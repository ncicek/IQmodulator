// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.11.3.469
// Netlist written on Sun Feb 07 01:50:57 2021
//
// Verilog Description of module top
//

module top (i_ref_clk, i_wbu_uart_rx, o_wbu_uart_tx, i_sw0, i_sw1, 
            o_dac_a, o_dac_b, dac_clk_p, dac_clk_n, o_dac_cw_b, i_clk_p, 
            i_clk_n, q_clk_p, q_clk_n) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(4[8:11])
    input i_ref_clk;   // d:/documents/git_local/fm_modulator/rtl/top.v(26[12:21])
    input i_wbu_uart_rx;   // d:/documents/git_local/fm_modulator/rtl/top.v(28[12:25])
    output o_wbu_uart_tx;   // d:/documents/git_local/fm_modulator/rtl/top.v(29[13:26])
    input i_sw0;   // d:/documents/git_local/fm_modulator/rtl/top.v(31[12:17])
    input i_sw1;   // d:/documents/git_local/fm_modulator/rtl/top.v(31[19:24])
    output [9:0]o_dac_a;   // d:/documents/git_local/fm_modulator/rtl/top.v(33[38:45])
    output [9:0]o_dac_b;   // d:/documents/git_local/fm_modulator/rtl/top.v(33[47:54])
    output dac_clk_p;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[49:58])
    output dac_clk_n;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[60:69])
    output o_dac_cw_b;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[71:81])
    output i_clk_p;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[13:20])
    output i_clk_n;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[22:29])
    output q_clk_p;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[31:38])
    output q_clk_n;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[40:47])
    
    wire i_ref_clk_c /* synthesis is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(26[12:21])
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[49:58])
    wire lo_pll_out /* synthesis is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(166[6:16])
    wire o_dac_b_c_15 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire o_dac_b_c_14 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire o_dac_b_c_13 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire o_dac_b_c_12 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire o_dac_b_c_11 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire o_dac_b_c_10 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire n3639 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire o_dac_b_c_8 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire o_dac_b_c_7 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire i_clk_2f_N_2268 /* synthesis is_inv_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/clock_phase_shifter.v(11[21:28])
    
    wire GND_net, VCC_net, i_wbu_uart_rx_c, o_wbu_uart_tx_c, i_sw0_c, 
        o_dac_a_c_9, o_dac_a_c_7, o_dac_a_c_6, o_dac_a_c_5, o_dac_a_c_4, 
        o_dac_a_c_3, o_dac_a_c_2, o_dac_a_c_1, o_dac_a_c_0, o_dac_b_c_9, 
        i_clk_p_c, q_clk_p_c, dac_clk_n_c, o_dac_cw_b_c, rx_stb;
    wire [7:0]rx_data;   // d:/documents/git_local/fm_modulator/rtl/top.v(61[12:19])
    
    wire tx_busy, wb_cyc, wb_stb, wb_we;
    wire [29:0]wb_addr;   // d:/documents/git_local/fm_modulator/rtl/top.v(78[13:20])
    wire [31:0]wb_odata;   // d:/documents/git_local/fm_modulator/rtl/top.v(79[13:21])
    
    wire wb_ack, wb_err;
    wire [31:0]wb_idata;   // d:/documents/git_local/fm_modulator/rtl/top.v(84[12:20])
    wire [29:0]bus_err_address;   // d:/documents/git_local/fm_modulator/rtl/top.v(108[12:27])
    
    wire wb_fm_ack;
    wire [31:0]wb_fm_data;   // d:/documents/git_local/fm_modulator/rtl/top.v(112[13:23])
    wire [31:0]wb_smpl_data;   // d:/documents/git_local/fm_modulator/rtl/top.v(115[12:24])
    
    wire wb_smpl_ack;
    wire [7:0]wb_lo_data;   // d:/documents/git_local/fm_modulator/rtl/top.v(144[12:22])
    
    wire wb_lo_ack, pll_clk, pll_rst, pll_stb, pll_we, pll_ack;
    wire [7:0]pll_data_i;   // d:/documents/git_local/fm_modulator/rtl/top.v(150[12:22])
    wire [7:0]pll_data_o;   // d:/documents/git_local/fm_modulator/rtl/top.v(150[24:34])
    wire [4:0]pll_addr;   // d:/documents/git_local/fm_modulator/rtl/top.v(151[12:20])
    wire [31:0]smpl_register;   // d:/documents/git_local/fm_modulator/rtl/top.v(210[13:26])
    wire [31:0]power_counter;   // d:/documents/git_local/fm_modulator/rtl/top.v(210[28:41])
    
    wire smpl_interrupt, none_sel, o_dac_a_9__N_1, wb_lo_data_7__N_96, 
        n21078, n7;
    wire [31:0]wb_smpl_data_31__N_64;
    wire [31:0]power_counter_31__N_232;
    wire [30:0]power_counter_31__N_201;
    wire [31:0]power_counter_31__N_129;
    
    wire wb_smpl_sel_N_310, wb_lo_sel_N_312;
    wire [31:0]wb_idata_31__N_266;
    wire [31:0]wb_idata_31__N_2;
    wire [23:0]chg_counter;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(97[17:28])
    
    wire chg_counter_23__N_405;
    wire [3:0]state_adj_3094;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(83[12:17])
    wire [7:0]lcl_data;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(84[12:20])
    
    wire zero_baud_counter, o_busy_N_535;
    wire [7:0]lcl_data_7__N_510;
    
    wire n2116, n2115, n27051, n2112, n2111, n2110, n2109, n2108, 
        n27058, n27059, n2104, n2102, n21592, n21586, n21590, 
        n17849, i_clk_n_c, q_clk_n_c, dac_clk_p_c_enable_297, n21102, 
        n2101, n2100, n2099, n2098, n17855, n17872, n17854, n21096, 
        n2117, n27380, n2, n2097, n2096, n2095, n27057, n2093, 
        n2092, n27050, n2119, n2120, n2121, n2122, dac_clk_p_c_enable_199, 
        n17860, n17871, n17853, n17847, n21088, n17870, n21546, 
        n17852, n17869, n17851, n17868, n27056, n27313, n17850, 
        n27304, n21044, n17867, n38, n17848, n34, n17866, n21032, 
        n17846, n21396, n21026, n18134, n27281, n10106, dac_clk_p_c_enable_224, 
        n17865, n17858, n21344, n21326, n4, n21320, n17845, n21540, 
        n4_adj_3041, n17864, n17857, n27184, n12753, n21248, n17863, 
        n17843, n17842, n27061, n27049, n17862, n17859, n17844, 
        n17861, dac_clk_p_c_enable_346, n21190, n21584, n27140, n21188, 
        n21186, n21176, n2_adj_3042, n1, n2_adj_3043, n1_adj_3044, 
        n2_adj_3045, n2_adj_3046, n1_adj_3047, n2_adj_3048, n1_adj_3049, 
        n2_adj_3050, n29969, n1_adj_3051, n2_adj_3052, n1_adj_3053, 
        n2_adj_3054, n1_adj_3055, n2_adj_3056, n1_adj_3057, n2_adj_3058, 
        n1_adj_3059, n2_adj_3060, n1_adj_3061, n2_adj_3062, n2_adj_3063, 
        n1_adj_3064, n2_adj_3065, n2_adj_3066, n2_adj_3067, n2_adj_3068, 
        n1_adj_3069, n2_adj_3070, n1_adj_3071, n2_adj_3072, n1_adj_3073, 
        n2_adj_3074, n1_adj_3075, n2_adj_3076, n21562, n1_adj_3077, 
        n2_adj_3078, n2_adj_3079, n2_adj_3080, n1_adj_3081, n2_adj_3082, 
        n1_adj_3083, n2_adj_3084, n1_adj_3085, n2_adj_3086, n2_adj_3087, 
        n1_adj_3088, n2_adj_3089, n1_adj_3090, n2_adj_3091, n1_adj_3092, 
        n17856, n27114, n27444, n21604, n21560, n21600, n29968;
    
    VHI i2 (.Z(VCC_net));
    GSR GSR_INST (.GSR(i_sw0_c)) /* synthesis syn_instantiated=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(41[6:29])
    LUT4 mux_434_Mux_22_i2_3_lut (.A(bus_err_address[20]), .B(power_counter[22]), 
         .C(wb_addr[0]), .Z(n2_adj_3058)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(228[3] 235[10])
    defparam mux_434_Mux_22_i2_3_lut.init = 16'hcaca;
    hbbus genbus (.dac_clk_p_c(dac_clk_p_c), .wb_cyc(wb_cyc), .wb_odata({wb_odata}), 
          .wb_we(wb_we), .wb_stb(wb_stb), .wb_err(wb_err), .wb_ack(wb_ack), 
          .\wb_idata[0] (wb_idata[0]), .wb_addr({wb_addr}), .\wb_idata[2] (wb_idata[2]), 
          .\wb_idata[3] (wb_idata[3]), .\wb_idata[4] (wb_idata[4]), .\wb_idata[5] (wb_idata[5]), 
          .\wb_idata[6] (wb_idata[6]), .\wb_idata[7] (wb_idata[7]), .\wb_idata[8] (wb_idata[8]), 
          .\wb_idata[9] (wb_idata[9]), .\wb_idata[10] (wb_idata[10]), .\wb_idata[11] (wb_idata[11]), 
          .\wb_idata[12] (wb_idata[12]), .\wb_idata[13] (wb_idata[13]), 
          .\wb_idata[14] (wb_idata[14]), .\wb_idata[15] (wb_idata[15]), 
          .\wb_idata[16] (wb_idata[16]), .\wb_idata[17] (wb_idata[17]), 
          .\wb_idata[18] (wb_idata[18]), .\wb_idata[19] (wb_idata[19]), 
          .\wb_idata[20] (wb_idata[20]), .\wb_idata[21] (wb_idata[21]), 
          .\wb_idata[22] (wb_idata[22]), .\wb_idata[23] (wb_idata[23]), 
          .\wb_idata[24] (wb_idata[24]), .\wb_idata[25] (wb_idata[25]), 
          .\wb_idata[26] (wb_idata[26]), .\wb_idata[27] (wb_idata[27]), 
          .\wb_idata[28] (wb_idata[28]), .\wb_idata[29] (wb_idata[29]), 
          .\wb_idata[30] (wb_idata[30]), .\wb_idata[31] (wb_idata[31]), 
          .n2(n2), .GND_net(GND_net), .n12753(n12753), .n29969(n29969), 
          .VCC_net(VCC_net), .rx_stb(rx_stb), .\rx_data[3] (rx_data[3]), 
          .\rx_data[6] (rx_data[6]), .\rx_data[2] (rx_data[2]), .\rx_data[4] (rx_data[4]), 
          .\rx_data[5] (rx_data[5]), .\rx_data[0] (rx_data[0]), .\rx_data[1] (rx_data[1]), 
          .tx_busy(tx_busy), .n27281(n27281), .\lcl_data[1] (lcl_data[1]), 
          .\lcl_data_7__N_510[0] (lcl_data_7__N_510[0]), .zero_baud_counter(zero_baud_counter), 
          .dac_clk_p_c_enable_346(dac_clk_p_c_enable_346), .\lcl_data[4] (lcl_data[4]), 
          .\lcl_data_7__N_510[3] (lcl_data_7__N_510[3]), .\lcl_data[7] (lcl_data[7]), 
          .\lcl_data_7__N_510[6] (lcl_data_7__N_510[6]), .\lcl_data[6] (lcl_data[6]), 
          .\lcl_data_7__N_510[5] (lcl_data_7__N_510[5]), .\lcl_data[5] (lcl_data[5]), 
          .\lcl_data_7__N_510[4] (lcl_data_7__N_510[4]), .\lcl_data[3] (lcl_data[3]), 
          .\lcl_data_7__N_510[2] (lcl_data_7__N_510[2]), .\lcl_data[2] (lcl_data[2]), 
          .\lcl_data_7__N_510[1] (lcl_data_7__N_510[1]), .o_busy_N_535(o_busy_N_535), 
          .\state[0] (state_adj_3094[0]), .n18134(n18134)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(87[7] 103[22])
    FD1S3AX power_counter_i0 (.D(power_counter_31__N_129[0]), .CK(dac_clk_p_c), 
            .Q(power_counter[0])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(239[9] 244[54])
    defparam power_counter_i0.GSR = "DISABLED";
    FD1S3AX wb_idata_i0 (.D(wb_idata_31__N_2[0]), .CK(dac_clk_p_c), .Q(wb_idata[0]));   // d:/documents/git_local/fm_modulator/rtl/top.v(280[9] 288[53])
    defparam wb_idata_i0.GSR = "DISABLED";
    FD1S3JX wb_ack_67 (.D(n4), .CK(dac_clk_p_c), .PD(wb_smpl_ack), .Q(wb_ack)) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(277[9] 278[57])
    defparam wb_ack_67.GSR = "DISABLED";
    FD1S3IX wb_smpl_ack_60 (.D(wb_stb), .CK(dac_clk_p_c), .CD(wb_smpl_sel_N_310), 
            .Q(wb_smpl_ack)) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(213[9] 214[44])
    defparam wb_smpl_ack_60.GSR = "DISABLED";
    \rxuartlite(CLOCKS_PER_BAUD=10000)  rxtransport (.\rx_data[0] (rx_data[0]), 
            .dac_clk_p_c(dac_clk_p_c), .rx_stb(rx_stb), .i_wbu_uart_rx_c(i_wbu_uart_rx_c), 
            .chg_counter({chg_counter}), .dac_clk_p_c_enable_199(dac_clk_p_c_enable_199), 
            .chg_counter_23__N_405(chg_counter_23__N_405), .GND_net(GND_net), 
            .\rx_data[6] (rx_data[6]), .\rx_data[5] (rx_data[5]), .\rx_data[4] (rx_data[4]), 
            .\rx_data[3] (rx_data[3]), .\rx_data[2] (rx_data[2]), .\rx_data[1] (rx_data[1])) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(63[57:105])
    PUR PUR_INST (.PUR(i_sw0_c)) /* synthesis syn_instantiated=1 */ ;
    defparam PUR_INST.RST_PULSE = 1;
    OB o_dac_a_pad_7 (.I(o_dac_a_c_7), .O(o_dac_a[7]));   // d:/documents/git_local/fm_modulator/rtl/top.v(33[38:45])
    \txuartlite(TIMING_BITS=24,CLOCKS_PER_BAUD=10000)  txtransport (.n27281(n27281), 
            .state({Open_0, Open_1, Open_2, state_adj_3094[0]}), .dac_clk_p_c(dac_clk_p_c), 
            .dac_clk_p_c_enable_346(dac_clk_p_c_enable_346), .\lcl_data_7__N_510[0] (lcl_data_7__N_510[0]), 
            .zero_baud_counter(zero_baud_counter), .o_wbu_uart_tx_c(o_wbu_uart_tx_c), 
            .\lcl_data[7] (lcl_data[7]), .n29969(n29969), .GND_net(GND_net), 
            .\lcl_data[6] (lcl_data[6]), .\lcl_data_7__N_510[6] (lcl_data_7__N_510[6]), 
            .\lcl_data[5] (lcl_data[5]), .\lcl_data_7__N_510[5] (lcl_data_7__N_510[5]), 
            .\lcl_data[4] (lcl_data[4]), .\lcl_data_7__N_510[4] (lcl_data_7__N_510[4]), 
            .\lcl_data[3] (lcl_data[3]), .\lcl_data_7__N_510[3] (lcl_data_7__N_510[3]), 
            .\lcl_data[2] (lcl_data[2]), .\lcl_data_7__N_510[2] (lcl_data_7__N_510[2]), 
            .\lcl_data[1] (lcl_data[1]), .\lcl_data_7__N_510[1] (lcl_data_7__N_510[1]), 
            .o_busy_N_535(o_busy_N_535), .tx_busy(tx_busy), .n18134(n18134)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(72[58:115])
    FD1P3AX smpl_register_i0_i0 (.D(wb_odata[0]), .SP(dac_clk_p_c_enable_297), 
            .CK(dac_clk_p_c), .Q(smpl_register[0]));   // d:/documents/git_local/fm_modulator/rtl/top.v(217[9] 225[6])
    defparam smpl_register_i0_i0.GSR = "DISABLED";
    FD1S3IX wb_err_65 (.D(none_sel), .CK(dac_clk_p_c), .CD(n2), .Q(wb_err));   // d:/documents/git_local/fm_modulator/rtl/top.v(266[9] 267[34])
    defparam wb_err_65.GSR = "DISABLED";
    PFUMX mux_434_Mux_3_i3 (.BLUT(n1_adj_3090), .ALUT(n2_adj_3089), .C0(wb_addr[1]), 
          .Z(n2120));
    OB o_dac_a_pad_8 (.I(n27380), .O(o_dac_a[8]));   // d:/documents/git_local/fm_modulator/rtl/top.v(33[38:45])
    OB o_dac_a_pad_9 (.I(o_dac_a_c_9), .O(o_dac_a[9]));   // d:/documents/git_local/fm_modulator/rtl/top.v(33[38:45])
    FD1P3AX bus_err_address_i0_i0 (.D(wb_addr[0]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[0])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[9] 272[31])
    defparam bus_err_address_i0_i0.GSR = "DISABLED";
    OB o_wbu_uart_tx_pad (.I(o_wbu_uart_tx_c), .O(o_wbu_uart_tx));   // d:/documents/git_local/fm_modulator/rtl/top.v(29[13:26])
    LUT4 mux_434_Mux_2_i2_3_lut (.A(bus_err_address[0]), .B(power_counter[2]), 
         .C(wb_addr[0]), .Z(n2_adj_3091)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(228[3] 235[10])
    defparam mux_434_Mux_2_i2_3_lut.init = 16'hcaca;
    CCU2D add_31_27 (.A0(power_counter[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17854), .COUT(n17855), .S0(power_counter_31__N_232[25]), 
          .S1(power_counter_31__N_232[26]));   // d:/documents/git_local/fm_modulator/rtl/top.v(242[21:41])
    defparam add_31_27.INIT0 = 16'h5aaa;
    defparam add_31_27.INIT1 = 16'h5aaa;
    defparam add_31_27.INJECT1_0 = "NO";
    defparam add_31_27.INJECT1_1 = "NO";
    PFUMX mux_434_Mux_23_i3 (.BLUT(n1_adj_3057), .ALUT(n2_adj_3056), .C0(wb_addr[1]), 
          .Z(n2100));
    LUT4 o_clk_q_I_0_1_lut (.A(q_clk_p_c), .Z(q_clk_n_c)) /* synthesis lut_function=(!(A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/clock_phase_shifter.v(18[16:24])
    defparam o_clk_q_I_0_1_lut.init = 16'h5555;
    LUT4 mux_434_Mux_26_i2_3_lut (.A(bus_err_address[24]), .B(power_counter[26]), 
         .C(wb_addr[0]), .Z(n2_adj_3050)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(228[3] 235[10])
    defparam mux_434_Mux_26_i2_3_lut.init = 16'hcaca;
    PFUMX mux_434_Mux_24_i3 (.BLUT(n1_adj_3055), .ALUT(n2_adj_3054), .C0(wb_addr[1]), 
          .Z(n2099));
    PFUMX mux_434_Mux_4_i3 (.BLUT(n1_adj_3088), .ALUT(n2_adj_3087), .C0(wb_addr[1]), 
          .Z(n2119));
    FD1P3AX smpl_interrupt_62 (.D(wb_odata[0]), .SP(dac_clk_p_c_enable_224), 
            .CK(dac_clk_p_c), .Q(smpl_interrupt)) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(217[9] 225[6])
    defparam smpl_interrupt_62.GSR = "DISABLED";
    LUT4 o_clk_i_I_0_1_lut (.A(i_clk_p_c), .Z(i_clk_n_c)) /* synthesis lut_function=(!(A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/clock_phase_shifter.v(14[16:24])
    defparam o_clk_i_I_0_1_lut.init = 16'h5555;
    PFUMX mux_434_Mux_6_i3 (.BLUT(n1_adj_3085), .ALUT(n2_adj_3084), .C0(wb_addr[1]), 
          .Z(n2117));
    PFUMX mux_434_Mux_7_i3 (.BLUT(n1_adj_3083), .ALUT(n2_adj_3082), .C0(wb_addr[1]), 
          .Z(n2116));
    LUT4 i1_2_lut_rep_475_3_lut (.A(wb_addr[12]), .B(wb_addr[8]), .C(wb_addr[1]), 
         .Z(n27140)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(256[23:49])
    defparam i1_2_lut_rep_475_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_3_lut_4_lut (.A(wb_addr[12]), .B(wb_addr[8]), .C(n27313), 
         .D(wb_addr[1]), .Z(n21078)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(256[23:49])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 wb_cyc_I_0_2_lut (.A(wb_cyc), .B(wb_lo_sel_N_312), .Z(wb_lo_data_7__N_96)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(191[13:36])
    defparam wb_cyc_I_0_2_lut.init = 16'h2222;
    LUT4 i1_4_lut (.A(n27184), .B(n21248), .C(wb_addr[9]), .D(wb_addr[8]), 
         .Z(wb_lo_sel_N_312)) /* synthesis lut_function=(A+(B+!(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(256[23:49])
    defparam i1_4_lut.init = 16'hefff;
    LUT4 i1_4_lut_adj_145 (.A(n38), .B(n4_adj_3041), .C(n21540), .D(n21032), 
         .Z(dac_clk_p_c_enable_297)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut_adj_145.init = 16'h0100;
    LUT4 i1_4_lut_adj_146 (.A(n27313), .B(n21026), .C(wb_addr[1]), .D(wb_addr[12]), 
         .Z(n21032)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_4_lut_adj_146.init = 16'h0004;
    LUT4 i1_3_lut_4_lut (.A(wb_addr[12]), .B(wb_addr[8]), .C(wb_addr[0]), 
         .D(n27313), .Z(n21044)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(256[23:49])
    defparam i1_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_3_lut_4_lut_adj_147 (.A(wb_addr[12]), .B(wb_addr[8]), .C(wb_addr[15]), 
         .D(n27313), .Z(n21344)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(256[23:49])
    defparam i1_3_lut_4_lut_adj_147.init = 16'hffef;
    PFUMX mux_434_Mux_8_i3 (.BLUT(n1_adj_3081), .ALUT(n2_adj_3080), .C0(wb_addr[1]), 
          .Z(n2115));
    PFUMX mux_434_Mux_2_i3 (.BLUT(n1_adj_3092), .ALUT(n2_adj_3091), .C0(wb_addr[1]), 
          .Z(n2121));
    PFUMX mux_434_Mux_25_i3 (.BLUT(n1_adj_3053), .ALUT(n2_adj_3052), .C0(wb_addr[1]), 
          .Z(n2098));
    LUT4 i18010_2_lut_rep_779 (.A(wb_addr[2]), .B(wb_addr[3]), .Z(n27444)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i18010_2_lut_rep_779.init = 16'heeee;
    LUT4 i19260_2_lut_3_lut (.A(wb_addr[2]), .B(wb_addr[3]), .C(n34), 
         .Z(n21540)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i19260_2_lut_3_lut.init = 16'hfefe;
    FD1P3AX smpl_register_i0_i31 (.D(wb_odata[31]), .SP(dac_clk_p_c_enable_297), 
            .CK(dac_clk_p_c), .Q(smpl_register[31]));   // d:/documents/git_local/fm_modulator/rtl/top.v(217[9] 225[6])
    defparam smpl_register_i0_i31.GSR = "DISABLED";
    LUT4 power_counter_31__I_0_74_i1_3_lut (.A(power_counter_31__N_232[0]), 
         .B(power_counter_31__N_201[0]), .C(power_counter[31]), .Z(power_counter_31__N_129[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[4:54])
    defparam power_counter_31__I_0_74_i1_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_148 (.A(wb_lo_sel_N_312), .B(wb_smpl_sel_N_310), .C(n27114), 
         .D(n21344), .Z(none_sel)) /* synthesis lut_function=(A (B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(262[20:68])
    defparam i1_4_lut_adj_148.init = 16'h8880;
    LUT4 i1_4_lut_adj_149 (.A(n21586), .B(n21604), .C(n21600), .D(chg_counter_23__N_405), 
         .Z(dac_clk_p_c_enable_199)) /* synthesis lut_function=((((D)+!C)+!B)+!A) */ ;
    defparam i1_4_lut_adj_149.init = 16'hff7f;
    LUT4 i19306_4_lut (.A(chg_counter[15]), .B(chg_counter[17]), .C(chg_counter[10]), 
         .D(chg_counter[9]), .Z(n21586)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i19306_4_lut.init = 16'h8000;
    LUT4 i19324_4_lut (.A(n21560), .B(n21592), .C(n21590), .D(n21562), 
         .Z(n21604)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i19324_4_lut.init = 16'h8000;
    LUT4 i19320_4_lut (.A(chg_counter[2]), .B(n21584), .C(n21546), .D(chg_counter[3]), 
         .Z(n21600)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i19320_4_lut.init = 16'h8000;
    LUT4 i19280_2_lut (.A(chg_counter[5]), .B(chg_counter[7]), .Z(n21560)) /* synthesis lut_function=(A (B)) */ ;
    defparam i19280_2_lut.init = 16'h8888;
    FD1P3AX smpl_register_i0_i30 (.D(wb_odata[30]), .SP(dac_clk_p_c_enable_297), 
            .CK(dac_clk_p_c), .Q(smpl_register[30]));   // d:/documents/git_local/fm_modulator/rtl/top.v(217[9] 225[6])
    defparam smpl_register_i0_i30.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i29 (.D(wb_odata[29]), .SP(dac_clk_p_c_enable_297), 
            .CK(dac_clk_p_c), .Q(smpl_register[29]));   // d:/documents/git_local/fm_modulator/rtl/top.v(217[9] 225[6])
    defparam smpl_register_i0_i29.GSR = "DISABLED";
    LUT4 i19312_4_lut (.A(chg_counter[20]), .B(chg_counter[22]), .C(chg_counter[16]), 
         .D(chg_counter[4]), .Z(n21592)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i19312_4_lut.init = 16'h8000;
    FD1P3AX smpl_register_i0_i28 (.D(wb_odata[28]), .SP(dac_clk_p_c_enable_297), 
            .CK(dac_clk_p_c), .Q(smpl_register[28]));   // d:/documents/git_local/fm_modulator/rtl/top.v(217[9] 225[6])
    defparam smpl_register_i0_i28.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i27 (.D(wb_odata[27]), .SP(dac_clk_p_c_enable_297), 
            .CK(dac_clk_p_c), .Q(smpl_register[27]));   // d:/documents/git_local/fm_modulator/rtl/top.v(217[9] 225[6])
    defparam smpl_register_i0_i27.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i26 (.D(wb_odata[26]), .SP(dac_clk_p_c_enable_297), 
            .CK(dac_clk_p_c), .Q(smpl_register[26]));   // d:/documents/git_local/fm_modulator/rtl/top.v(217[9] 225[6])
    defparam smpl_register_i0_i26.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i25 (.D(wb_odata[25]), .SP(dac_clk_p_c_enable_297), 
            .CK(dac_clk_p_c), .Q(smpl_register[25]));   // d:/documents/git_local/fm_modulator/rtl/top.v(217[9] 225[6])
    defparam smpl_register_i0_i25.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i24 (.D(wb_odata[24]), .SP(dac_clk_p_c_enable_297), 
            .CK(dac_clk_p_c), .Q(smpl_register[24]));   // d:/documents/git_local/fm_modulator/rtl/top.v(217[9] 225[6])
    defparam smpl_register_i0_i24.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i23 (.D(wb_odata[23]), .SP(dac_clk_p_c_enable_297), 
            .CK(dac_clk_p_c), .Q(smpl_register[23]));   // d:/documents/git_local/fm_modulator/rtl/top.v(217[9] 225[6])
    defparam smpl_register_i0_i23.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i22 (.D(wb_odata[22]), .SP(dac_clk_p_c_enable_297), 
            .CK(dac_clk_p_c), .Q(smpl_register[22]));   // d:/documents/git_local/fm_modulator/rtl/top.v(217[9] 225[6])
    defparam smpl_register_i0_i22.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i21 (.D(wb_odata[21]), .SP(dac_clk_p_c_enable_297), 
            .CK(dac_clk_p_c), .Q(smpl_register[21]));   // d:/documents/git_local/fm_modulator/rtl/top.v(217[9] 225[6])
    defparam smpl_register_i0_i21.GSR = "DISABLED";
    LUT4 i19310_4_lut (.A(chg_counter[18]), .B(chg_counter[8]), .C(chg_counter[1]), 
         .D(chg_counter[23]), .Z(n21590)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i19310_4_lut.init = 16'h8000;
    FD1P3AX smpl_register_i0_i20 (.D(wb_odata[20]), .SP(dac_clk_p_c_enable_297), 
            .CK(dac_clk_p_c), .Q(smpl_register[20]));   // d:/documents/git_local/fm_modulator/rtl/top.v(217[9] 225[6])
    defparam smpl_register_i0_i20.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i19 (.D(wb_odata[19]), .SP(dac_clk_p_c_enable_297), 
            .CK(dac_clk_p_c), .Q(smpl_register[19]));   // d:/documents/git_local/fm_modulator/rtl/top.v(217[9] 225[6])
    defparam smpl_register_i0_i19.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i18 (.D(wb_odata[18]), .SP(dac_clk_p_c_enable_297), 
            .CK(dac_clk_p_c), .Q(smpl_register[18]));   // d:/documents/git_local/fm_modulator/rtl/top.v(217[9] 225[6])
    defparam smpl_register_i0_i18.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i17 (.D(wb_odata[17]), .SP(dac_clk_p_c_enable_297), 
            .CK(dac_clk_p_c), .Q(smpl_register[17]));   // d:/documents/git_local/fm_modulator/rtl/top.v(217[9] 225[6])
    defparam smpl_register_i0_i17.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i16 (.D(wb_odata[16]), .SP(dac_clk_p_c_enable_297), 
            .CK(dac_clk_p_c), .Q(smpl_register[16]));   // d:/documents/git_local/fm_modulator/rtl/top.v(217[9] 225[6])
    defparam smpl_register_i0_i16.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i15 (.D(wb_odata[15]), .SP(dac_clk_p_c_enable_297), 
            .CK(dac_clk_p_c), .Q(smpl_register[15]));   // d:/documents/git_local/fm_modulator/rtl/top.v(217[9] 225[6])
    defparam smpl_register_i0_i15.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i14 (.D(wb_odata[14]), .SP(dac_clk_p_c_enable_297), 
            .CK(dac_clk_p_c), .Q(smpl_register[14]));   // d:/documents/git_local/fm_modulator/rtl/top.v(217[9] 225[6])
    defparam smpl_register_i0_i14.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i13 (.D(wb_odata[13]), .SP(dac_clk_p_c_enable_297), 
            .CK(dac_clk_p_c), .Q(smpl_register[13]));   // d:/documents/git_local/fm_modulator/rtl/top.v(217[9] 225[6])
    defparam smpl_register_i0_i13.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i12 (.D(wb_odata[12]), .SP(dac_clk_p_c_enable_297), 
            .CK(dac_clk_p_c), .Q(smpl_register[12]));   // d:/documents/git_local/fm_modulator/rtl/top.v(217[9] 225[6])
    defparam smpl_register_i0_i12.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i11 (.D(wb_odata[11]), .SP(dac_clk_p_c_enable_297), 
            .CK(dac_clk_p_c), .Q(smpl_register[11]));   // d:/documents/git_local/fm_modulator/rtl/top.v(217[9] 225[6])
    defparam smpl_register_i0_i11.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i10 (.D(wb_odata[10]), .SP(dac_clk_p_c_enable_297), 
            .CK(dac_clk_p_c), .Q(smpl_register[10]));   // d:/documents/git_local/fm_modulator/rtl/top.v(217[9] 225[6])
    defparam smpl_register_i0_i10.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i9 (.D(wb_odata[9]), .SP(dac_clk_p_c_enable_297), 
            .CK(dac_clk_p_c), .Q(smpl_register[9]));   // d:/documents/git_local/fm_modulator/rtl/top.v(217[9] 225[6])
    defparam smpl_register_i0_i9.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i8 (.D(wb_odata[8]), .SP(dac_clk_p_c_enable_297), 
            .CK(dac_clk_p_c), .Q(smpl_register[8]));   // d:/documents/git_local/fm_modulator/rtl/top.v(217[9] 225[6])
    defparam smpl_register_i0_i8.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i7 (.D(wb_odata[7]), .SP(dac_clk_p_c_enable_297), 
            .CK(dac_clk_p_c), .Q(smpl_register[7]));   // d:/documents/git_local/fm_modulator/rtl/top.v(217[9] 225[6])
    defparam smpl_register_i0_i7.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i6 (.D(wb_odata[6]), .SP(dac_clk_p_c_enable_297), 
            .CK(dac_clk_p_c), .Q(smpl_register[6]));   // d:/documents/git_local/fm_modulator/rtl/top.v(217[9] 225[6])
    defparam smpl_register_i0_i6.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i5 (.D(wb_odata[5]), .SP(dac_clk_p_c_enable_297), 
            .CK(dac_clk_p_c), .Q(smpl_register[5]));   // d:/documents/git_local/fm_modulator/rtl/top.v(217[9] 225[6])
    defparam smpl_register_i0_i5.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i4 (.D(wb_odata[4]), .SP(dac_clk_p_c_enable_297), 
            .CK(dac_clk_p_c), .Q(smpl_register[4]));   // d:/documents/git_local/fm_modulator/rtl/top.v(217[9] 225[6])
    defparam smpl_register_i0_i4.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i3 (.D(wb_odata[3]), .SP(dac_clk_p_c_enable_297), 
            .CK(dac_clk_p_c), .Q(smpl_register[3]));   // d:/documents/git_local/fm_modulator/rtl/top.v(217[9] 225[6])
    defparam smpl_register_i0_i3.GSR = "DISABLED";
    LUT4 i11436_2_lut (.A(smpl_register[26]), .B(wb_addr[0]), .Z(n1_adj_3051)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(228[3] 235[10])
    defparam i11436_2_lut.init = 16'h8888;
    LUT4 i19282_2_lut (.A(chg_counter[12]), .B(chg_counter[14]), .Z(n21562)) /* synthesis lut_function=(A (B)) */ ;
    defparam i19282_2_lut.init = 16'h8888;
    LUT4 i19304_4_lut (.A(chg_counter[19]), .B(chg_counter[13]), .C(chg_counter[21]), 
         .D(chg_counter[0]), .Z(n21584)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i19304_4_lut.init = 16'h8000;
    FD1P3AX smpl_register_i0_i2 (.D(wb_odata[2]), .SP(dac_clk_p_c_enable_297), 
            .CK(dac_clk_p_c), .Q(smpl_register[2]));   // d:/documents/git_local/fm_modulator/rtl/top.v(217[9] 225[6])
    defparam smpl_register_i0_i2.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i1 (.D(wb_odata[1]), .SP(dac_clk_p_c_enable_297), 
            .CK(dac_clk_p_c), .Q(smpl_register[1]));   // d:/documents/git_local/fm_modulator/rtl/top.v(217[9] 225[6])
    defparam smpl_register_i0_i1.GSR = "DISABLED";
    LUT4 i19266_2_lut (.A(chg_counter[6]), .B(chg_counter[11]), .Z(n21546)) /* synthesis lut_function=(A (B)) */ ;
    defparam i19266_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_150 (.A(n27313), .B(n38), .C(n34), .D(n21326), 
         .Z(o_dac_a_9__N_1)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut_adj_150.init = 16'h0100;
    LUT4 i1_4_lut_adj_151 (.A(wb_addr[12]), .B(wb_addr[8]), .C(n21320), 
         .D(wb_stb), .Z(n21326)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_4_lut_adj_151.init = 16'h1000;
    LUT4 i1_2_lut (.A(wb_addr[15]), .B(wb_addr[9]), .Z(n21320)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i11432_2_lut (.A(smpl_register[22]), .B(wb_addr[0]), .Z(n1_adj_3059)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(228[3] 235[10])
    defparam i11432_2_lut.init = 16'h8888;
    LUT4 mux_434_Mux_21_i2_3_lut (.A(bus_err_address[19]), .B(power_counter[21]), 
         .C(wb_addr[0]), .Z(n2_adj_3060)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(228[3] 235[10])
    defparam mux_434_Mux_21_i2_3_lut.init = 16'hcaca;
    PFUMX mux_434_Mux_26_i3 (.BLUT(n1_adj_3051), .ALUT(n2_adj_3050), .C0(wb_addr[1]), 
          .Z(n2097));
    LUT4 wb_idata_31__I_0_i1_3_lut (.A(wb_idata_31__N_266[0]), .B(wb_fm_data[0]), 
         .C(wb_fm_ack), .Z(wb_idata_31__N_2[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(283[8] 288[53])
    defparam wb_idata_31__I_0_i1_3_lut.init = 16'hcaca;
    LUT4 mux_56_i1_4_lut (.A(wb_lo_data[0]), .B(wb_smpl_data[0]), .C(wb_smpl_ack), 
         .D(wb_lo_ack), .Z(wb_idata_31__N_266[0])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(285[8] 288[53])
    defparam mux_56_i1_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i32_4_lut (.A(wb_smpl_data[31]), .B(wb_fm_data[31]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_2[31])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(283[8] 288[53])
    defparam wb_idata_31__I_0_i32_4_lut.init = 16'hcac0;
    LUT4 i11431_2_lut (.A(smpl_register[21]), .B(wb_addr[0]), .Z(n1_adj_3061)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(228[3] 235[10])
    defparam i11431_2_lut.init = 16'h8888;
    LUT4 mux_434_Mux_20_i2_3_lut (.A(bus_err_address[18]), .B(power_counter[20]), 
         .C(wb_addr[0]), .Z(n2_adj_3062)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(228[3] 235[10])
    defparam mux_434_Mux_20_i2_3_lut.init = 16'hcaca;
    LUT4 mux_434_Mux_19_i2_3_lut (.A(bus_err_address[17]), .B(power_counter[19]), 
         .C(wb_addr[0]), .Z(n2_adj_3063)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(228[3] 235[10])
    defparam mux_434_Mux_19_i2_3_lut.init = 16'hcaca;
    LUT4 i11429_2_lut (.A(smpl_register[19]), .B(wb_addr[0]), .Z(n1_adj_3064)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(228[3] 235[10])
    defparam i11429_2_lut.init = 16'h8888;
    LUT4 mux_434_Mux_18_i2_3_lut (.A(bus_err_address[16]), .B(power_counter[18]), 
         .C(wb_addr[0]), .Z(n2_adj_3065)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(228[3] 235[10])
    defparam mux_434_Mux_18_i2_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_152 (.A(wb_fm_ack), .B(wb_lo_ack), .Z(n4)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(278[13:56])
    defparam i1_2_lut_adj_152.init = 16'heeee;
    LUT4 mux_434_Mux_17_i2_3_lut (.A(bus_err_address[15]), .B(power_counter[17]), 
         .C(wb_addr[0]), .Z(n2_adj_3066)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(228[3] 235[10])
    defparam mux_434_Mux_17_i2_3_lut.init = 16'hcaca;
    LUT4 mux_434_Mux_16_i2_3_lut (.A(bus_err_address[14]), .B(power_counter[16]), 
         .C(wb_addr[0]), .Z(n2_adj_3067)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(228[3] 235[10])
    defparam mux_434_Mux_16_i2_3_lut.init = 16'hcaca;
    PFUMX mux_434_Mux_27_i3 (.BLUT(n1_adj_3049), .ALUT(n2_adj_3048), .C0(wb_addr[1]), 
          .Z(n2096));
    LUT4 i1_2_lut_adj_153 (.A(wb_addr[9]), .B(wb_addr[8]), .Z(n4_adj_3041)) /* synthesis lut_function=(A+!(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(256[23:49])
    defparam i1_2_lut_adj_153.init = 16'hbbbb;
    LUT4 i1_4_lut_adj_154 (.A(wb_addr[28]), .B(wb_addr[19]), .C(wb_addr[13]), 
         .D(wb_addr[29]), .Z(n34)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(256[23:49])
    defparam i1_4_lut_adj_154.init = 16'hfffe;
    LUT4 i1_4_lut_adj_155 (.A(n21186), .B(n21188), .C(n21190), .D(n21176), 
         .Z(n38)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(256[23:49])
    defparam i1_4_lut_adj_155.init = 16'hfffe;
    LUT4 i1_2_lut_adj_156 (.A(wb_addr[11]), .B(wb_addr[16]), .Z(n21186)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(256[23:49])
    defparam i1_2_lut_adj_156.init = 16'heeee;
    LUT4 i1_4_lut_adj_157 (.A(wb_addr[17]), .B(wb_addr[14]), .C(wb_addr[23]), 
         .D(wb_addr[20]), .Z(n21188)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(256[23:49])
    defparam i1_4_lut_adj_157.init = 16'hfffe;
    LUT4 i1_4_lut_adj_158 (.A(wb_addr[25]), .B(wb_addr[10]), .C(wb_addr[26]), 
         .D(wb_addr[21]), .Z(n21190)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(256[23:49])
    defparam i1_4_lut_adj_158.init = 16'hfffe;
    LUT4 i1_2_lut_adj_159 (.A(wb_addr[27]), .B(wb_addr[18]), .Z(n21176)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(256[23:49])
    defparam i1_2_lut_adj_159.init = 16'heeee;
    LUT4 i1_4_lut_adj_160 (.A(wb_addr[1]), .B(wb_addr[2]), .C(wb_addr[0]), 
         .D(wb_addr[3]), .Z(n7)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(222[4:8])
    defparam i1_4_lut_adj_160.init = 16'hfffb;
    LUT4 i11412_2_lut (.A(smpl_register[2]), .B(wb_addr[0]), .Z(n1_adj_3092)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(228[3] 235[10])
    defparam i11412_2_lut.init = 16'h8888;
    LUT4 mux_434_Mux_15_i2_3_lut (.A(bus_err_address[13]), .B(power_counter[15]), 
         .C(wb_addr[0]), .Z(n2_adj_3068)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(228[3] 235[10])
    defparam mux_434_Mux_15_i2_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_519 (.A(wb_addr[15]), .B(n34), .Z(n27184)) /* synthesis lut_function=((B)+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(256[23:49])
    defparam i1_2_lut_rep_519.init = 16'hdddd;
    LUT4 i1_3_lut_4_lut_adj_161 (.A(wb_addr[15]), .B(n34), .C(n4_adj_3041), 
         .D(n21248), .Z(wb_smpl_sel_N_310)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(256[23:49])
    defparam i1_3_lut_4_lut_adj_161.init = 16'hfffd;
    LUT4 i11425_2_lut (.A(smpl_register[15]), .B(wb_addr[0]), .Z(n1_adj_3069)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(228[3] 235[10])
    defparam i11425_2_lut.init = 16'h8888;
    PFUMX mux_434_Mux_11_i3 (.BLUT(n1_adj_3077), .ALUT(n2_adj_3076), .C0(wb_addr[1]), 
          .Z(n2112));
    PFUMX mux_434_Mux_12_i3 (.BLUT(n1_adj_3075), .ALUT(n2_adj_3074), .C0(wb_addr[1]), 
          .Z(n2111));
    LUT4 mux_434_Mux_14_i2_3_lut (.A(bus_err_address[12]), .B(power_counter[14]), 
         .C(wb_addr[0]), .Z(n2_adj_3070)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(228[3] 235[10])
    defparam mux_434_Mux_14_i2_3_lut.init = 16'hcaca;
    LUT4 mux_434_Mux_31_i2_3_lut (.A(bus_err_address[29]), .B(power_counter[31]), 
         .C(wb_addr[0]), .Z(n2_adj_3042)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(228[3] 235[10])
    defparam mux_434_Mux_31_i2_3_lut.init = 16'hcaca;
    LUT4 i11424_2_lut (.A(smpl_register[14]), .B(wb_addr[0]), .Z(n1_adj_3071)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(228[3] 235[10])
    defparam i11424_2_lut.init = 16'h8888;
    LUT4 i11441_2_lut (.A(smpl_register[31]), .B(wb_addr[0]), .Z(n1)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(228[3] 235[10])
    defparam i11441_2_lut.init = 16'h8888;
    LUT4 mux_434_Mux_30_i2_3_lut (.A(bus_err_address[28]), .B(power_counter[30]), 
         .C(wb_addr[0]), .Z(n2_adj_3043)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(228[3] 235[10])
    defparam mux_434_Mux_30_i2_3_lut.init = 16'hcaca;
    LUT4 i11440_2_lut (.A(smpl_register[30]), .B(wb_addr[0]), .Z(n1_adj_3044)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(228[3] 235[10])
    defparam i11440_2_lut.init = 16'h8888;
    LUT4 mux_434_Mux_29_i2_3_lut (.A(bus_err_address[27]), .B(power_counter[29]), 
         .C(wb_addr[0]), .Z(n2_adj_3045)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(228[3] 235[10])
    defparam mux_434_Mux_29_i2_3_lut.init = 16'hcaca;
    LUT4 mux_434_Mux_13_i2_3_lut (.A(bus_err_address[11]), .B(power_counter[13]), 
         .C(wb_addr[0]), .Z(n2_adj_3072)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(228[3] 235[10])
    defparam mux_434_Mux_13_i2_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_rep_449 (.A(n34), .B(n38), .C(wb_addr[9]), .Z(n27114)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(256[23:49])
    defparam i1_3_lut_rep_449.init = 16'hefef;
    LUT4 i1_2_lut_4_lut (.A(n34), .B(n38), .C(wb_addr[9]), .D(n27304), 
         .Z(n21088)) /* synthesis lut_function=(A+(B+!(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(256[23:49])
    defparam i1_2_lut_4_lut.init = 16'hefff;
    LUT4 i11423_2_lut (.A(smpl_register[13]), .B(wb_addr[0]), .Z(n1_adj_3073)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(228[3] 235[10])
    defparam i11423_2_lut.init = 16'h8888;
    LUT4 mux_434_Mux_28_i2_3_lut (.A(bus_err_address[26]), .B(power_counter[28]), 
         .C(wb_addr[0]), .Z(n2_adj_3046)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(228[3] 235[10])
    defparam mux_434_Mux_28_i2_3_lut.init = 16'hcaca;
    LUT4 i11438_2_lut (.A(smpl_register[28]), .B(wb_addr[0]), .Z(n1_adj_3047)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(228[3] 235[10])
    defparam i11438_2_lut.init = 16'h8888;
    LUT4 mux_434_Mux_27_i2_3_lut (.A(bus_err_address[25]), .B(power_counter[27]), 
         .C(wb_addr[0]), .Z(n2_adj_3048)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(228[3] 235[10])
    defparam mux_434_Mux_27_i2_3_lut.init = 16'hcaca;
    LUT4 mux_434_Mux_12_i2_3_lut (.A(bus_err_address[10]), .B(power_counter[12]), 
         .C(wb_addr[0]), .Z(n2_adj_3074)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(228[3] 235[10])
    defparam mux_434_Mux_12_i2_3_lut.init = 16'hcaca;
    PFUMX mux_434_Mux_28_i3 (.BLUT(n1_adj_3047), .ALUT(n2_adj_3046), .C0(wb_addr[1]), 
          .Z(n2095));
    LUT4 i11437_2_lut (.A(smpl_register[27]), .B(wb_addr[0]), .Z(n1_adj_3049)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(228[3] 235[10])
    defparam i11437_2_lut.init = 16'h8888;
    PFUMX mux_434_Mux_13_i3 (.BLUT(n1_adj_3073), .ALUT(n2_adj_3072), .C0(wb_addr[1]), 
          .Z(n2110));
    LUT4 i11422_2_lut (.A(smpl_register[12]), .B(wb_addr[0]), .Z(n1_adj_3075)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(228[3] 235[10])
    defparam i11422_2_lut.init = 16'h8888;
    LUT4 mux_434_Mux_11_i2_3_lut (.A(bus_err_address[9]), .B(power_counter[11]), 
         .C(wb_addr[0]), .Z(n2_adj_3076)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(228[3] 235[10])
    defparam mux_434_Mux_11_i2_3_lut.init = 16'hcaca;
    LUT4 i11421_2_lut (.A(smpl_register[11]), .B(wb_addr[0]), .Z(n1_adj_3077)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(228[3] 235[10])
    defparam i11421_2_lut.init = 16'h8888;
    LUT4 mux_434_Mux_10_i2_3_lut (.A(bus_err_address[8]), .B(power_counter[10]), 
         .C(wb_addr[0]), .Z(n2_adj_3078)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(228[3] 235[10])
    defparam mux_434_Mux_10_i2_3_lut.init = 16'hcaca;
    PFUMX mux_434_Mux_30_i3 (.BLUT(n1_adj_3044), .ALUT(n2_adj_3043), .C0(wb_addr[1]), 
          .Z(n2093));
    LUT4 wb_idata_31__I_0_i31_4_lut (.A(wb_smpl_data[30]), .B(wb_fm_data[30]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_2[30])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(283[8] 288[53])
    defparam wb_idata_31__I_0_i31_4_lut.init = 16'hcac0;
    LUT4 i10187_1_lut (.A(wb_idata[1]), .Z(n12753)) /* synthesis lut_function=(!(A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(280[9] 288[53])
    defparam i10187_1_lut.init = 16'h5555;
    LUT4 wb_idata_31__I_0_i30_4_lut (.A(wb_smpl_data[29]), .B(wb_fm_data[29]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_2[29])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(283[8] 288[53])
    defparam wb_idata_31__I_0_i30_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i29_4_lut (.A(wb_smpl_data[28]), .B(wb_fm_data[28]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_2[28])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(283[8] 288[53])
    defparam wb_idata_31__I_0_i29_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i28_4_lut (.A(wb_smpl_data[27]), .B(wb_fm_data[27]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_2[27])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(283[8] 288[53])
    defparam wb_idata_31__I_0_i28_4_lut.init = 16'hcac0;
    PFUMX mux_434_Mux_31_i3 (.BLUT(n1), .ALUT(n2_adj_3042), .C0(wb_addr[1]), 
          .Z(n2092));
    LUT4 mux_433_i1_4_lut (.A(smpl_interrupt), .B(n21396), .C(n7), .D(n10106), 
         .Z(wb_smpl_data_31__N_64[0])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(228[3] 235[10])
    defparam mux_433_i1_4_lut.init = 16'hca0a;
    LUT4 i1_3_lut (.A(wb_addr[3]), .B(wb_addr[2]), .C(wb_addr[0]), .Z(n21396)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_3_lut.init = 16'h1010;
    LUT4 i7685_3_lut (.A(smpl_register[0]), .B(power_counter[0]), .C(wb_addr[1]), 
         .Z(n10106)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(228[3] 235[10])
    defparam i7685_3_lut.init = 16'hcaca;
    LUT4 wb_idata_31__I_0_i27_4_lut (.A(wb_smpl_data[26]), .B(wb_fm_data[26]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_2[26])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(283[8] 288[53])
    defparam wb_idata_31__I_0_i27_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i26_4_lut (.A(wb_smpl_data[25]), .B(wb_fm_data[25]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_2[25])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(283[8] 288[53])
    defparam wb_idata_31__I_0_i26_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i25_4_lut (.A(wb_smpl_data[24]), .B(wb_fm_data[24]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_2[24])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(283[8] 288[53])
    defparam wb_idata_31__I_0_i25_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i24_4_lut (.A(wb_smpl_data[23]), .B(wb_fm_data[23]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_2[23])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(283[8] 288[53])
    defparam wb_idata_31__I_0_i24_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i23_4_lut (.A(wb_smpl_data[22]), .B(wb_fm_data[22]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_2[22])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(283[8] 288[53])
    defparam wb_idata_31__I_0_i23_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i22_4_lut (.A(wb_smpl_data[21]), .B(wb_fm_data[21]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_2[21])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(283[8] 288[53])
    defparam wb_idata_31__I_0_i22_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i21_4_lut (.A(wb_smpl_data[20]), .B(wb_fm_data[20]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_2[20])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(283[8] 288[53])
    defparam wb_idata_31__I_0_i21_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i20_4_lut (.A(wb_smpl_data[19]), .B(wb_fm_data[19]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_2[19])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(283[8] 288[53])
    defparam wb_idata_31__I_0_i20_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i19_4_lut (.A(wb_smpl_data[18]), .B(wb_fm_data[18]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_2[18])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(283[8] 288[53])
    defparam wb_idata_31__I_0_i19_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i18_4_lut (.A(wb_smpl_data[17]), .B(wb_fm_data[17]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_2[17])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(283[8] 288[53])
    defparam wb_idata_31__I_0_i18_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i17_4_lut (.A(wb_smpl_data[16]), .B(wb_fm_data[16]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_2[16])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(283[8] 288[53])
    defparam wb_idata_31__I_0_i17_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i16_4_lut (.A(wb_smpl_data[15]), .B(wb_fm_data[15]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_2[15])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(283[8] 288[53])
    defparam wb_idata_31__I_0_i16_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i15_4_lut (.A(wb_smpl_data[14]), .B(wb_fm_data[14]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_2[14])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(283[8] 288[53])
    defparam wb_idata_31__I_0_i15_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i14_4_lut (.A(wb_smpl_data[13]), .B(wb_fm_data[13]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_2[13])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(283[8] 288[53])
    defparam wb_idata_31__I_0_i14_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i13_4_lut (.A(wb_smpl_data[12]), .B(wb_fm_data[12]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_2[12])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(283[8] 288[53])
    defparam wb_idata_31__I_0_i13_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i12_4_lut (.A(wb_smpl_data[11]), .B(wb_fm_data[11]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_2[11])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(283[8] 288[53])
    defparam wb_idata_31__I_0_i12_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i11_4_lut (.A(wb_smpl_data[10]), .B(wb_fm_data[10]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_2[10])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(283[8] 288[53])
    defparam wb_idata_31__I_0_i11_4_lut.init = 16'hcac0;
    PFUMX mux_434_Mux_14_i3 (.BLUT(n1_adj_3071), .ALUT(n2_adj_3070), .C0(wb_addr[1]), 
          .Z(n2109));
    LUT4 wb_idata_31__I_0_i10_4_lut (.A(wb_smpl_data[9]), .B(wb_fm_data[9]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_2[9])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(283[8] 288[53])
    defparam wb_idata_31__I_0_i10_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i9_4_lut (.A(wb_smpl_data[8]), .B(wb_fm_data[8]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_2[8])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(283[8] 288[53])
    defparam wb_idata_31__I_0_i9_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i8_3_lut (.A(wb_idata_31__N_266[7]), .B(wb_fm_data[7]), 
         .C(wb_fm_ack), .Z(wb_idata_31__N_2[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(283[8] 288[53])
    defparam wb_idata_31__I_0_i8_3_lut.init = 16'hcaca;
    LUT4 mux_56_i8_4_lut (.A(wb_lo_data[7]), .B(wb_smpl_data[7]), .C(wb_smpl_ack), 
         .D(wb_lo_ack), .Z(wb_idata_31__N_266[7])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(285[8] 288[53])
    defparam mux_56_i8_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i7_3_lut (.A(wb_idata_31__N_266[6]), .B(wb_fm_data[6]), 
         .C(wb_fm_ack), .Z(wb_idata_31__N_2[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(283[8] 288[53])
    defparam wb_idata_31__I_0_i7_3_lut.init = 16'hcaca;
    LUT4 mux_56_i7_4_lut (.A(wb_lo_data[6]), .B(wb_smpl_data[6]), .C(wb_smpl_ack), 
         .D(wb_lo_ack), .Z(wb_idata_31__N_266[6])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(285[8] 288[53])
    defparam mux_56_i7_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i6_3_lut (.A(wb_idata_31__N_266[5]), .B(wb_fm_data[5]), 
         .C(wb_fm_ack), .Z(wb_idata_31__N_2[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(283[8] 288[53])
    defparam wb_idata_31__I_0_i6_3_lut.init = 16'hcaca;
    LUT4 mux_56_i6_4_lut (.A(wb_lo_data[5]), .B(wb_smpl_data[5]), .C(wb_smpl_ack), 
         .D(wb_lo_ack), .Z(wb_idata_31__N_266[5])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(285[8] 288[53])
    defparam mux_56_i6_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i5_3_lut (.A(wb_idata_31__N_266[4]), .B(wb_fm_data[4]), 
         .C(wb_fm_ack), .Z(wb_idata_31__N_2[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(283[8] 288[53])
    defparam wb_idata_31__I_0_i5_3_lut.init = 16'hcaca;
    LUT4 mux_56_i5_4_lut (.A(wb_lo_data[4]), .B(wb_smpl_data[4]), .C(wb_smpl_ack), 
         .D(wb_lo_ack), .Z(wb_idata_31__N_266[4])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(285[8] 288[53])
    defparam mux_56_i5_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i4_3_lut (.A(wb_idata_31__N_266[3]), .B(wb_fm_data[3]), 
         .C(wb_fm_ack), .Z(wb_idata_31__N_2[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(283[8] 288[53])
    defparam wb_idata_31__I_0_i4_3_lut.init = 16'hcaca;
    LUT4 mux_56_i4_4_lut (.A(wb_lo_data[3]), .B(wb_smpl_data[3]), .C(wb_smpl_ack), 
         .D(wb_lo_ack), .Z(wb_idata_31__N_266[3])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(285[8] 288[53])
    defparam mux_56_i4_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i3_3_lut (.A(wb_idata_31__N_266[2]), .B(wb_fm_data[2]), 
         .C(wb_fm_ack), .Z(wb_idata_31__N_2[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(283[8] 288[53])
    defparam wb_idata_31__I_0_i3_3_lut.init = 16'hcaca;
    LUT4 mux_56_i3_4_lut (.A(wb_lo_data[2]), .B(wb_smpl_data[2]), .C(wb_smpl_ack), 
         .D(wb_lo_ack), .Z(wb_idata_31__N_266[2])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(285[8] 288[53])
    defparam mux_56_i3_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i2_3_lut (.A(wb_idata_31__N_266[1]), .B(wb_fm_data[1]), 
         .C(wb_fm_ack), .Z(wb_idata_31__N_2[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(283[8] 288[53])
    defparam wb_idata_31__I_0_i2_3_lut.init = 16'hcaca;
    LUT4 mux_56_i2_4_lut (.A(wb_lo_data[1]), .B(wb_smpl_data[1]), .C(wb_smpl_ack), 
         .D(wb_lo_ack), .Z(wb_idata_31__N_266[1])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(285[8] 288[53])
    defparam mux_56_i2_4_lut.init = 16'hcac0;
    LUT4 power_counter_31__I_0_74_i31_3_lut (.A(power_counter_31__N_232[30]), 
         .B(power_counter_31__N_201[30]), .C(power_counter[31]), .Z(power_counter_31__N_129[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[4:54])
    defparam power_counter_31__I_0_74_i31_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_74_i30_3_lut (.A(power_counter_31__N_232[29]), 
         .B(power_counter_31__N_201[29]), .C(power_counter[31]), .Z(power_counter_31__N_129[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[4:54])
    defparam power_counter_31__I_0_74_i30_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_74_i29_3_lut (.A(power_counter_31__N_232[28]), 
         .B(power_counter_31__N_201[28]), .C(power_counter[31]), .Z(power_counter_31__N_129[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[4:54])
    defparam power_counter_31__I_0_74_i29_3_lut.init = 16'hcaca;
    CCU2D add_31_25 (.A0(power_counter[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17853), .COUT(n17854), .S0(power_counter_31__N_232[23]), 
          .S1(power_counter_31__N_232[24]));   // d:/documents/git_local/fm_modulator/rtl/top.v(242[21:41])
    defparam add_31_25.INIT0 = 16'h5aaa;
    defparam add_31_25.INIT1 = 16'h5aaa;
    defparam add_31_25.INJECT1_0 = "NO";
    defparam add_31_25.INJECT1_1 = "NO";
    LUT4 power_counter_31__I_0_74_i28_3_lut (.A(power_counter_31__N_232[27]), 
         .B(power_counter_31__N_201[27]), .C(power_counter[31]), .Z(power_counter_31__N_129[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[4:54])
    defparam power_counter_31__I_0_74_i28_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_74_i27_3_lut (.A(power_counter_31__N_232[26]), 
         .B(power_counter_31__N_201[26]), .C(power_counter[31]), .Z(power_counter_31__N_129[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[4:54])
    defparam power_counter_31__I_0_74_i27_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_74_i26_3_lut (.A(power_counter_31__N_232[25]), 
         .B(power_counter_31__N_201[25]), .C(power_counter[31]), .Z(power_counter_31__N_129[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[4:54])
    defparam power_counter_31__I_0_74_i26_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_74_i25_3_lut (.A(power_counter_31__N_232[24]), 
         .B(power_counter_31__N_201[24]), .C(power_counter[31]), .Z(power_counter_31__N_129[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[4:54])
    defparam power_counter_31__I_0_74_i25_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_74_i24_3_lut (.A(power_counter_31__N_232[23]), 
         .B(power_counter_31__N_201[23]), .C(power_counter[31]), .Z(power_counter_31__N_129[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[4:54])
    defparam power_counter_31__I_0_74_i24_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_74_i23_3_lut (.A(power_counter_31__N_232[22]), 
         .B(power_counter_31__N_201[22]), .C(power_counter[31]), .Z(power_counter_31__N_129[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[4:54])
    defparam power_counter_31__I_0_74_i23_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_74_i22_3_lut (.A(power_counter_31__N_232[21]), 
         .B(power_counter_31__N_201[21]), .C(power_counter[31]), .Z(power_counter_31__N_129[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[4:54])
    defparam power_counter_31__I_0_74_i22_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_74_i21_3_lut (.A(power_counter_31__N_232[20]), 
         .B(power_counter_31__N_201[20]), .C(power_counter[31]), .Z(power_counter_31__N_129[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[4:54])
    defparam power_counter_31__I_0_74_i21_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_74_i20_3_lut (.A(power_counter_31__N_232[19]), 
         .B(power_counter_31__N_201[19]), .C(power_counter[31]), .Z(power_counter_31__N_129[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[4:54])
    defparam power_counter_31__I_0_74_i20_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_74_i19_3_lut (.A(power_counter_31__N_232[18]), 
         .B(power_counter_31__N_201[18]), .C(power_counter[31]), .Z(power_counter_31__N_129[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[4:54])
    defparam power_counter_31__I_0_74_i19_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_74_i18_3_lut (.A(power_counter_31__N_232[17]), 
         .B(power_counter_31__N_201[17]), .C(power_counter[31]), .Z(power_counter_31__N_129[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[4:54])
    defparam power_counter_31__I_0_74_i18_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_74_i17_3_lut (.A(power_counter_31__N_232[16]), 
         .B(power_counter_31__N_201[16]), .C(power_counter[31]), .Z(power_counter_31__N_129[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[4:54])
    defparam power_counter_31__I_0_74_i17_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_74_i16_3_lut (.A(power_counter_31__N_232[15]), 
         .B(power_counter_31__N_201[15]), .C(power_counter[31]), .Z(power_counter_31__N_129[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[4:54])
    defparam power_counter_31__I_0_74_i16_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_74_i15_3_lut (.A(power_counter_31__N_232[14]), 
         .B(power_counter_31__N_201[14]), .C(power_counter[31]), .Z(power_counter_31__N_129[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[4:54])
    defparam power_counter_31__I_0_74_i15_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_74_i14_3_lut (.A(power_counter_31__N_232[13]), 
         .B(power_counter_31__N_201[13]), .C(power_counter[31]), .Z(power_counter_31__N_129[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[4:54])
    defparam power_counter_31__I_0_74_i14_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_74_i13_3_lut (.A(power_counter_31__N_232[12]), 
         .B(power_counter_31__N_201[12]), .C(power_counter[31]), .Z(power_counter_31__N_129[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[4:54])
    defparam power_counter_31__I_0_74_i13_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_74_i12_3_lut (.A(power_counter_31__N_232[11]), 
         .B(power_counter_31__N_201[11]), .C(power_counter[31]), .Z(power_counter_31__N_129[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[4:54])
    defparam power_counter_31__I_0_74_i12_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_74_i11_3_lut (.A(power_counter_31__N_232[10]), 
         .B(power_counter_31__N_201[10]), .C(power_counter[31]), .Z(power_counter_31__N_129[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[4:54])
    defparam power_counter_31__I_0_74_i11_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_74_i10_3_lut (.A(power_counter_31__N_232[9]), 
         .B(power_counter_31__N_201[9]), .C(power_counter[31]), .Z(power_counter_31__N_129[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[4:54])
    defparam power_counter_31__I_0_74_i10_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_74_i9_3_lut (.A(power_counter_31__N_232[8]), 
         .B(power_counter_31__N_201[8]), .C(power_counter[31]), .Z(power_counter_31__N_129[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[4:54])
    defparam power_counter_31__I_0_74_i9_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_74_i8_3_lut (.A(power_counter_31__N_232[7]), 
         .B(power_counter_31__N_201[7]), .C(power_counter[31]), .Z(power_counter_31__N_129[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[4:54])
    defparam power_counter_31__I_0_74_i8_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_74_i7_3_lut (.A(power_counter_31__N_232[6]), 
         .B(power_counter_31__N_201[6]), .C(power_counter[31]), .Z(power_counter_31__N_129[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[4:54])
    defparam power_counter_31__I_0_74_i7_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_74_i6_3_lut (.A(power_counter_31__N_232[5]), 
         .B(power_counter_31__N_201[5]), .C(power_counter[31]), .Z(power_counter_31__N_129[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[4:54])
    defparam power_counter_31__I_0_74_i6_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_74_i5_3_lut (.A(power_counter_31__N_232[4]), 
         .B(power_counter_31__N_201[4]), .C(power_counter[31]), .Z(power_counter_31__N_129[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[4:54])
    defparam power_counter_31__I_0_74_i5_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_74_i4_3_lut (.A(power_counter_31__N_232[3]), 
         .B(power_counter_31__N_201[3]), .C(power_counter[31]), .Z(power_counter_31__N_129[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[4:54])
    defparam power_counter_31__I_0_74_i4_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_74_i3_3_lut (.A(power_counter_31__N_232[2]), 
         .B(power_counter_31__N_201[2]), .C(power_counter[31]), .Z(power_counter_31__N_129[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[4:54])
    defparam power_counter_31__I_0_74_i3_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_74_i2_3_lut (.A(power_counter_31__N_232[1]), 
         .B(power_counter_31__N_201[1]), .C(power_counter[31]), .Z(power_counter_31__N_129[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[4:54])
    defparam power_counter_31__I_0_74_i2_3_lut.init = 16'hcaca;
    CCU2D add_32_31 (.A0(power_counter[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17872), .S0(power_counter_31__N_201[29]), 
          .S1(power_counter_31__N_201[30]));   // d:/documents/git_local/fm_modulator/rtl/top.v(244[27:53])
    defparam add_32_31.INIT0 = 16'h5aaa;
    defparam add_32_31.INIT1 = 16'h5aaa;
    defparam add_32_31.INJECT1_0 = "NO";
    defparam add_32_31.INJECT1_1 = "NO";
    PFUMX mux_434_Mux_15_i3 (.BLUT(n1_adj_3069), .ALUT(n2_adj_3068), .C0(wb_addr[1]), 
          .Z(n2108));
    CCU2D add_31_23 (.A0(power_counter[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17852), .COUT(n17853), .S0(power_counter_31__N_232[21]), 
          .S1(power_counter_31__N_232[22]));   // d:/documents/git_local/fm_modulator/rtl/top.v(242[21:41])
    defparam add_31_23.INIT0 = 16'h5aaa;
    defparam add_31_23.INIT1 = 16'h5aaa;
    defparam add_31_23.INJECT1_0 = "NO";
    defparam add_31_23.INJECT1_1 = "NO";
    CCU2D add_32_29 (.A0(power_counter[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17871), .COUT(n17872), .S0(power_counter_31__N_201[27]), 
          .S1(power_counter_31__N_201[28]));   // d:/documents/git_local/fm_modulator/rtl/top.v(244[27:53])
    defparam add_32_29.INIT0 = 16'h5aaa;
    defparam add_32_29.INIT1 = 16'h5aaa;
    defparam add_32_29.INJECT1_0 = "NO";
    defparam add_32_29.INJECT1_1 = "NO";
    LUT4 dac_clk_p_I_0_1_lut (.A(dac_clk_p_c), .Z(dac_clk_n_c)) /* synthesis lut_function=(!(A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(56[20:30])
    defparam dac_clk_p_I_0_1_lut.init = 16'h5555;
    LUT4 mux_434_Mux_25_i2_3_lut (.A(bus_err_address[23]), .B(power_counter[25]), 
         .C(wb_addr[0]), .Z(n2_adj_3052)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(228[3] 235[10])
    defparam mux_434_Mux_25_i2_3_lut.init = 16'hcaca;
    LUT4 mux_434_Mux_9_i2_3_lut (.A(bus_err_address[7]), .B(power_counter[9]), 
         .C(wb_addr[0]), .Z(n2_adj_3079)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(228[3] 235[10])
    defparam mux_434_Mux_9_i2_3_lut.init = 16'hcaca;
    LUT4 mux_434_Mux_8_i2_3_lut (.A(bus_err_address[6]), .B(power_counter[8]), 
         .C(wb_addr[0]), .Z(n2_adj_3080)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(228[3] 235[10])
    defparam mux_434_Mux_8_i2_3_lut.init = 16'hcaca;
    LUT4 i11435_2_lut (.A(smpl_register[25]), .B(wb_addr[0]), .Z(n1_adj_3053)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(228[3] 235[10])
    defparam i11435_2_lut.init = 16'h8888;
    LUT4 i11418_2_lut (.A(smpl_register[8]), .B(wb_addr[0]), .Z(n1_adj_3081)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(228[3] 235[10])
    defparam i11418_2_lut.init = 16'h8888;
    LUT4 mux_434_Mux_7_i2_3_lut (.A(bus_err_address[5]), .B(power_counter[7]), 
         .C(wb_addr[0]), .Z(n2_adj_3082)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(228[3] 235[10])
    defparam mux_434_Mux_7_i2_3_lut.init = 16'hcaca;
    LUT4 mux_434_Mux_24_i2_3_lut (.A(bus_err_address[22]), .B(power_counter[24]), 
         .C(wb_addr[0]), .Z(n2_adj_3054)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(228[3] 235[10])
    defparam mux_434_Mux_24_i2_3_lut.init = 16'hcaca;
    LUT4 i11417_2_lut (.A(smpl_register[7]), .B(wb_addr[0]), .Z(n1_adj_3083)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(228[3] 235[10])
    defparam i11417_2_lut.init = 16'h8888;
    VLO i1 (.Z(GND_net));
    FD1S3AX wb_idata_i31 (.D(wb_idata_31__N_2[31]), .CK(dac_clk_p_c), .Q(wb_idata[31]));   // d:/documents/git_local/fm_modulator/rtl/top.v(280[9] 288[53])
    defparam wb_idata_i31.GSR = "DISABLED";
    LUT4 i11434_2_lut (.A(smpl_register[24]), .B(wb_addr[0]), .Z(n1_adj_3055)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(228[3] 235[10])
    defparam i11434_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_rep_639 (.A(wb_stb), .B(wb_we), .Z(n27304)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(218[7:30])
    defparam i1_2_lut_rep_639.init = 16'h8888;
    LUT4 i1_3_lut_4_lut_adj_162 (.A(wb_stb), .B(wb_we), .C(wb_addr[15]), 
         .D(wb_addr[0]), .Z(n21026)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(218[7:30])
    defparam i1_3_lut_4_lut_adj_162.init = 16'h8000;
    LUT4 i23043_3_lut_4_lut (.A(wb_stb), .B(wb_we), .C(n7), .D(wb_smpl_sel_N_310), 
         .Z(dac_clk_p_c_enable_224)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(218[7:30])
    defparam i23043_3_lut_4_lut.init = 16'h0008;
    LUT4 i1_4_lut_adj_163 (.A(n27140), .B(n21096), .C(n34), .D(wb_addr[0]), 
         .Z(n21102)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(256[23:49])
    defparam i1_4_lut_adj_163.init = 16'hfffe;
    LUT4 mux_434_Mux_6_i2_3_lut (.A(bus_err_address[4]), .B(power_counter[6]), 
         .C(wb_addr[0]), .Z(n2_adj_3084)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(228[3] 235[10])
    defparam mux_434_Mux_6_i2_3_lut.init = 16'hcaca;
    LUT4 i11416_2_lut (.A(smpl_register[6]), .B(wb_addr[0]), .Z(n1_adj_3085)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(228[3] 235[10])
    defparam i11416_2_lut.init = 16'h8888;
    LUT4 mux_434_Mux_5_i2_3_lut (.A(bus_err_address[3]), .B(power_counter[5]), 
         .C(wb_addr[0]), .Z(n2_adj_3086)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(228[3] 235[10])
    defparam mux_434_Mux_5_i2_3_lut.init = 16'hcaca;
    LUT4 i6_2_lut_rep_648 (.A(wb_addr[22]), .B(wb_addr[24]), .Z(n27313)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(256[23:49])
    defparam i6_2_lut_rep_648.init = 16'heeee;
    LUT4 i1_2_lut_3_lut (.A(wb_addr[22]), .B(wb_addr[24]), .C(wb_addr[9]), 
         .Z(n21096)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(256[23:49])
    defparam i1_2_lut_3_lut.init = 16'hefef;
    LUT4 mux_434_Mux_4_i2_3_lut (.A(bus_err_address[2]), .B(power_counter[4]), 
         .C(wb_addr[0]), .Z(n2_adj_3087)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(228[3] 235[10])
    defparam mux_434_Mux_4_i2_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_4_lut_adj_164 (.A(wb_addr[22]), .B(wb_addr[24]), .C(wb_addr[12]), 
         .D(n38), .Z(n21248)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(256[23:49])
    defparam i1_3_lut_4_lut_adj_164.init = 16'hfffe;
    LUT4 i11414_2_lut (.A(smpl_register[4]), .B(wb_addr[0]), .Z(n1_adj_3088)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(228[3] 235[10])
    defparam i11414_2_lut.init = 16'h8888;
    PFUMX mux_434_Mux_19_i3 (.BLUT(n1_adj_3064), .ALUT(n2_adj_3063), .C0(wb_addr[1]), 
          .Z(n2104));
    PFUMX mux_434_Mux_21_i3 (.BLUT(n1_adj_3061), .ALUT(n2_adj_3060), .C0(wb_addr[1]), 
          .Z(n2102));
    LUT4 mux_434_Mux_3_i2_3_lut (.A(bus_err_address[1]), .B(power_counter[3]), 
         .C(wb_addr[0]), .Z(n2_adj_3089)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(228[3] 235[10])
    defparam mux_434_Mux_3_i2_3_lut.init = 16'hcaca;
    TSALL TSALL_INST (.TSALL(GND_net));
    LUT4 i11413_2_lut (.A(smpl_register[3]), .B(wb_addr[0]), .Z(n1_adj_3090)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(228[3] 235[10])
    defparam i11413_2_lut.init = 16'h8888;
    FD1S3AX wb_idata_i30 (.D(wb_idata_31__N_2[30]), .CK(dac_clk_p_c), .Q(wb_idata[30]));   // d:/documents/git_local/fm_modulator/rtl/top.v(280[9] 288[53])
    defparam wb_idata_i30.GSR = "DISABLED";
    FD1S3AX wb_idata_i29 (.D(wb_idata_31__N_2[29]), .CK(dac_clk_p_c), .Q(wb_idata[29]));   // d:/documents/git_local/fm_modulator/rtl/top.v(280[9] 288[53])
    defparam wb_idata_i29.GSR = "DISABLED";
    PFUMX mux_434_Mux_22_i3 (.BLUT(n1_adj_3059), .ALUT(n2_adj_3058), .C0(wb_addr[1]), 
          .Z(n2101));
    CCU2D add_31_21 (.A0(power_counter[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17851), .COUT(n17852), .S0(power_counter_31__N_232[19]), 
          .S1(power_counter_31__N_232[20]));   // d:/documents/git_local/fm_modulator/rtl/top.v(242[21:41])
    defparam add_31_21.INIT0 = 16'h5aaa;
    defparam add_31_21.INIT1 = 16'h5aaa;
    defparam add_31_21.INJECT1_0 = "NO";
    defparam add_31_21.INJECT1_1 = "NO";
    FD1S3AX wb_idata_i28 (.D(wb_idata_31__N_2[28]), .CK(dac_clk_p_c), .Q(wb_idata[28]));   // d:/documents/git_local/fm_modulator/rtl/top.v(280[9] 288[53])
    defparam wb_idata_i28.GSR = "DISABLED";
    LUT4 mux_434_Mux_23_i2_3_lut (.A(bus_err_address[21]), .B(power_counter[23]), 
         .C(wb_addr[0]), .Z(n2_adj_3056)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(228[3] 235[10])
    defparam mux_434_Mux_23_i2_3_lut.init = 16'hcaca;
    FD1S3AX wb_idata_i27 (.D(wb_idata_31__N_2[27]), .CK(dac_clk_p_c), .Q(wb_idata[27]));   // d:/documents/git_local/fm_modulator/rtl/top.v(280[9] 288[53])
    defparam wb_idata_i27.GSR = "DISABLED";
    LUT4 i11433_2_lut (.A(smpl_register[23]), .B(wb_addr[0]), .Z(n1_adj_3057)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(228[3] 235[10])
    defparam i11433_2_lut.init = 16'h8888;
    efb_inst wb_lo_data_7__I_0 (.dac_clk_p_c(dac_clk_p_c), .i_sw0_c(i_sw0_c), 
            .wb_cyc(wb_cyc), .wb_lo_data_7__N_96(wb_lo_data_7__N_96), .wb_we(wb_we), 
            .\wb_addr[7] (wb_addr[7]), .\wb_addr[6] (wb_addr[6]), .\wb_addr[5] (wb_addr[5]), 
            .\wb_addr[4] (wb_addr[4]), .\wb_addr[3] (wb_addr[3]), .\wb_addr[2] (wb_addr[2]), 
            .\wb_addr[1] (wb_addr[1]), .\wb_addr[0] (wb_addr[0]), .\wb_odata[7] (wb_odata[7]), 
            .\wb_odata[6] (wb_odata[6]), .\wb_odata[5] (wb_odata[5]), .\wb_odata[4] (wb_odata[4]), 
            .\wb_odata[3] (wb_odata[3]), .\wb_odata[2] (wb_odata[2]), .\wb_odata[1] (wb_odata[1]), 
            .\wb_odata[0] (wb_odata[0]), .pll_data_o({pll_data_o}), .pll_ack(pll_ack), 
            .wb_lo_data({wb_lo_data}), .wb_lo_ack(wb_lo_ack), .pll_clk(pll_clk), 
            .pll_rst(pll_rst), .pll_stb(pll_stb), .pll_we(pll_we), .pll_addr({pll_addr}), 
            .pll_data_i({pll_data_i}), .GND_net(GND_net), .VCC_net(VCC_net)) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(187[11] 199[4])
    clock_phase_shifter clock_phase_shifter_inst (.q_clk_p_c(q_clk_p_c), .i_clk_2f_N_2268(i_clk_2f_N_2268), 
            .q_clk_n_c(q_clk_n_c), .i_clk_p_c(i_clk_p_c), .lo_pll_out(lo_pll_out), 
            .i_clk_n_c(i_clk_n_c)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(167[21] 171[2])
    FD1S3AX wb_smpl_data_i0 (.D(wb_smpl_data_31__N_64[0]), .CK(dac_clk_p_c), 
            .Q(wb_smpl_data[0]));   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 235[10])
    defparam wb_smpl_data_i0.GSR = "DISABLED";
    CCU2D add_32_27 (.A0(power_counter[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17870), .COUT(n17871), .S0(power_counter_31__N_201[25]), 
          .S1(power_counter_31__N_201[26]));   // d:/documents/git_local/fm_modulator/rtl/top.v(244[27:53])
    defparam add_32_27.INIT0 = 16'h5aaa;
    defparam add_32_27.INIT1 = 16'h5aaa;
    defparam add_32_27.INJECT1_0 = "NO";
    defparam add_32_27.INJECT1_1 = "NO";
    CCU2D add_31_19 (.A0(power_counter[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17850), .COUT(n17851), .S0(power_counter_31__N_232[17]), 
          .S1(power_counter_31__N_232[18]));   // d:/documents/git_local/fm_modulator/rtl/top.v(242[21:41])
    defparam add_31_19.INIT0 = 16'h5aaa;
    defparam add_31_19.INIT1 = 16'h5aaa;
    defparam add_31_19.INJECT1_0 = "NO";
    defparam add_31_19.INJECT1_1 = "NO";
    CCU2D add_32_25 (.A0(power_counter[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17869), .COUT(n17870), .S0(power_counter_31__N_201[23]), 
          .S1(power_counter_31__N_201[24]));   // d:/documents/git_local/fm_modulator/rtl/top.v(244[27:53])
    defparam add_32_25.INIT0 = 16'h5aaa;
    defparam add_32_25.INIT1 = 16'h5aaa;
    defparam add_32_25.INJECT1_0 = "NO";
    defparam add_32_25.INJECT1_1 = "NO";
    CCU2D add_31_17 (.A0(power_counter[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17849), .COUT(n17850), .S0(power_counter_31__N_232[15]), 
          .S1(power_counter_31__N_232[16]));   // d:/documents/git_local/fm_modulator/rtl/top.v(242[21:41])
    defparam add_31_17.INIT0 = 16'h5aaa;
    defparam add_31_17.INIT1 = 16'h5aaa;
    defparam add_31_17.INJECT1_0 = "NO";
    defparam add_31_17.INJECT1_1 = "NO";
    CCU2D add_32_23 (.A0(power_counter[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17868), .COUT(n17869), .S0(power_counter_31__N_201[21]), 
          .S1(power_counter_31__N_201[22]));   // d:/documents/git_local/fm_modulator/rtl/top.v(244[27:53])
    defparam add_32_23.INIT0 = 16'h5aaa;
    defparam add_32_23.INIT1 = 16'h5aaa;
    defparam add_32_23.INJECT1_0 = "NO";
    defparam add_32_23.INJECT1_1 = "NO";
    CCU2D add_31_15 (.A0(power_counter[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17848), .COUT(n17849), .S0(power_counter_31__N_232[13]), 
          .S1(power_counter_31__N_232[14]));   // d:/documents/git_local/fm_modulator/rtl/top.v(242[21:41])
    defparam add_31_15.INIT0 = 16'h5aaa;
    defparam add_31_15.INIT1 = 16'h5aaa;
    defparam add_31_15.INJECT1_0 = "NO";
    defparam add_31_15.INJECT1_1 = "NO";
    CCU2D add_32_21 (.A0(power_counter[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17867), .COUT(n17868), .S0(power_counter_31__N_201[19]), 
          .S1(power_counter_31__N_201[20]));   // d:/documents/git_local/fm_modulator/rtl/top.v(244[27:53])
    defparam add_32_21.INIT0 = 16'h5aaa;
    defparam add_32_21.INIT1 = 16'h5aaa;
    defparam add_32_21.INJECT1_0 = "NO";
    defparam add_32_21.INJECT1_1 = "NO";
    CCU2D add_31_5 (.A0(power_counter[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17843), .COUT(n17844), .S0(power_counter_31__N_232[3]), 
          .S1(power_counter_31__N_232[4]));   // d:/documents/git_local/fm_modulator/rtl/top.v(242[21:41])
    defparam add_31_5.INIT0 = 16'h5aaa;
    defparam add_31_5.INIT1 = 16'h5aaa;
    defparam add_31_5.INJECT1_0 = "NO";
    defparam add_31_5.INJECT1_1 = "NO";
    CCU2D add_32_19 (.A0(power_counter[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17866), .COUT(n17867), .S0(power_counter_31__N_201[17]), 
          .S1(power_counter_31__N_201[18]));   // d:/documents/git_local/fm_modulator/rtl/top.v(244[27:53])
    defparam add_32_19.INIT0 = 16'h5aaa;
    defparam add_32_19.INIT1 = 16'h5aaa;
    defparam add_32_19.INJECT1_0 = "NO";
    defparam add_32_19.INJECT1_1 = "NO";
    CCU2D add_32_17 (.A0(power_counter[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17865), .COUT(n17866), .S0(power_counter_31__N_201[15]), 
          .S1(power_counter_31__N_201[16]));   // d:/documents/git_local/fm_modulator/rtl/top.v(244[27:53])
    defparam add_32_17.INIT0 = 16'h5aaa;
    defparam add_32_17.INIT1 = 16'h5aaa;
    defparam add_32_17.INJECT1_0 = "NO";
    defparam add_32_17.INJECT1_1 = "NO";
    CCU2D add_32_15 (.A0(power_counter[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17864), .COUT(n17865), .S0(power_counter_31__N_201[13]), 
          .S1(power_counter_31__N_201[14]));   // d:/documents/git_local/fm_modulator/rtl/top.v(244[27:53])
    defparam add_32_15.INIT0 = 16'h5aaa;
    defparam add_32_15.INIT1 = 16'h5aaa;
    defparam add_32_15.INJECT1_0 = "NO";
    defparam add_32_15.INJECT1_1 = "NO";
    CCU2D add_32_13 (.A0(power_counter[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17863), .COUT(n17864), .S0(power_counter_31__N_201[11]), 
          .S1(power_counter_31__N_201[12]));   // d:/documents/git_local/fm_modulator/rtl/top.v(244[27:53])
    defparam add_32_13.INIT0 = 16'h5aaa;
    defparam add_32_13.INIT1 = 16'h5aaa;
    defparam add_32_13.INJECT1_0 = "NO";
    defparam add_32_13.INJECT1_1 = "NO";
    CCU2D add_31_9 (.A0(power_counter[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17845), .COUT(n17846), .S0(power_counter_31__N_232[7]), 
          .S1(power_counter_31__N_232[8]));   // d:/documents/git_local/fm_modulator/rtl/top.v(242[21:41])
    defparam add_31_9.INIT0 = 16'h5aaa;
    defparam add_31_9.INIT1 = 16'h5aaa;
    defparam add_31_9.INJECT1_0 = "NO";
    defparam add_31_9.INJECT1_1 = "NO";
    CCU2D add_32_11 (.A0(power_counter[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17862), .COUT(n17863), .S0(power_counter_31__N_201[9]), 
          .S1(power_counter_31__N_201[10]));   // d:/documents/git_local/fm_modulator/rtl/top.v(244[27:53])
    defparam add_32_11.INIT0 = 16'h5aaa;
    defparam add_32_11.INIT1 = 16'h5aaa;
    defparam add_32_11.INJECT1_0 = "NO";
    defparam add_32_11.INJECT1_1 = "NO";
    CCU2D add_32_9 (.A0(power_counter[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17861), .COUT(n17862), .S0(power_counter_31__N_201[7]), 
          .S1(power_counter_31__N_201[8]));   // d:/documents/git_local/fm_modulator/rtl/top.v(244[27:53])
    defparam add_32_9.INIT0 = 16'h5aaa;
    defparam add_32_9.INIT1 = 16'h5aaa;
    defparam add_32_9.INJECT1_0 = "NO";
    defparam add_32_9.INJECT1_1 = "NO";
    CCU2D add_31_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(power_counter[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n17842), .S1(power_counter_31__N_232[0]));   // d:/documents/git_local/fm_modulator/rtl/top.v(242[21:41])
    defparam add_31_1.INIT0 = 16'hF000;
    defparam add_31_1.INIT1 = 16'h5555;
    defparam add_31_1.INJECT1_0 = "NO";
    defparam add_31_1.INJECT1_1 = "NO";
    CCU2D add_32_7 (.A0(power_counter[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17860), .COUT(n17861), .S0(power_counter_31__N_201[5]), 
          .S1(power_counter_31__N_201[6]));   // d:/documents/git_local/fm_modulator/rtl/top.v(244[27:53])
    defparam add_32_7.INIT0 = 16'h5aaa;
    defparam add_32_7.INIT1 = 16'h5aaa;
    defparam add_32_7.INJECT1_0 = "NO";
    defparam add_32_7.INJECT1_1 = "NO";
    CCU2D add_32_5 (.A0(power_counter[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17859), .COUT(n17860), .S0(power_counter_31__N_201[3]), 
          .S1(power_counter_31__N_201[4]));   // d:/documents/git_local/fm_modulator/rtl/top.v(244[27:53])
    defparam add_32_5.INIT0 = 16'h5aaa;
    defparam add_32_5.INIT1 = 16'h5aaa;
    defparam add_32_5.INJECT1_0 = "NO";
    defparam add_32_5.INJECT1_1 = "NO";
    CCU2D add_31_3 (.A0(power_counter[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17842), .COUT(n17843), .S0(power_counter_31__N_232[1]), 
          .S1(power_counter_31__N_232[2]));   // d:/documents/git_local/fm_modulator/rtl/top.v(242[21:41])
    defparam add_31_3.INIT0 = 16'h5aaa;
    defparam add_31_3.INIT1 = 16'h5aaa;
    defparam add_31_3.INJECT1_0 = "NO";
    defparam add_31_3.INJECT1_1 = "NO";
    CCU2D add_32_3 (.A0(power_counter[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17858), .COUT(n17859), .S0(power_counter_31__N_201[1]), 
          .S1(power_counter_31__N_201[2]));   // d:/documents/git_local/fm_modulator/rtl/top.v(244[27:53])
    defparam add_32_3.INIT0 = 16'h5aaa;
    defparam add_32_3.INIT1 = 16'h5aaa;
    defparam add_32_3.INJECT1_0 = "NO";
    defparam add_32_3.INJECT1_1 = "NO";
    CCU2D add_31_13 (.A0(power_counter[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17847), .COUT(n17848), .S0(power_counter_31__N_232[11]), 
          .S1(power_counter_31__N_232[12]));   // d:/documents/git_local/fm_modulator/rtl/top.v(242[21:41])
    defparam add_31_13.INIT0 = 16'h5aaa;
    defparam add_31_13.INIT1 = 16'h5aaa;
    defparam add_31_13.INJECT1_0 = "NO";
    defparam add_31_13.INJECT1_1 = "NO";
    CCU2D add_32_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(power_counter[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n17858), .S1(power_counter_31__N_201[0]));   // d:/documents/git_local/fm_modulator/rtl/top.v(244[27:53])
    defparam add_32_1.INIT0 = 16'hF000;
    defparam add_32_1.INIT1 = 16'h5555;
    defparam add_32_1.INJECT1_0 = "NO";
    defparam add_32_1.INJECT1_1 = "NO";
    CCU2D add_31_7 (.A0(power_counter[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17844), .COUT(n17845), .S0(power_counter_31__N_232[5]), 
          .S1(power_counter_31__N_232[6]));   // d:/documents/git_local/fm_modulator/rtl/top.v(242[21:41])
    defparam add_31_7.INIT0 = 16'h5aaa;
    defparam add_31_7.INIT1 = 16'h5aaa;
    defparam add_31_7.INJECT1_0 = "NO";
    defparam add_31_7.INJECT1_1 = "NO";
    CCU2D add_31_33 (.A0(power_counter[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n17857), .S0(power_counter_31__N_232[31]));   // d:/documents/git_local/fm_modulator/rtl/top.v(242[21:41])
    defparam add_31_33.INIT0 = 16'h5aaa;
    defparam add_31_33.INIT1 = 16'h0000;
    defparam add_31_33.INJECT1_0 = "NO";
    defparam add_31_33.INJECT1_1 = "NO";
    OB o_dac_a_pad_6 (.I(o_dac_a_c_6), .O(o_dac_a[6]));   // d:/documents/git_local/fm_modulator/rtl/top.v(33[38:45])
    FD1S3AX wb_idata_i26 (.D(wb_idata_31__N_2[26]), .CK(dac_clk_p_c), .Q(wb_idata[26]));   // d:/documents/git_local/fm_modulator/rtl/top.v(280[9] 288[53])
    defparam wb_idata_i26.GSR = "DISABLED";
    FD1S3AX wb_idata_i25 (.D(wb_idata_31__N_2[25]), .CK(dac_clk_p_c), .Q(wb_idata[25]));   // d:/documents/git_local/fm_modulator/rtl/top.v(280[9] 288[53])
    defparam wb_idata_i25.GSR = "DISABLED";
    FD1S3AX wb_idata_i24 (.D(wb_idata_31__N_2[24]), .CK(dac_clk_p_c), .Q(wb_idata[24]));   // d:/documents/git_local/fm_modulator/rtl/top.v(280[9] 288[53])
    defparam wb_idata_i24.GSR = "DISABLED";
    FD1S3AX wb_idata_i23 (.D(wb_idata_31__N_2[23]), .CK(dac_clk_p_c), .Q(wb_idata[23]));   // d:/documents/git_local/fm_modulator/rtl/top.v(280[9] 288[53])
    defparam wb_idata_i23.GSR = "DISABLED";
    FD1S3AX wb_idata_i22 (.D(wb_idata_31__N_2[22]), .CK(dac_clk_p_c), .Q(wb_idata[22]));   // d:/documents/git_local/fm_modulator/rtl/top.v(280[9] 288[53])
    defparam wb_idata_i22.GSR = "DISABLED";
    FD1S3AX wb_idata_i21 (.D(wb_idata_31__N_2[21]), .CK(dac_clk_p_c), .Q(wb_idata[21]));   // d:/documents/git_local/fm_modulator/rtl/top.v(280[9] 288[53])
    defparam wb_idata_i21.GSR = "DISABLED";
    FD1S3AX wb_idata_i20 (.D(wb_idata_31__N_2[20]), .CK(dac_clk_p_c), .Q(wb_idata[20]));   // d:/documents/git_local/fm_modulator/rtl/top.v(280[9] 288[53])
    defparam wb_idata_i20.GSR = "DISABLED";
    FD1S3AX wb_idata_i19 (.D(wb_idata_31__N_2[19]), .CK(dac_clk_p_c), .Q(wb_idata[19]));   // d:/documents/git_local/fm_modulator/rtl/top.v(280[9] 288[53])
    defparam wb_idata_i19.GSR = "DISABLED";
    FD1S3AX wb_idata_i18 (.D(wb_idata_31__N_2[18]), .CK(dac_clk_p_c), .Q(wb_idata[18]));   // d:/documents/git_local/fm_modulator/rtl/top.v(280[9] 288[53])
    defparam wb_idata_i18.GSR = "DISABLED";
    FD1S3AX wb_idata_i17 (.D(wb_idata_31__N_2[17]), .CK(dac_clk_p_c), .Q(wb_idata[17]));   // d:/documents/git_local/fm_modulator/rtl/top.v(280[9] 288[53])
    defparam wb_idata_i17.GSR = "DISABLED";
    FD1S3AX wb_idata_i16 (.D(wb_idata_31__N_2[16]), .CK(dac_clk_p_c), .Q(wb_idata[16]));   // d:/documents/git_local/fm_modulator/rtl/top.v(280[9] 288[53])
    defparam wb_idata_i16.GSR = "DISABLED";
    FD1S3AX wb_idata_i15 (.D(wb_idata_31__N_2[15]), .CK(dac_clk_p_c), .Q(wb_idata[15]));   // d:/documents/git_local/fm_modulator/rtl/top.v(280[9] 288[53])
    defparam wb_idata_i15.GSR = "DISABLED";
    FD1S3AX wb_idata_i14 (.D(wb_idata_31__N_2[14]), .CK(dac_clk_p_c), .Q(wb_idata[14]));   // d:/documents/git_local/fm_modulator/rtl/top.v(280[9] 288[53])
    defparam wb_idata_i14.GSR = "DISABLED";
    FD1S3AX wb_idata_i13 (.D(wb_idata_31__N_2[13]), .CK(dac_clk_p_c), .Q(wb_idata[13]));   // d:/documents/git_local/fm_modulator/rtl/top.v(280[9] 288[53])
    defparam wb_idata_i13.GSR = "DISABLED";
    FD1S3AX wb_idata_i12 (.D(wb_idata_31__N_2[12]), .CK(dac_clk_p_c), .Q(wb_idata[12]));   // d:/documents/git_local/fm_modulator/rtl/top.v(280[9] 288[53])
    defparam wb_idata_i12.GSR = "DISABLED";
    FD1S3AX wb_idata_i11 (.D(wb_idata_31__N_2[11]), .CK(dac_clk_p_c), .Q(wb_idata[11]));   // d:/documents/git_local/fm_modulator/rtl/top.v(280[9] 288[53])
    defparam wb_idata_i11.GSR = "DISABLED";
    FD1S3AX wb_idata_i10 (.D(wb_idata_31__N_2[10]), .CK(dac_clk_p_c), .Q(wb_idata[10]));   // d:/documents/git_local/fm_modulator/rtl/top.v(280[9] 288[53])
    defparam wb_idata_i10.GSR = "DISABLED";
    FD1S3AX wb_idata_i9 (.D(wb_idata_31__N_2[9]), .CK(dac_clk_p_c), .Q(wb_idata[9]));   // d:/documents/git_local/fm_modulator/rtl/top.v(280[9] 288[53])
    defparam wb_idata_i9.GSR = "DISABLED";
    FD1S3AX wb_idata_i8 (.D(wb_idata_31__N_2[8]), .CK(dac_clk_p_c), .Q(wb_idata[8]));   // d:/documents/git_local/fm_modulator/rtl/top.v(280[9] 288[53])
    defparam wb_idata_i8.GSR = "DISABLED";
    FD1S3AX wb_idata_i7 (.D(wb_idata_31__N_2[7]), .CK(dac_clk_p_c), .Q(wb_idata[7]));   // d:/documents/git_local/fm_modulator/rtl/top.v(280[9] 288[53])
    defparam wb_idata_i7.GSR = "DISABLED";
    FD1S3AX wb_idata_i6 (.D(wb_idata_31__N_2[6]), .CK(dac_clk_p_c), .Q(wb_idata[6]));   // d:/documents/git_local/fm_modulator/rtl/top.v(280[9] 288[53])
    defparam wb_idata_i6.GSR = "DISABLED";
    FD1S3AX wb_idata_i5 (.D(wb_idata_31__N_2[5]), .CK(dac_clk_p_c), .Q(wb_idata[5]));   // d:/documents/git_local/fm_modulator/rtl/top.v(280[9] 288[53])
    defparam wb_idata_i5.GSR = "DISABLED";
    FD1S3AX wb_idata_i4 (.D(wb_idata_31__N_2[4]), .CK(dac_clk_p_c), .Q(wb_idata[4]));   // d:/documents/git_local/fm_modulator/rtl/top.v(280[9] 288[53])
    defparam wb_idata_i4.GSR = "DISABLED";
    FD1S3AX wb_idata_i3 (.D(wb_idata_31__N_2[3]), .CK(dac_clk_p_c), .Q(wb_idata[3]));   // d:/documents/git_local/fm_modulator/rtl/top.v(280[9] 288[53])
    defparam wb_idata_i3.GSR = "DISABLED";
    FD1S3AX wb_idata_i2 (.D(wb_idata_31__N_2[2]), .CK(dac_clk_p_c), .Q(wb_idata[2]));   // d:/documents/git_local/fm_modulator/rtl/top.v(280[9] 288[53])
    defparam wb_idata_i2.GSR = "DISABLED";
    FD1S3AX wb_idata_i1 (.D(wb_idata_31__N_2[1]), .CK(dac_clk_p_c), .Q(wb_idata[1]));   // d:/documents/git_local/fm_modulator/rtl/top.v(280[9] 288[53])
    defparam wb_idata_i1.GSR = "DISABLED";
    sys_clk sys_clk_inst (.i_ref_clk_c(i_ref_clk_c), .dac_clk_p_c(dac_clk_p_c), 
            .GND_net(GND_net)) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(47[10:54])
    CCU2D add_31_31 (.A0(power_counter[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17856), .COUT(n17857), .S0(power_counter_31__N_232[29]), 
          .S1(power_counter_31__N_232[30]));   // d:/documents/git_local/fm_modulator/rtl/top.v(242[21:41])
    defparam add_31_31.INIT0 = 16'h5aaa;
    defparam add_31_31.INIT1 = 16'h5aaa;
    defparam add_31_31.INJECT1_0 = "NO";
    defparam add_31_31.INJECT1_1 = "NO";
    CCU2D add_31_11 (.A0(power_counter[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17846), .COUT(n17847), .S0(power_counter_31__N_232[9]), 
          .S1(power_counter_31__N_232[10]));   // d:/documents/git_local/fm_modulator/rtl/top.v(242[21:41])
    defparam add_31_11.INIT0 = 16'h5aaa;
    defparam add_31_11.INIT1 = 16'h5aaa;
    defparam add_31_11.INJECT1_0 = "NO";
    defparam add_31_11.INJECT1_1 = "NO";
    CCU2D add_31_29 (.A0(power_counter[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17855), .COUT(n17856), .S0(power_counter_31__N_232[27]), 
          .S1(power_counter_31__N_232[28]));   // d:/documents/git_local/fm_modulator/rtl/top.v(242[21:41])
    defparam add_31_29.INIT0 = 16'h5aaa;
    defparam add_31_29.INIT1 = 16'h5aaa;
    defparam add_31_29.INJECT1_0 = "NO";
    defparam add_31_29.INJECT1_1 = "NO";
    LUT4 m1_lut (.Z(n29969)) /* synthesis lut_function=1, syn_instantiated=1 */ ;
    defparam m1_lut.init = 16'hffff;
    FD1P3AX power_counter_i31 (.D(n29969), .SP(power_counter_31__N_232[31]), 
            .CK(dac_clk_p_c), .Q(power_counter[31])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(239[9] 244[54])
    defparam power_counter_i31.GSR = "DISABLED";
    FD1S3AX power_counter_i30 (.D(power_counter_31__N_129[30]), .CK(dac_clk_p_c), 
            .Q(power_counter[30])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(239[9] 244[54])
    defparam power_counter_i30.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i29 (.D(wb_addr[29]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[29])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[9] 272[31])
    defparam bus_err_address_i0_i29.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i28 (.D(wb_addr[28]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[28])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[9] 272[31])
    defparam bus_err_address_i0_i28.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i27 (.D(wb_addr[27]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[27])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[9] 272[31])
    defparam bus_err_address_i0_i27.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i26 (.D(wb_addr[26]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[26])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[9] 272[31])
    defparam bus_err_address_i0_i26.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i25 (.D(wb_addr[25]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[25])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[9] 272[31])
    defparam bus_err_address_i0_i25.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i24 (.D(wb_addr[24]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[24])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[9] 272[31])
    defparam bus_err_address_i0_i24.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i23 (.D(wb_addr[23]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[23])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[9] 272[31])
    defparam bus_err_address_i0_i23.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i22 (.D(wb_addr[22]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[22])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[9] 272[31])
    defparam bus_err_address_i0_i22.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i21 (.D(wb_addr[21]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[21])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[9] 272[31])
    defparam bus_err_address_i0_i21.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i20 (.D(wb_addr[20]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[20])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[9] 272[31])
    defparam bus_err_address_i0_i20.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i19 (.D(wb_addr[19]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[19])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[9] 272[31])
    defparam bus_err_address_i0_i19.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i18 (.D(wb_addr[18]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[18])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[9] 272[31])
    defparam bus_err_address_i0_i18.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i17 (.D(wb_addr[17]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[17])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[9] 272[31])
    defparam bus_err_address_i0_i17.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i16 (.D(wb_addr[16]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[16])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[9] 272[31])
    defparam bus_err_address_i0_i16.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i15 (.D(wb_addr[15]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[15])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[9] 272[31])
    defparam bus_err_address_i0_i15.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i14 (.D(wb_addr[14]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[14])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[9] 272[31])
    defparam bus_err_address_i0_i14.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i13 (.D(wb_addr[13]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[13])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[9] 272[31])
    defparam bus_err_address_i0_i13.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i12 (.D(wb_addr[12]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[12])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[9] 272[31])
    defparam bus_err_address_i0_i12.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i11 (.D(wb_addr[11]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[11])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[9] 272[31])
    defparam bus_err_address_i0_i11.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i10 (.D(wb_addr[10]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[10])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[9] 272[31])
    defparam bus_err_address_i0_i10.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i9 (.D(wb_addr[9]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[9])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[9] 272[31])
    defparam bus_err_address_i0_i9.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i8 (.D(wb_addr[8]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[8])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[9] 272[31])
    defparam bus_err_address_i0_i8.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i7 (.D(wb_addr[7]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[7])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[9] 272[31])
    defparam bus_err_address_i0_i7.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i6 (.D(wb_addr[6]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[6])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[9] 272[31])
    defparam bus_err_address_i0_i6.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i5 (.D(wb_addr[5]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[5])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[9] 272[31])
    defparam bus_err_address_i0_i5.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i4 (.D(wb_addr[4]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[4])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[9] 272[31])
    defparam bus_err_address_i0_i4.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i3 (.D(wb_addr[3]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[3])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[9] 272[31])
    defparam bus_err_address_i0_i3.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i2 (.D(wb_addr[2]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[2])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[9] 272[31])
    defparam bus_err_address_i0_i2.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i1 (.D(wb_addr[1]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[1])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[9] 272[31])
    defparam bus_err_address_i0_i1.GSR = "DISABLED";
    FD1S3AX power_counter_i29 (.D(power_counter_31__N_129[29]), .CK(dac_clk_p_c), 
            .Q(power_counter[29])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(239[9] 244[54])
    defparam power_counter_i29.GSR = "DISABLED";
    FD1S3AX power_counter_i28 (.D(power_counter_31__N_129[28]), .CK(dac_clk_p_c), 
            .Q(power_counter[28])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(239[9] 244[54])
    defparam power_counter_i28.GSR = "DISABLED";
    FD1S3AX power_counter_i27 (.D(power_counter_31__N_129[27]), .CK(dac_clk_p_c), 
            .Q(power_counter[27])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(239[9] 244[54])
    defparam power_counter_i27.GSR = "DISABLED";
    FD1S3AX power_counter_i26 (.D(power_counter_31__N_129[26]), .CK(dac_clk_p_c), 
            .Q(power_counter[26])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(239[9] 244[54])
    defparam power_counter_i26.GSR = "DISABLED";
    FD1S3AX power_counter_i25 (.D(power_counter_31__N_129[25]), .CK(dac_clk_p_c), 
            .Q(power_counter[25])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(239[9] 244[54])
    defparam power_counter_i25.GSR = "DISABLED";
    FD1S3AX power_counter_i24 (.D(power_counter_31__N_129[24]), .CK(dac_clk_p_c), 
            .Q(power_counter[24])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(239[9] 244[54])
    defparam power_counter_i24.GSR = "DISABLED";
    FD1S3AX power_counter_i23 (.D(power_counter_31__N_129[23]), .CK(dac_clk_p_c), 
            .Q(power_counter[23])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(239[9] 244[54])
    defparam power_counter_i23.GSR = "DISABLED";
    FD1S3AX power_counter_i22 (.D(power_counter_31__N_129[22]), .CK(dac_clk_p_c), 
            .Q(power_counter[22])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(239[9] 244[54])
    defparam power_counter_i22.GSR = "DISABLED";
    FD1S3AX power_counter_i21 (.D(power_counter_31__N_129[21]), .CK(dac_clk_p_c), 
            .Q(power_counter[21])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(239[9] 244[54])
    defparam power_counter_i21.GSR = "DISABLED";
    FD1S3AX power_counter_i20 (.D(power_counter_31__N_129[20]), .CK(dac_clk_p_c), 
            .Q(power_counter[20])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(239[9] 244[54])
    defparam power_counter_i20.GSR = "DISABLED";
    FD1S3AX power_counter_i19 (.D(power_counter_31__N_129[19]), .CK(dac_clk_p_c), 
            .Q(power_counter[19])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(239[9] 244[54])
    defparam power_counter_i19.GSR = "DISABLED";
    FD1S3AX power_counter_i18 (.D(power_counter_31__N_129[18]), .CK(dac_clk_p_c), 
            .Q(power_counter[18])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(239[9] 244[54])
    defparam power_counter_i18.GSR = "DISABLED";
    FD1S3AX power_counter_i17 (.D(power_counter_31__N_129[17]), .CK(dac_clk_p_c), 
            .Q(power_counter[17])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(239[9] 244[54])
    defparam power_counter_i17.GSR = "DISABLED";
    FD1S3AX power_counter_i16 (.D(power_counter_31__N_129[16]), .CK(dac_clk_p_c), 
            .Q(power_counter[16])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(239[9] 244[54])
    defparam power_counter_i16.GSR = "DISABLED";
    FD1S3AX power_counter_i15 (.D(power_counter_31__N_129[15]), .CK(dac_clk_p_c), 
            .Q(power_counter[15])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(239[9] 244[54])
    defparam power_counter_i15.GSR = "DISABLED";
    FD1S3AX power_counter_i14 (.D(power_counter_31__N_129[14]), .CK(dac_clk_p_c), 
            .Q(power_counter[14])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(239[9] 244[54])
    defparam power_counter_i14.GSR = "DISABLED";
    FD1S3AX power_counter_i13 (.D(power_counter_31__N_129[13]), .CK(dac_clk_p_c), 
            .Q(power_counter[13])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(239[9] 244[54])
    defparam power_counter_i13.GSR = "DISABLED";
    FD1S3AX power_counter_i12 (.D(power_counter_31__N_129[12]), .CK(dac_clk_p_c), 
            .Q(power_counter[12])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(239[9] 244[54])
    defparam power_counter_i12.GSR = "DISABLED";
    FD1S3AX power_counter_i11 (.D(power_counter_31__N_129[11]), .CK(dac_clk_p_c), 
            .Q(power_counter[11])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(239[9] 244[54])
    defparam power_counter_i11.GSR = "DISABLED";
    FD1S3AX power_counter_i10 (.D(power_counter_31__N_129[10]), .CK(dac_clk_p_c), 
            .Q(power_counter[10])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(239[9] 244[54])
    defparam power_counter_i10.GSR = "DISABLED";
    FD1S3AX power_counter_i9 (.D(power_counter_31__N_129[9]), .CK(dac_clk_p_c), 
            .Q(power_counter[9])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(239[9] 244[54])
    defparam power_counter_i9.GSR = "DISABLED";
    FD1S3AX power_counter_i8 (.D(power_counter_31__N_129[8]), .CK(dac_clk_p_c), 
            .Q(power_counter[8])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(239[9] 244[54])
    defparam power_counter_i8.GSR = "DISABLED";
    FD1S3AX power_counter_i7 (.D(power_counter_31__N_129[7]), .CK(dac_clk_p_c), 
            .Q(power_counter[7])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(239[9] 244[54])
    defparam power_counter_i7.GSR = "DISABLED";
    FD1S3AX power_counter_i6 (.D(power_counter_31__N_129[6]), .CK(dac_clk_p_c), 
            .Q(power_counter[6])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(239[9] 244[54])
    defparam power_counter_i6.GSR = "DISABLED";
    FD1S3AX power_counter_i5 (.D(power_counter_31__N_129[5]), .CK(dac_clk_p_c), 
            .Q(power_counter[5])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(239[9] 244[54])
    defparam power_counter_i5.GSR = "DISABLED";
    FD1S3AX power_counter_i4 (.D(power_counter_31__N_129[4]), .CK(dac_clk_p_c), 
            .Q(power_counter[4])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(239[9] 244[54])
    defparam power_counter_i4.GSR = "DISABLED";
    FD1S3AX power_counter_i3 (.D(power_counter_31__N_129[3]), .CK(dac_clk_p_c), 
            .Q(power_counter[3])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(239[9] 244[54])
    defparam power_counter_i3.GSR = "DISABLED";
    FD1S3AX power_counter_i2 (.D(power_counter_31__N_129[2]), .CK(dac_clk_p_c), 
            .Q(power_counter[2])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(239[9] 244[54])
    defparam power_counter_i2.GSR = "DISABLED";
    FD1S3AX power_counter_i1 (.D(power_counter_31__N_129[1]), .CK(dac_clk_p_c), 
            .Q(power_counter[1])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(239[9] 244[54])
    defparam power_counter_i1.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i31 (.D(n2092), .CK(dac_clk_p_c), .CD(n27444), 
            .Q(wb_smpl_data[31]));   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 235[10])
    defparam wb_smpl_data_i31.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i30 (.D(n2093), .CK(dac_clk_p_c), .CD(n27444), 
            .Q(wb_smpl_data[30]));   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 235[10])
    defparam wb_smpl_data_i30.GSR = "DISABLED";
    dynamic_pll lo_gen (.i_clk_2f_N_2268(i_clk_2f_N_2268), .lo_pll_out(lo_pll_out), 
            .i_ref_clk_c(i_ref_clk_c), .pll_clk(pll_clk), .pll_rst(pll_rst), 
            .pll_stb(pll_stb), .pll_we(pll_we), .pll_data_i({pll_data_i}), 
            .pll_addr({pll_addr}), .pll_data_o({pll_data_o}), .pll_ack(pll_ack), 
            .GND_net(GND_net)) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(174[14] 185[5])
    LUT4 m0_lut (.Z(n29968)) /* synthesis lut_function=0, syn_instantiated=1 */ ;
    defparam m0_lut.init = 16'h0000;
    OB o_dac_a_pad_5 (.I(o_dac_a_c_5), .O(o_dac_a[5]));   // d:/documents/git_local/fm_modulator/rtl/top.v(33[38:45])
    OB o_dac_a_pad_4 (.I(o_dac_a_c_4), .O(o_dac_a[4]));   // d:/documents/git_local/fm_modulator/rtl/top.v(33[38:45])
    OB o_dac_a_pad_3 (.I(o_dac_a_c_3), .O(o_dac_a[3]));   // d:/documents/git_local/fm_modulator/rtl/top.v(33[38:45])
    OB o_dac_a_pad_2 (.I(o_dac_a_c_2), .O(o_dac_a[2]));   // d:/documents/git_local/fm_modulator/rtl/top.v(33[38:45])
    OB o_dac_a_pad_1 (.I(o_dac_a_c_1), .O(o_dac_a[1]));   // d:/documents/git_local/fm_modulator/rtl/top.v(33[38:45])
    OB o_dac_a_pad_0 (.I(o_dac_a_c_0), .O(o_dac_a[0]));   // d:/documents/git_local/fm_modulator/rtl/top.v(33[38:45])
    OB o_dac_b_pad_9 (.I(o_dac_b_c_9), .O(o_dac_b[9]));   // d:/documents/git_local/fm_modulator/rtl/top.v(33[47:54])
    OB o_dac_b_pad_8 (.I(o_dac_b_c_15), .O(o_dac_b[8]));   // d:/documents/git_local/fm_modulator/rtl/top.v(33[47:54])
    OB o_dac_b_pad_7 (.I(o_dac_b_c_14), .O(o_dac_b[7]));   // d:/documents/git_local/fm_modulator/rtl/top.v(33[47:54])
    OB o_dac_b_pad_6 (.I(o_dac_b_c_13), .O(o_dac_b[6]));   // d:/documents/git_local/fm_modulator/rtl/top.v(33[47:54])
    OB o_dac_b_pad_5 (.I(o_dac_b_c_12), .O(o_dac_b[5]));   // d:/documents/git_local/fm_modulator/rtl/top.v(33[47:54])
    OB o_dac_b_pad_4 (.I(o_dac_b_c_11), .O(o_dac_b[4]));   // d:/documents/git_local/fm_modulator/rtl/top.v(33[47:54])
    OB o_dac_b_pad_3 (.I(o_dac_b_c_10), .O(o_dac_b[3]));   // d:/documents/git_local/fm_modulator/rtl/top.v(33[47:54])
    OB o_dac_b_pad_2 (.I(n3639), .O(o_dac_b[2]));   // d:/documents/git_local/fm_modulator/rtl/top.v(33[47:54])
    OB o_dac_b_pad_1 (.I(o_dac_b_c_8), .O(o_dac_b[1]));   // d:/documents/git_local/fm_modulator/rtl/top.v(33[47:54])
    OB o_dac_b_pad_0 (.I(o_dac_b_c_7), .O(o_dac_b[0]));   // d:/documents/git_local/fm_modulator/rtl/top.v(33[47:54])
    OB dac_clk_p_pad (.I(dac_clk_p_c), .O(dac_clk_p));   // d:/documents/git_local/fm_modulator/rtl/top.v(34[49:58])
    OB dac_clk_n_pad (.I(dac_clk_n_c), .O(dac_clk_n));   // d:/documents/git_local/fm_modulator/rtl/top.v(34[60:69])
    OB o_dac_cw_b_pad (.I(o_dac_cw_b_c), .O(o_dac_cw_b));   // d:/documents/git_local/fm_modulator/rtl/top.v(34[71:81])
    OB i_clk_p_pad (.I(i_clk_p_c), .O(i_clk_p));   // d:/documents/git_local/fm_modulator/rtl/top.v(34[13:20])
    OB i_clk_n_pad (.I(i_clk_n_c), .O(i_clk_n));   // d:/documents/git_local/fm_modulator/rtl/top.v(34[22:29])
    OB q_clk_p_pad (.I(q_clk_p_c), .O(q_clk_p));   // d:/documents/git_local/fm_modulator/rtl/top.v(34[31:38])
    OB q_clk_n_pad (.I(q_clk_n_c), .O(q_clk_n));   // d:/documents/git_local/fm_modulator/rtl/top.v(34[40:47])
    IB i_ref_clk_pad (.I(i_ref_clk), .O(i_ref_clk_c));   // d:/documents/git_local/fm_modulator/rtl/top.v(26[12:21])
    IB i_wbu_uart_rx_pad (.I(i_wbu_uart_rx), .O(i_wbu_uart_rx_c));   // d:/documents/git_local/fm_modulator/rtl/top.v(28[12:25])
    IB i_sw0_pad (.I(i_sw0), .O(i_sw0_c));   // d:/documents/git_local/fm_modulator/rtl/top.v(31[12:17])
    FD1S3IX wb_smpl_data_i11 (.D(n2112), .CK(dac_clk_p_c), .CD(n27444), 
            .Q(wb_smpl_data[11]));   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 235[10])
    defparam wb_smpl_data_i11.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i29 (.D(n27056), .CK(dac_clk_p_c), .CD(n27444), 
            .Q(wb_smpl_data[29]));   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 235[10])
    defparam wb_smpl_data_i29.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i10 (.D(n27051), .CK(dac_clk_p_c), .CD(n27444), 
            .Q(wb_smpl_data[10]));   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 235[10])
    defparam wb_smpl_data_i10.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i28 (.D(n2095), .CK(dac_clk_p_c), .CD(n27444), 
            .Q(wb_smpl_data[28]));   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 235[10])
    defparam wb_smpl_data_i28.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i9 (.D(n27050), .CK(dac_clk_p_c), .CD(n27444), 
            .Q(wb_smpl_data[9]));   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 235[10])
    defparam wb_smpl_data_i9.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i27 (.D(n2096), .CK(dac_clk_p_c), .CD(n27444), 
            .Q(wb_smpl_data[27]));   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 235[10])
    defparam wb_smpl_data_i27.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i8 (.D(n2115), .CK(dac_clk_p_c), .CD(n27444), 
            .Q(wb_smpl_data[8]));   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 235[10])
    defparam wb_smpl_data_i8.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i26 (.D(n2097), .CK(dac_clk_p_c), .CD(n27444), 
            .Q(wb_smpl_data[26]));   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 235[10])
    defparam wb_smpl_data_i26.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i7 (.D(n2116), .CK(dac_clk_p_c), .CD(n27444), 
            .Q(wb_smpl_data[7]));   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 235[10])
    defparam wb_smpl_data_i7.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i25 (.D(n2098), .CK(dac_clk_p_c), .CD(n27444), 
            .Q(wb_smpl_data[25]));   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 235[10])
    defparam wb_smpl_data_i25.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i6 (.D(n2117), .CK(dac_clk_p_c), .CD(n27444), 
            .Q(wb_smpl_data[6]));   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 235[10])
    defparam wb_smpl_data_i6.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i24 (.D(n2099), .CK(dac_clk_p_c), .CD(n27444), 
            .Q(wb_smpl_data[24]));   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 235[10])
    defparam wb_smpl_data_i24.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i5 (.D(n27049), .CK(dac_clk_p_c), .CD(n27444), 
            .Q(wb_smpl_data[5]));   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 235[10])
    defparam wb_smpl_data_i5.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i23 (.D(n2100), .CK(dac_clk_p_c), .CD(n27444), 
            .Q(wb_smpl_data[23]));   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 235[10])
    defparam wb_smpl_data_i23.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i4 (.D(n2119), .CK(dac_clk_p_c), .CD(n27444), 
            .Q(wb_smpl_data[4]));   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 235[10])
    defparam wb_smpl_data_i4.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i22 (.D(n2101), .CK(dac_clk_p_c), .CD(n27444), 
            .Q(wb_smpl_data[22]));   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 235[10])
    defparam wb_smpl_data_i22.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i3 (.D(n2120), .CK(dac_clk_p_c), .CD(n27444), 
            .Q(wb_smpl_data[3]));   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 235[10])
    defparam wb_smpl_data_i3.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i21 (.D(n2102), .CK(dac_clk_p_c), .CD(n27444), 
            .Q(wb_smpl_data[21]));   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 235[10])
    defparam wb_smpl_data_i21.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i2 (.D(n2121), .CK(dac_clk_p_c), .CD(n27444), 
            .Q(wb_smpl_data[2]));   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 235[10])
    defparam wb_smpl_data_i2.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i20 (.D(n27061), .CK(dac_clk_p_c), .CD(n27444), 
            .Q(wb_smpl_data[20]));   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 235[10])
    defparam wb_smpl_data_i20.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i1 (.D(n2122), .CK(dac_clk_p_c), .CD(n27444), 
            .Q(wb_smpl_data[1]));   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 235[10])
    defparam wb_smpl_data_i1.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i19 (.D(n2104), .CK(dac_clk_p_c), .CD(n27444), 
            .Q(wb_smpl_data[19]));   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 235[10])
    defparam wb_smpl_data_i19.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i18 (.D(n27059), .CK(dac_clk_p_c), .CD(n27444), 
            .Q(wb_smpl_data[18]));   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 235[10])
    defparam wb_smpl_data_i18.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i17 (.D(n27058), .CK(dac_clk_p_c), .CD(n27444), 
            .Q(wb_smpl_data[17]));   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 235[10])
    defparam wb_smpl_data_i17.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i16 (.D(n27057), .CK(dac_clk_p_c), .CD(n27444), 
            .Q(wb_smpl_data[16]));   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 235[10])
    defparam wb_smpl_data_i16.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i15 (.D(n2108), .CK(dac_clk_p_c), .CD(n27444), 
            .Q(wb_smpl_data[15]));   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 235[10])
    defparam wb_smpl_data_i15.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i14 (.D(n2109), .CK(dac_clk_p_c), .CD(n27444), 
            .Q(wb_smpl_data[14]));   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 235[10])
    defparam wb_smpl_data_i14.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i13 (.D(n2110), .CK(dac_clk_p_c), .CD(n27444), 
            .Q(wb_smpl_data[13]));   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 235[10])
    defparam wb_smpl_data_i13.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i12 (.D(n2111), .CK(dac_clk_p_c), .CD(n27444), 
            .Q(wb_smpl_data[12]));   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 235[10])
    defparam wb_smpl_data_i12.GSR = "DISABLED";
    fm_generator_wb_slave o_dac_a_9__I_0 (.dac_clk_p_c(dac_clk_p_c), .wb_odata({wb_odata}), 
            .i_sw0_c(i_sw0_c), .wb_fm_data({wb_fm_data}), .wb_fm_ack(wb_fm_ack), 
            .o_dac_a_9__N_1(o_dac_a_9__N_1), .\wb_addr[0] (wb_addr[0]), 
            .\wb_addr[1] (wb_addr[1]), .\power_counter[1] (power_counter[1]), 
            .\smpl_register[1] (smpl_register[1]), .n2122(n2122), .n27114(n27114), 
            .n27304(n27304), .n27313(n27313), .\wb_addr[15] (wb_addr[15]), 
            .\wb_addr[8] (wb_addr[8]), .\wb_addr[12] (wb_addr[12]), .GND_net(GND_net), 
            .o_dac_a_c_7(o_dac_a_c_7), .o_dac_a_c_6(o_dac_a_c_6), .o_dac_a_c_5(o_dac_a_c_5), 
            .o_dac_a_c_4(o_dac_a_c_4), .o_dac_a_c_3(o_dac_a_c_3), .o_dac_a_c_2(o_dac_a_c_2), 
            .o_dac_a_c_1(o_dac_a_c_1), .o_dac_a_c_0(o_dac_a_c_0), .o_dac_b_c_15(o_dac_b_c_15), 
            .o_dac_b_c_9(o_dac_b_c_9), .o_dac_cw_b_c(o_dac_cw_b_c), .n27380(n27380), 
            .o_dac_a_c_9(o_dac_a_c_9), .n21102(n21102), .n38(n38), .n2(n2_adj_3086), 
            .\smpl_register[5] (smpl_register[5]), .n27049(n27049), .n2_adj_1(n2_adj_3062), 
            .\smpl_register[20] (smpl_register[20]), .n27061(n27061), .n2_adj_2(n2_adj_3065), 
            .\smpl_register[18] (smpl_register[18]), .n27059(n27059), .n2_adj_3(n2_adj_3066), 
            .\smpl_register[17] (smpl_register[17]), .n27058(n27058), .n2_adj_4(n2_adj_3067), 
            .\smpl_register[16] (smpl_register[16]), .n27057(n27057), .n2_adj_5(n2_adj_3045), 
            .\smpl_register[29] (smpl_register[29]), .n27056(n27056), .n2_adj_6(n2_adj_3078), 
            .\smpl_register[10] (smpl_register[10]), .n27051(n27051), .n2_adj_7(n2_adj_3079), 
            .\smpl_register[9] (smpl_register[9]), .n27050(n27050), .n21088(n21088), 
            .n21078(n21078), .n21044(n21044), .n29969(n29969), .o_dac_b_c_7(o_dac_b_c_7), 
            .n29968(n29968), .o_dac_b_c_14(o_dac_b_c_14), .o_dac_b_c_13(o_dac_b_c_13), 
            .o_dac_b_c_12(o_dac_b_c_12), .o_dac_b_c_11(o_dac_b_c_11), .o_dac_b_c_10(o_dac_b_c_10), 
            .n3639(n3639), .o_dac_b_c_8(o_dac_b_c_8)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(129[2] 141[2])
    
endmodule
//
// Verilog Description of module hbbus
//

module hbbus (dac_clk_p_c, wb_cyc, wb_odata, wb_we, wb_stb, wb_err, 
            wb_ack, \wb_idata[0] , wb_addr, \wb_idata[2] , \wb_idata[3] , 
            \wb_idata[4] , \wb_idata[5] , \wb_idata[6] , \wb_idata[7] , 
            \wb_idata[8] , \wb_idata[9] , \wb_idata[10] , \wb_idata[11] , 
            \wb_idata[12] , \wb_idata[13] , \wb_idata[14] , \wb_idata[15] , 
            \wb_idata[16] , \wb_idata[17] , \wb_idata[18] , \wb_idata[19] , 
            \wb_idata[20] , \wb_idata[21] , \wb_idata[22] , \wb_idata[23] , 
            \wb_idata[24] , \wb_idata[25] , \wb_idata[26] , \wb_idata[27] , 
            \wb_idata[28] , \wb_idata[29] , \wb_idata[30] , \wb_idata[31] , 
            n2, GND_net, n12753, n29969, VCC_net, rx_stb, \rx_data[3] , 
            \rx_data[6] , \rx_data[2] , \rx_data[4] , \rx_data[5] , 
            \rx_data[0] , \rx_data[1] , tx_busy, n27281, \lcl_data[1] , 
            \lcl_data_7__N_510[0] , zero_baud_counter, dac_clk_p_c_enable_346, 
            \lcl_data[4] , \lcl_data_7__N_510[3] , \lcl_data[7] , \lcl_data_7__N_510[6] , 
            \lcl_data[6] , \lcl_data_7__N_510[5] , \lcl_data[5] , \lcl_data_7__N_510[4] , 
            \lcl_data[3] , \lcl_data_7__N_510[2] , \lcl_data[2] , \lcl_data_7__N_510[1] , 
            o_busy_N_535, \state[0] , n18134) /* synthesis syn_module_defined=1 */ ;
    input dac_clk_p_c;
    output wb_cyc;
    output [31:0]wb_odata;
    output wb_we;
    output wb_stb;
    input wb_err;
    input wb_ack;
    input \wb_idata[0] ;
    output [29:0]wb_addr;
    input \wb_idata[2] ;
    input \wb_idata[3] ;
    input \wb_idata[4] ;
    input \wb_idata[5] ;
    input \wb_idata[6] ;
    input \wb_idata[7] ;
    input \wb_idata[8] ;
    input \wb_idata[9] ;
    input \wb_idata[10] ;
    input \wb_idata[11] ;
    input \wb_idata[12] ;
    input \wb_idata[13] ;
    input \wb_idata[14] ;
    input \wb_idata[15] ;
    input \wb_idata[16] ;
    input \wb_idata[17] ;
    input \wb_idata[18] ;
    input \wb_idata[19] ;
    input \wb_idata[20] ;
    input \wb_idata[21] ;
    input \wb_idata[22] ;
    input \wb_idata[23] ;
    input \wb_idata[24] ;
    input \wb_idata[25] ;
    input \wb_idata[26] ;
    input \wb_idata[27] ;
    input \wb_idata[28] ;
    input \wb_idata[29] ;
    input \wb_idata[30] ;
    input \wb_idata[31] ;
    output n2;
    input GND_net;
    input n12753;
    input n29969;
    input VCC_net;
    input rx_stb;
    input \rx_data[3] ;
    input \rx_data[6] ;
    input \rx_data[2] ;
    input \rx_data[4] ;
    input \rx_data[5] ;
    input \rx_data[0] ;
    input \rx_data[1] ;
    input tx_busy;
    output n27281;
    input \lcl_data[1] ;
    output \lcl_data_7__N_510[0] ;
    input zero_baud_counter;
    output dac_clk_p_c_enable_346;
    input \lcl_data[4] ;
    output \lcl_data_7__N_510[3] ;
    input \lcl_data[7] ;
    output \lcl_data_7__N_510[6] ;
    input \lcl_data[6] ;
    output \lcl_data_7__N_510[5] ;
    input \lcl_data[5] ;
    output \lcl_data_7__N_510[4] ;
    input \lcl_data[3] ;
    output \lcl_data_7__N_510[2] ;
    input \lcl_data[2] ;
    output \lcl_data_7__N_510[1] ;
    input o_busy_N_535;
    input \state[0] ;
    output n18134;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[49:58])
    
    wire newaddr_N_989;
    wire [33:0]iw_word;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(71[14:21])
    
    wire inc, dac_clk_p_c_enable_138, ow_stb;
    wire [33:0]ow_word;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(73[14:21])
    
    wire n30028, i_cmd_wr, n22542, n30027, n17754, n27423, n27443, 
        dac_clk_p_c_enable_471, dac_clk_p_c_enable_332;
    wire [4:0]hb_bits;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(79[13:20])
    
    wire dac_clk_p_c_enable_219;
    wire [33:0]idl_word;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(77[14:22])
    
    wire hb_busy, w_reset, idl_stb, n27258, nl_busy, hx_stb, dac_clk_p_c_enable_405;
    wire [4:0]dec_bits;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(69[13:21])
    
    wire o_pck_stb_N_764, cmd_loaded, dac_clk_p_c_enable_222, cmd_loaded_N_767, 
        dac_clk_p_c_enable_374;
    wire [33:0]n14;
    wire [7:0]w_gx_char;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbgenhex.v(80[12:21])
    
    wire n11763;
    wire [33:0]int_word;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(75[14:22])
    
    wire dac_clk_p_c_enable_442, n12767, n27315, n27249, int_stb;
    
    hbexec wbexec (.dac_clk_p_c(dac_clk_p_c), .wb_cyc(wb_cyc), .newaddr_N_989(newaddr_N_989), 
           .wb_odata({wb_odata}), .\iw_word[0] (iw_word[0]), .inc(inc), 
           .dac_clk_p_c_enable_138(dac_clk_p_c_enable_138), .ow_stb(ow_stb), 
           .ow_word({ow_word}), .n30028(n30028), .wb_we(wb_we), .i_cmd_wr(i_cmd_wr), 
           .wb_stb(wb_stb), .n22542(n22542), .\iw_word[31] (iw_word[31]), 
           .\iw_word[1] (iw_word[1]), .\iw_word[30] (iw_word[30]), .\iw_word[28] (iw_word[28]), 
           .\iw_word[29] (iw_word[29]), .\iw_word[26] (iw_word[26]), .\iw_word[27] (iw_word[27]), 
           .\iw_word[24] (iw_word[24]), .\iw_word[25] (iw_word[25]), .\iw_word[22] (iw_word[22]), 
           .\iw_word[23] (iw_word[23]), .\iw_word[20] (iw_word[20]), .\iw_word[21] (iw_word[21]), 
           .\iw_word[18] (iw_word[18]), .\iw_word[19] (iw_word[19]), .\iw_word[16] (iw_word[16]), 
           .\iw_word[17] (iw_word[17]), .wb_err(wb_err), .n30027(n30027), 
           .wb_ack(wb_ack), .\iw_word[14] (iw_word[14]), .\iw_word[15] (iw_word[15]), 
           .\wb_idata[0] (\wb_idata[0] ), .wb_addr({wb_addr}), .\wb_idata[2] (\wb_idata[2] ), 
           .\wb_idata[3] (\wb_idata[3] ), .\wb_idata[4] (\wb_idata[4] ), 
           .\wb_idata[5] (\wb_idata[5] ), .\wb_idata[6] (\wb_idata[6] ), 
           .\wb_idata[7] (\wb_idata[7] ), .\wb_idata[8] (\wb_idata[8] ), 
           .\wb_idata[9] (\wb_idata[9] ), .\wb_idata[10] (\wb_idata[10] ), 
           .\wb_idata[11] (\wb_idata[11] ), .\wb_idata[12] (\wb_idata[12] ), 
           .\wb_idata[13] (\wb_idata[13] ), .\wb_idata[14] (\wb_idata[14] ), 
           .\wb_idata[15] (\wb_idata[15] ), .\wb_idata[16] (\wb_idata[16] ), 
           .\wb_idata[17] (\wb_idata[17] ), .\wb_idata[18] (\wb_idata[18] ), 
           .\wb_idata[19] (\wb_idata[19] ), .\iw_word[12] (iw_word[12]), 
           .\iw_word[13] (iw_word[13]), .\wb_idata[20] (\wb_idata[20] ), 
           .\wb_idata[21] (\wb_idata[21] ), .\wb_idata[22] (\wb_idata[22] ), 
           .\wb_idata[23] (\wb_idata[23] ), .\wb_idata[24] (\wb_idata[24] ), 
           .\wb_idata[25] (\wb_idata[25] ), .\wb_idata[26] (\wb_idata[26] ), 
           .\iw_word[10] (iw_word[10]), .\iw_word[11] (iw_word[11]), .\wb_idata[27] (\wb_idata[27] ), 
           .\wb_idata[28] (\wb_idata[28] ), .\wb_idata[29] (\wb_idata[29] ), 
           .\wb_idata[30] (\wb_idata[30] ), .\wb_idata[31] (\wb_idata[31] ), 
           .\iw_word[8] (iw_word[8]), .\iw_word[9] (iw_word[9]), .\iw_word[6] (iw_word[6]), 
           .\iw_word[7] (iw_word[7]), .\iw_word[5] (iw_word[5]), .\iw_word[4] (iw_word[4]), 
           .\iw_word[3] (iw_word[3]), .\iw_word[2] (iw_word[2]), .n2(n2), 
           .n17754(n17754), .GND_net(GND_net), .n27423(n27423), .\iw_word[32] (iw_word[32]), 
           .n27443(n27443), .dac_clk_p_c_enable_471(dac_clk_p_c_enable_471), 
           .n12753(n12753)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(105[15] 109[15])
    hbdeword unpackx (.dac_clk_p_c(dac_clk_p_c), .dac_clk_p_c_enable_332(dac_clk_p_c_enable_332), 
            .hb_bits({hb_bits}), .dac_clk_p_c_enable_219(dac_clk_p_c_enable_219), 
            .n30028(n30028), .idl_word({idl_word}), .n29969(n29969), .hb_busy(hb_busy), 
            .w_reset(w_reset), .idl_stb(idl_stb), .n27258(n27258), .nl_busy(nl_busy), 
            .hx_stb(hx_stb), .n30027(n30027)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(127[11] 129[29])
    hbpack packxi (.iw_word({Open_3, iw_word[32], Open_4, Open_5, Open_6, 
           Open_7, Open_8, Open_9, Open_10, Open_11, Open_12, Open_13, 
           Open_14, Open_15, Open_16, Open_17, Open_18, Open_19, 
           Open_20, Open_21, Open_22, Open_23, Open_24, Open_25, 
           Open_26, Open_27, Open_28, Open_29, Open_30, Open_31, 
           Open_32, Open_33, Open_34, iw_word[0]}), .n27423(n27423), 
           .wb_stb(wb_stb), .wb_cyc(wb_cyc), .dac_clk_p_c_enable_471(dac_clk_p_c_enable_471), 
           .dac_clk_p_c(dac_clk_p_c), .dac_clk_p_c_enable_405(dac_clk_p_c_enable_405), 
           .n30028(n30028), .\dec_bits[1] (dec_bits[1]), .\dec_bits[4] (dec_bits[4]), 
           .w_reset(w_reset), .o_pck_stb_N_764(o_pck_stb_N_764), .cmd_loaded(cmd_loaded), 
           .dac_clk_p_c_enable_222(dac_clk_p_c_enable_222), .cmd_loaded_N_767(cmd_loaded_N_767), 
           .n27443(n27443), .i_cmd_wr(i_cmd_wr), .n22542(n22542), .\iw_word[2] (iw_word[2]), 
           .inc(inc), .n17754(n17754), .\iw_word[31] (iw_word[31]), .\iw_word[30] (iw_word[30]), 
           .\iw_word[29] (iw_word[29]), .\iw_word[28] (iw_word[28]), .\iw_word[27] (iw_word[27]), 
           .\iw_word[26] (iw_word[26]), .\iw_word[25] (iw_word[25]), .\iw_word[24] (iw_word[24]), 
           .\iw_word[23] (iw_word[23]), .\iw_word[22] (iw_word[22]), .\iw_word[21] (iw_word[21]), 
           .\iw_word[20] (iw_word[20]), .\iw_word[19] (iw_word[19]), .\iw_word[18] (iw_word[18]), 
           .\iw_word[17] (iw_word[17]), .\iw_word[16] (iw_word[16]), .\iw_word[15] (iw_word[15]), 
           .\iw_word[14] (iw_word[14]), .\iw_word[13] (iw_word[13]), .\iw_word[12] (iw_word[12]), 
           .\iw_word[11] (iw_word[11]), .\iw_word[10] (iw_word[10]), .\iw_word[9] (iw_word[9]), 
           .\iw_word[8] (iw_word[8]), .\iw_word[7] (iw_word[7]), .\iw_word[6] (iw_word[6]), 
           .\iw_word[5] (iw_word[5]), .\iw_word[4] (iw_word[4]), .\iw_word[3] (iw_word[3]), 
           .\iw_word[1] (iw_word[1]), .\dec_bits[0] (dec_bits[0]), .dac_clk_p_c_enable_374(dac_clk_p_c_enable_374), 
           .n45(n14[3]), .n46(n14[2]), .dac_clk_p_c_enable_138(dac_clk_p_c_enable_138), 
           .n30027(n30027), .newaddr_N_989(newaddr_N_989)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(99[9] 100[38])
    hbgenhex genhex (.hx_stb(hx_stb), .dac_clk_p_c(dac_clk_p_c), .n30028(n30028), 
            .hb_busy(hb_busy), .hb_bits({hb_bits}), .\w_gx_char[0] (w_gx_char[0]), 
            .\w_gx_char[1] (w_gx_char[1]), .\w_gx_char[2] (w_gx_char[2]), 
            .\w_gx_char[3] (w_gx_char[3]), .\w_gx_char[4] (w_gx_char[4]), 
            .\w_gx_char[5] (w_gx_char[5]), .\w_gx_char[6] (w_gx_char[6]), 
            .dac_clk_p_c_enable_332(dac_clk_p_c_enable_332), .GND_net(GND_net), 
            .VCC_net(VCC_net), .n11763(n11763), .nl_busy(nl_busy), .n30027(n30027), 
            .n27258(n27258), .dac_clk_p_c_enable_219(dac_clk_p_c_enable_219)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(132[11] 133[29])
    hbdechex dechxi (.dac_clk_p_c(dac_clk_p_c), .dec_bits({dec_bits[4], 
            Open_35, Open_36, Open_37, Open_38}), .n45(n14[3]), .\dec_bits[0] (dec_bits[0]), 
            .w_reset(w_reset), .n46(n14[2]), .rx_stb(rx_stb), .\rx_data[3] (\rx_data[3] ), 
            .\rx_data[6] (\rx_data[6] ), .\rx_data[2] (\rx_data[2] ), .\rx_data[4] (\rx_data[4] ), 
            .\rx_data[5] (\rx_data[5] ), .\rx_data[0] (\rx_data[0] ), .\rx_data[1] (\rx_data[1] ), 
            .n30028(n30028), .\dec_bits[1] (dec_bits[1]), .n30027(n30027), 
            .cmd_loaded(cmd_loaded), .o_pck_stb_N_764(o_pck_stb_N_764), 
            .dac_clk_p_c_enable_222(dac_clk_p_c_enable_222), .cmd_loaded_N_767(cmd_loaded_N_767), 
            .dac_clk_p_c_enable_405(dac_clk_p_c_enable_405), .dac_clk_p_c_enable_374(dac_clk_p_c_enable_374)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(93[11] 95[30])
    hbnewline addnl (.dac_clk_p_c(dac_clk_p_c), .n30028(n30028), .w_reset(w_reset), 
            .hx_stb(hx_stb), .tx_busy(tx_busy), .nl_busy(nl_busy), .\w_gx_char[2] (w_gx_char[2]), 
            .\w_gx_char[0] (w_gx_char[0]), .\w_gx_char[4] (w_gx_char[4]), 
            .n30027(n30027), .\w_gx_char[3] (w_gx_char[3]), .\w_gx_char[5] (w_gx_char[5]), 
            .\w_gx_char[1] (w_gx_char[1]), .\w_gx_char[6] (w_gx_char[6]), 
            .n11763(n11763), .n27281(n27281), .\lcl_data[1] (\lcl_data[1] ), 
            .\lcl_data_7__N_510[0] (\lcl_data_7__N_510[0] ), .zero_baud_counter(zero_baud_counter), 
            .dac_clk_p_c_enable_346(dac_clk_p_c_enable_346), .\lcl_data[4] (\lcl_data[4] ), 
            .\lcl_data_7__N_510[3] (\lcl_data_7__N_510[3] ), .\lcl_data[7] (\lcl_data[7] ), 
            .\lcl_data_7__N_510[6] (\lcl_data_7__N_510[6] ), .\lcl_data[6] (\lcl_data[6] ), 
            .\lcl_data_7__N_510[5] (\lcl_data_7__N_510[5] ), .\lcl_data[5] (\lcl_data[5] ), 
            .\lcl_data_7__N_510[4] (\lcl_data_7__N_510[4] ), .\lcl_data[3] (\lcl_data[3] ), 
            .\lcl_data_7__N_510[2] (\lcl_data_7__N_510[2] ), .\lcl_data[2] (\lcl_data[2] ), 
            .\lcl_data_7__N_510[1] (\lcl_data_7__N_510[1] ), .o_busy_N_535(o_busy_N_535), 
            .\state[0] (\state[0] ), .n18134(n18134)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(138[12] 139[40])
    hbints addints (.int_word({int_word}), .dac_clk_p_c(dac_clk_p_c), .dac_clk_p_c_enable_442(dac_clk_p_c_enable_442), 
           .n12767(n12767), .ow_word({ow_word}), .n30027(n30027), .n27315(n27315), 
           .n27249(n27249), .int_stb(int_stb), .ow_stb(ow_stb), .n30028(n30028)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(114[9] 116[32])
    hbidle addidles (.idl_word({idl_word}), .dac_clk_p_c(dac_clk_p_c), .int_word({int_word}), 
           .idl_stb(idl_stb), .w_reset(w_reset), .hb_busy(hb_busy), .int_stb(int_stb), 
           .n27249(n27249), .n30027(n30027), .n27315(n27315), .dac_clk_p_c_enable_442(dac_clk_p_c_enable_442), 
           .n12767(n12767)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(121[9] 123[31])
    
endmodule
//
// Verilog Description of module hbexec
//

module hbexec (dac_clk_p_c, wb_cyc, newaddr_N_989, wb_odata, \iw_word[0] , 
            inc, dac_clk_p_c_enable_138, ow_stb, ow_word, n30028, 
            wb_we, i_cmd_wr, wb_stb, n22542, \iw_word[31] , \iw_word[1] , 
            \iw_word[30] , \iw_word[28] , \iw_word[29] , \iw_word[26] , 
            \iw_word[27] , \iw_word[24] , \iw_word[25] , \iw_word[22] , 
            \iw_word[23] , \iw_word[20] , \iw_word[21] , \iw_word[18] , 
            \iw_word[19] , \iw_word[16] , \iw_word[17] , wb_err, n30027, 
            wb_ack, \iw_word[14] , \iw_word[15] , \wb_idata[0] , wb_addr, 
            \wb_idata[2] , \wb_idata[3] , \wb_idata[4] , \wb_idata[5] , 
            \wb_idata[6] , \wb_idata[7] , \wb_idata[8] , \wb_idata[9] , 
            \wb_idata[10] , \wb_idata[11] , \wb_idata[12] , \wb_idata[13] , 
            \wb_idata[14] , \wb_idata[15] , \wb_idata[16] , \wb_idata[17] , 
            \wb_idata[18] , \wb_idata[19] , \iw_word[12] , \iw_word[13] , 
            \wb_idata[20] , \wb_idata[21] , \wb_idata[22] , \wb_idata[23] , 
            \wb_idata[24] , \wb_idata[25] , \wb_idata[26] , \iw_word[10] , 
            \iw_word[11] , \wb_idata[27] , \wb_idata[28] , \wb_idata[29] , 
            \wb_idata[30] , \wb_idata[31] , \iw_word[8] , \iw_word[9] , 
            \iw_word[6] , \iw_word[7] , \iw_word[5] , \iw_word[4] , 
            \iw_word[3] , \iw_word[2] , n2, n17754, GND_net, n27423, 
            \iw_word[32] , n27443, dac_clk_p_c_enable_471, n12753) /* synthesis syn_module_defined=1 */ ;
    input dac_clk_p_c;
    output wb_cyc;
    input newaddr_N_989;
    output [31:0]wb_odata;
    input \iw_word[0] ;
    output inc;
    input dac_clk_p_c_enable_138;
    output ow_stb;
    output [33:0]ow_word;
    input n30028;
    output wb_we;
    input i_cmd_wr;
    output wb_stb;
    input n22542;
    input \iw_word[31] ;
    input \iw_word[1] ;
    input \iw_word[30] ;
    input \iw_word[28] ;
    input \iw_word[29] ;
    input \iw_word[26] ;
    input \iw_word[27] ;
    input \iw_word[24] ;
    input \iw_word[25] ;
    input \iw_word[22] ;
    input \iw_word[23] ;
    input \iw_word[20] ;
    input \iw_word[21] ;
    input \iw_word[18] ;
    input \iw_word[19] ;
    input \iw_word[16] ;
    input \iw_word[17] ;
    input wb_err;
    input n30027;
    input wb_ack;
    input \iw_word[14] ;
    input \iw_word[15] ;
    input \wb_idata[0] ;
    output [29:0]wb_addr;
    input \wb_idata[2] ;
    input \wb_idata[3] ;
    input \wb_idata[4] ;
    input \wb_idata[5] ;
    input \wb_idata[6] ;
    input \wb_idata[7] ;
    input \wb_idata[8] ;
    input \wb_idata[9] ;
    input \wb_idata[10] ;
    input \wb_idata[11] ;
    input \wb_idata[12] ;
    input \wb_idata[13] ;
    input \wb_idata[14] ;
    input \wb_idata[15] ;
    input \wb_idata[16] ;
    input \wb_idata[17] ;
    input \wb_idata[18] ;
    input \wb_idata[19] ;
    input \iw_word[12] ;
    input \iw_word[13] ;
    input \wb_idata[20] ;
    input \wb_idata[21] ;
    input \wb_idata[22] ;
    input \wb_idata[23] ;
    input \wb_idata[24] ;
    input \wb_idata[25] ;
    input \wb_idata[26] ;
    input \iw_word[10] ;
    input \iw_word[11] ;
    input \wb_idata[27] ;
    input \wb_idata[28] ;
    input \wb_idata[29] ;
    input \wb_idata[30] ;
    input \wb_idata[31] ;
    input \iw_word[8] ;
    input \iw_word[9] ;
    input \iw_word[6] ;
    input \iw_word[7] ;
    input \iw_word[5] ;
    input \iw_word[4] ;
    input \iw_word[3] ;
    input \iw_word[2] ;
    output n2;
    input n17754;
    input GND_net;
    input n27423;
    input \iw_word[32] ;
    input n27443;
    input dac_clk_p_c_enable_471;
    input n12753;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[49:58])
    
    wire newaddr, i_cmd_word_0__N_994, n9811, o_rsp_stb_N_986;
    wire [33:0]n338;
    wire [33:0]o_rsp_word_33__N_950;
    
    wire o_cmd_busy_N_930, n20129, n18012, n17699, n17697;
    wire [29:0]n125;
    
    wire n18011, n17703, n17701, n18010, n17707, n17705, n18009, 
        n17711, n17709, n18008, n17715, n17713, n18007, n17719, 
        n17717, n18006, n17723, n17721, n18005, n17727, n17725, 
        n18004, n17731, n17729, n18003, n17735, n17733, n18002, 
        n17739, n17737;
    wire [32:0]n2210;
    
    wire n18001, n17743, n17741, n18000, n17747, n17745, n17999, 
        n17751, n17749, n17998, n17753, n3, n20752, o_cmd_busy_N_940, 
        o_cmd_busy_N_932, dac_clk_p_c_enable_438;
    
    FD1S3IX newaddr_72 (.D(newaddr_N_989), .CK(dac_clk_p_c), .CD(wb_cyc), 
            .Q(newaddr)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(192[9] 236[5])
    defparam newaddr_72.GSR = "DISABLED";
    FD1S3AX o_wb_data_i0 (.D(\iw_word[0] ), .CK(dac_clk_p_c), .Q(wb_odata[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i0.GSR = "DISABLED";
    FD1P3AX inc_71 (.D(i_cmd_word_0__N_994), .SP(dac_clk_p_c_enable_138), 
            .CK(dac_clk_p_c), .Q(inc)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(192[9] 236[5])
    defparam inc_71.GSR = "DISABLED";
    FD1S3JX o_rsp_stb_74 (.D(o_rsp_stb_N_986), .CK(dac_clk_p_c), .PD(n9811), 
            .Q(ow_stb)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_stb_74.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i0 (.D(n338[0]), .CK(dac_clk_p_c), .CD(n9811), 
            .Q(ow_word[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i0.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i2 (.D(n338[2]), .CK(dac_clk_p_c), .CD(n9811), 
            .Q(ow_word[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i2.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i3 (.D(n338[3]), .CK(dac_clk_p_c), .CD(n9811), 
            .Q(ow_word[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i3.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i4 (.D(n338[4]), .CK(dac_clk_p_c), .CD(n9811), 
            .Q(ow_word[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i4.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i5 (.D(n338[5]), .CK(dac_clk_p_c), .CD(n9811), 
            .Q(ow_word[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i5.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i6 (.D(n338[6]), .CK(dac_clk_p_c), .CD(n9811), 
            .Q(ow_word[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i6.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i7 (.D(n338[7]), .CK(dac_clk_p_c), .CD(n9811), 
            .Q(ow_word[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i7.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i8 (.D(n338[8]), .CK(dac_clk_p_c), .CD(n9811), 
            .Q(ow_word[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i8.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i9 (.D(n338[9]), .CK(dac_clk_p_c), .CD(n9811), 
            .Q(ow_word[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i9.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i10 (.D(n338[10]), .CK(dac_clk_p_c), .CD(n9811), 
            .Q(ow_word[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i10.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i11 (.D(n338[11]), .CK(dac_clk_p_c), .CD(n9811), 
            .Q(ow_word[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i11.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i12 (.D(n338[12]), .CK(dac_clk_p_c), .CD(n9811), 
            .Q(ow_word[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i12.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i13 (.D(n338[13]), .CK(dac_clk_p_c), .CD(n9811), 
            .Q(ow_word[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i13.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i14 (.D(n338[14]), .CK(dac_clk_p_c), .CD(n9811), 
            .Q(ow_word[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i14.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i15 (.D(n338[15]), .CK(dac_clk_p_c), .CD(n9811), 
            .Q(ow_word[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i15.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i16 (.D(n338[16]), .CK(dac_clk_p_c), .CD(n9811), 
            .Q(ow_word[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i16.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i17 (.D(n338[17]), .CK(dac_clk_p_c), .CD(n9811), 
            .Q(ow_word[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i17.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i18 (.D(n338[18]), .CK(dac_clk_p_c), .CD(n9811), 
            .Q(ow_word[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i18.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i19 (.D(n338[19]), .CK(dac_clk_p_c), .CD(n9811), 
            .Q(ow_word[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i19.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i20 (.D(n338[20]), .CK(dac_clk_p_c), .CD(n9811), 
            .Q(ow_word[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i20.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i21 (.D(n338[21]), .CK(dac_clk_p_c), .CD(n9811), 
            .Q(ow_word[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i21.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i22 (.D(n338[22]), .CK(dac_clk_p_c), .CD(n9811), 
            .Q(ow_word[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i22.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i23 (.D(n338[23]), .CK(dac_clk_p_c), .CD(n9811), 
            .Q(ow_word[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i23.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i24 (.D(n338[24]), .CK(dac_clk_p_c), .CD(n9811), 
            .Q(ow_word[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i24.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i25 (.D(n338[25]), .CK(dac_clk_p_c), .CD(n9811), 
            .Q(ow_word[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i25.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i26 (.D(n338[26]), .CK(dac_clk_p_c), .CD(n9811), 
            .Q(ow_word[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i26.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i27 (.D(n338[27]), .CK(dac_clk_p_c), .CD(n9811), 
            .Q(ow_word[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i27.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i28 (.D(n338[28]), .CK(dac_clk_p_c), .CD(n9811), 
            .Q(ow_word[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i28.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i29 (.D(o_rsp_word_33__N_950[29]), .CK(dac_clk_p_c), 
            .CD(n30028), .Q(ow_word[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i29.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i30 (.D(n338[30]), .CK(dac_clk_p_c), .CD(n9811), 
            .Q(ow_word[30])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i30.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i31 (.D(n338[31]), .CK(dac_clk_p_c), .CD(n9811), 
            .Q(ow_word[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i31.GSR = "DISABLED";
    FD1S3JX o_rsp_word_i32 (.D(n338[32]), .CK(dac_clk_p_c), .PD(n9811), 
            .Q(ow_word[32])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i32.GSR = "DISABLED";
    FD1S3JX o_rsp_word_i33 (.D(o_cmd_busy_N_930), .CK(dac_clk_p_c), .PD(n9811), 
            .Q(ow_word[33])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i33.GSR = "DISABLED";
    FD1P3AX o_wb_we_69 (.D(i_cmd_wr), .SP(o_cmd_busy_N_930), .CK(dac_clk_p_c), 
            .Q(wb_we)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(184[9] 186[26])
    defparam o_wb_we_69.GSR = "DISABLED";
    FD1P3IX o_wb_stb_68 (.D(n22542), .SP(o_cmd_busy_N_930), .CD(n20129), 
            .CK(dac_clk_p_c), .Q(wb_stb)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(121[9] 168[5])
    defparam o_wb_stb_68.GSR = "DISABLED";
    FD1S3AX o_wb_data_i31 (.D(\iw_word[31] ), .CK(dac_clk_p_c), .Q(wb_odata[31])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i31.GSR = "DISABLED";
    CCU2D o_wb_addr_598_add_4_31 (.A0(n17699), .B0(\iw_word[1] ), .C0(dac_clk_p_c_enable_138), 
          .D0(\iw_word[30] ), .A1(n17697), .B1(\iw_word[1] ), .C1(dac_clk_p_c_enable_138), 
          .D1(\iw_word[31] ), .CIN(n18012), .S0(n125[28]), .S1(n125[29]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_598_add_4_31.INIT0 = 16'h5aaa;
    defparam o_wb_addr_598_add_4_31.INIT1 = 16'h5aaa;
    defparam o_wb_addr_598_add_4_31.INJECT1_0 = "NO";
    defparam o_wb_addr_598_add_4_31.INJECT1_1 = "NO";
    CCU2D o_wb_addr_598_add_4_29 (.A0(n17703), .B0(\iw_word[1] ), .C0(dac_clk_p_c_enable_138), 
          .D0(\iw_word[28] ), .A1(n17701), .B1(\iw_word[1] ), .C1(dac_clk_p_c_enable_138), 
          .D1(\iw_word[29] ), .CIN(n18011), .COUT(n18012), .S0(n125[26]), 
          .S1(n125[27]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_598_add_4_29.INIT0 = 16'h5aaa;
    defparam o_wb_addr_598_add_4_29.INIT1 = 16'h5aaa;
    defparam o_wb_addr_598_add_4_29.INJECT1_0 = "NO";
    defparam o_wb_addr_598_add_4_29.INJECT1_1 = "NO";
    CCU2D o_wb_addr_598_add_4_27 (.A0(n17707), .B0(\iw_word[1] ), .C0(dac_clk_p_c_enable_138), 
          .D0(\iw_word[26] ), .A1(n17705), .B1(\iw_word[1] ), .C1(dac_clk_p_c_enable_138), 
          .D1(\iw_word[27] ), .CIN(n18010), .COUT(n18011), .S0(n125[24]), 
          .S1(n125[25]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_598_add_4_27.INIT0 = 16'h5aaa;
    defparam o_wb_addr_598_add_4_27.INIT1 = 16'h5aaa;
    defparam o_wb_addr_598_add_4_27.INJECT1_0 = "NO";
    defparam o_wb_addr_598_add_4_27.INJECT1_1 = "NO";
    CCU2D o_wb_addr_598_add_4_25 (.A0(n17711), .B0(\iw_word[1] ), .C0(dac_clk_p_c_enable_138), 
          .D0(\iw_word[24] ), .A1(n17709), .B1(\iw_word[1] ), .C1(dac_clk_p_c_enable_138), 
          .D1(\iw_word[25] ), .CIN(n18009), .COUT(n18010), .S0(n125[22]), 
          .S1(n125[23]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_598_add_4_25.INIT0 = 16'h5aaa;
    defparam o_wb_addr_598_add_4_25.INIT1 = 16'h5aaa;
    defparam o_wb_addr_598_add_4_25.INJECT1_0 = "NO";
    defparam o_wb_addr_598_add_4_25.INJECT1_1 = "NO";
    CCU2D o_wb_addr_598_add_4_23 (.A0(n17715), .B0(\iw_word[1] ), .C0(dac_clk_p_c_enable_138), 
          .D0(\iw_word[22] ), .A1(n17713), .B1(\iw_word[1] ), .C1(dac_clk_p_c_enable_138), 
          .D1(\iw_word[23] ), .CIN(n18008), .COUT(n18009), .S0(n125[20]), 
          .S1(n125[21]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_598_add_4_23.INIT0 = 16'h5aaa;
    defparam o_wb_addr_598_add_4_23.INIT1 = 16'h5aaa;
    defparam o_wb_addr_598_add_4_23.INJECT1_0 = "NO";
    defparam o_wb_addr_598_add_4_23.INJECT1_1 = "NO";
    CCU2D o_wb_addr_598_add_4_21 (.A0(n17719), .B0(\iw_word[1] ), .C0(dac_clk_p_c_enable_138), 
          .D0(\iw_word[20] ), .A1(n17717), .B1(\iw_word[1] ), .C1(dac_clk_p_c_enable_138), 
          .D1(\iw_word[21] ), .CIN(n18007), .COUT(n18008), .S0(n125[18]), 
          .S1(n125[19]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_598_add_4_21.INIT0 = 16'h5aaa;
    defparam o_wb_addr_598_add_4_21.INIT1 = 16'h5aaa;
    defparam o_wb_addr_598_add_4_21.INJECT1_0 = "NO";
    defparam o_wb_addr_598_add_4_21.INJECT1_1 = "NO";
    CCU2D o_wb_addr_598_add_4_19 (.A0(n17723), .B0(\iw_word[1] ), .C0(dac_clk_p_c_enable_138), 
          .D0(\iw_word[18] ), .A1(n17721), .B1(\iw_word[1] ), .C1(dac_clk_p_c_enable_138), 
          .D1(\iw_word[19] ), .CIN(n18006), .COUT(n18007), .S0(n125[16]), 
          .S1(n125[17]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_598_add_4_19.INIT0 = 16'h5aaa;
    defparam o_wb_addr_598_add_4_19.INIT1 = 16'h5aaa;
    defparam o_wb_addr_598_add_4_19.INJECT1_0 = "NO";
    defparam o_wb_addr_598_add_4_19.INJECT1_1 = "NO";
    CCU2D o_wb_addr_598_add_4_17 (.A0(n17727), .B0(\iw_word[1] ), .C0(dac_clk_p_c_enable_138), 
          .D0(\iw_word[16] ), .A1(n17725), .B1(\iw_word[1] ), .C1(dac_clk_p_c_enable_138), 
          .D1(\iw_word[17] ), .CIN(n18005), .COUT(n18006), .S0(n125[14]), 
          .S1(n125[15]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_598_add_4_17.INIT0 = 16'h5aaa;
    defparam o_wb_addr_598_add_4_17.INIT1 = 16'h5aaa;
    defparam o_wb_addr_598_add_4_17.INJECT1_0 = "NO";
    defparam o_wb_addr_598_add_4_17.INJECT1_1 = "NO";
    LUT4 i_cmd_word_0__I_0_1_lut (.A(\iw_word[0] ), .Z(i_cmd_word_0__N_994)) /* synthesis lut_function=(!(A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(214[11:25])
    defparam i_cmd_word_0__I_0_1_lut.init = 16'h5555;
    LUT4 i7390_2_lut (.A(wb_err), .B(n30027), .Z(n9811)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(283[11] 309[5])
    defparam i7390_2_lut.init = 16'heeee;
    LUT4 newaddr_I_0_3_lut (.A(newaddr), .B(wb_ack), .C(wb_cyc), .Z(o_rsp_stb_N_986)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam newaddr_I_0_3_lut.init = 16'hcaca;
    CCU2D o_wb_addr_598_add_4_15 (.A0(n17731), .B0(\iw_word[1] ), .C0(dac_clk_p_c_enable_138), 
          .D0(\iw_word[14] ), .A1(n17729), .B1(\iw_word[1] ), .C1(dac_clk_p_c_enable_138), 
          .D1(\iw_word[15] ), .CIN(n18004), .COUT(n18005), .S0(n125[12]), 
          .S1(n125[13]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_598_add_4_15.INIT0 = 16'h5aaa;
    defparam o_wb_addr_598_add_4_15.INIT1 = 16'h5aaa;
    defparam o_wb_addr_598_add_4_15.INJECT1_0 = "NO";
    defparam o_wb_addr_598_add_4_15.INJECT1_1 = "NO";
    LUT4 mux_59_i1_4_lut (.A(inc), .B(\wb_idata[0] ), .C(wb_cyc), .D(wb_we), 
         .Z(n338[0])) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A (B (C (D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i1_4_lut.init = 16'h05c5;
    LUT4 mux_59_i3_4_lut (.A(wb_addr[0]), .B(\wb_idata[2] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[2])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i3_4_lut.init = 16'h0aca;
    LUT4 mux_59_i4_4_lut (.A(wb_addr[1]), .B(\wb_idata[3] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[3])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i4_4_lut.init = 16'h0aca;
    LUT4 mux_59_i5_4_lut (.A(wb_addr[2]), .B(\wb_idata[4] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[4])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i5_4_lut.init = 16'h0aca;
    LUT4 mux_59_i6_4_lut (.A(wb_addr[3]), .B(\wb_idata[5] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[5])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i6_4_lut.init = 16'h0aca;
    LUT4 mux_59_i7_4_lut (.A(wb_addr[4]), .B(\wb_idata[6] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[6])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i7_4_lut.init = 16'h0aca;
    LUT4 mux_59_i8_4_lut (.A(wb_addr[5]), .B(\wb_idata[7] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[7])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i8_4_lut.init = 16'h0aca;
    LUT4 mux_59_i9_4_lut (.A(wb_addr[6]), .B(\wb_idata[8] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[8])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i9_4_lut.init = 16'h0aca;
    LUT4 mux_59_i10_4_lut (.A(wb_addr[7]), .B(\wb_idata[9] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[9])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i10_4_lut.init = 16'h0aca;
    LUT4 mux_59_i11_4_lut (.A(wb_addr[8]), .B(\wb_idata[10] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[10])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i11_4_lut.init = 16'h0aca;
    LUT4 mux_59_i12_4_lut (.A(wb_addr[9]), .B(\wb_idata[11] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[11])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i12_4_lut.init = 16'h0aca;
    LUT4 mux_59_i13_4_lut (.A(wb_addr[10]), .B(\wb_idata[12] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[12])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i13_4_lut.init = 16'h0aca;
    LUT4 mux_59_i14_4_lut (.A(wb_addr[11]), .B(\wb_idata[13] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[13])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i14_4_lut.init = 16'h0aca;
    LUT4 mux_59_i15_4_lut (.A(wb_addr[12]), .B(\wb_idata[14] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[14])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i15_4_lut.init = 16'h0aca;
    LUT4 mux_59_i16_4_lut (.A(wb_addr[13]), .B(\wb_idata[15] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[15])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i16_4_lut.init = 16'h0aca;
    LUT4 mux_59_i17_4_lut (.A(wb_addr[14]), .B(\wb_idata[16] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[16])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i17_4_lut.init = 16'h0aca;
    LUT4 mux_59_i18_4_lut (.A(wb_addr[15]), .B(\wb_idata[17] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[17])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i18_4_lut.init = 16'h0aca;
    LUT4 mux_59_i19_4_lut (.A(wb_addr[16]), .B(\wb_idata[18] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[18])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i19_4_lut.init = 16'h0aca;
    LUT4 mux_59_i20_4_lut (.A(wb_addr[17]), .B(\wb_idata[19] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[19])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i20_4_lut.init = 16'h0aca;
    CCU2D o_wb_addr_598_add_4_13 (.A0(n17735), .B0(\iw_word[1] ), .C0(dac_clk_p_c_enable_138), 
          .D0(\iw_word[12] ), .A1(n17733), .B1(\iw_word[1] ), .C1(dac_clk_p_c_enable_138), 
          .D1(\iw_word[13] ), .CIN(n18003), .COUT(n18004), .S0(n125[10]), 
          .S1(n125[11]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_598_add_4_13.INIT0 = 16'h5aaa;
    defparam o_wb_addr_598_add_4_13.INIT1 = 16'h5aaa;
    defparam o_wb_addr_598_add_4_13.INJECT1_0 = "NO";
    defparam o_wb_addr_598_add_4_13.INJECT1_1 = "NO";
    LUT4 mux_59_i21_4_lut (.A(wb_addr[18]), .B(\wb_idata[20] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[20])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i21_4_lut.init = 16'h0aca;
    LUT4 mux_59_i22_4_lut (.A(wb_addr[19]), .B(\wb_idata[21] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[21])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i22_4_lut.init = 16'h0aca;
    LUT4 mux_59_i23_4_lut (.A(wb_addr[20]), .B(\wb_idata[22] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[22])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i23_4_lut.init = 16'h0aca;
    LUT4 mux_59_i24_4_lut (.A(wb_addr[21]), .B(\wb_idata[23] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[23])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i24_4_lut.init = 16'h0aca;
    LUT4 mux_59_i25_4_lut (.A(wb_addr[22]), .B(\wb_idata[24] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[24])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i25_4_lut.init = 16'h0aca;
    LUT4 mux_59_i26_4_lut (.A(wb_addr[23]), .B(\wb_idata[25] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[25])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i26_4_lut.init = 16'h0aca;
    LUT4 mux_59_i27_4_lut (.A(wb_addr[24]), .B(\wb_idata[26] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[26])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i27_4_lut.init = 16'h0aca;
    CCU2D o_wb_addr_598_add_4_11 (.A0(n17739), .B0(\iw_word[1] ), .C0(dac_clk_p_c_enable_138), 
          .D0(\iw_word[10] ), .A1(n17737), .B1(\iw_word[1] ), .C1(dac_clk_p_c_enable_138), 
          .D1(\iw_word[11] ), .CIN(n18002), .COUT(n18003), .S0(n125[8]), 
          .S1(n125[9]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_598_add_4_11.INIT0 = 16'h5aaa;
    defparam o_wb_addr_598_add_4_11.INIT1 = 16'h5aaa;
    defparam o_wb_addr_598_add_4_11.INJECT1_0 = "NO";
    defparam o_wb_addr_598_add_4_11.INJECT1_1 = "NO";
    LUT4 mux_59_i28_4_lut (.A(wb_addr[25]), .B(\wb_idata[27] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[27])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i28_4_lut.init = 16'h0aca;
    LUT4 mux_59_i29_4_lut (.A(wb_addr[26]), .B(\wb_idata[28] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[28])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i29_4_lut.init = 16'h0aca;
    LUT4 i11681_4_lut (.A(wb_addr[27]), .B(wb_err), .C(n2210[29]), .D(wb_cyc), 
         .Z(o_rsp_word_33__N_950[29])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(287[11] 309[5])
    defparam i11681_4_lut.init = 16'hfcee;
    LUT4 i11730_2_lut (.A(\wb_idata[29] ), .B(wb_we), .Z(n2210[29])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(299[4:47])
    defparam i11730_2_lut.init = 16'h2222;
    LUT4 mux_59_i31_4_lut (.A(wb_addr[28]), .B(\wb_idata[30] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[30])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i31_4_lut.init = 16'h0aca;
    LUT4 mux_59_i32_4_lut (.A(wb_addr[29]), .B(\wb_idata[31] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[31])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i32_4_lut.init = 16'h0aca;
    LUT4 i11683_2_lut (.A(wb_we), .B(wb_cyc), .Z(n338[32])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam i11683_2_lut.init = 16'h8888;
    LUT4 o_cmd_busy_I_0_1_lut (.A(wb_cyc), .Z(o_cmd_busy_N_930)) /* synthesis lut_function=(!(A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(194[21:34])
    defparam o_cmd_busy_I_0_1_lut.init = 16'h5555;
    CCU2D o_wb_addr_598_add_4_9 (.A0(n17743), .B0(\iw_word[1] ), .C0(dac_clk_p_c_enable_138), 
          .D0(\iw_word[8] ), .A1(n17741), .B1(\iw_word[1] ), .C1(dac_clk_p_c_enable_138), 
          .D1(\iw_word[9] ), .CIN(n18001), .COUT(n18002), .S0(n125[6]), 
          .S1(n125[7]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_598_add_4_9.INIT0 = 16'h5aaa;
    defparam o_wb_addr_598_add_4_9.INIT1 = 16'h5aaa;
    defparam o_wb_addr_598_add_4_9.INJECT1_0 = "NO";
    defparam o_wb_addr_598_add_4_9.INJECT1_1 = "NO";
    CCU2D o_wb_addr_598_add_4_7 (.A0(n17747), .B0(\iw_word[1] ), .C0(dac_clk_p_c_enable_138), 
          .D0(\iw_word[6] ), .A1(n17745), .B1(\iw_word[1] ), .C1(dac_clk_p_c_enable_138), 
          .D1(\iw_word[7] ), .CIN(n18000), .COUT(n18001), .S0(n125[4]), 
          .S1(n125[5]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_598_add_4_7.INIT0 = 16'h5aaa;
    defparam o_wb_addr_598_add_4_7.INIT1 = 16'h5aaa;
    defparam o_wb_addr_598_add_4_7.INJECT1_0 = "NO";
    defparam o_wb_addr_598_add_4_7.INJECT1_1 = "NO";
    FD1S3AX o_wb_data_i30 (.D(\iw_word[30] ), .CK(dac_clk_p_c), .Q(wb_odata[30])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i30.GSR = "DISABLED";
    FD1S3AX o_wb_data_i29 (.D(\iw_word[29] ), .CK(dac_clk_p_c), .Q(wb_odata[29])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i29.GSR = "DISABLED";
    FD1S3AX o_wb_data_i28 (.D(\iw_word[28] ), .CK(dac_clk_p_c), .Q(wb_odata[28])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i28.GSR = "DISABLED";
    FD1S3AX o_wb_data_i27 (.D(\iw_word[27] ), .CK(dac_clk_p_c), .Q(wb_odata[27])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i27.GSR = "DISABLED";
    FD1S3AX o_wb_data_i26 (.D(\iw_word[26] ), .CK(dac_clk_p_c), .Q(wb_odata[26])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i26.GSR = "DISABLED";
    FD1S3AX o_wb_data_i25 (.D(\iw_word[25] ), .CK(dac_clk_p_c), .Q(wb_odata[25])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i25.GSR = "DISABLED";
    FD1S3AX o_wb_data_i24 (.D(\iw_word[24] ), .CK(dac_clk_p_c), .Q(wb_odata[24])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i24.GSR = "DISABLED";
    FD1S3AX o_wb_data_i23 (.D(\iw_word[23] ), .CK(dac_clk_p_c), .Q(wb_odata[23])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i23.GSR = "DISABLED";
    FD1S3AX o_wb_data_i22 (.D(\iw_word[22] ), .CK(dac_clk_p_c), .Q(wb_odata[22])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i22.GSR = "DISABLED";
    FD1S3AX o_wb_data_i21 (.D(\iw_word[21] ), .CK(dac_clk_p_c), .Q(wb_odata[21])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i21.GSR = "DISABLED";
    FD1S3AX o_wb_data_i20 (.D(\iw_word[20] ), .CK(dac_clk_p_c), .Q(wb_odata[20])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i20.GSR = "DISABLED";
    FD1S3AX o_wb_data_i19 (.D(\iw_word[19] ), .CK(dac_clk_p_c), .Q(wb_odata[19])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i19.GSR = "DISABLED";
    FD1S3AX o_wb_data_i18 (.D(\iw_word[18] ), .CK(dac_clk_p_c), .Q(wb_odata[18])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i18.GSR = "DISABLED";
    FD1S3AX o_wb_data_i17 (.D(\iw_word[17] ), .CK(dac_clk_p_c), .Q(wb_odata[17])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i17.GSR = "DISABLED";
    FD1S3AX o_wb_data_i16 (.D(\iw_word[16] ), .CK(dac_clk_p_c), .Q(wb_odata[16])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i16.GSR = "DISABLED";
    FD1S3AX o_wb_data_i15 (.D(\iw_word[15] ), .CK(dac_clk_p_c), .Q(wb_odata[15])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i15.GSR = "DISABLED";
    FD1S3AX o_wb_data_i14 (.D(\iw_word[14] ), .CK(dac_clk_p_c), .Q(wb_odata[14])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i14.GSR = "DISABLED";
    FD1S3AX o_wb_data_i13 (.D(\iw_word[13] ), .CK(dac_clk_p_c), .Q(wb_odata[13])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i13.GSR = "DISABLED";
    FD1S3AX o_wb_data_i12 (.D(\iw_word[12] ), .CK(dac_clk_p_c), .Q(wb_odata[12])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i12.GSR = "DISABLED";
    FD1S3AX o_wb_data_i11 (.D(\iw_word[11] ), .CK(dac_clk_p_c), .Q(wb_odata[11])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i11.GSR = "DISABLED";
    FD1S3AX o_wb_data_i10 (.D(\iw_word[10] ), .CK(dac_clk_p_c), .Q(wb_odata[10])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i10.GSR = "DISABLED";
    FD1S3AX o_wb_data_i9 (.D(\iw_word[9] ), .CK(dac_clk_p_c), .Q(wb_odata[9])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i9.GSR = "DISABLED";
    FD1S3AX o_wb_data_i8 (.D(\iw_word[8] ), .CK(dac_clk_p_c), .Q(wb_odata[8])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i8.GSR = "DISABLED";
    FD1S3AX o_wb_data_i7 (.D(\iw_word[7] ), .CK(dac_clk_p_c), .Q(wb_odata[7])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i7.GSR = "DISABLED";
    FD1S3AX o_wb_data_i6 (.D(\iw_word[6] ), .CK(dac_clk_p_c), .Q(wb_odata[6])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i6.GSR = "DISABLED";
    FD1S3AX o_wb_data_i5 (.D(\iw_word[5] ), .CK(dac_clk_p_c), .Q(wb_odata[5])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i5.GSR = "DISABLED";
    FD1S3AX o_wb_data_i4 (.D(\iw_word[4] ), .CK(dac_clk_p_c), .Q(wb_odata[4])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i4.GSR = "DISABLED";
    FD1S3AX o_wb_data_i3 (.D(\iw_word[3] ), .CK(dac_clk_p_c), .Q(wb_odata[3])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i3.GSR = "DISABLED";
    FD1S3AX o_wb_data_i2 (.D(\iw_word[2] ), .CK(dac_clk_p_c), .Q(wb_odata[2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i2.GSR = "DISABLED";
    FD1S3AX o_wb_data_i1 (.D(\iw_word[1] ), .CK(dac_clk_p_c), .Q(wb_odata[1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i1.GSR = "DISABLED";
    LUT4 i2_1_lut (.A(wb_stb), .Z(n2)) /* synthesis lut_function=(!(A)) */ ;
    defparam i2_1_lut.init = 16'h5555;
    CCU2D o_wb_addr_598_add_4_5 (.A0(n17751), .B0(\iw_word[1] ), .C0(dac_clk_p_c_enable_138), 
          .D0(\iw_word[4] ), .A1(n17749), .B1(\iw_word[1] ), .C1(dac_clk_p_c_enable_138), 
          .D1(\iw_word[5] ), .CIN(n17999), .COUT(n18000), .S0(n125[2]), 
          .S1(n125[3]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_598_add_4_5.INIT0 = 16'h5aaa;
    defparam o_wb_addr_598_add_4_5.INIT1 = 16'h5aaa;
    defparam o_wb_addr_598_add_4_5.INJECT1_0 = "NO";
    defparam o_wb_addr_598_add_4_5.INJECT1_1 = "NO";
    CCU2D o_wb_addr_598_add_4_3 (.A0(n17754), .B0(dac_clk_p_c_enable_138), 
          .C0(\iw_word[1] ), .D0(wb_addr[0]), .A1(n17753), .B1(\iw_word[1] ), 
          .C1(dac_clk_p_c_enable_138), .D1(\iw_word[3] ), .CIN(n17998), 
          .COUT(n17999), .S0(n125[0]), .S1(n125[1]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_598_add_4_3.INIT0 = 16'h59aa;
    defparam o_wb_addr_598_add_4_3.INIT1 = 16'h5aaa;
    defparam o_wb_addr_598_add_4_3.INJECT1_0 = "NO";
    defparam o_wb_addr_598_add_4_3.INJECT1_1 = "NO";
    CCU2D o_wb_addr_598_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\iw_word[1] ), .B1(dac_clk_p_c_enable_138), 
          .C1(GND_net), .D1(GND_net), .COUT(n17998));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_598_add_4_1.INIT0 = 16'hF000;
    defparam o_wb_addr_598_add_4_1.INIT1 = 16'hffff;
    defparam o_wb_addr_598_add_4_1.INJECT1_0 = "NO";
    defparam o_wb_addr_598_add_4_1.INJECT1_1 = "NO";
    LUT4 i15960_2_lut (.A(wb_addr[28]), .B(n3), .Z(n17699)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15960_2_lut.init = 16'h8888;
    LUT4 i15961_2_lut (.A(wb_addr[29]), .B(n3), .Z(n17697)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15961_2_lut.init = 16'h8888;
    LUT4 i1_4_lut (.A(\iw_word[1] ), .B(n27423), .C(wb_cyc), .D(\iw_word[32] ), 
         .Z(n3)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;
    defparam i1_4_lut.init = 16'hfffb;
    LUT4 i15958_2_lut (.A(wb_addr[26]), .B(n3), .Z(n17703)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15958_2_lut.init = 16'h8888;
    LUT4 i15959_2_lut (.A(wb_addr[27]), .B(n3), .Z(n17701)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15959_2_lut.init = 16'h8888;
    LUT4 i15956_2_lut (.A(wb_addr[24]), .B(n3), .Z(n17707)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15956_2_lut.init = 16'h8888;
    LUT4 i15957_2_lut (.A(wb_addr[25]), .B(n3), .Z(n17705)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15957_2_lut.init = 16'h8888;
    LUT4 i15937_2_lut (.A(wb_addr[22]), .B(n3), .Z(n17711)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15937_2_lut.init = 16'h8888;
    LUT4 i15947_2_lut (.A(wb_addr[23]), .B(n3), .Z(n17709)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15947_2_lut.init = 16'h8888;
    LUT4 i15909_2_lut (.A(wb_addr[20]), .B(n3), .Z(n17715)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15909_2_lut.init = 16'h8888;
    LUT4 i15963_2_lut (.A(wb_addr[21]), .B(n3), .Z(n17713)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15963_2_lut.init = 16'h8888;
    LUT4 i15912_2_lut (.A(wb_addr[18]), .B(n3), .Z(n17719)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15912_2_lut.init = 16'h8888;
    LUT4 i15941_2_lut (.A(wb_addr[19]), .B(n3), .Z(n17717)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15941_2_lut.init = 16'h8888;
    LUT4 i15929_2_lut (.A(wb_addr[16]), .B(n3), .Z(n17723)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15929_2_lut.init = 16'h8888;
    LUT4 i15962_2_lut (.A(wb_addr[17]), .B(n3), .Z(n17721)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15962_2_lut.init = 16'h8888;
    LUT4 i15911_2_lut (.A(wb_addr[14]), .B(n3), .Z(n17727)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15911_2_lut.init = 16'h8888;
    LUT4 i15923_2_lut (.A(wb_addr[15]), .B(n3), .Z(n17725)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15923_2_lut.init = 16'h8888;
    LUT4 i15949_2_lut (.A(wb_addr[12]), .B(n3), .Z(n17731)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15949_2_lut.init = 16'h8888;
    LUT4 i15966_2_lut (.A(wb_addr[13]), .B(n3), .Z(n17729)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15966_2_lut.init = 16'h8888;
    LUT4 i15942_2_lut (.A(wb_addr[10]), .B(n3), .Z(n17735)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15942_2_lut.init = 16'h8888;
    LUT4 i15943_2_lut (.A(wb_addr[11]), .B(n3), .Z(n17733)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15943_2_lut.init = 16'h8888;
    LUT4 i15928_2_lut (.A(wb_addr[8]), .B(n3), .Z(n17739)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15928_2_lut.init = 16'h8888;
    LUT4 i15930_2_lut (.A(wb_addr[9]), .B(n3), .Z(n17737)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15930_2_lut.init = 16'h8888;
    LUT4 i15922_2_lut (.A(wb_addr[6]), .B(n3), .Z(n17743)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15922_2_lut.init = 16'h8888;
    LUT4 i15924_2_lut (.A(wb_addr[7]), .B(n3), .Z(n17741)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15924_2_lut.init = 16'h8888;
    LUT4 i15914_2_lut (.A(wb_addr[4]), .B(n3), .Z(n17747)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15914_2_lut.init = 16'h8888;
    LUT4 i15915_2_lut (.A(wb_addr[5]), .B(n3), .Z(n17745)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15915_2_lut.init = 16'h8888;
    LUT4 i15910_2_lut (.A(wb_addr[2]), .B(n3), .Z(n17751)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15910_2_lut.init = 16'h8888;
    LUT4 i15913_2_lut (.A(wb_addr[3]), .B(n3), .Z(n17749)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15913_2_lut.init = 16'h8888;
    LUT4 i15908_2_lut (.A(wb_addr[1]), .B(n3), .Z(n17753)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15908_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_143 (.A(wb_err), .B(n30027), .C(wb_we), .D(wb_cyc), 
         .Z(n20752)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut_adj_143.init = 16'h0100;
    LUT4 i1_4_lut_adj_144 (.A(n27443), .B(o_cmd_busy_N_940), .C(wb_ack), 
         .D(o_cmd_busy_N_932), .Z(dac_clk_p_c_enable_438)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+!((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(122[6:41])
    defparam i1_4_lut_adj_144.init = 16'heefc;
    LUT4 i23168_2_lut (.A(wb_cyc), .B(wb_stb), .Z(o_cmd_busy_N_932)) /* synthesis lut_function=(!(A+(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(149[11] 168[5])
    defparam i23168_2_lut.init = 16'h1111;
    FD1P3AX o_wb_addr_598__i0 (.D(n125[0]), .SP(dac_clk_p_c_enable_471), 
            .CK(dac_clk_p_c), .Q(wb_addr[0])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_598__i0.GSR = "DISABLED";
    LUT4 i1_2_lut_3_lut_4_lut (.A(wb_err), .B(wb_cyc), .C(wb_stb), .D(n30027), 
         .Z(n20129)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(122[17:41])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfff8;
    LUT4 i1_2_lut_rep_566_3_lut (.A(wb_err), .B(wb_cyc), .C(n30027), .Z(o_cmd_busy_N_940)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(122[17:41])
    defparam i1_2_lut_rep_566_3_lut.init = 16'hf8f8;
    FD1S3IX o_rsp_word_i1 (.D(n20752), .CK(dac_clk_p_c), .CD(n12753), 
            .Q(ow_word[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i1.GSR = "DISABLED";
    FD1P3IX o_wb_cyc_67 (.D(o_cmd_busy_N_932), .SP(dac_clk_p_c_enable_438), 
            .CD(o_cmd_busy_N_940), .CK(dac_clk_p_c), .Q(wb_cyc)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(121[9] 168[5])
    defparam o_wb_cyc_67.GSR = "DISABLED";
    FD1P3AX o_wb_addr_598__i29 (.D(n125[29]), .SP(dac_clk_p_c_enable_471), 
            .CK(dac_clk_p_c), .Q(wb_addr[29])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_598__i29.GSR = "DISABLED";
    FD1P3AX o_wb_addr_598__i28 (.D(n125[28]), .SP(dac_clk_p_c_enable_471), 
            .CK(dac_clk_p_c), .Q(wb_addr[28])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_598__i28.GSR = "DISABLED";
    FD1P3AX o_wb_addr_598__i27 (.D(n125[27]), .SP(dac_clk_p_c_enable_471), 
            .CK(dac_clk_p_c), .Q(wb_addr[27])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_598__i27.GSR = "DISABLED";
    FD1P3AX o_wb_addr_598__i26 (.D(n125[26]), .SP(dac_clk_p_c_enable_471), 
            .CK(dac_clk_p_c), .Q(wb_addr[26])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_598__i26.GSR = "DISABLED";
    FD1P3AX o_wb_addr_598__i25 (.D(n125[25]), .SP(dac_clk_p_c_enable_471), 
            .CK(dac_clk_p_c), .Q(wb_addr[25])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_598__i25.GSR = "DISABLED";
    FD1P3AX o_wb_addr_598__i24 (.D(n125[24]), .SP(dac_clk_p_c_enable_471), 
            .CK(dac_clk_p_c), .Q(wb_addr[24])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_598__i24.GSR = "DISABLED";
    FD1P3AX o_wb_addr_598__i23 (.D(n125[23]), .SP(dac_clk_p_c_enable_471), 
            .CK(dac_clk_p_c), .Q(wb_addr[23])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_598__i23.GSR = "DISABLED";
    FD1P3AX o_wb_addr_598__i22 (.D(n125[22]), .SP(dac_clk_p_c_enable_471), 
            .CK(dac_clk_p_c), .Q(wb_addr[22])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_598__i22.GSR = "DISABLED";
    FD1P3AX o_wb_addr_598__i21 (.D(n125[21]), .SP(dac_clk_p_c_enable_471), 
            .CK(dac_clk_p_c), .Q(wb_addr[21])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_598__i21.GSR = "DISABLED";
    FD1P3AX o_wb_addr_598__i20 (.D(n125[20]), .SP(dac_clk_p_c_enable_471), 
            .CK(dac_clk_p_c), .Q(wb_addr[20])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_598__i20.GSR = "DISABLED";
    FD1P3AX o_wb_addr_598__i19 (.D(n125[19]), .SP(dac_clk_p_c_enable_471), 
            .CK(dac_clk_p_c), .Q(wb_addr[19])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_598__i19.GSR = "DISABLED";
    FD1P3AX o_wb_addr_598__i18 (.D(n125[18]), .SP(dac_clk_p_c_enable_471), 
            .CK(dac_clk_p_c), .Q(wb_addr[18])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_598__i18.GSR = "DISABLED";
    FD1P3AX o_wb_addr_598__i17 (.D(n125[17]), .SP(dac_clk_p_c_enable_471), 
            .CK(dac_clk_p_c), .Q(wb_addr[17])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_598__i17.GSR = "DISABLED";
    FD1P3AX o_wb_addr_598__i16 (.D(n125[16]), .SP(dac_clk_p_c_enable_471), 
            .CK(dac_clk_p_c), .Q(wb_addr[16])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_598__i16.GSR = "DISABLED";
    FD1P3AX o_wb_addr_598__i15 (.D(n125[15]), .SP(dac_clk_p_c_enable_471), 
            .CK(dac_clk_p_c), .Q(wb_addr[15])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_598__i15.GSR = "DISABLED";
    FD1P3AX o_wb_addr_598__i14 (.D(n125[14]), .SP(dac_clk_p_c_enable_471), 
            .CK(dac_clk_p_c), .Q(wb_addr[14])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_598__i14.GSR = "DISABLED";
    FD1P3AX o_wb_addr_598__i13 (.D(n125[13]), .SP(dac_clk_p_c_enable_471), 
            .CK(dac_clk_p_c), .Q(wb_addr[13])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_598__i13.GSR = "DISABLED";
    FD1P3AX o_wb_addr_598__i12 (.D(n125[12]), .SP(dac_clk_p_c_enable_471), 
            .CK(dac_clk_p_c), .Q(wb_addr[12])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_598__i12.GSR = "DISABLED";
    FD1P3AX o_wb_addr_598__i11 (.D(n125[11]), .SP(dac_clk_p_c_enable_471), 
            .CK(dac_clk_p_c), .Q(wb_addr[11])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_598__i11.GSR = "DISABLED";
    FD1P3AX o_wb_addr_598__i10 (.D(n125[10]), .SP(dac_clk_p_c_enable_471), 
            .CK(dac_clk_p_c), .Q(wb_addr[10])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_598__i10.GSR = "DISABLED";
    FD1P3AX o_wb_addr_598__i9 (.D(n125[9]), .SP(dac_clk_p_c_enable_471), 
            .CK(dac_clk_p_c), .Q(wb_addr[9])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_598__i9.GSR = "DISABLED";
    FD1P3AX o_wb_addr_598__i8 (.D(n125[8]), .SP(dac_clk_p_c_enable_471), 
            .CK(dac_clk_p_c), .Q(wb_addr[8])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_598__i8.GSR = "DISABLED";
    FD1P3AX o_wb_addr_598__i7 (.D(n125[7]), .SP(dac_clk_p_c_enable_471), 
            .CK(dac_clk_p_c), .Q(wb_addr[7])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_598__i7.GSR = "DISABLED";
    FD1P3AX o_wb_addr_598__i6 (.D(n125[6]), .SP(dac_clk_p_c_enable_471), 
            .CK(dac_clk_p_c), .Q(wb_addr[6])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_598__i6.GSR = "DISABLED";
    FD1P3AX o_wb_addr_598__i5 (.D(n125[5]), .SP(dac_clk_p_c_enable_471), 
            .CK(dac_clk_p_c), .Q(wb_addr[5])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_598__i5.GSR = "DISABLED";
    FD1P3AX o_wb_addr_598__i4 (.D(n125[4]), .SP(dac_clk_p_c_enable_471), 
            .CK(dac_clk_p_c), .Q(wb_addr[4])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_598__i4.GSR = "DISABLED";
    FD1P3AX o_wb_addr_598__i3 (.D(n125[3]), .SP(dac_clk_p_c_enable_471), 
            .CK(dac_clk_p_c), .Q(wb_addr[3])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_598__i3.GSR = "DISABLED";
    FD1P3AX o_wb_addr_598__i2 (.D(n125[2]), .SP(dac_clk_p_c_enable_471), 
            .CK(dac_clk_p_c), .Q(wb_addr[2])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_598__i2.GSR = "DISABLED";
    FD1P3AX o_wb_addr_598__i1 (.D(n125[1]), .SP(dac_clk_p_c_enable_471), 
            .CK(dac_clk_p_c), .Q(wb_addr[1])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_598__i1.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module hbdeword
//

module hbdeword (dac_clk_p_c, dac_clk_p_c_enable_332, hb_bits, dac_clk_p_c_enable_219, 
            n30028, idl_word, n29969, hb_busy, w_reset, idl_stb, 
            n27258, nl_busy, hx_stb, n30027) /* synthesis syn_module_defined=1 */ ;
    input dac_clk_p_c;
    input dac_clk_p_c_enable_332;
    output [4:0]hb_bits;
    input dac_clk_p_c_enable_219;
    input n30028;
    input [33:0]idl_word;
    input n29969;
    output hb_busy;
    input w_reset;
    input idl_stb;
    output n27258;
    input nl_busy;
    input hx_stb;
    input n30027;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[49:58])
    wire [3:0]r_len;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(58[12:17])
    
    wire n27141;
    wire [3:0]n13;
    
    wire dac_clk_p_c_enable_261;
    wire [4:0]o_dw_bits_4__N_1187;
    wire [31:0]r_word;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(59[13:19])
    wire [31:0]r_word_31__N_1196;
    wire [3:0]r_len_3__N_1228;
    
    wire n12840, o_dw_busy_N_1268, n11587, n27259;
    wire [4:0]o_dw_bits_4__N_1278;
    
    wire n26614, n20553, n11583, n26931;
    
    FD1P3IX r_len__i0 (.D(n13[0]), .SP(dac_clk_p_c_enable_332), .CD(n27141), 
            .CK(dac_clk_p_c), .Q(r_len[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(64[9] 81[6])
    defparam r_len__i0.GSR = "DISABLED";
    FD1P3AX o_dw_bits_i0 (.D(o_dw_bits_4__N_1187[0]), .SP(dac_clk_p_c_enable_261), 
            .CK(dac_clk_p_c), .Q(hb_bits[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(95[9] 103[41])
    defparam o_dw_bits_i0.GSR = "DISABLED";
    FD1P3AX o_dw_bits_i3 (.D(o_dw_bits_4__N_1187[3]), .SP(dac_clk_p_c_enable_261), 
            .CK(dac_clk_p_c), .Q(hb_bits[3])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(95[9] 103[41])
    defparam o_dw_bits_i3.GSR = "DISABLED";
    FD1P3AX o_dw_bits_i2 (.D(o_dw_bits_4__N_1187[2]), .SP(dac_clk_p_c_enable_261), 
            .CK(dac_clk_p_c), .Q(hb_bits[2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(95[9] 103[41])
    defparam o_dw_bits_i2.GSR = "DISABLED";
    FD1P3AX o_dw_bits_i1 (.D(o_dw_bits_4__N_1187[1]), .SP(dac_clk_p_c_enable_261), 
            .CK(dac_clk_p_c), .Q(hb_bits[1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(95[9] 103[41])
    defparam o_dw_bits_i1.GSR = "DISABLED";
    FD1P3AX r_word_i31 (.D(r_word_31__N_1196[31]), .SP(dac_clk_p_c_enable_261), 
            .CK(dac_clk_p_c), .Q(r_word[31])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i31.GSR = "DISABLED";
    FD1P3IX r_len__i3 (.D(r_len_3__N_1228[3]), .SP(dac_clk_p_c_enable_219), 
            .CD(n30028), .CK(dac_clk_p_c), .Q(r_len[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(64[9] 81[6])
    defparam r_len__i3.GSR = "DISABLED";
    FD1P3IX r_word_i1 (.D(idl_word[1]), .SP(dac_clk_p_c_enable_261), .CD(n12840), 
            .CK(dac_clk_p_c), .Q(r_word[1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i1.GSR = "DISABLED";
    FD1P3IX r_word_i2 (.D(idl_word[2]), .SP(dac_clk_p_c_enable_261), .CD(n12840), 
            .CK(dac_clk_p_c), .Q(r_word[2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i2.GSR = "DISABLED";
    FD1P3IX r_word_i3 (.D(idl_word[3]), .SP(dac_clk_p_c_enable_261), .CD(n12840), 
            .CK(dac_clk_p_c), .Q(r_word[3])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i3.GSR = "DISABLED";
    FD1P3IX o_dw_bits_i4 (.D(n29969), .SP(dac_clk_p_c_enable_261), .CD(n12840), 
            .CK(dac_clk_p_c), .Q(hb_bits[4])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(95[9] 103[41])
    defparam o_dw_bits_i4.GSR = "DISABLED";
    FD1P3IX o_dw_stb_36 (.D(o_dw_busy_N_1268), .SP(dac_clk_p_c_enable_219), 
            .CD(w_reset), .CK(dac_clk_p_c), .Q(hb_busy)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(64[9] 81[6])
    defparam o_dw_stb_36.GSR = "DISABLED";
    FD1P3IX r_word_i0 (.D(idl_word[0]), .SP(dac_clk_p_c_enable_261), .CD(n12840), 
            .CK(dac_clk_p_c), .Q(r_word[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i0.GSR = "DISABLED";
    FD1P3AX r_word_i30 (.D(r_word_31__N_1196[30]), .SP(dac_clk_p_c_enable_261), 
            .CK(dac_clk_p_c), .Q(r_word[30])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i30.GSR = "DISABLED";
    FD1P3AX r_word_i29 (.D(r_word_31__N_1196[29]), .SP(dac_clk_p_c_enable_261), 
            .CK(dac_clk_p_c), .Q(r_word[29])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i29.GSR = "DISABLED";
    FD1P3AX r_word_i28 (.D(r_word_31__N_1196[28]), .SP(dac_clk_p_c_enable_261), 
            .CK(dac_clk_p_c), .Q(r_word[28])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i28.GSR = "DISABLED";
    FD1P3AX r_word_i27 (.D(r_word_31__N_1196[27]), .SP(dac_clk_p_c_enable_261), 
            .CK(dac_clk_p_c), .Q(r_word[27])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i27.GSR = "DISABLED";
    FD1P3AX r_word_i26 (.D(r_word_31__N_1196[26]), .SP(dac_clk_p_c_enable_261), 
            .CK(dac_clk_p_c), .Q(r_word[26])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i26.GSR = "DISABLED";
    FD1P3AX r_word_i25 (.D(r_word_31__N_1196[25]), .SP(dac_clk_p_c_enable_261), 
            .CK(dac_clk_p_c), .Q(r_word[25])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i25.GSR = "DISABLED";
    FD1P3AX r_word_i24 (.D(r_word_31__N_1196[24]), .SP(dac_clk_p_c_enable_261), 
            .CK(dac_clk_p_c), .Q(r_word[24])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i24.GSR = "DISABLED";
    FD1P3AX r_word_i23 (.D(r_word_31__N_1196[23]), .SP(dac_clk_p_c_enable_261), 
            .CK(dac_clk_p_c), .Q(r_word[23])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i23.GSR = "DISABLED";
    FD1P3AX r_word_i22 (.D(r_word_31__N_1196[22]), .SP(dac_clk_p_c_enable_261), 
            .CK(dac_clk_p_c), .Q(r_word[22])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i22.GSR = "DISABLED";
    FD1P3AX r_word_i21 (.D(r_word_31__N_1196[21]), .SP(dac_clk_p_c_enable_261), 
            .CK(dac_clk_p_c), .Q(r_word[21])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i21.GSR = "DISABLED";
    FD1P3AX r_word_i20 (.D(r_word_31__N_1196[20]), .SP(dac_clk_p_c_enable_261), 
            .CK(dac_clk_p_c), .Q(r_word[20])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i20.GSR = "DISABLED";
    FD1P3AX r_word_i19 (.D(r_word_31__N_1196[19]), .SP(dac_clk_p_c_enable_261), 
            .CK(dac_clk_p_c), .Q(r_word[19])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i19.GSR = "DISABLED";
    FD1P3AX r_word_i18 (.D(r_word_31__N_1196[18]), .SP(dac_clk_p_c_enable_261), 
            .CK(dac_clk_p_c), .Q(r_word[18])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i18.GSR = "DISABLED";
    FD1P3AX r_word_i17 (.D(r_word_31__N_1196[17]), .SP(dac_clk_p_c_enable_261), 
            .CK(dac_clk_p_c), .Q(r_word[17])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i17.GSR = "DISABLED";
    FD1P3AX r_word_i16 (.D(r_word_31__N_1196[16]), .SP(dac_clk_p_c_enable_261), 
            .CK(dac_clk_p_c), .Q(r_word[16])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i16.GSR = "DISABLED";
    FD1P3AX r_word_i15 (.D(r_word_31__N_1196[15]), .SP(dac_clk_p_c_enable_261), 
            .CK(dac_clk_p_c), .Q(r_word[15])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i15.GSR = "DISABLED";
    FD1P3AX r_word_i14 (.D(r_word_31__N_1196[14]), .SP(dac_clk_p_c_enable_261), 
            .CK(dac_clk_p_c), .Q(r_word[14])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i14.GSR = "DISABLED";
    FD1P3AX r_word_i13 (.D(r_word_31__N_1196[13]), .SP(dac_clk_p_c_enable_261), 
            .CK(dac_clk_p_c), .Q(r_word[13])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i13.GSR = "DISABLED";
    FD1P3AX r_word_i12 (.D(r_word_31__N_1196[12]), .SP(dac_clk_p_c_enable_261), 
            .CK(dac_clk_p_c), .Q(r_word[12])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i12.GSR = "DISABLED";
    FD1P3AX r_word_i11 (.D(r_word_31__N_1196[11]), .SP(dac_clk_p_c_enable_261), 
            .CK(dac_clk_p_c), .Q(r_word[11])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i11.GSR = "DISABLED";
    FD1P3AX r_word_i10 (.D(r_word_31__N_1196[10]), .SP(dac_clk_p_c_enable_261), 
            .CK(dac_clk_p_c), .Q(r_word[10])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i10.GSR = "DISABLED";
    FD1P3AX r_word_i9 (.D(r_word_31__N_1196[9]), .SP(dac_clk_p_c_enable_261), 
            .CK(dac_clk_p_c), .Q(r_word[9])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i9.GSR = "DISABLED";
    FD1P3AX r_word_i8 (.D(r_word_31__N_1196[8]), .SP(dac_clk_p_c_enable_261), 
            .CK(dac_clk_p_c), .Q(r_word[8])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i8.GSR = "DISABLED";
    FD1P3AX r_word_i7 (.D(r_word_31__N_1196[7]), .SP(dac_clk_p_c_enable_261), 
            .CK(dac_clk_p_c), .Q(r_word[7])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i7.GSR = "DISABLED";
    FD1P3AX r_word_i6 (.D(r_word_31__N_1196[6]), .SP(dac_clk_p_c_enable_261), 
            .CK(dac_clk_p_c), .Q(r_word[6])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i6.GSR = "DISABLED";
    FD1P3AX r_word_i5 (.D(r_word_31__N_1196[5]), .SP(dac_clk_p_c_enable_261), 
            .CK(dac_clk_p_c), .Q(r_word[5])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i5.GSR = "DISABLED";
    FD1P3AX r_word_i4 (.D(r_word_31__N_1196[4]), .SP(dac_clk_p_c_enable_261), 
            .CK(dac_clk_p_c), .Q(r_word[4])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i4.GSR = "DISABLED";
    LUT4 i1_3_lut_4_lut_3_lut_4_lut (.A(r_len[0]), .B(r_len[1]), .C(r_len[2]), 
         .D(r_len[3]), .Z(n11587)) /* synthesis lut_function=(A (B)+!A !(B+!(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(80[14:26])
    defparam i1_3_lut_4_lut_3_lut_4_lut.init = 16'h9998;
    LUT4 i_stb_I_0_2_lut_rep_593 (.A(idl_stb), .B(hb_busy), .Z(n27258)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam i_stb_I_0_2_lut_rep_593.init = 16'h2222;
    LUT4 i11341_2_lut_3_lut (.A(idl_stb), .B(hb_busy), .C(n27259), .Z(o_dw_busy_N_1268)) /* synthesis lut_function=(A ((C)+!B)+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam i11341_2_lut_3_lut.init = 16'hf2f2;
    LUT4 i1_2_lut_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(nl_busy), 
         .D(hx_stb), .Z(dac_clk_p_c_enable_261)) /* synthesis lut_function=(!(A (B (C (D)))+!A (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h2fff;
    LUT4 i11334_2_lut (.A(idl_word[32]), .B(idl_word[33]), .Z(o_dw_bits_4__N_1278[3])) /* synthesis lut_function=(A (B)) */ ;
    defparam i11334_2_lut.init = 16'h8888;
    LUT4 o_dw_bits_4__I_0_i4_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(o_dw_bits_4__N_1278[3]), 
         .D(r_word[31]), .Z(o_dw_bits_4__N_1187[3])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam o_dw_bits_4__I_0_i4_3_lut_4_lut.init = 16'hfd20;
    LUT4 i1_2_lut_rep_476_3_lut (.A(idl_stb), .B(hb_busy), .C(n30027), 
         .Z(n27141)) /* synthesis lut_function=(A ((C)+!B)+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam i1_2_lut_rep_476_3_lut.init = 16'hf2f2;
    LUT4 r_word_31__I_0_i32_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[31]), 
         .D(r_word[27]), .Z(r_word_31__N_1196[31])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i32_3_lut_4_lut.init = 16'hfd20;
    LUT4 i23052_2_lut_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(nl_busy), 
         .D(hx_stb), .Z(n12840)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam i23052_2_lut_3_lut_4_lut.init = 16'h0ddd;
    LUT4 r_word_29__bdd_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(n26614), 
         .D(r_word[29]), .Z(o_dw_bits_4__N_1187[1])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_29__bdd_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i31_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[30]), 
         .D(r_word[26]), .Z(r_word_31__N_1196[30])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i31_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i30_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[29]), 
         .D(r_word[25]), .Z(r_word_31__N_1196[29])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i30_3_lut_4_lut.init = 16'hfd20;
    LUT4 o_dw_bits_4__I_0_i3_4_lut (.A(r_word[30]), .B(idl_word[31]), .C(n27258), 
         .D(o_dw_bits_4__N_1278[3]), .Z(o_dw_bits_4__N_1187[2])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(102[12] 103[41])
    defparam o_dw_bits_4__I_0_i3_4_lut.init = 16'hca0a;
    LUT4 mux_15_i4_4_lut (.A(r_len[3]), .B(o_dw_bits_4__N_1278[3]), .C(n27258), 
         .D(n20553), .Z(r_len_3__N_1228[3])) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(76[12] 81[6])
    defparam mux_15_i4_4_lut.init = 16'h3a35;
    LUT4 r_word_31__I_0_i29_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[28]), 
         .D(r_word[24]), .Z(r_word_31__N_1196[28])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i29_3_lut_4_lut.init = 16'hfd20;
    FD1P3IX r_len__i2 (.D(n11583), .SP(dac_clk_p_c_enable_332), .CD(n27141), 
            .CK(dac_clk_p_c), .Q(r_len[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(64[9] 81[6])
    defparam r_len__i2.GSR = "DISABLED";
    FD1P3IX r_len__i1 (.D(n11587), .SP(dac_clk_p_c_enable_332), .CD(n27141), 
            .CK(dac_clk_p_c), .Q(r_len[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(64[9] 81[6])
    defparam r_len__i1.GSR = "DISABLED";
    LUT4 r_word_31__I_0_i28_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[27]), 
         .D(r_word[23]), .Z(r_word_31__N_1196[27])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i28_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i27_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[26]), 
         .D(r_word[22]), .Z(r_word_31__N_1196[26])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i27_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i26_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[25]), 
         .D(r_word[21]), .Z(r_word_31__N_1196[25])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i26_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i25_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[24]), 
         .D(r_word[20]), .Z(r_word_31__N_1196[24])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i25_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i24_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[23]), 
         .D(r_word[19]), .Z(r_word_31__N_1196[23])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i24_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i23_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[22]), 
         .D(r_word[18]), .Z(r_word_31__N_1196[22])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i23_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_29__bdd_3_lut_24797 (.A(idl_word[30]), .B(idl_word[33]), 
         .C(idl_word[32]), .Z(n26614)) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam r_word_29__bdd_3_lut_24797.init = 16'h8c8c;
    LUT4 r_word_31__I_0_i22_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[21]), 
         .D(r_word[17]), .Z(r_word_31__N_1196[21])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i22_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i21_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[20]), 
         .D(r_word[16]), .Z(r_word_31__N_1196[20])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i21_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i20_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[19]), 
         .D(r_word[15]), .Z(r_word_31__N_1196[19])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i20_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i19_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[18]), 
         .D(r_word[14]), .Z(r_word_31__N_1196[18])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i19_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i18_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[17]), 
         .D(r_word[13]), .Z(r_word_31__N_1196[17])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i18_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i17_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[16]), 
         .D(r_word[12]), .Z(r_word_31__N_1196[16])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i17_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i16_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[15]), 
         .D(r_word[11]), .Z(r_word_31__N_1196[15])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i16_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_28__bdd_3_lut_25053 (.A(idl_word[29]), .B(idl_word[32]), 
         .C(idl_word[33]), .Z(n26931)) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam r_word_28__bdd_3_lut_25053.init = 16'h8c8c;
    LUT4 r_word_31__I_0_i15_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[14]), 
         .D(r_word[10]), .Z(r_word_31__N_1196[14])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i15_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i14_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[13]), 
         .D(r_word[9]), .Z(r_word_31__N_1196[13])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i14_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i13_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[12]), 
         .D(r_word[8]), .Z(r_word_31__N_1196[12])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i13_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i12_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[11]), 
         .D(r_word[7]), .Z(r_word_31__N_1196[11])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i12_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i11_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[10]), 
         .D(r_word[6]), .Z(r_word_31__N_1196[10])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i11_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i10_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[9]), 
         .D(r_word[5]), .Z(r_word_31__N_1196[9])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i10_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i9_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[8]), 
         .D(r_word[4]), .Z(r_word_31__N_1196[8])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i9_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i8_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[7]), 
         .D(r_word[3]), .Z(r_word_31__N_1196[7])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i8_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i7_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[6]), 
         .D(r_word[2]), .Z(r_word_31__N_1196[6])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i7_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i6_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[5]), 
         .D(r_word[1]), .Z(r_word_31__N_1196[5])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i6_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i5_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[4]), 
         .D(r_word[0]), .Z(r_word_31__N_1196[4])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i5_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_28__bdd_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(n26931), 
         .D(r_word[28]), .Z(o_dw_bits_4__N_1187[0])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_28__bdd_3_lut_4_lut.init = 16'hfd20;
    LUT4 i3_4_lut_rep_594 (.A(r_len[0]), .B(r_len[1]), .C(r_len[2]), .D(r_len[3]), 
         .Z(n27259)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(78[16:31])
    defparam i3_4_lut_rep_594.init = 16'hfffe;
    LUT4 i1_2_lut_4_lut (.A(r_len[0]), .B(r_len[1]), .C(r_len[2]), .D(r_len[3]), 
         .Z(n13[0])) /* synthesis lut_function=(!(A+!(B+(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(78[16:31])
    defparam i1_2_lut_4_lut.init = 16'h5554;
    LUT4 i1_3_lut_3_lut_4_lut (.A(r_len[0]), .B(r_len[1]), .C(r_len[3]), 
         .D(r_len[2]), .Z(n11583)) /* synthesis lut_function=(A (D)+!A (B (D)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(80[14:26])
    defparam i1_3_lut_3_lut_4_lut.init = 16'hee10;
    LUT4 i1_4_lut_4_lut (.A(r_len[0]), .B(r_len[1]), .C(r_len[3]), .D(r_len[2]), 
         .Z(n20553)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(80[14:26])
    defparam i1_4_lut_4_lut.init = 16'hffef;
    
endmodule
//
// Verilog Description of module hbpack
//

module hbpack (iw_word, n27423, wb_stb, wb_cyc, dac_clk_p_c_enable_471, 
            dac_clk_p_c, dac_clk_p_c_enable_405, n30028, \dec_bits[1] , 
            \dec_bits[4] , w_reset, o_pck_stb_N_764, cmd_loaded, dac_clk_p_c_enable_222, 
            cmd_loaded_N_767, n27443, i_cmd_wr, n22542, \iw_word[2] , 
            inc, n17754, \iw_word[31] , \iw_word[30] , \iw_word[29] , 
            \iw_word[28] , \iw_word[27] , \iw_word[26] , \iw_word[25] , 
            \iw_word[24] , \iw_word[23] , \iw_word[22] , \iw_word[21] , 
            \iw_word[20] , \iw_word[19] , \iw_word[18] , \iw_word[17] , 
            \iw_word[16] , \iw_word[15] , \iw_word[14] , \iw_word[13] , 
            \iw_word[12] , \iw_word[11] , \iw_word[10] , \iw_word[9] , 
            \iw_word[8] , \iw_word[7] , \iw_word[6] , \iw_word[5] , 
            \iw_word[4] , \iw_word[3] , \iw_word[1] , \dec_bits[0] , 
            dac_clk_p_c_enable_374, n45, n46, dac_clk_p_c_enable_138, 
            n30027, newaddr_N_989) /* synthesis syn_module_defined=1 */ ;
    output [33:0]iw_word;
    output n27423;
    input wb_stb;
    input wb_cyc;
    output dac_clk_p_c_enable_471;
    input dac_clk_p_c;
    input dac_clk_p_c_enable_405;
    input n30028;
    input \dec_bits[1] ;
    input \dec_bits[4] ;
    input w_reset;
    input o_pck_stb_N_764;
    output cmd_loaded;
    input dac_clk_p_c_enable_222;
    input cmd_loaded_N_767;
    output n27443;
    output i_cmd_wr;
    output n22542;
    output \iw_word[2] ;
    input inc;
    output n17754;
    output \iw_word[31] ;
    output \iw_word[30] ;
    output \iw_word[29] ;
    output \iw_word[28] ;
    output \iw_word[27] ;
    output \iw_word[26] ;
    output \iw_word[25] ;
    output \iw_word[24] ;
    output \iw_word[23] ;
    output \iw_word[22] ;
    output \iw_word[21] ;
    output \iw_word[20] ;
    output \iw_word[19] ;
    output \iw_word[18] ;
    output \iw_word[17] ;
    output \iw_word[16] ;
    output \iw_word[15] ;
    output \iw_word[14] ;
    output \iw_word[13] ;
    output \iw_word[12] ;
    output \iw_word[11] ;
    output \iw_word[10] ;
    output \iw_word[9] ;
    output \iw_word[8] ;
    output \iw_word[7] ;
    output \iw_word[6] ;
    output \iw_word[5] ;
    output \iw_word[4] ;
    output \iw_word[3] ;
    output \iw_word[1] ;
    input \dec_bits[0] ;
    input dac_clk_p_c_enable_374;
    input n45;
    input n46;
    output dac_clk_p_c_enable_138;
    input n30027;
    output newaddr_N_989;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[49:58])
    wire [33:0]r_word;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(71[13:19])
    wire [33:0]n14;
    
    wire iw_stb;
    wire [33:0]iw_word_c;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(71[14:21])
    
    wire n27235;
    
    LUT4 i11393_2_lut_3_lut_4_lut (.A(iw_word[32]), .B(n27423), .C(wb_stb), 
         .D(wb_cyc), .Z(dac_clk_p_c_enable_471)) /* synthesis lut_function=(A (C)+!A (B (C+!(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(83[9] 84[65])
    defparam i11393_2_lut_3_lut_4_lut.init = 16'hf0f4;
    FD1P3IX r_word__i0 (.D(n14[0]), .SP(dac_clk_p_c_enable_405), .CD(n30028), 
            .CK(dac_clk_p_c), .Q(r_word[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i0.GSR = "DISABLED";
    FD1P3IX o_pck_word__i0 (.D(r_word[0]), .SP(dac_clk_p_c_enable_405), 
            .CD(n30028), .CK(dac_clk_p_c), .Q(iw_word[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i0.GSR = "DISABLED";
    LUT4 i11719_2_lut (.A(\dec_bits[1] ), .B(\dec_bits[4] ), .Z(n14[1])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11719_2_lut.init = 16'h2222;
    FD1S3IX o_pck_stb_24 (.D(o_pck_stb_N_764), .CK(dac_clk_p_c), .CD(w_reset), 
            .Q(iw_stb)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(83[9] 84[65])
    defparam o_pck_stb_24.GSR = "DISABLED";
    FD1P3IX cmd_loaded_23 (.D(cmd_loaded_N_767), .SP(dac_clk_p_c_enable_222), 
            .CD(n30028), .CK(dac_clk_p_c), .Q(cmd_loaded)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(74[9] 80[23])
    defparam cmd_loaded_23.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_778 (.A(iw_stb), .B(iw_word_c[33]), .Z(n27443)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(83[9] 84[65])
    defparam i1_2_lut_rep_778.init = 16'h2222;
    LUT4 i1_2_lut_3_lut (.A(iw_stb), .B(iw_word_c[33]), .C(iw_word[32]), 
         .Z(i_cmd_wr)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(83[9] 84[65])
    defparam i1_2_lut_3_lut.init = 16'h2020;
    LUT4 i20187_3_lut_3_lut (.A(iw_stb), .B(iw_word_c[33]), .C(wb_stb), 
         .Z(n22542)) /* synthesis lut_function=(A ((C)+!B)+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(83[9] 84[65])
    defparam i20187_3_lut_3_lut.init = 16'hf2f2;
    LUT4 i15965_3_lut_4_lut (.A(wb_cyc), .B(n27235), .C(\iw_word[2] ), 
         .D(inc), .Z(n17754)) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(83[9] 84[65])
    defparam i15965_3_lut_4_lut.init = 16'hfb40;
    FD1P3IX o_pck_word__i33 (.D(r_word[33]), .SP(dac_clk_p_c_enable_405), 
            .CD(w_reset), .CK(dac_clk_p_c), .Q(iw_word_c[33])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i33.GSR = "DISABLED";
    FD1P3IX o_pck_word__i32 (.D(r_word[32]), .SP(dac_clk_p_c_enable_405), 
            .CD(w_reset), .CK(dac_clk_p_c), .Q(iw_word[32])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i32.GSR = "DISABLED";
    FD1P3IX o_pck_word__i31 (.D(r_word[31]), .SP(dac_clk_p_c_enable_405), 
            .CD(w_reset), .CK(dac_clk_p_c), .Q(\iw_word[31] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i31.GSR = "DISABLED";
    FD1P3IX o_pck_word__i30 (.D(r_word[30]), .SP(dac_clk_p_c_enable_405), 
            .CD(w_reset), .CK(dac_clk_p_c), .Q(\iw_word[30] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i30.GSR = "DISABLED";
    FD1P3IX o_pck_word__i29 (.D(r_word[29]), .SP(dac_clk_p_c_enable_405), 
            .CD(w_reset), .CK(dac_clk_p_c), .Q(\iw_word[29] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i29.GSR = "DISABLED";
    FD1P3IX o_pck_word__i28 (.D(r_word[28]), .SP(dac_clk_p_c_enable_405), 
            .CD(w_reset), .CK(dac_clk_p_c), .Q(\iw_word[28] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i28.GSR = "DISABLED";
    FD1P3IX o_pck_word__i27 (.D(r_word[27]), .SP(dac_clk_p_c_enable_405), 
            .CD(w_reset), .CK(dac_clk_p_c), .Q(\iw_word[27] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i27.GSR = "DISABLED";
    FD1P3IX o_pck_word__i26 (.D(r_word[26]), .SP(dac_clk_p_c_enable_405), 
            .CD(w_reset), .CK(dac_clk_p_c), .Q(\iw_word[26] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i26.GSR = "DISABLED";
    FD1P3IX o_pck_word__i25 (.D(r_word[25]), .SP(dac_clk_p_c_enable_405), 
            .CD(w_reset), .CK(dac_clk_p_c), .Q(\iw_word[25] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i25.GSR = "DISABLED";
    FD1P3IX o_pck_word__i24 (.D(r_word[24]), .SP(dac_clk_p_c_enable_405), 
            .CD(w_reset), .CK(dac_clk_p_c), .Q(\iw_word[24] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i24.GSR = "DISABLED";
    FD1P3IX o_pck_word__i23 (.D(r_word[23]), .SP(dac_clk_p_c_enable_405), 
            .CD(n30028), .CK(dac_clk_p_c), .Q(\iw_word[23] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i23.GSR = "DISABLED";
    FD1P3IX o_pck_word__i22 (.D(r_word[22]), .SP(dac_clk_p_c_enable_405), 
            .CD(w_reset), .CK(dac_clk_p_c), .Q(\iw_word[22] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i22.GSR = "DISABLED";
    FD1P3IX o_pck_word__i21 (.D(r_word[21]), .SP(dac_clk_p_c_enable_405), 
            .CD(n30028), .CK(dac_clk_p_c), .Q(\iw_word[21] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i21.GSR = "DISABLED";
    FD1P3IX o_pck_word__i20 (.D(r_word[20]), .SP(dac_clk_p_c_enable_405), 
            .CD(n30028), .CK(dac_clk_p_c), .Q(\iw_word[20] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i20.GSR = "DISABLED";
    FD1P3IX o_pck_word__i19 (.D(r_word[19]), .SP(dac_clk_p_c_enable_405), 
            .CD(n30028), .CK(dac_clk_p_c), .Q(\iw_word[19] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i19.GSR = "DISABLED";
    FD1P3IX o_pck_word__i18 (.D(r_word[18]), .SP(dac_clk_p_c_enable_405), 
            .CD(n30028), .CK(dac_clk_p_c), .Q(\iw_word[18] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i18.GSR = "DISABLED";
    FD1P3IX o_pck_word__i17 (.D(r_word[17]), .SP(dac_clk_p_c_enable_405), 
            .CD(n30028), .CK(dac_clk_p_c), .Q(\iw_word[17] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i17.GSR = "DISABLED";
    FD1P3IX o_pck_word__i16 (.D(r_word[16]), .SP(dac_clk_p_c_enable_405), 
            .CD(n30028), .CK(dac_clk_p_c), .Q(\iw_word[16] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i16.GSR = "DISABLED";
    FD1P3IX o_pck_word__i15 (.D(r_word[15]), .SP(dac_clk_p_c_enable_405), 
            .CD(n30028), .CK(dac_clk_p_c), .Q(\iw_word[15] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i15.GSR = "DISABLED";
    FD1P3IX o_pck_word__i14 (.D(r_word[14]), .SP(dac_clk_p_c_enable_405), 
            .CD(n30028), .CK(dac_clk_p_c), .Q(\iw_word[14] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i14.GSR = "DISABLED";
    FD1P3IX o_pck_word__i13 (.D(r_word[13]), .SP(dac_clk_p_c_enable_405), 
            .CD(n30028), .CK(dac_clk_p_c), .Q(\iw_word[13] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i13.GSR = "DISABLED";
    FD1P3IX o_pck_word__i12 (.D(r_word[12]), .SP(dac_clk_p_c_enable_405), 
            .CD(n30028), .CK(dac_clk_p_c), .Q(\iw_word[12] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i12.GSR = "DISABLED";
    FD1P3IX o_pck_word__i11 (.D(r_word[11]), .SP(dac_clk_p_c_enable_405), 
            .CD(n30028), .CK(dac_clk_p_c), .Q(\iw_word[11] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i11.GSR = "DISABLED";
    FD1P3IX o_pck_word__i10 (.D(r_word[10]), .SP(dac_clk_p_c_enable_405), 
            .CD(n30028), .CK(dac_clk_p_c), .Q(\iw_word[10] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i10.GSR = "DISABLED";
    FD1P3IX o_pck_word__i9 (.D(r_word[9]), .SP(dac_clk_p_c_enable_405), 
            .CD(n30028), .CK(dac_clk_p_c), .Q(\iw_word[9] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i9.GSR = "DISABLED";
    FD1P3IX o_pck_word__i8 (.D(r_word[8]), .SP(dac_clk_p_c_enable_405), 
            .CD(n30028), .CK(dac_clk_p_c), .Q(\iw_word[8] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i8.GSR = "DISABLED";
    FD1P3IX o_pck_word__i7 (.D(r_word[7]), .SP(dac_clk_p_c_enable_405), 
            .CD(n30028), .CK(dac_clk_p_c), .Q(\iw_word[7] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i7.GSR = "DISABLED";
    FD1P3IX o_pck_word__i6 (.D(r_word[6]), .SP(dac_clk_p_c_enable_405), 
            .CD(n30028), .CK(dac_clk_p_c), .Q(\iw_word[6] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i6.GSR = "DISABLED";
    FD1P3IX o_pck_word__i5 (.D(r_word[5]), .SP(dac_clk_p_c_enable_405), 
            .CD(n30028), .CK(dac_clk_p_c), .Q(\iw_word[5] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i5.GSR = "DISABLED";
    FD1P3IX o_pck_word__i4 (.D(r_word[4]), .SP(dac_clk_p_c_enable_405), 
            .CD(n30028), .CK(dac_clk_p_c), .Q(\iw_word[4] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i4.GSR = "DISABLED";
    FD1P3IX o_pck_word__i3 (.D(r_word[3]), .SP(dac_clk_p_c_enable_405), 
            .CD(n30028), .CK(dac_clk_p_c), .Q(\iw_word[3] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i3.GSR = "DISABLED";
    FD1P3IX o_pck_word__i2 (.D(r_word[2]), .SP(dac_clk_p_c_enable_405), 
            .CD(n30028), .CK(dac_clk_p_c), .Q(\iw_word[2] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i2.GSR = "DISABLED";
    FD1P3IX o_pck_word__i1 (.D(r_word[1]), .SP(dac_clk_p_c_enable_405), 
            .CD(n30028), .CK(dac_clk_p_c), .Q(\iw_word[1] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i1.GSR = "DISABLED";
    LUT4 i11329_2_lut (.A(\dec_bits[0] ), .B(\dec_bits[4] ), .Z(n14[0])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11329_2_lut.init = 16'h2222;
    LUT4 i11691_2_lut (.A(r_word[27]), .B(\dec_bits[4] ), .Z(n14[31])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11691_2_lut.init = 16'h2222;
    LUT4 i11692_2_lut (.A(r_word[26]), .B(\dec_bits[4] ), .Z(n14[30])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11692_2_lut.init = 16'h2222;
    LUT4 i11693_2_lut (.A(r_word[25]), .B(\dec_bits[4] ), .Z(n14[29])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11693_2_lut.init = 16'h2222;
    LUT4 i11694_2_lut (.A(r_word[24]), .B(\dec_bits[4] ), .Z(n14[28])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11694_2_lut.init = 16'h2222;
    LUT4 i11695_2_lut (.A(r_word[23]), .B(\dec_bits[4] ), .Z(n14[27])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11695_2_lut.init = 16'h2222;
    LUT4 i11696_2_lut (.A(r_word[22]), .B(\dec_bits[4] ), .Z(n14[26])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11696_2_lut.init = 16'h2222;
    LUT4 i11697_2_lut (.A(r_word[21]), .B(\dec_bits[4] ), .Z(n14[25])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11697_2_lut.init = 16'h2222;
    LUT4 i11698_2_lut (.A(r_word[20]), .B(\dec_bits[4] ), .Z(n14[24])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11698_2_lut.init = 16'h2222;
    LUT4 i11699_2_lut (.A(r_word[19]), .B(\dec_bits[4] ), .Z(n14[23])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11699_2_lut.init = 16'h2222;
    LUT4 i11700_2_lut (.A(r_word[18]), .B(\dec_bits[4] ), .Z(n14[22])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11700_2_lut.init = 16'h2222;
    LUT4 i11701_2_lut (.A(r_word[17]), .B(\dec_bits[4] ), .Z(n14[21])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11701_2_lut.init = 16'h2222;
    LUT4 i11702_2_lut (.A(r_word[16]), .B(\dec_bits[4] ), .Z(n14[20])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11702_2_lut.init = 16'h2222;
    LUT4 i11703_2_lut (.A(r_word[15]), .B(\dec_bits[4] ), .Z(n14[19])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11703_2_lut.init = 16'h2222;
    LUT4 i11704_2_lut (.A(r_word[14]), .B(\dec_bits[4] ), .Z(n14[18])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11704_2_lut.init = 16'h2222;
    LUT4 i11705_2_lut (.A(r_word[13]), .B(\dec_bits[4] ), .Z(n14[17])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11705_2_lut.init = 16'h2222;
    LUT4 i11706_2_lut (.A(r_word[12]), .B(\dec_bits[4] ), .Z(n14[16])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11706_2_lut.init = 16'h2222;
    LUT4 i11707_2_lut (.A(r_word[11]), .B(\dec_bits[4] ), .Z(n14[15])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11707_2_lut.init = 16'h2222;
    LUT4 i11708_2_lut (.A(r_word[10]), .B(\dec_bits[4] ), .Z(n14[14])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11708_2_lut.init = 16'h2222;
    LUT4 i11709_2_lut (.A(r_word[9]), .B(\dec_bits[4] ), .Z(n14[13])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11709_2_lut.init = 16'h2222;
    LUT4 i11710_2_lut (.A(r_word[8]), .B(\dec_bits[4] ), .Z(n14[12])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11710_2_lut.init = 16'h2222;
    LUT4 i11711_2_lut (.A(r_word[7]), .B(\dec_bits[4] ), .Z(n14[11])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11711_2_lut.init = 16'h2222;
    LUT4 i11712_2_lut (.A(r_word[6]), .B(\dec_bits[4] ), .Z(n14[10])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11712_2_lut.init = 16'h2222;
    LUT4 i11713_2_lut (.A(r_word[5]), .B(\dec_bits[4] ), .Z(n14[9])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11713_2_lut.init = 16'h2222;
    LUT4 i11714_2_lut (.A(r_word[4]), .B(\dec_bits[4] ), .Z(n14[8])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11714_2_lut.init = 16'h2222;
    LUT4 i11715_2_lut (.A(r_word[3]), .B(\dec_bits[4] ), .Z(n14[7])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11715_2_lut.init = 16'h2222;
    LUT4 i11716_2_lut (.A(r_word[2]), .B(\dec_bits[4] ), .Z(n14[6])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11716_2_lut.init = 16'h2222;
    LUT4 i11717_2_lut (.A(r_word[1]), .B(\dec_bits[4] ), .Z(n14[5])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11717_2_lut.init = 16'h2222;
    LUT4 i11718_2_lut (.A(r_word[0]), .B(\dec_bits[4] ), .Z(n14[4])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11718_2_lut.init = 16'h2222;
    FD1P3IX r_word__i33 (.D(\dec_bits[1] ), .SP(dac_clk_p_c_enable_374), 
            .CD(n30028), .CK(dac_clk_p_c), .Q(r_word[33])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i33.GSR = "DISABLED";
    FD1P3IX r_word__i32 (.D(\dec_bits[0] ), .SP(dac_clk_p_c_enable_374), 
            .CD(n30028), .CK(dac_clk_p_c), .Q(r_word[32])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i32.GSR = "DISABLED";
    FD1P3IX r_word__i31 (.D(n14[31]), .SP(dac_clk_p_c_enable_405), .CD(n30028), 
            .CK(dac_clk_p_c), .Q(r_word[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i31.GSR = "DISABLED";
    FD1P3IX r_word__i30 (.D(n14[30]), .SP(dac_clk_p_c_enable_405), .CD(n30028), 
            .CK(dac_clk_p_c), .Q(r_word[30])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i30.GSR = "DISABLED";
    FD1P3IX r_word__i29 (.D(n14[29]), .SP(dac_clk_p_c_enable_405), .CD(n30028), 
            .CK(dac_clk_p_c), .Q(r_word[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i29.GSR = "DISABLED";
    FD1P3IX r_word__i28 (.D(n14[28]), .SP(dac_clk_p_c_enable_405), .CD(n30028), 
            .CK(dac_clk_p_c), .Q(r_word[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i28.GSR = "DISABLED";
    FD1P3IX r_word__i27 (.D(n14[27]), .SP(dac_clk_p_c_enable_405), .CD(n30028), 
            .CK(dac_clk_p_c), .Q(r_word[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i27.GSR = "DISABLED";
    FD1P3IX r_word__i26 (.D(n14[26]), .SP(dac_clk_p_c_enable_405), .CD(n30028), 
            .CK(dac_clk_p_c), .Q(r_word[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i26.GSR = "DISABLED";
    FD1P3IX r_word__i25 (.D(n14[25]), .SP(dac_clk_p_c_enable_405), .CD(n30028), 
            .CK(dac_clk_p_c), .Q(r_word[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i25.GSR = "DISABLED";
    FD1P3IX r_word__i24 (.D(n14[24]), .SP(dac_clk_p_c_enable_405), .CD(n30028), 
            .CK(dac_clk_p_c), .Q(r_word[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i24.GSR = "DISABLED";
    FD1P3IX r_word__i23 (.D(n14[23]), .SP(dac_clk_p_c_enable_405), .CD(n30028), 
            .CK(dac_clk_p_c), .Q(r_word[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i23.GSR = "DISABLED";
    FD1P3IX r_word__i22 (.D(n14[22]), .SP(dac_clk_p_c_enable_405), .CD(n30028), 
            .CK(dac_clk_p_c), .Q(r_word[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i22.GSR = "DISABLED";
    FD1P3IX r_word__i21 (.D(n14[21]), .SP(dac_clk_p_c_enable_405), .CD(n30028), 
            .CK(dac_clk_p_c), .Q(r_word[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i21.GSR = "DISABLED";
    FD1P3IX r_word__i20 (.D(n14[20]), .SP(dac_clk_p_c_enable_405), .CD(n30028), 
            .CK(dac_clk_p_c), .Q(r_word[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i20.GSR = "DISABLED";
    FD1P3IX r_word__i19 (.D(n14[19]), .SP(dac_clk_p_c_enable_405), .CD(n30028), 
            .CK(dac_clk_p_c), .Q(r_word[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i19.GSR = "DISABLED";
    FD1P3IX r_word__i18 (.D(n14[18]), .SP(dac_clk_p_c_enable_405), .CD(n30028), 
            .CK(dac_clk_p_c), .Q(r_word[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i18.GSR = "DISABLED";
    FD1P3IX r_word__i17 (.D(n14[17]), .SP(dac_clk_p_c_enable_405), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i17.GSR = "DISABLED";
    FD1P3IX r_word__i16 (.D(n14[16]), .SP(dac_clk_p_c_enable_405), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i16.GSR = "DISABLED";
    FD1P3IX r_word__i15 (.D(n14[15]), .SP(dac_clk_p_c_enable_405), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i15.GSR = "DISABLED";
    FD1P3IX r_word__i14 (.D(n14[14]), .SP(dac_clk_p_c_enable_405), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i14.GSR = "DISABLED";
    FD1P3IX r_word__i13 (.D(n14[13]), .SP(dac_clk_p_c_enable_405), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i13.GSR = "DISABLED";
    FD1P3IX r_word__i12 (.D(n14[12]), .SP(dac_clk_p_c_enable_405), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i12.GSR = "DISABLED";
    FD1P3IX r_word__i11 (.D(n14[11]), .SP(dac_clk_p_c_enable_405), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i11.GSR = "DISABLED";
    FD1P3IX r_word__i10 (.D(n14[10]), .SP(dac_clk_p_c_enable_405), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i10.GSR = "DISABLED";
    FD1P3IX r_word__i9 (.D(n14[9]), .SP(dac_clk_p_c_enable_405), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i9.GSR = "DISABLED";
    FD1P3IX r_word__i8 (.D(n14[8]), .SP(dac_clk_p_c_enable_405), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i8.GSR = "DISABLED";
    FD1P3IX r_word__i7 (.D(n14[7]), .SP(dac_clk_p_c_enable_405), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i7.GSR = "DISABLED";
    FD1P3IX r_word__i6 (.D(n14[6]), .SP(dac_clk_p_c_enable_405), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i6.GSR = "DISABLED";
    FD1P3IX r_word__i5 (.D(n14[5]), .SP(dac_clk_p_c_enable_405), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i5.GSR = "DISABLED";
    FD1P3IX r_word__i4 (.D(n14[4]), .SP(dac_clk_p_c_enable_405), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i4.GSR = "DISABLED";
    FD1P3IX r_word__i3 (.D(n45), .SP(dac_clk_p_c_enable_405), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i3.GSR = "DISABLED";
    FD1P3IX r_word__i2 (.D(n46), .SP(dac_clk_p_c_enable_405), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i2.GSR = "DISABLED";
    FD1P3IX r_word__i1 (.D(n14[1]), .SP(dac_clk_p_c_enable_405), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i1.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_758 (.A(iw_word_c[33]), .B(iw_stb), .Z(n27423)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(83[9] 84[65])
    defparam i1_2_lut_rep_758.init = 16'h8888;
    LUT4 i1_2_lut_rep_469_3_lut_4_lut (.A(iw_word_c[33]), .B(iw_stb), .C(wb_cyc), 
         .D(iw_word[32]), .Z(dac_clk_p_c_enable_138)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(83[9] 84[65])
    defparam i1_2_lut_rep_469_3_lut_4_lut.init = 16'h0008;
    LUT4 i2_2_lut_rep_570_3_lut (.A(iw_word_c[33]), .B(iw_stb), .C(iw_word[32]), 
         .Z(n27235)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(83[9] 84[65])
    defparam i2_2_lut_rep_570_3_lut.init = 16'h0808;
    LUT4 i1_2_lut_3_lut_4_lut (.A(iw_word_c[33]), .B(iw_stb), .C(n30027), 
         .D(iw_word[32]), .Z(newaddr_N_989)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(83[9] 84[65])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0008;
    
endmodule
//
// Verilog Description of module hbgenhex
//

module hbgenhex (hx_stb, dac_clk_p_c, n30028, hb_busy, hb_bits, \w_gx_char[0] , 
            \w_gx_char[1] , \w_gx_char[2] , \w_gx_char[3] , \w_gx_char[4] , 
            \w_gx_char[5] , \w_gx_char[6] , dac_clk_p_c_enable_332, GND_net, 
            VCC_net, n11763, nl_busy, n30027, n27258, dac_clk_p_c_enable_219) /* synthesis syn_module_defined=1 */ ;
    output hx_stb;
    input dac_clk_p_c;
    input n30028;
    input hb_busy;
    input [4:0]hb_bits;
    output \w_gx_char[0] ;
    output \w_gx_char[1] ;
    output \w_gx_char[2] ;
    output \w_gx_char[3] ;
    output \w_gx_char[4] ;
    output \w_gx_char[5] ;
    output \w_gx_char[6] ;
    output dac_clk_p_c_enable_332;
    input GND_net;
    input VCC_net;
    output n11763;
    input nl_busy;
    input n30027;
    input n27258;
    output dac_clk_p_c_enable_219;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[49:58])
    
    wire dac_clk_p_c_enable_1, n20902;
    
    FD1P3IX o_gx_stb_13 (.D(hb_busy), .SP(dac_clk_p_c_enable_1), .CD(n30028), 
            .CK(dac_clk_p_c), .Q(hx_stb)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=132, LSE_RLINE=133 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbgenhex.v(74[9] 78[21])
    defparam o_gx_stb_13.GSR = "DISABLED";
    SP8KC mux_98 (.DI0(GND_net), .DI1(GND_net), .DI2(GND_net), .DI3(GND_net), 
          .DI4(GND_net), .DI5(GND_net), .DI6(GND_net), .DI7(GND_net), 
          .DI8(GND_net), .AD0(GND_net), .AD1(GND_net), .AD2(GND_net), 
          .AD3(hb_bits[0]), .AD4(hb_bits[1]), .AD5(hb_bits[2]), .AD6(hb_bits[3]), 
          .AD7(hb_bits[4]), .AD8(GND_net), .AD9(GND_net), .AD10(GND_net), 
          .AD11(GND_net), .AD12(GND_net), .CE(dac_clk_p_c_enable_332), 
          .OCE(VCC_net), .CLK(dac_clk_p_c), .WE(GND_net), .CS0(GND_net), 
          .CS1(GND_net), .CS2(GND_net), .RST(GND_net), .DO0(\w_gx_char[0] ), 
          .DO1(\w_gx_char[1] ), .DO2(\w_gx_char[2] ), .DO3(\w_gx_char[3] ), 
          .DO4(\w_gx_char[4] ), .DO5(\w_gx_char[5] ), .DO6(\w_gx_char[6] ));
    defparam mux_98.DATA_WIDTH = 9;
    defparam mux_98.REGMODE = "NOREG";
    defparam mux_98.CSDECODE = "0b000";
    defparam mux_98.WRITEMODE = "NORMAL";
    defparam mux_98.GSR = "DISABLED";
    defparam mux_98.RESETMODE = "ASYNC";
    defparam mux_98.ASYNC_RESET_RELEASE = "SYNC";
    defparam mux_98.INIT_DATA = "STATIC";
    defparam mux_98.INITVAL_00 = "0x01A0D01A0D0B44908A5401A0D01A0D0A641096520CC650C8630C4610723806E3606A340663206230";
    defparam mux_98.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_98.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_98.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_98.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_98.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_98.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_98.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_98.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_98.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_98.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_98.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_98.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_98.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_98.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_98.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_98.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_98.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_98.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_98.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_98.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_98.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_98.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_98.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_98.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_98.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_98.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_98.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_98.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_98.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_98.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_98.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    LUT4 i1_4_lut (.A(\w_gx_char[3] ), .B(\w_gx_char[0] ), .C(\w_gx_char[2] ), 
         .D(n20902), .Z(n11763)) /* synthesis lut_function=((((D)+!C)+!B)+!A) */ ;
    defparam i1_4_lut.init = 16'hff7f;
    LUT4 i1_4_lut_adj_142 (.A(\w_gx_char[1] ), .B(\w_gx_char[6] ), .C(\w_gx_char[4] ), 
         .D(\w_gx_char[5] ), .Z(n20902)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_142.init = 16'hfffe;
    LUT4 i23038_2_lut_rep_565 (.A(hx_stb), .B(nl_busy), .Z(dac_clk_p_c_enable_332)) /* synthesis lut_function=(!(A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(76[16:26])
    defparam i23038_2_lut_rep_565.init = 16'h7777;
    LUT4 i690_2_lut_3_lut (.A(hx_stb), .B(nl_busy), .C(n30027), .Z(dac_clk_p_c_enable_1)) /* synthesis lut_function=(((C)+!B)+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(76[16:26])
    defparam i690_2_lut_3_lut.init = 16'hf7f7;
    LUT4 i1_2_lut_3_lut_4_lut (.A(hx_stb), .B(nl_busy), .C(n30027), .D(n27258), 
         .Z(dac_clk_p_c_enable_219)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(76[16:26])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfff7;
    
endmodule
//
// Verilog Description of module hbdechex
//

module hbdechex (dac_clk_p_c, dec_bits, n45, \dec_bits[0] , w_reset, 
            n46, rx_stb, \rx_data[3] , \rx_data[6] , \rx_data[2] , 
            \rx_data[4] , \rx_data[5] , \rx_data[0] , \rx_data[1] , 
            n30028, \dec_bits[1] , n30027, cmd_loaded, o_pck_stb_N_764, 
            dac_clk_p_c_enable_222, cmd_loaded_N_767, dac_clk_p_c_enable_405, 
            dac_clk_p_c_enable_374) /* synthesis syn_module_defined=1 */ ;
    input dac_clk_p_c;
    output [4:0]dec_bits;
    output n45;
    output \dec_bits[0] ;
    output w_reset;
    output n46;
    input rx_stb;
    input \rx_data[3] ;
    input \rx_data[6] ;
    input \rx_data[2] ;
    input \rx_data[4] ;
    input \rx_data[5] ;
    input \rx_data[0] ;
    input \rx_data[1] ;
    output n30028;
    output \dec_bits[1] ;
    output n30027;
    input cmd_loaded;
    output o_pck_stb_N_764;
    output dac_clk_p_c_enable_222;
    output cmd_loaded_N_767;
    output dac_clk_p_c_enable_405;
    output dac_clk_p_c_enable_374;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[49:58])
    
    wire dec_stb, o_dh_stb_N_622;
    wire [4:0]dec_bits_c;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(69[13:21])
    wire [4:0]o_dh_bits_4__N_595;
    
    wire o_reset_N_624, n21302, n20095, n21300, n20272, n20844, 
        n35, n29910, n50, n20160, n20702, n47, n9, n50_adj_3039, 
        n27445, n27244, n27447, n52, n27982, n27983, n20978, n27986, 
        n20988, n20826, n27984, n4, n27448, n20097, n27245, n26373, 
        n26376, n28999, n29909, n41, n20832, n27135, n20850, n49, 
        n20974, n42, n33, n35_adj_3040, n20982;
    
    FD1S3AX o_dh_stb_35 (.D(o_dh_stb_N_622), .CK(dac_clk_p_c), .Q(dec_stb)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=30, LSE_LLINE=93, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(57[9] 58[47])
    defparam o_dh_stb_35.GSR = "DISABLED";
    LUT4 i1_2_lut (.A(dec_bits[4]), .B(dec_bits_c[3]), .Z(n45)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(60[9] 100[5])
    defparam i1_2_lut.init = 16'h4444;
    FD1S3AX o_dh_bits_i0 (.D(o_dh_bits_4__N_595[0]), .CK(dac_clk_p_c), .Q(\dec_bits[0] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=30, LSE_LLINE=93, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(60[9] 100[5])
    defparam o_dh_bits_i0.GSR = "DISABLED";
    FD1S3AY o_reset_34 (.D(o_reset_N_624), .CK(dac_clk_p_c), .Q(w_reset)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=30, LSE_LLINE=93, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(53[9] 54[46])
    defparam o_reset_34.GSR = "DISABLED";
    LUT4 i1_2_lut_adj_123 (.A(dec_bits[4]), .B(dec_bits_c[2]), .Z(n46)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(60[9] 100[5])
    defparam i1_2_lut_adj_123.init = 16'h4444;
    LUT4 i_stb_I_0_58_4_lut (.A(rx_stb), .B(n21302), .C(n20095), .D(n21300), 
         .Z(o_dh_stb_N_622)) /* synthesis lut_function=(!((B (C (D)))+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(58[15:46])
    defparam i_stb_I_0_58_4_lut.init = 16'h2aaa;
    LUT4 i1_3_lut (.A(\rx_data[3] ), .B(\rx_data[6] ), .C(\rx_data[2] ), 
         .Z(n21302)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_adj_124 (.A(\rx_data[4] ), .B(\rx_data[5] ), .Z(n20095)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_124.init = 16'h8888;
    LUT4 i1_2_lut_adj_125 (.A(\rx_data[0] ), .B(\rx_data[1] ), .Z(n21300)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_125.init = 16'h8888;
    LUT4 i1_4_lut (.A(n20272), .B(\rx_data[6] ), .C(n20844), .D(n35), 
         .Z(o_dh_bits_4__N_595[0])) /* synthesis lut_function=((B (C+(D))+!B (C))+!A) */ ;
    defparam i1_4_lut.init = 16'hfdf5;
    LUT4 i1_4_lut_adj_126 (.A(n29910), .B(\rx_data[6] ), .C(n50), .D(n20160), 
         .Z(n20844)) /* synthesis lut_function=(A+(B (C)+!B (C+!(D)))) */ ;
    defparam i1_4_lut_adj_126.init = 16'hfafb;
    LUT4 i1_4_lut_adj_127 (.A(\rx_data[5] ), .B(\rx_data[4] ), .C(\rx_data[6] ), 
         .D(\rx_data[3] ), .Z(n20702)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(87[3:8])
    defparam i1_4_lut_adj_127.init = 16'hfff7;
    LUT4 i1_3_lut_adj_128 (.A(\rx_data[4] ), .B(\rx_data[3] ), .C(n47), 
         .Z(n35)) /* synthesis lut_function=(A (B+!(C))+!A (B)) */ ;
    defparam i1_3_lut_adj_128.init = 16'hcece;
    LUT4 i1_4_lut_adj_129 (.A(\rx_data[5] ), .B(\rx_data[2] ), .C(\rx_data[1] ), 
         .D(\rx_data[0] ), .Z(n47)) /* synthesis lut_function=(!(A+!(B (C (D)+!C !(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(65[3] 99[10])
    defparam i1_4_lut_adj_129.init = 16'h5014;
    LUT4 i1_3_lut_adj_130 (.A(\rx_data[0] ), .B(\rx_data[2] ), .C(\rx_data[1] ), 
         .Z(n9)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(72[3:8])
    defparam i1_3_lut_adj_130.init = 16'hfbfb;
    FD1S3AY o_reset_34_rep_833 (.D(o_reset_N_624), .CK(dac_clk_p_c), .Q(n30028)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=30, LSE_LLINE=93, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(53[9] 54[46])
    defparam o_reset_34_rep_833.GSR = "DISABLED";
    LUT4 i1_4_lut_4_lut (.A(\rx_data[5] ), .B(\rx_data[2] ), .C(\rx_data[1] ), 
         .D(\rx_data[0] ), .Z(n50_adj_3039)) /* synthesis lut_function=(!((B (C (D))+!B !(C+(D)))+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(65[3] 99[10])
    defparam i1_4_lut_4_lut.init = 16'h2aa8;
    LUT4 i1_2_lut_rep_780 (.A(\rx_data[5] ), .B(\rx_data[3] ), .Z(n27445)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_780.init = 16'heeee;
    LUT4 i1_3_lut_rep_579_4_lut (.A(\rx_data[5] ), .B(\rx_data[3] ), .C(\rx_data[4] ), 
         .D(\rx_data[6] ), .Z(n27244)) /* synthesis lut_function=(A+(B+!(C (D)))) */ ;
    defparam i1_3_lut_rep_579_4_lut.init = 16'hefff;
    LUT4 i_stb_I_0_2_lut_3_lut (.A(n9), .B(n27244), .C(rx_stb), .Z(o_reset_N_624)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(54[23:45])
    defparam i_stb_I_0_2_lut_3_lut.init = 16'h1010;
    LUT4 i18056_3_lut_4_lut (.A(n27447), .B(n50_adj_3039), .C(\rx_data[6] ), 
         .D(\rx_data[4] ), .Z(n20272)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(65[3] 99[10])
    defparam i18056_3_lut_4_lut.init = 16'hffe0;
    LUT4 i82_3_lut_4_lut (.A(n27447), .B(n50_adj_3039), .C(\rx_data[4] ), 
         .D(n47), .Z(n52)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(65[3] 99[10])
    defparam i82_3_lut_4_lut.init = 16'hfe0e;
    LUT4 rx_data_0__bdd_3_lut_25499 (.A(\rx_data[0] ), .B(\rx_data[6] ), 
         .C(\rx_data[4] ), .Z(n27982)) /* synthesis lut_function=(!(A (B+!(C))+!A ((C)+!B))) */ ;
    defparam rx_data_0__bdd_3_lut_25499.init = 16'h2424;
    LUT4 rx_data_0__bdd_4_lut_26220 (.A(\rx_data[0] ), .B(\rx_data[1] ), 
         .C(\rx_data[6] ), .D(\rx_data[4] ), .Z(n27983)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (((D)+!C)+!B))) */ ;
    defparam rx_data_0__bdd_4_lut_26220.init = 16'h0840;
    LUT4 i1_2_lut_3_lut (.A(\rx_data[5] ), .B(\rx_data[3] ), .C(\rx_data[4] ), 
         .Z(n20978)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_3_lut.init = 16'hfefe;
    LUT4 rx_data_0__bdd_3_lut_26787 (.A(\rx_data[0] ), .B(\rx_data[1] ), 
         .C(\rx_data[4] ), .Z(n27986)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam rx_data_0__bdd_3_lut_26787.init = 16'h8080;
    LUT4 i1_4_lut_4_lut_adj_131 (.A(\rx_data[1] ), .B(\rx_data[2] ), .C(n20988), 
         .D(n20702), .Z(n20826)) /* synthesis lut_function=((B (C (D))+!B (D))+!A) */ ;
    defparam i1_4_lut_4_lut_adj_131.init = 16'hf755;
    FD1S3AX o_dh_bits_i4 (.D(o_dh_bits_4__N_595[4]), .CK(dac_clk_p_c), .Q(dec_bits[4])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=30, LSE_LLINE=93, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(60[9] 100[5])
    defparam o_dh_bits_i4.GSR = "DISABLED";
    LUT4 n27984_bdd_4_lut (.A(n27984), .B(\rx_data[3] ), .C(n27986), .D(\rx_data[5] ), 
         .Z(n29910)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A ((D)+!C))) */ ;
    defparam n27984_bdd_4_lut.init = 16'h22f0;
    LUT4 i1_3_lut_4_lut_3_lut (.A(\rx_data[1] ), .B(\rx_data[2] ), .C(\rx_data[0] ), 
         .Z(n4)) /* synthesis lut_function=(!(A ((C)+!B))) */ ;
    defparam i1_3_lut_4_lut_3_lut.init = 16'h5d5d;
    LUT4 i1_3_lut_rep_782 (.A(\rx_data[1] ), .B(\rx_data[2] ), .C(\rx_data[0] ), 
         .Z(n27447)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_3_lut_rep_782.init = 16'h1010;
    LUT4 i1_2_lut_rep_783 (.A(\rx_data[2] ), .B(\rx_data[1] ), .Z(n27448)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(65[3] 99[10])
    defparam i1_2_lut_rep_783.init = 16'heeee;
    FD1S3AX o_dh_bits_i3 (.D(o_dh_bits_4__N_595[3]), .CK(dac_clk_p_c), .Q(dec_bits_c[3])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=30, LSE_LLINE=93, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(60[9] 100[5])
    defparam o_dh_bits_i3.GSR = "DISABLED";
    FD1S3AX o_dh_bits_i2 (.D(o_dh_bits_4__N_595[2]), .CK(dac_clk_p_c), .Q(dec_bits_c[2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=30, LSE_LLINE=93, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(60[9] 100[5])
    defparam o_dh_bits_i2.GSR = "DISABLED";
    FD1S3AX o_dh_bits_i1 (.D(o_dh_bits_4__N_595[1]), .CK(dac_clk_p_c), .Q(\dec_bits[1] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=30, LSE_LLINE=93, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(60[9] 100[5])
    defparam o_dh_bits_i1.GSR = "DISABLED";
    FD1S3AY o_reset_34_rep_832 (.D(o_reset_N_624), .CK(dac_clk_p_c), .Q(n30027)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=30, LSE_LLINE=93, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(53[9] 54[46])
    defparam o_reset_34_rep_832.GSR = "DISABLED";
    LUT4 i1_2_lut_3_lut_4_lut (.A(\rx_data[2] ), .B(\rx_data[1] ), .C(n20095), 
         .D(\rx_data[3] ), .Z(n20097)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(65[3] 99[10])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h10f0;
    LUT4 i_byte_6__I_0_38_i9_2_lut_rep_580_3_lut (.A(\rx_data[2] ), .B(\rx_data[1] ), 
         .C(\rx_data[0] ), .Z(n27245)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(65[3] 99[10])
    defparam i_byte_6__I_0_38_i9_2_lut_rep_580_3_lut.init = 16'hefef;
    LUT4 n26375_bdd_2_lut_3_lut_4_lut (.A(n26373), .B(\rx_data[4] ), .C(\rx_data[3] ), 
         .D(\rx_data[6] ), .Z(n26376)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;
    defparam n26375_bdd_2_lut_3_lut_4_lut.init = 16'hfeff;
    LUT4 rx_data_0__bdd_4_lut_26788 (.A(\rx_data[0] ), .B(\rx_data[4] ), 
         .C(\rx_data[1] ), .D(\rx_data[2] ), .Z(n28999)) /* synthesis lut_function=(!(A (B (C)+!B !(C+(D)))+!A !((C (D)+!C !(D))+!B))) */ ;
    defparam rx_data_0__bdd_4_lut_26788.init = 16'h7b3d;
    LUT4 n29002_bdd_2_lut (.A(n29909), .B(\rx_data[3] ), .Z(o_dh_bits_4__N_595[3])) /* synthesis lut_function=(A+(B)) */ ;
    defparam n29002_bdd_2_lut.init = 16'heeee;
    LUT4 rx_data_0__bdd_4_lut_24716 (.A(\rx_data[0] ), .B(\rx_data[5] ), 
         .C(\rx_data[1] ), .D(\rx_data[2] ), .Z(n26373)) /* synthesis lut_function=(A (B (C)+!B (C+(D)))+!A (((D)+!C)+!B)) */ ;
    defparam rx_data_0__bdd_4_lut_24716.init = 16'hf7b5;
    LUT4 i17953_2_lut_3_lut_4_lut (.A(\rx_data[2] ), .B(\rx_data[1] ), .C(\rx_data[5] ), 
         .D(\rx_data[3] ), .Z(n20160)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(65[3] 99[10])
    defparam i17953_2_lut_3_lut_4_lut.init = 16'h10f0;
    LUT4 i23156_4_lut (.A(n27244), .B(n41), .C(n20832), .D(n4), .Z(o_dh_bits_4__N_595[4])) /* synthesis lut_function=(!(A (B (C))+!A (B (C (D))))) */ ;
    defparam i23156_4_lut.init = 16'h3f7f;
    LUT4 i1_4_lut_adj_132 (.A(n27135), .B(\rx_data[6] ), .C(n27245), .D(n20978), 
         .Z(n20832)) /* synthesis lut_function=(A ((C+(D))+!B)) */ ;
    defparam i1_4_lut_adj_132.init = 16'haaa2;
    LUT4 i1_4_lut_adj_133 (.A(n20850), .B(n20160), .C(n35), .D(\rx_data[6] ), 
         .Z(o_dh_bits_4__N_595[2])) /* synthesis lut_function=(A+(B (C (D))+!B (C+!(D)))) */ ;
    defparam i1_4_lut_adj_133.init = 16'hfabb;
    LUT4 i1_4_lut_adj_134 (.A(n20272), .B(n49), .C(n20974), .D(n42), 
         .Z(n20850)) /* synthesis lut_function=((B+(C (D)))+!A) */ ;
    defparam i1_4_lut_adj_134.init = 16'hfddd;
    LUT4 i1_4_lut_adj_135 (.A(\rx_data[2] ), .B(n20702), .C(\rx_data[1] ), 
         .D(n33), .Z(n49)) /* synthesis lut_function=(!((B (C+!(D)))+!A)) */ ;
    defparam i1_4_lut_adj_135.init = 16'h2a22;
    LUT4 i23159_4_lut (.A(n26376), .B(n41), .C(n35_adj_3040), .D(n20826), 
         .Z(o_dh_bits_4__N_595[1])) /* synthesis lut_function=(((C+!(D))+!B)+!A) */ ;
    defparam i23159_4_lut.init = 16'hf7ff;
    LUT4 i1_4_lut_adj_136 (.A(n27244), .B(n21300), .C(n9), .D(\rx_data[2] ), 
         .Z(n35_adj_3040)) /* synthesis lut_function=(!(A+(B (C (D))+!B (C)))) */ ;
    defparam i1_4_lut_adj_136.init = 16'h0545;
    LUT4 i1_4_lut_adj_137 (.A(\rx_data[5] ), .B(\rx_data[6] ), .C(n20982), 
         .D(\rx_data[4] ), .Z(n20988)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;
    defparam i1_4_lut_adj_137.init = 16'hfff7;
    LUT4 i1_2_lut_adj_138 (.A(\rx_data[0] ), .B(\rx_data[3] ), .Z(n20982)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_138.init = 16'heeee;
    LUT4 n28999_bdd_4_lut_4_lut (.A(\rx_data[4] ), .B(\rx_data[5] ), .C(\rx_data[6] ), 
         .D(n28999), .Z(n29909)) /* synthesis lut_function=(A (B (C)+!B ((D)+!C))+!A (B+((D)+!C))) */ ;
    defparam n28999_bdd_4_lut_4_lut.init = 16'hf7c7;
    LUT4 i_byte_6__I_0_57_i13_2_lut_rep_470_4_lut (.A(\rx_data[6] ), .B(\rx_data[4] ), 
         .C(n27445), .D(n9), .Z(n27135)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(93[3:8])
    defparam i_byte_6__I_0_57_i13_2_lut_rep_470_4_lut.init = 16'hfff7;
    LUT4 i1_3_lut_4_lut (.A(\rx_data[0] ), .B(n27448), .C(\rx_data[3] ), 
         .D(n20702), .Z(n50)) /* synthesis lut_function=(!((B+!(C+!(D)))+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(69[3:8])
    defparam i1_3_lut_4_lut.init = 16'h2022;
    LUT4 i1_2_lut_3_lut_adj_139 (.A(dec_stb), .B(dec_bits[4]), .C(cmd_loaded), 
         .Z(o_pck_stb_N_764)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(60[9] 100[5])
    defparam i1_2_lut_3_lut_adj_139.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_140 (.A(dec_stb), .B(dec_bits[4]), .C(n30027), 
         .Z(dac_clk_p_c_enable_222)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(60[9] 100[5])
    defparam i1_2_lut_3_lut_adj_140.init = 16'hf8f8;
    LUT4 i2_3_lut_4_lut (.A(dec_stb), .B(dec_bits[4]), .C(dec_bits_c[2]), 
         .D(dec_bits_c[3]), .Z(cmd_loaded_N_767)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(60[9] 100[5])
    defparam i2_3_lut_4_lut.init = 16'h0008;
    LUT4 i1_3_lut_4_lut_adj_141 (.A(\rx_data[5] ), .B(\rx_data[4] ), .C(\rx_data[0] ), 
         .D(n20974), .Z(n33)) /* synthesis lut_function=(A (D)+!A (B ((D)+!C)+!B (D))) */ ;
    defparam i1_3_lut_4_lut_adj_141.init = 16'hff04;
    LUT4 i66_3_lut_3_lut (.A(\rx_data[2] ), .B(\rx_data[1] ), .C(\rx_data[0] ), 
         .Z(n42)) /* synthesis lut_function=(!(A (C)+!A !(B (C)))) */ ;
    defparam i66_3_lut_3_lut.init = 16'h4a4a;
    LUT4 rx_data_4__bdd_3_lut_4_lut (.A(\rx_data[6] ), .B(\rx_data[5] ), 
         .C(\rx_data[3] ), .D(\rx_data[4] ), .Z(n20974)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam rx_data_4__bdd_3_lut_4_lut.init = 16'h0008;
    LUT4 i83_4_lut_4_lut (.A(\rx_data[3] ), .B(n52), .C(\rx_data[6] ), 
         .D(n20097), .Z(n41)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(58[24:46])
    defparam i83_4_lut_4_lut.init = 16'h4f40;
    LUT4 i1_2_lut_rep_647 (.A(n30027), .B(dec_stb), .Z(dac_clk_p_c_enable_405)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(53[9] 54[46])
    defparam i1_2_lut_rep_647.init = 16'heeee;
    LUT4 i7017_2_lut_3_lut (.A(n30027), .B(dec_stb), .C(dec_bits[4]), 
         .Z(dac_clk_p_c_enable_374)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(53[9] 54[46])
    defparam i7017_2_lut_3_lut.init = 16'he0e0;
    PFUMX i25497 (.BLUT(n27983), .ALUT(n27982), .C0(\rx_data[2] ), .Z(n27984));
    
endmodule
//
// Verilog Description of module hbnewline
//

module hbnewline (dac_clk_p_c, n30028, w_reset, hx_stb, tx_busy, nl_busy, 
            \w_gx_char[2] , \w_gx_char[0] , \w_gx_char[4] , n30027, 
            \w_gx_char[3] , \w_gx_char[5] , \w_gx_char[1] , \w_gx_char[6] , 
            n11763, n27281, \lcl_data[1] , \lcl_data_7__N_510[0] , zero_baud_counter, 
            dac_clk_p_c_enable_346, \lcl_data[4] , \lcl_data_7__N_510[3] , 
            \lcl_data[7] , \lcl_data_7__N_510[6] , \lcl_data[6] , \lcl_data_7__N_510[5] , 
            \lcl_data[5] , \lcl_data_7__N_510[4] , \lcl_data[3] , \lcl_data_7__N_510[2] , 
            \lcl_data[2] , \lcl_data_7__N_510[1] , o_busy_N_535, \state[0] , 
            n18134) /* synthesis syn_module_defined=1 */ ;
    input dac_clk_p_c;
    input n30028;
    input w_reset;
    input hx_stb;
    input tx_busy;
    output nl_busy;
    input \w_gx_char[2] ;
    input \w_gx_char[0] ;
    input \w_gx_char[4] ;
    input n30027;
    input \w_gx_char[3] ;
    input \w_gx_char[5] ;
    input \w_gx_char[1] ;
    input \w_gx_char[6] ;
    input n11763;
    output n27281;
    input \lcl_data[1] ;
    output \lcl_data_7__N_510[0] ;
    input zero_baud_counter;
    output dac_clk_p_c_enable_346;
    input \lcl_data[4] ;
    output \lcl_data_7__N_510[3] ;
    input \lcl_data[7] ;
    output \lcl_data_7__N_510[6] ;
    input \lcl_data[6] ;
    output \lcl_data_7__N_510[5] ;
    input \lcl_data[5] ;
    output \lcl_data_7__N_510[4] ;
    input \lcl_data[3] ;
    output \lcl_data_7__N_510[2] ;
    input \lcl_data[2] ;
    output \lcl_data_7__N_510[1] ;
    input o_busy_N_535;
    input \state[0] ;
    output n18134;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[49:58])
    
    wire tx_stb, o_nl_stb_N_1314, last_cr, last_cr_N_1322;
    wire [7:0]tx_data;   // d:/documents/git_local/fm_modulator/rtl/top.v(69[12:19])
    
    wire dac_clk_p_c_enable_225;
    wire [6:0]o_nl_byte_6__N_1301;
    wire [6:0]o_nl_byte_6__N_1294;
    
    wire cr_state, cr_state_N_1330, loaded, n27115, n27555, n27556, 
        n25095, n25094;
    wire [6:0]n32;
    
    wire n27234;
    
    FD1S3IX o_nl_stb_46 (.D(o_nl_stb_N_1314), .CK(dac_clk_p_c), .CD(n30028), 
            .Q(tx_stb)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=12, LSE_RCOL=40, LSE_LLINE=138, LSE_RLINE=139 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam o_nl_stb_46.GSR = "DISABLED";
    FD1S3JX last_cr_45 (.D(last_cr_N_1322), .CK(dac_clk_p_c), .PD(n30028), 
            .Q(last_cr)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=12, LSE_RCOL=40, LSE_LLINE=138, LSE_RLINE=139 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam last_cr_45.GSR = "DISABLED";
    FD1P3JX o_nl_byte_i2 (.D(o_nl_byte_6__N_1301[1]), .SP(dac_clk_p_c_enable_225), 
            .PD(w_reset), .CK(dac_clk_p_c), .Q(tx_data[1])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=12, LSE_RCOL=40, LSE_LLINE=138, LSE_RLINE=139 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam o_nl_byte_i2.GSR = "DISABLED";
    FD1P3JX o_nl_byte_i3 (.D(o_nl_byte_6__N_1301[2]), .SP(dac_clk_p_c_enable_225), 
            .PD(w_reset), .CK(dac_clk_p_c), .Q(tx_data[2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=12, LSE_RCOL=40, LSE_LLINE=138, LSE_RLINE=139 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam o_nl_byte_i3.GSR = "DISABLED";
    FD1P3AY o_nl_byte_i4 (.D(o_nl_byte_6__N_1294[3]), .SP(dac_clk_p_c_enable_225), 
            .CK(dac_clk_p_c), .Q(tx_data[3])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=12, LSE_RCOL=40, LSE_LLINE=138, LSE_RLINE=139 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam o_nl_byte_i4.GSR = "DISABLED";
    FD1P3JX o_nl_byte_i5 (.D(o_nl_byte_6__N_1301[4]), .SP(dac_clk_p_c_enable_225), 
            .PD(w_reset), .CK(dac_clk_p_c), .Q(tx_data[4])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=12, LSE_RCOL=40, LSE_LLINE=138, LSE_RLINE=139 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam o_nl_byte_i5.GSR = "DISABLED";
    FD1P3JX o_nl_byte_i6 (.D(o_nl_byte_6__N_1301[5]), .SP(dac_clk_p_c_enable_225), 
            .PD(w_reset), .CK(dac_clk_p_c), .Q(tx_data[5])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=12, LSE_RCOL=40, LSE_LLINE=138, LSE_RLINE=139 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam o_nl_byte_i6.GSR = "DISABLED";
    FD1P3JX o_nl_byte_i7 (.D(o_nl_byte_6__N_1301[6]), .SP(dac_clk_p_c_enable_225), 
            .PD(w_reset), .CK(dac_clk_p_c), .Q(tx_data[6])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=12, LSE_RCOL=40, LSE_LLINE=138, LSE_RLINE=139 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam o_nl_byte_i7.GSR = "DISABLED";
    FD1P3IX cr_state_44 (.D(cr_state_N_1330), .SP(dac_clk_p_c_enable_225), 
            .CD(w_reset), .CK(dac_clk_p_c), .Q(cr_state)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=12, LSE_RCOL=40, LSE_LLINE=138, LSE_RLINE=139 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam cr_state_44.GSR = "DISABLED";
    FD1P3IX loaded_47 (.D(n27115), .SP(dac_clk_p_c_enable_225), .CD(n30028), 
            .CK(dac_clk_p_c), .Q(loaded)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=12, LSE_RCOL=40, LSE_LLINE=138, LSE_RLINE=139 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam loaded_47.GSR = "DISABLED";
    FD1P3JX o_nl_byte_i1 (.D(o_nl_byte_6__N_1301[0]), .SP(dac_clk_p_c_enable_225), 
            .PD(n30028), .CK(dac_clk_p_c), .Q(tx_data[0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=12, LSE_RCOL=40, LSE_LLINE=138, LSE_RLINE=139 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam o_nl_byte_i1.GSR = "DISABLED";
    PFUMX i25208 (.BLUT(n27555), .ALUT(n27556), .C0(last_cr), .Z(last_cr_N_1322));
    LUT4 tx_stb_bdd_3_lut (.A(hx_stb), .B(last_cr), .C(cr_state), .Z(n25095)) /* synthesis lut_function=(A (B+!(C))+!A ((C)+!B)) */ ;
    defparam tx_stb_bdd_3_lut.init = 16'hdbdb;
    LUT4 tx_stb_bdd_2_lut (.A(tx_stb), .B(hx_stb), .Z(n25094)) /* synthesis lut_function=(A+(B)) */ ;
    defparam tx_stb_bdd_2_lut.init = 16'heeee;
    LUT4 i21484_4_lut (.A(cr_state), .B(tx_stb), .C(tx_busy), .D(loaded), 
         .Z(nl_busy)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(123[21] 124[30])
    defparam i21484_4_lut.init = 16'hca0a;
    LUT4 i1_2_lut (.A(last_cr), .B(cr_state), .Z(n32[4])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam i1_2_lut.init = 16'h2222;
    LUT4 i1_3_lut_4_lut (.A(last_cr), .B(n27234), .C(cr_state), .D(\w_gx_char[2] ), 
         .Z(o_nl_byte_6__N_1301[2])) /* synthesis lut_function=(A (B (D)+!B !(C))+!A ((D)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(97[12] 120[6])
    defparam i1_3_lut_4_lut.init = 16'hdf13;
    LUT4 i1_3_lut_4_lut_adj_120 (.A(last_cr), .B(n27234), .C(cr_state), 
         .D(\w_gx_char[0] ), .Z(o_nl_byte_6__N_1301[0])) /* synthesis lut_function=(A (B (D)+!B !(C))+!A ((D)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(97[12] 120[6])
    defparam i1_3_lut_4_lut_adj_120.init = 16'hdf13;
    LUT4 i_stb_I_0_2_lut_rep_569 (.A(hx_stb), .B(nl_busy), .Z(n27234)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(90[16:37])
    defparam i_stb_I_0_2_lut_rep_569.init = 16'h2222;
    LUT4 mux_24_i5_3_lut_4_lut (.A(hx_stb), .B(nl_busy), .C(\w_gx_char[4] ), 
         .D(n32[4]), .Z(o_nl_byte_6__N_1301[4])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(90[16:37])
    defparam mux_24_i5_3_lut_4_lut.init = 16'hfd20;
    LUT4 i1_3_lut_4_lut_adj_121 (.A(hx_stb), .B(nl_busy), .C(n30027), 
         .D(\w_gx_char[3] ), .Z(o_nl_byte_6__N_1294[3])) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(90[16:37])
    defparam i1_3_lut_4_lut_adj_121.init = 16'hfffd;
    LUT4 i1_3_lut_4_lut_adj_122 (.A(hx_stb), .B(nl_busy), .C(n30027), 
         .D(tx_busy), .Z(dac_clk_p_c_enable_225)) /* synthesis lut_function=(A ((C+!(D))+!B)+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(90[16:37])
    defparam i1_3_lut_4_lut_adj_122.init = 16'hf2ff;
    LUT4 i11343_3_lut_rep_450_4_lut (.A(hx_stb), .B(nl_busy), .C(cr_state), 
         .D(last_cr), .Z(n27115)) /* synthesis lut_function=(A ((C (D))+!B)+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(90[16:37])
    defparam i11343_3_lut_rep_450_4_lut.init = 16'hf222;
    LUT4 i11029_3_lut_4_lut (.A(hx_stb), .B(nl_busy), .C(\w_gx_char[5] ), 
         .D(n32[4]), .Z(o_nl_byte_6__N_1301[5])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(90[16:37])
    defparam i11029_3_lut_4_lut.init = 16'hfd20;
    LUT4 i11032_3_lut_4_lut (.A(hx_stb), .B(nl_busy), .C(\w_gx_char[1] ), 
         .D(last_cr), .Z(o_nl_byte_6__N_1301[1])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(90[16:37])
    defparam i11032_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_24_i7_3_lut_4_lut (.A(hx_stb), .B(nl_busy), .C(\w_gx_char[6] ), 
         .D(n32[4]), .Z(o_nl_byte_6__N_1301[6])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(90[16:37])
    defparam mux_24_i7_3_lut_4_lut.init = 16'hfd20;
    LUT4 cr_state_I_41_3_lut_4_lut (.A(hx_stb), .B(nl_busy), .C(n11763), 
         .D(last_cr), .Z(cr_state_N_1330)) /* synthesis lut_function=(!(A (B (D)+!B (C))+!A (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(90[16:37])
    defparam cr_state_I_41_3_lut_4_lut.init = 16'h02df;
    LUT4 i1_2_lut_rep_616 (.A(tx_stb), .B(tx_busy), .Z(n27281)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam i1_2_lut_rep_616.init = 16'h2222;
    LUT4 lcl_data_7__I_0_i1_3_lut_4_lut (.A(tx_stb), .B(tx_busy), .C(tx_data[0]), 
         .D(\lcl_data[1] ), .Z(\lcl_data_7__N_510[0] )) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam lcl_data_7__I_0_i1_3_lut_4_lut.init = 16'hfd20;
    LUT4 i611_2_lut_3_lut (.A(tx_stb), .B(tx_busy), .C(zero_baud_counter), 
         .Z(dac_clk_p_c_enable_346)) /* synthesis lut_function=(A ((C)+!B)+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam i611_2_lut_3_lut.init = 16'hf2f2;
    LUT4 lcl_data_7__I_0_i4_3_lut_4_lut (.A(tx_stb), .B(tx_busy), .C(tx_data[3]), 
         .D(\lcl_data[4] ), .Z(\lcl_data_7__N_510[3] )) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam lcl_data_7__I_0_i4_3_lut_4_lut.init = 16'hfd20;
    LUT4 lcl_data_7__I_0_i7_3_lut_4_lut (.A(tx_stb), .B(tx_busy), .C(tx_data[6]), 
         .D(\lcl_data[7] ), .Z(\lcl_data_7__N_510[6] )) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam lcl_data_7__I_0_i7_3_lut_4_lut.init = 16'hfd20;
    LUT4 lcl_data_7__I_0_i6_3_lut_4_lut (.A(tx_stb), .B(tx_busy), .C(tx_data[5]), 
         .D(\lcl_data[6] ), .Z(\lcl_data_7__N_510[5] )) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam lcl_data_7__I_0_i6_3_lut_4_lut.init = 16'hfd20;
    LUT4 lcl_data_7__I_0_i5_3_lut_4_lut (.A(tx_stb), .B(tx_busy), .C(tx_data[4]), 
         .D(\lcl_data[5] ), .Z(\lcl_data_7__N_510[4] )) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam lcl_data_7__I_0_i5_3_lut_4_lut.init = 16'hfd20;
    LUT4 lcl_data_7__I_0_i3_3_lut_4_lut (.A(tx_stb), .B(tx_busy), .C(tx_data[2]), 
         .D(\lcl_data[3] ), .Z(\lcl_data_7__N_510[2] )) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam lcl_data_7__I_0_i3_3_lut_4_lut.init = 16'hfd20;
    LUT4 lcl_data_7__I_0_i2_3_lut_4_lut (.A(tx_stb), .B(tx_busy), .C(tx_data[1]), 
         .D(\lcl_data[2] ), .Z(\lcl_data_7__N_510[1] )) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam lcl_data_7__I_0_i2_3_lut_4_lut.init = 16'hfd20;
    LUT4 state_596_mux_6_i1_3_lut_4_lut (.A(tx_stb), .B(tx_busy), .C(o_busy_N_535), 
         .D(\state[0] ), .Z(n18134)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam state_596_mux_6_i1_3_lut_4_lut.init = 16'hd0df;
    LUT4 last_cr_I_39_4_lut_then_3_lut (.A(n11763), .B(hx_stb), .C(nl_busy), 
         .Z(n27556)) /* synthesis lut_function=(((C)+!B)+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(97[12] 120[6])
    defparam last_cr_I_39_4_lut_then_3_lut.init = 16'hf7f7;
    LUT4 last_cr_I_39_4_lut_else_3_lut (.A(n11763), .B(tx_busy), .C(hx_stb), 
         .D(nl_busy), .Z(n27555)) /* synthesis lut_function=(!(A (B+(C))+!A (B ((D)+!C)+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(97[12] 120[6])
    defparam last_cr_I_39_4_lut_else_3_lut.init = 16'h0353;
    PFUMX i23464 (.BLUT(n25095), .ALUT(n25094), .C0(tx_busy), .Z(o_nl_stb_N_1314));
    
endmodule
//
// Verilog Description of module hbints
//

module hbints (int_word, dac_clk_p_c, dac_clk_p_c_enable_442, n12767, 
            ow_word, n30027, n27315, n27249, int_stb, ow_stb, n30028) /* synthesis syn_module_defined=1 */ ;
    output [33:0]int_word;
    input dac_clk_p_c;
    input dac_clk_p_c_enable_442;
    input n12767;
    input [33:0]ow_word;
    input n30027;
    output n27315;
    input n27249;
    output int_stb;
    input ow_stb;
    input n30028;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[49:58])
    
    wire dac_clk_p_c_enable_437, loaded, dac_clk_p_c_enable_434;
    
    FD1P3IX o_int_word_i9 (.D(ow_word[9]), .SP(dac_clk_p_c_enable_442), 
            .CD(n12767), .CK(dac_clk_p_c), .Q(int_word[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i9.GSR = "DISABLED";
    FD1P3JX o_int_word_i33 (.D(ow_word[33]), .SP(dac_clk_p_c_enable_442), 
            .PD(n12767), .CK(dac_clk_p_c), .Q(int_word[33])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i33.GSR = "DISABLED";
    FD1P3JX o_int_word_i32 (.D(ow_word[32]), .SP(dac_clk_p_c_enable_442), 
            .PD(n12767), .CK(dac_clk_p_c), .Q(int_word[32])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i32.GSR = "DISABLED";
    LUT4 i1_2_lut_3_lut_4_lut (.A(n30027), .B(n27315), .C(n27249), .D(int_stb), 
         .Z(dac_clk_p_c_enable_437)) /* synthesis lut_function=(A+(B+!(C+!(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'hefee;
    LUT4 i1_3_lut_4_lut (.A(n30027), .B(n27315), .C(loaded), .D(n27249), 
         .Z(dac_clk_p_c_enable_434)) /* synthesis lut_function=(A+(B+!(C (D)))) */ ;
    defparam i1_3_lut_4_lut.init = 16'hefff;
    FD1P3IX o_int_word_i31 (.D(ow_word[31]), .SP(dac_clk_p_c_enable_442), 
            .CD(n12767), .CK(dac_clk_p_c), .Q(int_word[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i31.GSR = "DISABLED";
    FD1P3IX o_int_word_i8 (.D(ow_word[8]), .SP(dac_clk_p_c_enable_442), 
            .CD(n12767), .CK(dac_clk_p_c), .Q(int_word[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i8.GSR = "DISABLED";
    FD1P3JX o_int_word_i30 (.D(ow_word[30]), .SP(dac_clk_p_c_enable_442), 
            .PD(n12767), .CK(dac_clk_p_c), .Q(int_word[30])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i30.GSR = "DISABLED";
    FD1P3IX o_int_word_i29 (.D(ow_word[29]), .SP(dac_clk_p_c_enable_442), 
            .CD(n12767), .CK(dac_clk_p_c), .Q(int_word[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i29.GSR = "DISABLED";
    FD1P3IX o_int_word_i28 (.D(ow_word[28]), .SP(dac_clk_p_c_enable_442), 
            .CD(n12767), .CK(dac_clk_p_c), .Q(int_word[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i28.GSR = "DISABLED";
    FD1P3IX o_int_word_i27 (.D(ow_word[27]), .SP(dac_clk_p_c_enable_442), 
            .CD(n12767), .CK(dac_clk_p_c), .Q(int_word[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i27.GSR = "DISABLED";
    FD1P3IX o_int_word_i7 (.D(ow_word[7]), .SP(dac_clk_p_c_enable_442), 
            .CD(n12767), .CK(dac_clk_p_c), .Q(int_word[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i7.GSR = "DISABLED";
    FD1P3IX o_int_word_i26 (.D(ow_word[26]), .SP(dac_clk_p_c_enable_442), 
            .CD(n12767), .CK(dac_clk_p_c), .Q(int_word[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i26.GSR = "DISABLED";
    FD1P3IX o_int_word_i6 (.D(ow_word[6]), .SP(dac_clk_p_c_enable_442), 
            .CD(n12767), .CK(dac_clk_p_c), .Q(int_word[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i6.GSR = "DISABLED";
    FD1P3IX o_int_word_i25 (.D(ow_word[25]), .SP(dac_clk_p_c_enable_442), 
            .CD(n12767), .CK(dac_clk_p_c), .Q(int_word[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i25.GSR = "DISABLED";
    FD1P3IX o_int_word_i5 (.D(ow_word[5]), .SP(dac_clk_p_c_enable_442), 
            .CD(n12767), .CK(dac_clk_p_c), .Q(int_word[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i5.GSR = "DISABLED";
    FD1P3IX o_int_word_i24 (.D(ow_word[24]), .SP(dac_clk_p_c_enable_442), 
            .CD(n12767), .CK(dac_clk_p_c), .Q(int_word[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i24.GSR = "DISABLED";
    LUT4 i_stb_I_0_3_lut_rep_650 (.A(ow_stb), .B(int_stb), .C(loaded), 
         .Z(n27315)) /* synthesis lut_function=(!((B (C))+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(93[12:34])
    defparam i_stb_I_0_3_lut_rep_650.init = 16'h2a2a;
    FD1P3IX o_int_word_i4 (.D(ow_word[4]), .SP(dac_clk_p_c_enable_442), 
            .CD(n12767), .CK(dac_clk_p_c), .Q(int_word[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i4.GSR = "DISABLED";
    FD1P3IX o_int_word_i3 (.D(ow_word[3]), .SP(dac_clk_p_c_enable_442), 
            .CD(n12767), .CK(dac_clk_p_c), .Q(int_word[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i3.GSR = "DISABLED";
    FD1P3IX o_int_word_i23 (.D(ow_word[23]), .SP(dac_clk_p_c_enable_442), 
            .CD(n12767), .CK(dac_clk_p_c), .Q(int_word[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i23.GSR = "DISABLED";
    FD1P3IX o_int_word_i2 (.D(ow_word[2]), .SP(dac_clk_p_c_enable_442), 
            .CD(n12767), .CK(dac_clk_p_c), .Q(int_word[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i2.GSR = "DISABLED";
    FD1P3IX o_int_word_i22 (.D(ow_word[22]), .SP(dac_clk_p_c_enable_442), 
            .CD(n12767), .CK(dac_clk_p_c), .Q(int_word[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i22.GSR = "DISABLED";
    FD1P3IX o_int_word_i1 (.D(ow_word[1]), .SP(dac_clk_p_c_enable_442), 
            .CD(n12767), .CK(dac_clk_p_c), .Q(int_word[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i1.GSR = "DISABLED";
    FD1P3IX o_int_word_i0 (.D(ow_word[0]), .SP(dac_clk_p_c_enable_442), 
            .CD(n12767), .CK(dac_clk_p_c), .Q(int_word[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i0.GSR = "DISABLED";
    FD1P3IX o_int_word_i21 (.D(ow_word[21]), .SP(dac_clk_p_c_enable_442), 
            .CD(n12767), .CK(dac_clk_p_c), .Q(int_word[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i21.GSR = "DISABLED";
    FD1P3IX o_int_word_i20 (.D(ow_word[20]), .SP(dac_clk_p_c_enable_442), 
            .CD(n12767), .CK(dac_clk_p_c), .Q(int_word[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i20.GSR = "DISABLED";
    FD1P3IX o_int_word_i19 (.D(ow_word[19]), .SP(dac_clk_p_c_enable_442), 
            .CD(n12767), .CK(dac_clk_p_c), .Q(int_word[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i19.GSR = "DISABLED";
    FD1P3IX o_int_word_i18 (.D(ow_word[18]), .SP(dac_clk_p_c_enable_442), 
            .CD(n12767), .CK(dac_clk_p_c), .Q(int_word[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i18.GSR = "DISABLED";
    FD1P3IX o_int_word_i17 (.D(ow_word[17]), .SP(dac_clk_p_c_enable_442), 
            .CD(n12767), .CK(dac_clk_p_c), .Q(int_word[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i17.GSR = "DISABLED";
    FD1P3IX o_int_word_i16 (.D(ow_word[16]), .SP(dac_clk_p_c_enable_442), 
            .CD(n12767), .CK(dac_clk_p_c), .Q(int_word[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i16.GSR = "DISABLED";
    FD1P3IX o_int_word_i15 (.D(ow_word[15]), .SP(dac_clk_p_c_enable_442), 
            .CD(n12767), .CK(dac_clk_p_c), .Q(int_word[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i15.GSR = "DISABLED";
    FD1P3IX o_int_stb_58 (.D(n27315), .SP(dac_clk_p_c_enable_434), .CD(n30028), 
            .CK(dac_clk_p_c), .Q(int_stb)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(90[9] 98[22])
    defparam o_int_stb_58.GSR = "DISABLED";
    FD1P3IX o_int_word_i14 (.D(ow_word[14]), .SP(dac_clk_p_c_enable_442), 
            .CD(n12767), .CK(dac_clk_p_c), .Q(int_word[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i14.GSR = "DISABLED";
    FD1P3IX o_int_word_i13 (.D(ow_word[13]), .SP(dac_clk_p_c_enable_442), 
            .CD(n12767), .CK(dac_clk_p_c), .Q(int_word[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i13.GSR = "DISABLED";
    FD1P3IX loaded_57 (.D(n27315), .SP(dac_clk_p_c_enable_437), .CD(n30028), 
            .CK(dac_clk_p_c), .Q(loaded)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(81[9] 87[19])
    defparam loaded_57.GSR = "DISABLED";
    FD1P3IX o_int_word_i12 (.D(ow_word[12]), .SP(dac_clk_p_c_enable_442), 
            .CD(n12767), .CK(dac_clk_p_c), .Q(int_word[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i12.GSR = "DISABLED";
    FD1P3IX o_int_word_i11 (.D(ow_word[11]), .SP(dac_clk_p_c_enable_442), 
            .CD(n12767), .CK(dac_clk_p_c), .Q(int_word[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i11.GSR = "DISABLED";
    FD1P3IX o_int_word_i10 (.D(ow_word[10]), .SP(dac_clk_p_c_enable_442), 
            .CD(n12767), .CK(dac_clk_p_c), .Q(int_word[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i10.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module hbidle
//

module hbidle (idl_word, dac_clk_p_c, int_word, idl_stb, w_reset, 
            hb_busy, int_stb, n27249, n30027, n27315, dac_clk_p_c_enable_442, 
            n12767) /* synthesis syn_module_defined=1 */ ;
    output [33:0]idl_word;
    input dac_clk_p_c;
    input [33:0]int_word;
    output idl_stb;
    input w_reset;
    input hb_busy;
    input int_stb;
    output n27249;
    input n30027;
    input n27315;
    output dac_clk_p_c_enable_442;
    output n12767;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[49:58])
    
    wire dac_clk_p_c_enable_429, n12797, dac_clk_p_c_enable_221, n27137;
    
    FD1P3IX o_idl_word_i11 (.D(int_word[11]), .SP(dac_clk_p_c_enable_429), 
            .CD(n12797), .CK(dac_clk_p_c), .Q(idl_word[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i11.GSR = "DISABLED";
    FD1P3IX o_idl_word_i10 (.D(int_word[10]), .SP(dac_clk_p_c_enable_429), 
            .CD(n12797), .CK(dac_clk_p_c), .Q(idl_word[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i10.GSR = "DISABLED";
    FD1P3IX o_idl_word_i9 (.D(int_word[9]), .SP(dac_clk_p_c_enable_429), 
            .CD(n12797), .CK(dac_clk_p_c), .Q(idl_word[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i9.GSR = "DISABLED";
    FD1P3IX o_idl_word_i8 (.D(int_word[8]), .SP(dac_clk_p_c_enable_429), 
            .CD(n12797), .CK(dac_clk_p_c), .Q(idl_word[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i8.GSR = "DISABLED";
    FD1P3IX o_idl_word_i7 (.D(int_word[7]), .SP(dac_clk_p_c_enable_429), 
            .CD(n12797), .CK(dac_clk_p_c), .Q(idl_word[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i7.GSR = "DISABLED";
    FD1P3IX o_idl_word_i6 (.D(int_word[6]), .SP(dac_clk_p_c_enable_429), 
            .CD(n12797), .CK(dac_clk_p_c), .Q(idl_word[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i6.GSR = "DISABLED";
    FD1P3IX o_idl_word_i5 (.D(int_word[5]), .SP(dac_clk_p_c_enable_429), 
            .CD(n12797), .CK(dac_clk_p_c), .Q(idl_word[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i5.GSR = "DISABLED";
    FD1P3IX o_idl_word_i4 (.D(int_word[4]), .SP(dac_clk_p_c_enable_429), 
            .CD(n12797), .CK(dac_clk_p_c), .Q(idl_word[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i4.GSR = "DISABLED";
    FD1P3IX o_idl_stb_28 (.D(n27137), .SP(dac_clk_p_c_enable_221), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(idl_stb)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(80[9] 88[22])
    defparam o_idl_stb_28.GSR = "DISABLED";
    FD1P3JX o_idl_word_i33 (.D(int_word[33]), .SP(dac_clk_p_c_enable_429), 
            .PD(n12797), .CK(dac_clk_p_c), .Q(idl_word[33])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i33.GSR = "DISABLED";
    FD1P3JX o_idl_word_i32 (.D(int_word[32]), .SP(dac_clk_p_c_enable_429), 
            .PD(n12797), .CK(dac_clk_p_c), .Q(idl_word[32])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i32.GSR = "DISABLED";
    FD1P3IX o_idl_word_i31 (.D(int_word[31]), .SP(dac_clk_p_c_enable_429), 
            .CD(n12797), .CK(dac_clk_p_c), .Q(idl_word[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i31.GSR = "DISABLED";
    FD1P3JX o_idl_word_i30 (.D(int_word[30]), .SP(dac_clk_p_c_enable_429), 
            .PD(n12797), .CK(dac_clk_p_c), .Q(idl_word[30])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i30.GSR = "DISABLED";
    FD1P3JX o_idl_word_i29 (.D(int_word[29]), .SP(dac_clk_p_c_enable_429), 
            .PD(n12797), .CK(dac_clk_p_c), .Q(idl_word[29])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i29.GSR = "DISABLED";
    FD1P3IX o_idl_word_i28 (.D(int_word[28]), .SP(dac_clk_p_c_enable_429), 
            .CD(n12797), .CK(dac_clk_p_c), .Q(idl_word[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i28.GSR = "DISABLED";
    FD1P3IX o_idl_word_i27 (.D(int_word[27]), .SP(dac_clk_p_c_enable_429), 
            .CD(n12797), .CK(dac_clk_p_c), .Q(idl_word[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i27.GSR = "DISABLED";
    FD1P3IX o_idl_word_i3 (.D(int_word[3]), .SP(dac_clk_p_c_enable_429), 
            .CD(n12797), .CK(dac_clk_p_c), .Q(idl_word[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i3.GSR = "DISABLED";
    LUT4 i23069_2_lut (.A(hb_busy), .B(int_stb), .Z(n12797)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i23069_2_lut.init = 16'h1111;
    FD1P3IX o_idl_word_i2 (.D(int_word[2]), .SP(dac_clk_p_c_enable_429), 
            .CD(n12797), .CK(dac_clk_p_c), .Q(idl_word[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i2.GSR = "DISABLED";
    FD1P3IX o_idl_word_i1 (.D(int_word[1]), .SP(dac_clk_p_c_enable_429), 
            .CD(n12797), .CK(dac_clk_p_c), .Q(idl_word[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i1.GSR = "DISABLED";
    FD1P3IX o_idl_word_i0 (.D(int_word[0]), .SP(dac_clk_p_c_enable_429), 
            .CD(n12797), .CK(dac_clk_p_c), .Q(idl_word[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i0.GSR = "DISABLED";
    FD1P3IX o_idl_word_i14 (.D(int_word[14]), .SP(dac_clk_p_c_enable_429), 
            .CD(n12797), .CK(dac_clk_p_c), .Q(idl_word[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i14.GSR = "DISABLED";
    FD1P3IX o_idl_word_i26 (.D(int_word[26]), .SP(dac_clk_p_c_enable_429), 
            .CD(n12797), .CK(dac_clk_p_c), .Q(idl_word[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i26.GSR = "DISABLED";
    FD1P3IX o_idl_word_i25 (.D(int_word[25]), .SP(dac_clk_p_c_enable_429), 
            .CD(n12797), .CK(dac_clk_p_c), .Q(idl_word[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i25.GSR = "DISABLED";
    FD1P3IX o_idl_word_i24 (.D(int_word[24]), .SP(dac_clk_p_c_enable_429), 
            .CD(n12797), .CK(dac_clk_p_c), .Q(idl_word[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i24.GSR = "DISABLED";
    FD1P3IX o_idl_word_i23 (.D(int_word[23]), .SP(dac_clk_p_c_enable_429), 
            .CD(n12797), .CK(dac_clk_p_c), .Q(idl_word[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i23.GSR = "DISABLED";
    FD1P3IX o_idl_word_i22 (.D(int_word[22]), .SP(dac_clk_p_c_enable_429), 
            .CD(n12797), .CK(dac_clk_p_c), .Q(idl_word[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i22.GSR = "DISABLED";
    FD1P3IX o_idl_word_i21 (.D(int_word[21]), .SP(dac_clk_p_c_enable_429), 
            .CD(n12797), .CK(dac_clk_p_c), .Q(idl_word[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i21.GSR = "DISABLED";
    FD1P3IX o_idl_word_i20 (.D(int_word[20]), .SP(dac_clk_p_c_enable_429), 
            .CD(n12797), .CK(dac_clk_p_c), .Q(idl_word[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i20.GSR = "DISABLED";
    FD1P3IX o_idl_word_i19 (.D(int_word[19]), .SP(dac_clk_p_c_enable_429), 
            .CD(n12797), .CK(dac_clk_p_c), .Q(idl_word[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i19.GSR = "DISABLED";
    FD1P3IX o_idl_word_i18 (.D(int_word[18]), .SP(dac_clk_p_c_enable_429), 
            .CD(n12797), .CK(dac_clk_p_c), .Q(idl_word[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i18.GSR = "DISABLED";
    FD1P3IX o_idl_word_i17 (.D(int_word[17]), .SP(dac_clk_p_c_enable_429), 
            .CD(n12797), .CK(dac_clk_p_c), .Q(idl_word[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i17.GSR = "DISABLED";
    FD1P3IX o_idl_word_i16 (.D(int_word[16]), .SP(dac_clk_p_c_enable_429), 
            .CD(n12797), .CK(dac_clk_p_c), .Q(idl_word[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i16.GSR = "DISABLED";
    FD1P3IX o_idl_word_i15 (.D(int_word[15]), .SP(dac_clk_p_c_enable_429), 
            .CD(n12797), .CK(dac_clk_p_c), .Q(idl_word[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i15.GSR = "DISABLED";
    FD1P3IX o_idl_word_i13 (.D(int_word[13]), .SP(dac_clk_p_c_enable_429), 
            .CD(n12797), .CK(dac_clk_p_c), .Q(idl_word[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i13.GSR = "DISABLED";
    FD1P3IX o_idl_word_i12 (.D(int_word[12]), .SP(dac_clk_p_c_enable_429), 
            .CD(n12797), .CK(dac_clk_p_c), .Q(idl_word[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i12.GSR = "DISABLED";
    LUT4 o_idl_stb_I_0_30_2_lut_rep_584 (.A(idl_stb), .B(hb_busy), .Z(n27249)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(97[22:43])
    defparam o_idl_stb_I_0_30_2_lut_rep_584.init = 16'h8888;
    LUT4 o_int_stb_I_0_66_2_lut_rep_472_3_lut (.A(idl_stb), .B(hb_busy), 
         .C(int_stb), .Z(n27137)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(97[22:43])
    defparam o_int_stb_I_0_66_2_lut_rep_472_3_lut.init = 16'h7070;
    LUT4 i1_3_lut_4_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(n30027), .D(int_stb), 
         .Z(dac_clk_p_c_enable_221)) /* synthesis lut_function=(A ((C)+!B)+!A ((C+(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(97[22:43])
    defparam i1_3_lut_4_lut_4_lut.init = 16'hf7f3;
    LUT4 i1_2_lut_3_lut_3_lut (.A(idl_stb), .B(hb_busy), .C(int_stb), 
         .Z(dac_clk_p_c_enable_429)) /* synthesis lut_function=(!(A (B)+!A !((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(97[22:43])
    defparam i1_2_lut_3_lut_3_lut.init = 16'h7373;
    LUT4 i1_2_lut_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(n27315), .D(int_stb), 
         .Z(dac_clk_p_c_enable_442)) /* synthesis lut_function=(((C+!(D))+!B)+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(97[22:43])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hf7ff;
    LUT4 i23034_2_lut_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(n27315), 
         .D(int_stb), .Z(n12767)) /* synthesis lut_function=(!(A (B (C+(D))+!B (C))+!A (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(97[22:43])
    defparam i23034_2_lut_3_lut_4_lut.init = 16'h070f;
    
endmodule
//
// Verilog Description of module \rxuartlite(CLOCKS_PER_BAUD=10000) 
//

module \rxuartlite(CLOCKS_PER_BAUD=10000)  (\rx_data[0] , dac_clk_p_c, rx_stb, 
            i_wbu_uart_rx_c, chg_counter, dac_clk_p_c_enable_199, chg_counter_23__N_405, 
            GND_net, \rx_data[6] , \rx_data[5] , \rx_data[4] , \rx_data[3] , 
            \rx_data[2] , \rx_data[1] ) /* synthesis syn_module_defined=1 */ ;
    output \rx_data[0] ;
    input dac_clk_p_c;
    output rx_stb;
    input i_wbu_uart_rx_c;
    output [23:0]chg_counter;
    input dac_clk_p_c_enable_199;
    output chg_counter_23__N_405;
    input GND_net;
    output \rx_data[6] ;
    output \rx_data[5] ;
    output \rx_data[4] ;
    output \rx_data[3] ;
    output \rx_data[2] ;
    output \rx_data[1] ;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[49:58])
    
    wire o_data_7__N_417;
    wire [7:0]data_reg;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(142[12:20])
    
    wire qq_uart, q_uart, ck_uart;
    wire [3:0]state;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(75[13:18])
    
    wire dac_clk_p_c_enable_372;
    wire [3:0]state_3__N_321;
    
    wire half_baud_time, half_baud_time_N_456;
    wire [23:0]baud_counter;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(78[17:29])
    
    wire dac_clk_p_c_enable_440, baud_counter_23__N_444;
    wire [23:0]baud_counter_23__N_420;
    wire [23:0]n8;
    
    wire zero_baud_counter, dac_clk_p_c_enable_146, n14846, n27199, 
        n17946, n17947, n17945, n17944, n17943, n17942, n17941, 
        n17940, n17939, n17938;
    wire [23:0]n254;
    
    wire n17937, n17936, n17935, n17934, n17933, n17932, n17931, 
        n17885, n17884, n17930, n17883, n17882, n17929, n17928, 
        n17927, zero_baud_counter_N_453, n11702, state_3__N_414, n27133, 
        n20817, n21436, n21598, n21596, n21582, n21580, n21528, 
        n21574, n21532, n164, n27496, n17881, n171, n27495, n17880, 
        n17879, n17878, n27319, half_baud_time_N_457, n17877, data_reg_7__N_415, 
        n17876, n26513, n26512, n17875, dac_clk_p_c_enable_368;
    wire [3:0]n174;
    
    wire n17874, n17950, n17949, n17948;
    
    FD1P3AX o_data__i1 (.D(data_reg[0]), .SP(o_data_7__N_417), .CK(dac_clk_p_c), 
            .Q(\rx_data[0] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(155[9] 161[18])
    defparam o_data__i1.GSR = "DISABLED";
    FD1S3AY qq_uart_70 (.D(q_uart), .CK(dac_clk_p_c), .Q(qq_uart)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(90[9] 91[66])
    defparam qq_uart_70.GSR = "DISABLED";
    FD1S3AY ck_uart_71 (.D(qq_uart), .CK(dac_clk_p_c), .Q(ck_uart)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(90[9] 91[66])
    defparam ck_uart_71.GSR = "DISABLED";
    FD1P3AY state_i0 (.D(state_3__N_321[0]), .SP(dac_clk_p_c_enable_372), 
            .CK(dac_clk_p_c), .Q(state[0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(116[9] 134[5])
    defparam state_i0.GSR = "DISABLED";
    FD1S3AX half_baud_time_73 (.D(half_baud_time_N_456), .CK(dac_clk_p_c), 
            .Q(half_baud_time)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(111[9] 112[70])
    defparam half_baud_time_73.GSR = "DISABLED";
    FD1S3AX o_wr_76 (.D(o_data_7__N_417), .CK(dac_clk_p_c), .Q(rx_stb)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(155[9] 161[18])
    defparam o_wr_76.GSR = "DISABLED";
    FD1S3AY q_uart_69 (.D(i_wbu_uart_rx_c), .CK(dac_clk_p_c), .Q(q_uart)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(90[9] 91[66])
    defparam q_uart_69.GSR = "DISABLED";
    FD1P3JX baud_counter_i1 (.D(baud_counter_23__N_420[1]), .SP(dac_clk_p_c_enable_440), 
            .PD(baud_counter_23__N_444), .CK(dac_clk_p_c), .Q(baud_counter[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i1.GSR = "DISABLED";
    FD1P3IX chg_counter__i0 (.D(n8[0]), .SP(dac_clk_p_c_enable_199), .CD(chg_counter_23__N_405), 
            .CK(dac_clk_p_c), .Q(chg_counter[0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i0.GSR = "DISABLED";
    FD1P3AY zero_baud_counter_79 (.D(n14846), .SP(dac_clk_p_c_enable_146), 
            .CK(dac_clk_p_c), .Q(zero_baud_counter)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(187[9] 195[29])
    defparam zero_baud_counter_79.GSR = "DISABLED";
    LUT4 i1_3_lut_4_lut (.A(state[0]), .B(n27199), .C(ck_uart), .D(zero_baud_counter), 
         .Z(o_data_7__N_417)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(144[27:48])
    defparam i1_3_lut_4_lut.init = 16'h1000;
    CCU2D sub_435_add_2_18 (.A0(chg_counter[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17946), .COUT(n17947));
    defparam sub_435_add_2_18.INIT0 = 16'h5555;
    defparam sub_435_add_2_18.INIT1 = 16'h5555;
    defparam sub_435_add_2_18.INJECT1_0 = "NO";
    defparam sub_435_add_2_18.INJECT1_1 = "NO";
    CCU2D sub_435_add_2_16 (.A0(chg_counter[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17945), .COUT(n17946));
    defparam sub_435_add_2_16.INIT0 = 16'h5555;
    defparam sub_435_add_2_16.INIT1 = 16'h5555;
    defparam sub_435_add_2_16.INJECT1_0 = "NO";
    defparam sub_435_add_2_16.INJECT1_1 = "NO";
    FD1P3IX chg_counter__i23 (.D(n8[23]), .SP(dac_clk_p_c_enable_199), .CD(chg_counter_23__N_405), 
            .CK(dac_clk_p_c), .Q(chg_counter[23])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i23.GSR = "DISABLED";
    CCU2D sub_435_add_2_14 (.A0(chg_counter[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17944), .COUT(n17945));
    defparam sub_435_add_2_14.INIT0 = 16'h5aaa;
    defparam sub_435_add_2_14.INIT1 = 16'h5555;
    defparam sub_435_add_2_14.INJECT1_0 = "NO";
    defparam sub_435_add_2_14.INJECT1_1 = "NO";
    FD1P3JX baud_counter_i2 (.D(baud_counter_23__N_420[2]), .SP(dac_clk_p_c_enable_440), 
            .PD(baud_counter_23__N_444), .CK(dac_clk_p_c), .Q(baud_counter[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i2.GSR = "DISABLED";
    FD1P3JX baud_counter_i3 (.D(baud_counter_23__N_420[3]), .SP(dac_clk_p_c_enable_440), 
            .PD(baud_counter_23__N_444), .CK(dac_clk_p_c), .Q(baud_counter[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i3.GSR = "DISABLED";
    FD1P3JX baud_counter_i8 (.D(baud_counter_23__N_420[8]), .SP(dac_clk_p_c_enable_440), 
            .PD(baud_counter_23__N_444), .CK(dac_clk_p_c), .Q(baud_counter[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i8.GSR = "DISABLED";
    CCU2D sub_435_add_2_12 (.A0(chg_counter[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17943), .COUT(n17944));
    defparam sub_435_add_2_12.INIT0 = 16'h5555;
    defparam sub_435_add_2_12.INIT1 = 16'h5555;
    defparam sub_435_add_2_12.INJECT1_0 = "NO";
    defparam sub_435_add_2_12.INJECT1_1 = "NO";
    FD1P3IX chg_counter__i22 (.D(n8[22]), .SP(dac_clk_p_c_enable_199), .CD(chg_counter_23__N_405), 
            .CK(dac_clk_p_c), .Q(chg_counter[22])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i22.GSR = "DISABLED";
    FD1P3IX chg_counter__i21 (.D(n8[21]), .SP(dac_clk_p_c_enable_199), .CD(chg_counter_23__N_405), 
            .CK(dac_clk_p_c), .Q(chg_counter[21])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i21.GSR = "DISABLED";
    FD1P3IX chg_counter__i20 (.D(n8[20]), .SP(dac_clk_p_c_enable_199), .CD(chg_counter_23__N_405), 
            .CK(dac_clk_p_c), .Q(chg_counter[20])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i20.GSR = "DISABLED";
    FD1P3IX chg_counter__i19 (.D(n8[19]), .SP(dac_clk_p_c_enable_199), .CD(chg_counter_23__N_405), 
            .CK(dac_clk_p_c), .Q(chg_counter[19])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i19.GSR = "DISABLED";
    FD1P3IX chg_counter__i18 (.D(n8[18]), .SP(dac_clk_p_c_enable_199), .CD(chg_counter_23__N_405), 
            .CK(dac_clk_p_c), .Q(chg_counter[18])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i18.GSR = "DISABLED";
    FD1P3IX chg_counter__i17 (.D(n8[17]), .SP(dac_clk_p_c_enable_199), .CD(chg_counter_23__N_405), 
            .CK(dac_clk_p_c), .Q(chg_counter[17])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i17.GSR = "DISABLED";
    FD1P3IX chg_counter__i16 (.D(n8[16]), .SP(dac_clk_p_c_enable_199), .CD(chg_counter_23__N_405), 
            .CK(dac_clk_p_c), .Q(chg_counter[16])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i16.GSR = "DISABLED";
    FD1P3IX chg_counter__i15 (.D(n8[15]), .SP(dac_clk_p_c_enable_199), .CD(chg_counter_23__N_405), 
            .CK(dac_clk_p_c), .Q(chg_counter[15])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i15.GSR = "DISABLED";
    FD1P3IX chg_counter__i14 (.D(n8[14]), .SP(dac_clk_p_c_enable_199), .CD(chg_counter_23__N_405), 
            .CK(dac_clk_p_c), .Q(chg_counter[14])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i14.GSR = "DISABLED";
    FD1P3IX chg_counter__i13 (.D(n8[13]), .SP(dac_clk_p_c_enable_199), .CD(chg_counter_23__N_405), 
            .CK(dac_clk_p_c), .Q(chg_counter[13])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i13.GSR = "DISABLED";
    FD1P3IX chg_counter__i12 (.D(n8[12]), .SP(dac_clk_p_c_enable_199), .CD(chg_counter_23__N_405), 
            .CK(dac_clk_p_c), .Q(chg_counter[12])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i12.GSR = "DISABLED";
    FD1P3IX chg_counter__i11 (.D(n8[11]), .SP(dac_clk_p_c_enable_199), .CD(chg_counter_23__N_405), 
            .CK(dac_clk_p_c), .Q(chg_counter[11])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i11.GSR = "DISABLED";
    FD1P3IX chg_counter__i10 (.D(n8[10]), .SP(dac_clk_p_c_enable_199), .CD(chg_counter_23__N_405), 
            .CK(dac_clk_p_c), .Q(chg_counter[10])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i10.GSR = "DISABLED";
    FD1P3IX chg_counter__i9 (.D(n8[9]), .SP(dac_clk_p_c_enable_199), .CD(chg_counter_23__N_405), 
            .CK(dac_clk_p_c), .Q(chg_counter[9])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i9.GSR = "DISABLED";
    FD1P3IX chg_counter__i8 (.D(n8[8]), .SP(dac_clk_p_c_enable_199), .CD(chg_counter_23__N_405), 
            .CK(dac_clk_p_c), .Q(chg_counter[8])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i8.GSR = "DISABLED";
    FD1P3IX chg_counter__i7 (.D(n8[7]), .SP(dac_clk_p_c_enable_199), .CD(chg_counter_23__N_405), 
            .CK(dac_clk_p_c), .Q(chg_counter[7])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i7.GSR = "DISABLED";
    FD1P3IX chg_counter__i6 (.D(n8[6]), .SP(dac_clk_p_c_enable_199), .CD(chg_counter_23__N_405), 
            .CK(dac_clk_p_c), .Q(chg_counter[6])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i6.GSR = "DISABLED";
    FD1P3IX chg_counter__i5 (.D(n8[5]), .SP(dac_clk_p_c_enable_199), .CD(chg_counter_23__N_405), 
            .CK(dac_clk_p_c), .Q(chg_counter[5])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i5.GSR = "DISABLED";
    FD1P3IX chg_counter__i4 (.D(n8[4]), .SP(dac_clk_p_c_enable_199), .CD(chg_counter_23__N_405), 
            .CK(dac_clk_p_c), .Q(chg_counter[4])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i4.GSR = "DISABLED";
    FD1P3IX chg_counter__i3 (.D(n8[3]), .SP(dac_clk_p_c_enable_199), .CD(chg_counter_23__N_405), 
            .CK(dac_clk_p_c), .Q(chg_counter[3])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i3.GSR = "DISABLED";
    FD1P3IX chg_counter__i2 (.D(n8[2]), .SP(dac_clk_p_c_enable_199), .CD(chg_counter_23__N_405), 
            .CK(dac_clk_p_c), .Q(chg_counter[2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i2.GSR = "DISABLED";
    FD1P3IX chg_counter__i1 (.D(n8[1]), .SP(dac_clk_p_c_enable_199), .CD(chg_counter_23__N_405), 
            .CK(dac_clk_p_c), .Q(chg_counter[1])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i1.GSR = "DISABLED";
    FD1P3JX baud_counter_i9 (.D(baud_counter_23__N_420[9]), .SP(dac_clk_p_c_enable_440), 
            .PD(baud_counter_23__N_444), .CK(dac_clk_p_c), .Q(baud_counter[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i9.GSR = "DISABLED";
    FD1P3JX baud_counter_i10 (.D(baud_counter_23__N_420[10]), .SP(dac_clk_p_c_enable_440), 
            .PD(baud_counter_23__N_444), .CK(dac_clk_p_c), .Q(baud_counter[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i10.GSR = "DISABLED";
    FD1P3JX baud_counter_i13 (.D(baud_counter_23__N_420[13]), .SP(dac_clk_p_c_enable_440), 
            .PD(baud_counter_23__N_444), .CK(dac_clk_p_c), .Q(baud_counter[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i13.GSR = "DISABLED";
    CCU2D sub_435_add_2_10 (.A0(chg_counter[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17942), .COUT(n17943));
    defparam sub_435_add_2_10.INIT0 = 16'h5aaa;
    defparam sub_435_add_2_10.INIT1 = 16'h5aaa;
    defparam sub_435_add_2_10.INJECT1_0 = "NO";
    defparam sub_435_add_2_10.INJECT1_1 = "NO";
    CCU2D sub_435_add_2_8 (.A0(chg_counter[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17941), .COUT(n17942));
    defparam sub_435_add_2_8.INIT0 = 16'h5555;
    defparam sub_435_add_2_8.INIT1 = 16'h5aaa;
    defparam sub_435_add_2_8.INJECT1_0 = "NO";
    defparam sub_435_add_2_8.INJECT1_1 = "NO";
    CCU2D sub_435_add_2_6 (.A0(chg_counter[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17940), .COUT(n17941));
    defparam sub_435_add_2_6.INIT0 = 16'h5555;
    defparam sub_435_add_2_6.INIT1 = 16'h5555;
    defparam sub_435_add_2_6.INJECT1_0 = "NO";
    defparam sub_435_add_2_6.INJECT1_1 = "NO";
    CCU2D sub_435_add_2_4 (.A0(chg_counter[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17939), .COUT(n17940));
    defparam sub_435_add_2_4.INIT0 = 16'h5aaa;
    defparam sub_435_add_2_4.INIT1 = 16'h5555;
    defparam sub_435_add_2_4.INJECT1_0 = "NO";
    defparam sub_435_add_2_4.INJECT1_1 = "NO";
    CCU2D sub_435_add_2_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(chg_counter[1]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n17939));
    defparam sub_435_add_2_2.INIT0 = 16'h0000;
    defparam sub_435_add_2_2.INIT1 = 16'h5aaa;
    defparam sub_435_add_2_2.INJECT1_0 = "NO";
    defparam sub_435_add_2_2.INJECT1_1 = "NO";
    CCU2D sub_49_add_2_25 (.A0(baud_counter[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n17938), .S0(n254[23]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_25.INIT0 = 16'h5555;
    defparam sub_49_add_2_25.INIT1 = 16'h0000;
    defparam sub_49_add_2_25.INJECT1_0 = "NO";
    defparam sub_49_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_49_add_2_23 (.A0(baud_counter[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17937), .COUT(n17938), .S0(n254[21]), 
          .S1(n254[22]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_23.INIT0 = 16'h5555;
    defparam sub_49_add_2_23.INIT1 = 16'h5555;
    defparam sub_49_add_2_23.INJECT1_0 = "NO";
    defparam sub_49_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_49_add_2_21 (.A0(baud_counter[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17936), .COUT(n17937), .S0(n254[19]), 
          .S1(n254[20]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_21.INIT0 = 16'h5555;
    defparam sub_49_add_2_21.INIT1 = 16'h5555;
    defparam sub_49_add_2_21.INJECT1_0 = "NO";
    defparam sub_49_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_49_add_2_19 (.A0(baud_counter[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17935), .COUT(n17936), .S0(n254[17]), 
          .S1(n254[18]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_19.INIT0 = 16'h5555;
    defparam sub_49_add_2_19.INIT1 = 16'h5555;
    defparam sub_49_add_2_19.INJECT1_0 = "NO";
    defparam sub_49_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_49_add_2_17 (.A0(baud_counter[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17934), .COUT(n17935), .S0(n254[15]), 
          .S1(n254[16]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_17.INIT0 = 16'h5555;
    defparam sub_49_add_2_17.INIT1 = 16'h5555;
    defparam sub_49_add_2_17.INJECT1_0 = "NO";
    defparam sub_49_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_49_add_2_15 (.A0(baud_counter[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17933), .COUT(n17934), .S0(n254[13]), 
          .S1(n254[14]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_15.INIT0 = 16'h5555;
    defparam sub_49_add_2_15.INIT1 = 16'h5555;
    defparam sub_49_add_2_15.INJECT1_0 = "NO";
    defparam sub_49_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_49_add_2_13 (.A0(baud_counter[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17932), .COUT(n17933), .S0(n254[11]), 
          .S1(n254[12]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_13.INIT0 = 16'h5555;
    defparam sub_49_add_2_13.INIT1 = 16'h5555;
    defparam sub_49_add_2_13.INJECT1_0 = "NO";
    defparam sub_49_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_49_add_2_11 (.A0(baud_counter[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17931), .COUT(n17932), .S0(n254[9]), .S1(n254[10]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_11.INIT0 = 16'h5555;
    defparam sub_49_add_2_11.INIT1 = 16'h5555;
    defparam sub_49_add_2_11.INJECT1_0 = "NO";
    defparam sub_49_add_2_11.INJECT1_1 = "NO";
    CCU2D add_8_25 (.A0(chg_counter[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n17885), .S0(n8[23]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:36])
    defparam add_8_25.INIT0 = 16'h5aaa;
    defparam add_8_25.INIT1 = 16'h0000;
    defparam add_8_25.INJECT1_0 = "NO";
    defparam add_8_25.INJECT1_1 = "NO";
    CCU2D add_8_23 (.A0(chg_counter[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17884), .COUT(n17885), .S0(n8[21]), .S1(n8[22]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:36])
    defparam add_8_23.INIT0 = 16'h5aaa;
    defparam add_8_23.INIT1 = 16'h5aaa;
    defparam add_8_23.INJECT1_0 = "NO";
    defparam add_8_23.INJECT1_1 = "NO";
    CCU2D sub_49_add_2_9 (.A0(baud_counter[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17930), .COUT(n17931), .S0(n254[7]), .S1(n254[8]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_9.INIT0 = 16'h5555;
    defparam sub_49_add_2_9.INIT1 = 16'h5555;
    defparam sub_49_add_2_9.INJECT1_0 = "NO";
    defparam sub_49_add_2_9.INJECT1_1 = "NO";
    CCU2D add_8_21 (.A0(chg_counter[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17883), .COUT(n17884), .S0(n8[19]), .S1(n8[20]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:36])
    defparam add_8_21.INIT0 = 16'h5aaa;
    defparam add_8_21.INIT1 = 16'h5aaa;
    defparam add_8_21.INJECT1_0 = "NO";
    defparam add_8_21.INJECT1_1 = "NO";
    CCU2D add_8_19 (.A0(chg_counter[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17882), .COUT(n17883), .S0(n8[17]), .S1(n8[18]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:36])
    defparam add_8_19.INIT0 = 16'h5aaa;
    defparam add_8_19.INIT1 = 16'h5aaa;
    defparam add_8_19.INJECT1_0 = "NO";
    defparam add_8_19.INJECT1_1 = "NO";
    CCU2D sub_49_add_2_7 (.A0(baud_counter[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17929), .COUT(n17930), .S0(n254[5]), .S1(n254[6]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_7.INIT0 = 16'h5555;
    defparam sub_49_add_2_7.INIT1 = 16'h5555;
    defparam sub_49_add_2_7.INJECT1_0 = "NO";
    defparam sub_49_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_49_add_2_5 (.A0(baud_counter[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17928), .COUT(n17929), .S0(n254[3]), .S1(n254[4]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_5.INIT0 = 16'h5555;
    defparam sub_49_add_2_5.INIT1 = 16'h5555;
    defparam sub_49_add_2_5.INJECT1_0 = "NO";
    defparam sub_49_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_49_add_2_3 (.A0(baud_counter[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17927), .COUT(n17928), .S0(n254[1]), .S1(n254[2]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_3.INIT0 = 16'h5555;
    defparam sub_49_add_2_3.INIT1 = 16'h5555;
    defparam sub_49_add_2_3.INJECT1_0 = "NO";
    defparam sub_49_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_49_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(baud_counter[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n17927), .S1(n254[0]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_1.INIT0 = 16'hF000;
    defparam sub_49_add_2_1.INIT1 = 16'h5555;
    defparam sub_49_add_2_1.INJECT1_0 = "NO";
    defparam sub_49_add_2_1.INJECT1_1 = "NO";
    LUT4 i11830_3_lut_4_lut (.A(state[0]), .B(n27199), .C(zero_baud_counter_N_453), 
         .D(n254[1]), .Z(baud_counter_23__N_420[1])) /* synthesis lut_function=(A (B (C+(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(144[27:48])
    defparam i11830_3_lut_4_lut.init = 16'hddd0;
    LUT4 i1_2_lut_3_lut_4_lut (.A(state[0]), .B(n27199), .C(zero_baud_counter_N_453), 
         .D(baud_counter_23__N_444), .Z(n11702)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(144[27:48])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfff2;
    LUT4 i23030_3_lut_4_lut (.A(state[0]), .B(n27199), .C(baud_counter_23__N_444), 
         .D(zero_baud_counter_N_453), .Z(n14846)) /* synthesis lut_function=(!(A (B (C+(D))+!B (C))+!A (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(144[27:48])
    defparam i23030_3_lut_4_lut.init = 16'h020f;
    LUT4 i11829_3_lut_4_lut (.A(state[0]), .B(n27199), .C(zero_baud_counter_N_453), 
         .D(n254[2]), .Z(baud_counter_23__N_420[2])) /* synthesis lut_function=(A (B (C+(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(144[27:48])
    defparam i11829_3_lut_4_lut.init = 16'hddd0;
    LUT4 i11828_3_lut_4_lut (.A(state[0]), .B(n27199), .C(zero_baud_counter_N_453), 
         .D(n254[3]), .Z(baud_counter_23__N_420[3])) /* synthesis lut_function=(A (B (C+(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(144[27:48])
    defparam i11828_3_lut_4_lut.init = 16'hddd0;
    LUT4 i11827_3_lut_4_lut (.A(state[0]), .B(n27199), .C(zero_baud_counter_N_453), 
         .D(n254[8]), .Z(baud_counter_23__N_420[8])) /* synthesis lut_function=(A (B (C+(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(144[27:48])
    defparam i11827_3_lut_4_lut.init = 16'hddd0;
    LUT4 i11826_3_lut_4_lut (.A(state[0]), .B(n27199), .C(zero_baud_counter_N_453), 
         .D(n254[9]), .Z(baud_counter_23__N_420[9])) /* synthesis lut_function=(A (B (C+(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(144[27:48])
    defparam i11826_3_lut_4_lut.init = 16'hddd0;
    LUT4 i11825_3_lut_4_lut (.A(state[0]), .B(n27199), .C(zero_baud_counter_N_453), 
         .D(n254[10]), .Z(baud_counter_23__N_420[10])) /* synthesis lut_function=(A (B (C+(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(144[27:48])
    defparam i11825_3_lut_4_lut.init = 16'hddd0;
    LUT4 i11824_3_lut_4_lut (.A(state[0]), .B(n27199), .C(zero_baud_counter_N_453), 
         .D(n254[13]), .Z(baud_counter_23__N_420[13])) /* synthesis lut_function=(A (B (C+(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(144[27:48])
    defparam i11824_3_lut_4_lut.init = 16'hddd0;
    LUT4 i11314_3_lut_4_lut (.A(state[0]), .B(n27199), .C(zero_baud_counter_N_453), 
         .D(n254[0]), .Z(baud_counter_23__N_420[0])) /* synthesis lut_function=(A (B (C+(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(144[27:48])
    defparam i11314_3_lut_4_lut.init = 16'hddd0;
    LUT4 i1_3_lut (.A(ck_uart), .B(state_3__N_414), .C(half_baud_time), 
         .Z(baud_counter_23__N_444)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(171[6:57])
    defparam i1_3_lut.init = 16'h4040;
    LUT4 zero_baud_counter_I_0_2_lut (.A(zero_baud_counter), .B(state[3]), 
         .Z(zero_baud_counter_N_453)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(175[11:52])
    defparam zero_baud_counter_I_0_2_lut.init = 16'h2222;
    LUT4 qq_uart_I_0_2_lut (.A(qq_uart), .B(ck_uart), .Z(chg_counter_23__N_405)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(100[6:24])
    defparam qq_uart_I_0_2_lut.init = 16'h6666;
    LUT4 i1_4_lut (.A(zero_baud_counter_N_453), .B(n27133), .C(baud_counter_23__N_444), 
         .D(n20817), .Z(dac_clk_p_c_enable_146)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;
    defparam i1_4_lut.init = 16'hfffb;
    LUT4 i1_4_lut_adj_114 (.A(n21436), .B(n21598), .C(n21596), .D(n21582), 
         .Z(n20817)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_4_lut_adj_114.init = 16'h0002;
    LUT4 i1_4_lut_adj_115 (.A(baud_counter[3]), .B(baud_counter[2]), .C(baud_counter[16]), 
         .D(baud_counter[0]), .Z(n21436)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut_adj_115.init = 16'h0100;
    LUT4 i19318_4_lut (.A(baud_counter[23]), .B(n21580), .C(n21528), .D(baud_counter[11]), 
         .Z(n21598)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i19318_4_lut.init = 16'hfffe;
    LUT4 i19316_4_lut (.A(baud_counter[10]), .B(n21574), .C(n21532), .D(baud_counter[17]), 
         .Z(n21596)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i19316_4_lut.init = 16'hfffe;
    LUT4 i19302_4_lut (.A(baud_counter[22]), .B(baud_counter[8]), .C(baud_counter[15]), 
         .D(baud_counter[5]), .Z(n21582)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i19302_4_lut.init = 16'hfffe;
    LUT4 i19300_4_lut (.A(baud_counter[20]), .B(baud_counter[9]), .C(baud_counter[13]), 
         .D(baud_counter[19]), .Z(n21580)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i19300_4_lut.init = 16'hfffe;
    LUT4 i19248_2_lut (.A(baud_counter[7]), .B(baud_counter[4]), .Z(n21528)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i19248_2_lut.init = 16'heeee;
    LUT4 i19294_4_lut (.A(baud_counter[21]), .B(baud_counter[14]), .C(baud_counter[1]), 
         .D(baud_counter[18]), .Z(n21574)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i19294_4_lut.init = 16'hfffe;
    LUT4 i19252_2_lut (.A(baud_counter[6]), .B(baud_counter[12]), .Z(n21532)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i19252_2_lut.init = 16'heeee;
    LUT4 state_3__I_0_80_i4_4_lut_then_4_lut (.A(n164), .B(state[0]), .C(state[2]), 
         .D(state[1]), .Z(n27496)) /* synthesis lut_function=(!(A (B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(125[11] 134[5])
    defparam state_3__I_0_80_i4_4_lut_then_4_lut.init = 16'h7fff;
    CCU2D add_8_17 (.A0(chg_counter[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17881), .COUT(n17882), .S0(n8[15]), .S1(n8[16]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:36])
    defparam add_8_17.INIT0 = 16'h5aaa;
    defparam add_8_17.INIT1 = 16'h5aaa;
    defparam add_8_17.INJECT1_0 = "NO";
    defparam add_8_17.INJECT1_1 = "NO";
    LUT4 state_3__I_0_80_i4_4_lut_else_4_lut (.A(state[0]), .B(n171), .C(state[2]), 
         .D(state[1]), .Z(n27495)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(125[11] 134[5])
    defparam state_3__I_0_80_i4_4_lut_else_4_lut.init = 16'heccc;
    CCU2D add_8_15 (.A0(chg_counter[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17880), .COUT(n17881), .S0(n8[13]), .S1(n8[14]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:36])
    defparam add_8_15.INIT0 = 16'h5aaa;
    defparam add_8_15.INIT1 = 16'h5aaa;
    defparam add_8_15.INJECT1_0 = "NO";
    defparam add_8_15.INJECT1_1 = "NO";
    CCU2D add_8_13 (.A0(chg_counter[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17879), .COUT(n17880), .S0(n8[11]), .S1(n8[12]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:36])
    defparam add_8_13.INIT0 = 16'h5aaa;
    defparam add_8_13.INIT1 = 16'h5aaa;
    defparam add_8_13.INJECT1_0 = "NO";
    defparam add_8_13.INJECT1_1 = "NO";
    CCU2D add_8_11 (.A0(chg_counter[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(chg_counter[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n17878), .COUT(n17879), .S0(n8[9]), .S1(n8[10]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:36])
    defparam add_8_11.INIT0 = 16'h5aaa;
    defparam add_8_11.INIT1 = 16'h5aaa;
    defparam add_8_11.INJECT1_0 = "NO";
    defparam add_8_11.INJECT1_1 = "NO";
    LUT4 i1_3_lut_4_lut_adj_116 (.A(state[0]), .B(n27319), .C(ck_uart), 
         .D(state[3]), .Z(n171)) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(144[27:48])
    defparam i1_3_lut_4_lut_adj_116.init = 16'he000;
    LUT4 i1_3_lut_adj_117 (.A(state_3__N_414), .B(n171), .C(zero_baud_counter), 
         .Z(dac_clk_p_c_enable_372)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_3_lut_adj_117.init = 16'hfefe;
    LUT4 i21_2_lut (.A(ck_uart), .B(half_baud_time), .Z(n164)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(121[7:35])
    defparam i21_2_lut.init = 16'h4444;
    LUT4 i1_4_lut_adj_118 (.A(state[0]), .B(state[2]), .C(state[3]), .D(state[1]), 
         .Z(state_3__N_414)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_118.init = 16'h8000;
    LUT4 ck_uart_N_447_I_0_2_lut (.A(ck_uart), .B(half_baud_time_N_457), 
         .Z(half_baud_time_N_456)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(112[21:69])
    defparam ck_uart_N_447_I_0_2_lut.init = 16'h4444;
    CCU2D add_8_9 (.A0(chg_counter[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(chg_counter[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n17877), .COUT(n17878), .S0(n8[7]), .S1(n8[8]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:36])
    defparam add_8_9.INIT0 = 16'h5aaa;
    defparam add_8_9.INIT1 = 16'h5aaa;
    defparam add_8_9.INJECT1_0 = "NO";
    defparam add_8_9.INJECT1_1 = "NO";
    LUT4 zero_baud_counter_I_0_82_2_lut_3_lut_4_lut (.A(state[3]), .B(n27319), 
         .C(zero_baud_counter), .D(state[0]), .Z(data_reg_7__N_415)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(144[27:48])
    defparam zero_baud_counter_I_0_82_2_lut_3_lut_4_lut.init = 16'hf0d0;
    CCU2D add_8_7 (.A0(chg_counter[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(chg_counter[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n17876), .COUT(n17877), .S0(n8[5]), .S1(n8[6]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:36])
    defparam add_8_7.INIT0 = 16'h5aaa;
    defparam add_8_7.INIT1 = 16'h5aaa;
    defparam add_8_7.INJECT1_0 = "NO";
    defparam add_8_7.INJECT1_1 = "NO";
    LUT4 state_3__N_414_bdd_4_lut (.A(state[0]), .B(state[3]), .C(n27319), 
         .D(ck_uart), .Z(n26513)) /* synthesis lut_function=(A (B)+!A (((D)+!C)+!B)) */ ;
    defparam state_3__N_414_bdd_4_lut.init = 16'hdd9d;
    LUT4 state_3__N_414_bdd_2_lut (.A(half_baud_time), .B(ck_uart), .Z(n26512)) /* synthesis lut_function=((B)+!A) */ ;
    defparam state_3__N_414_bdd_2_lut.init = 16'hdddd;
    CCU2D add_8_5 (.A0(chg_counter[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(chg_counter[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n17875), .COUT(n17876), .S0(n8[3]), .S1(n8[4]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:36])
    defparam add_8_5.INIT0 = 16'h5aaa;
    defparam add_8_5.INIT1 = 16'h5aaa;
    defparam add_8_5.INJECT1_0 = "NO";
    defparam add_8_5.INJECT1_1 = "NO";
    LUT4 i1_3_lut_4_lut_adj_119 (.A(baud_counter_23__N_444), .B(n27133), 
         .C(state[3]), .D(zero_baud_counter), .Z(dac_clk_p_c_enable_440)) /* synthesis lut_function=(A+!(B (C (D)))) */ ;
    defparam i1_3_lut_4_lut_adj_119.init = 16'hbfff;
    FD1P3IX baud_counter_i23 (.D(n254[23]), .SP(dac_clk_p_c_enable_368), 
            .CD(n11702), .CK(dac_clk_p_c), .Q(baud_counter[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i23.GSR = "DISABLED";
    LUT4 i9727_1_lut (.A(zero_baud_counter), .Z(dac_clk_p_c_enable_368)) /* synthesis lut_function=(!(A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(187[9] 195[29])
    defparam i9727_1_lut.init = 16'h5555;
    LUT4 state_3__I_0_80_i3_4_lut (.A(n164), .B(n174[2]), .C(state_3__N_414), 
         .D(n171), .Z(state_3__N_321[2])) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A !(B+(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(125[11] 134[5])
    defparam state_3__I_0_80_i3_4_lut.init = 16'h5f5c;
    LUT4 state_3__I_0_80_i2_4_lut (.A(n164), .B(n174[1]), .C(state_3__N_414), 
         .D(n171), .Z(state_3__N_321[1])) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A !(B+(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(125[11] 134[5])
    defparam state_3__I_0_80_i2_4_lut.init = 16'h5f5c;
    FD1P3IX baud_counter_i22 (.D(n254[22]), .SP(dac_clk_p_c_enable_368), 
            .CD(n11702), .CK(dac_clk_p_c), .Q(baud_counter[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i22.GSR = "DISABLED";
    FD1P3IX baud_counter_i21 (.D(n254[21]), .SP(dac_clk_p_c_enable_368), 
            .CD(n11702), .CK(dac_clk_p_c), .Q(baud_counter[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i21.GSR = "DISABLED";
    FD1P3IX baud_counter_i20 (.D(n254[20]), .SP(dac_clk_p_c_enable_368), 
            .CD(n11702), .CK(dac_clk_p_c), .Q(baud_counter[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i20.GSR = "DISABLED";
    FD1P3IX baud_counter_i19 (.D(n254[19]), .SP(dac_clk_p_c_enable_368), 
            .CD(n11702), .CK(dac_clk_p_c), .Q(baud_counter[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i19.GSR = "DISABLED";
    FD1P3IX baud_counter_i18 (.D(n254[18]), .SP(dac_clk_p_c_enable_368), 
            .CD(n11702), .CK(dac_clk_p_c), .Q(baud_counter[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i18.GSR = "DISABLED";
    FD1P3IX baud_counter_i17 (.D(n254[17]), .SP(dac_clk_p_c_enable_368), 
            .CD(n11702), .CK(dac_clk_p_c), .Q(baud_counter[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i17.GSR = "DISABLED";
    FD1P3IX baud_counter_i16 (.D(n254[16]), .SP(dac_clk_p_c_enable_368), 
            .CD(n11702), .CK(dac_clk_p_c), .Q(baud_counter[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i16.GSR = "DISABLED";
    FD1P3IX baud_counter_i15 (.D(n254[15]), .SP(dac_clk_p_c_enable_368), 
            .CD(n11702), .CK(dac_clk_p_c), .Q(baud_counter[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i15.GSR = "DISABLED";
    FD1P3IX baud_counter_i14 (.D(n254[14]), .SP(dac_clk_p_c_enable_368), 
            .CD(n11702), .CK(dac_clk_p_c), .Q(baud_counter[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i14.GSR = "DISABLED";
    FD1P3IX baud_counter_i12 (.D(n254[12]), .SP(dac_clk_p_c_enable_368), 
            .CD(n11702), .CK(dac_clk_p_c), .Q(baud_counter[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i12.GSR = "DISABLED";
    FD1P3IX baud_counter_i11 (.D(n254[11]), .SP(dac_clk_p_c_enable_368), 
            .CD(n11702), .CK(dac_clk_p_c), .Q(baud_counter[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i11.GSR = "DISABLED";
    FD1P3IX baud_counter_i7 (.D(n254[7]), .SP(dac_clk_p_c_enable_368), .CD(n11702), 
            .CK(dac_clk_p_c), .Q(baud_counter[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i7.GSR = "DISABLED";
    FD1P3IX baud_counter_i6 (.D(n254[6]), .SP(dac_clk_p_c_enable_368), .CD(n11702), 
            .CK(dac_clk_p_c), .Q(baud_counter[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i6.GSR = "DISABLED";
    FD1P3IX baud_counter_i5 (.D(n254[5]), .SP(dac_clk_p_c_enable_368), .CD(n11702), 
            .CK(dac_clk_p_c), .Q(baud_counter[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i5.GSR = "DISABLED";
    FD1P3IX baud_counter_i4 (.D(n254[4]), .SP(dac_clk_p_c_enable_368), .CD(n11702), 
            .CK(dac_clk_p_c), .Q(baud_counter[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i4.GSR = "DISABLED";
    LUT4 i822_2_lut_3_lut (.A(state[0]), .B(state[3]), .C(state[1]), .Z(n174[1])) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(133[13:25])
    defparam i822_2_lut_3_lut.init = 16'hd2d2;
    FD1P3AY state_i3 (.D(state_3__N_321[3]), .SP(dac_clk_p_c_enable_372), 
            .CK(dac_clk_p_c), .Q(state[3])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(116[9] 134[5])
    defparam state_i3.GSR = "DISABLED";
    LUT4 i829_2_lut_3_lut_4_lut (.A(state[0]), .B(state[3]), .C(state[2]), 
         .D(state[1]), .Z(n174[2])) /* synthesis lut_function=(A (B (C)+!B !(C (D)+!C !(D)))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(133[13:25])
    defparam i829_2_lut_3_lut_4_lut.init = 16'hd2f0;
    FD1P3AY state_i2 (.D(state_3__N_321[2]), .SP(dac_clk_p_c_enable_372), 
            .CK(dac_clk_p_c), .Q(state[2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(116[9] 134[5])
    defparam state_i2.GSR = "DISABLED";
    FD1P3AY state_i1 (.D(state_3__N_321[1]), .SP(dac_clk_p_c_enable_372), 
            .CK(dac_clk_p_c), .Q(state[1])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(116[9] 134[5])
    defparam state_i1.GSR = "DISABLED";
    CCU2D add_8_3 (.A0(chg_counter[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(chg_counter[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n17874), .COUT(n17875), .S0(n8[1]), .S1(n8[2]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:36])
    defparam add_8_3.INIT0 = 16'h5aaa;
    defparam add_8_3.INIT1 = 16'h5aaa;
    defparam add_8_3.INJECT1_0 = "NO";
    defparam add_8_3.INJECT1_1 = "NO";
    CCU2D add_8_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(chg_counter[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n17874), .S1(n8[0]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:36])
    defparam add_8_1.INIT0 = 16'hF000;
    defparam add_8_1.INIT1 = 16'h5555;
    defparam add_8_1.INJECT1_0 = "NO";
    defparam add_8_1.INJECT1_1 = "NO";
    PFUMX i24714 (.BLUT(n26513), .ALUT(n26512), .C0(state_3__N_414), .Z(state_3__N_321[0]));
    FD1P3AX o_data__i7 (.D(data_reg[6]), .SP(o_data_7__N_417), .CK(dac_clk_p_c), 
            .Q(\rx_data[6] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(155[9] 161[18])
    defparam o_data__i7.GSR = "DISABLED";
    FD1P3AX o_data__i6 (.D(data_reg[5]), .SP(o_data_7__N_417), .CK(dac_clk_p_c), 
            .Q(\rx_data[5] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(155[9] 161[18])
    defparam o_data__i6.GSR = "DISABLED";
    FD1P3AX o_data__i5 (.D(data_reg[4]), .SP(o_data_7__N_417), .CK(dac_clk_p_c), 
            .Q(\rx_data[4] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(155[9] 161[18])
    defparam o_data__i5.GSR = "DISABLED";
    FD1P3AX o_data__i4 (.D(data_reg[3]), .SP(o_data_7__N_417), .CK(dac_clk_p_c), 
            .Q(\rx_data[3] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(155[9] 161[18])
    defparam o_data__i4.GSR = "DISABLED";
    FD1P3AX o_data__i3 (.D(data_reg[2]), .SP(o_data_7__N_417), .CK(dac_clk_p_c), 
            .Q(\rx_data[2] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(155[9] 161[18])
    defparam o_data__i3.GSR = "DISABLED";
    FD1P3AX o_data__i2 (.D(data_reg[1]), .SP(o_data_7__N_417), .CK(dac_clk_p_c), 
            .Q(\rx_data[1] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(155[9] 161[18])
    defparam o_data__i2.GSR = "DISABLED";
    PFUMX i25167 (.BLUT(n27495), .ALUT(n27496), .C0(state[3]), .Z(state_3__N_321[3]));
    FD1P3JX baud_counter_i0 (.D(baud_counter_23__N_420[0]), .SP(dac_clk_p_c_enable_440), 
            .PD(baud_counter_23__N_444), .CK(dac_clk_p_c), .Q(baud_counter[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i0.GSR = "DISABLED";
    CCU2D sub_435_add_2_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n17950), .S0(half_baud_time_N_457));
    defparam sub_435_add_2_cout.INIT0 = 16'h0000;
    defparam sub_435_add_2_cout.INIT1 = 16'h0000;
    defparam sub_435_add_2_cout.INJECT1_0 = "NO";
    defparam sub_435_add_2_cout.INJECT1_1 = "NO";
    LUT4 i6742_2_lut_rep_654 (.A(state[1]), .B(state[2]), .Z(n27319)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(129[7:26])
    defparam i6742_2_lut_rep_654.init = 16'heeee;
    LUT4 i1_2_lut_rep_534_3_lut (.A(state[1]), .B(state[2]), .C(state[3]), 
         .Z(n27199)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(129[7:26])
    defparam i1_2_lut_rep_534_3_lut.init = 16'hefef;
    LUT4 i1_2_lut_rep_468_3_lut_4_lut (.A(state[1]), .B(state[2]), .C(state[0]), 
         .D(state[3]), .Z(n27133)) /* synthesis lut_function=(A+(B+!(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(129[7:26])
    defparam i1_2_lut_rep_468_3_lut_4_lut.init = 16'hefff;
    CCU2D sub_435_add_2_24 (.A0(chg_counter[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17949), .COUT(n17950));
    defparam sub_435_add_2_24.INIT0 = 16'h5555;
    defparam sub_435_add_2_24.INIT1 = 16'h5555;
    defparam sub_435_add_2_24.INJECT1_0 = "NO";
    defparam sub_435_add_2_24.INJECT1_1 = "NO";
    CCU2D sub_435_add_2_22 (.A0(chg_counter[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17948), .COUT(n17949));
    defparam sub_435_add_2_22.INIT0 = 16'h5555;
    defparam sub_435_add_2_22.INIT1 = 16'h5555;
    defparam sub_435_add_2_22.INJECT1_0 = "NO";
    defparam sub_435_add_2_22.INJECT1_1 = "NO";
    CCU2D sub_435_add_2_20 (.A0(chg_counter[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17947), .COUT(n17948));
    defparam sub_435_add_2_20.INIT0 = 16'h5555;
    defparam sub_435_add_2_20.INIT1 = 16'h5555;
    defparam sub_435_add_2_20.INJECT1_0 = "NO";
    defparam sub_435_add_2_20.INJECT1_1 = "NO";
    FD1P3AX data_reg_i0_i7 (.D(qq_uart), .SP(data_reg_7__N_415), .CK(dac_clk_p_c), 
            .Q(data_reg[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(143[9] 145[42])
    defparam data_reg_i0_i7.GSR = "DISABLED";
    FD1P3AX data_reg_i0_i6 (.D(data_reg[7]), .SP(data_reg_7__N_415), .CK(dac_clk_p_c), 
            .Q(data_reg[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(143[9] 145[42])
    defparam data_reg_i0_i6.GSR = "DISABLED";
    FD1P3AX data_reg_i0_i5 (.D(data_reg[6]), .SP(data_reg_7__N_415), .CK(dac_clk_p_c), 
            .Q(data_reg[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(143[9] 145[42])
    defparam data_reg_i0_i5.GSR = "DISABLED";
    FD1P3AX data_reg_i0_i4 (.D(data_reg[5]), .SP(data_reg_7__N_415), .CK(dac_clk_p_c), 
            .Q(data_reg[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(143[9] 145[42])
    defparam data_reg_i0_i4.GSR = "DISABLED";
    FD1P3AX data_reg_i0_i3 (.D(data_reg[4]), .SP(data_reg_7__N_415), .CK(dac_clk_p_c), 
            .Q(data_reg[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(143[9] 145[42])
    defparam data_reg_i0_i3.GSR = "DISABLED";
    FD1P3AX data_reg_i0_i2 (.D(data_reg[3]), .SP(data_reg_7__N_415), .CK(dac_clk_p_c), 
            .Q(data_reg[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(143[9] 145[42])
    defparam data_reg_i0_i2.GSR = "DISABLED";
    FD1P3AX data_reg_i0_i1 (.D(data_reg[2]), .SP(data_reg_7__N_415), .CK(dac_clk_p_c), 
            .Q(data_reg[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(143[9] 145[42])
    defparam data_reg_i0_i1.GSR = "DISABLED";
    FD1P3AX data_reg_i0_i0 (.D(data_reg[1]), .SP(data_reg_7__N_415), .CK(dac_clk_p_c), 
            .Q(data_reg[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(143[9] 145[42])
    defparam data_reg_i0_i0.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module \txuartlite(TIMING_BITS=24,CLOCKS_PER_BAUD=10000) 
//

module \txuartlite(TIMING_BITS=24,CLOCKS_PER_BAUD=10000)  (n27281, state, 
            dac_clk_p_c, dac_clk_p_c_enable_346, \lcl_data_7__N_510[0] , 
            zero_baud_counter, o_wbu_uart_tx_c, \lcl_data[7] , n29969, 
            GND_net, \lcl_data[6] , \lcl_data_7__N_510[6] , \lcl_data[5] , 
            \lcl_data_7__N_510[5] , \lcl_data[4] , \lcl_data_7__N_510[4] , 
            \lcl_data[3] , \lcl_data_7__N_510[3] , \lcl_data[2] , \lcl_data_7__N_510[2] , 
            \lcl_data[1] , \lcl_data_7__N_510[1] , o_busy_N_535, tx_busy, 
            n18134) /* synthesis syn_module_defined=1 */ ;
    input n27281;
    output [3:0]state;
    input dac_clk_p_c;
    input dac_clk_p_c_enable_346;
    input \lcl_data_7__N_510[0] ;
    output zero_baud_counter;
    output o_wbu_uart_tx_c;
    output \lcl_data[7] ;
    input n29969;
    input GND_net;
    output \lcl_data[6] ;
    input \lcl_data_7__N_510[6] ;
    output \lcl_data[5] ;
    input \lcl_data_7__N_510[5] ;
    output \lcl_data[4] ;
    input \lcl_data_7__N_510[4] ;
    output \lcl_data[3] ;
    input \lcl_data_7__N_510[3] ;
    output \lcl_data[2] ;
    input \lcl_data_7__N_510[2] ;
    output \lcl_data[1] ;
    input \lcl_data_7__N_510[1] ;
    output o_busy_N_535;
    output tx_busy;
    input n18134;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[49:58])
    wire [3:0]state_c;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(83[12:17])
    
    wire n27483;
    wire [7:0]lcl_data;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(84[12:20])
    
    wire zero_baud_counter_N_524;
    wire [23:0]baud_counter;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(82[17:29])
    wire [23:0]baud_counter_23__N_482;
    
    wire n27482, n27484, n27261, n11549, n27485;
    wire [23:0]n108;
    wire [23:0]n133;
    
    wire n27142, zero_baud_counter_N_527, n27486, n20747, n21146, 
        n21154, n21152, n21144, n21130, n21140, n21142, n21132, 
        n17970, n17969, n17968, n17967, n17966, n8982, n17965;
    wire [3:0]n27;
    
    wire n17964, n17963, n17962, n17961, n17960, n17959, n27487;
    
    LUT4 state_596_mux_6_i3_4_lut_then_4_lut (.A(n27281), .B(state[0]), 
         .C(state_c[1]), .D(state_c[3]), .Z(n27483)) /* synthesis lut_function=(!(A (B (C+(D))+!B (D))+!A !(((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(110[14:26])
    defparam state_596_mux_6_i3_4_lut_then_4_lut.init = 16'h553f;
    FD1P3AY lcl_data_i0 (.D(\lcl_data_7__N_510[0] ), .SP(dac_clk_p_c_enable_346), 
            .CK(dac_clk_p_c), .Q(lcl_data[0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(139[9] 143[40])
    defparam lcl_data_i0.GSR = "DISABLED";
    FD1S3AY zero_baud_counter_49 (.D(zero_baud_counter_N_524), .CK(dac_clk_p_c), 
            .Q(zero_baud_counter)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam zero_baud_counter_49.GSR = "DISABLED";
    FD1S3AX baud_counter_i0 (.D(baud_counter_23__N_482[0]), .CK(dac_clk_p_c), 
            .Q(baud_counter[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i0.GSR = "DISABLED";
    PFUMX i25160 (.BLUT(n27482), .ALUT(n27483), .C0(state_c[2]), .Z(n27484));
    LUT4 state_596_mux_6_i3_4_lut_else_4_lut (.A(n27281), .B(state[0]), 
         .C(state_c[1]), .D(state_c[3]), .Z(n27482)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A !(B (C+(D))+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(110[14:26])
    defparam state_596_mux_6_i3_4_lut_else_4_lut.init = 16'h54c0;
    FD1P3IX o_uart_tx_48 (.D(lcl_data[0]), .SP(dac_clk_p_c_enable_346), 
            .CD(n27281), .CK(dac_clk_p_c), .Q(o_wbu_uart_tx_c)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(154[9] 158[29])
    defparam o_uart_tx_48.GSR = "DISABLED";
    LUT4 i1_2_lut_4_lut (.A(state_c[2]), .B(n27261), .C(state_c[1]), .D(zero_baud_counter), 
         .Z(n11549)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(110[14:26])
    defparam i1_2_lut_4_lut.init = 16'hff80;
    LUT4 state_596_mux_6_i4_4_lut_else_4_lut (.A(state_c[2]), .B(state[0]), 
         .C(state_c[1]), .Z(n27485)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(110[14:26])
    defparam state_596_mux_6_i4_4_lut_else_4_lut.init = 16'h8080;
    FD1S3IX baud_counter_i23 (.D(n108[23]), .CK(dac_clk_p_c), .CD(n11549), 
            .Q(baud_counter[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i23.GSR = "DISABLED";
    LUT4 baud_counter_23__I_10_i1_4_lut (.A(n27281), .B(n133[0]), .C(n27142), 
         .D(zero_baud_counter_N_527), .Z(baud_counter_23__N_482[0])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((C+(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(217[12] 224[43])
    defparam baud_counter_23__I_10_i1_4_lut.init = 16'ha0ac;
    LUT4 state_596_mux_6_i4_4_lut_then_4_lut (.A(n27281), .B(state_c[2]), 
         .C(state[0]), .D(state_c[1]), .Z(n27486)) /* synthesis lut_function=(!(A (B+(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(110[14:26])
    defparam state_596_mux_6_i4_4_lut_then_4_lut.init = 16'h5557;
    FD1S3IX baud_counter_i22 (.D(n108[22]), .CK(dac_clk_p_c), .CD(n11549), 
            .Q(baud_counter[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i22.GSR = "DISABLED";
    FD1S3IX baud_counter_i21 (.D(n108[21]), .CK(dac_clk_p_c), .CD(n11549), 
            .Q(baud_counter[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i21.GSR = "DISABLED";
    FD1S3IX baud_counter_i20 (.D(n108[20]), .CK(dac_clk_p_c), .CD(n11549), 
            .Q(baud_counter[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i20.GSR = "DISABLED";
    FD1S3IX baud_counter_i19 (.D(n108[19]), .CK(dac_clk_p_c), .CD(n11549), 
            .Q(baud_counter[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i19.GSR = "DISABLED";
    FD1S3IX baud_counter_i18 (.D(n108[18]), .CK(dac_clk_p_c), .CD(n11549), 
            .Q(baud_counter[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i18.GSR = "DISABLED";
    FD1S3IX baud_counter_i17 (.D(n108[17]), .CK(dac_clk_p_c), .CD(n11549), 
            .Q(baud_counter[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i17.GSR = "DISABLED";
    LUT4 zero_baud_counter_I_0_51_4_lut (.A(n27281), .B(n20747), .C(n27142), 
         .D(zero_baud_counter_N_527), .Z(zero_baud_counter_N_524)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C))+!A !((C+(D))+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(217[12] 224[43])
    defparam zero_baud_counter_I_0_51_4_lut.init = 16'h5f53;
    FD1S3IX baud_counter_i16 (.D(n108[16]), .CK(dac_clk_p_c), .CD(n11549), 
            .Q(baud_counter[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i16.GSR = "DISABLED";
    FD1S3IX baud_counter_i15 (.D(n108[15]), .CK(dac_clk_p_c), .CD(n11549), 
            .Q(baud_counter[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i15.GSR = "DISABLED";
    FD1S3IX baud_counter_i14 (.D(n108[14]), .CK(dac_clk_p_c), .CD(n11549), 
            .Q(baud_counter[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i14.GSR = "DISABLED";
    FD1S3AX baud_counter_i13 (.D(baud_counter_23__N_482[13]), .CK(dac_clk_p_c), 
            .Q(baud_counter[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i13.GSR = "DISABLED";
    FD1S3IX baud_counter_i12 (.D(n108[12]), .CK(dac_clk_p_c), .CD(n11549), 
            .Q(baud_counter[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i12.GSR = "DISABLED";
    FD1S3IX baud_counter_i11 (.D(n108[11]), .CK(dac_clk_p_c), .CD(n11549), 
            .Q(baud_counter[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i11.GSR = "DISABLED";
    FD1S3AX baud_counter_i10 (.D(baud_counter_23__N_482[10]), .CK(dac_clk_p_c), 
            .Q(baud_counter[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i10.GSR = "DISABLED";
    FD1S3AX baud_counter_i9 (.D(baud_counter_23__N_482[9]), .CK(dac_clk_p_c), 
            .Q(baud_counter[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i9.GSR = "DISABLED";
    FD1S3AX baud_counter_i8 (.D(baud_counter_23__N_482[8]), .CK(dac_clk_p_c), 
            .Q(baud_counter[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i8.GSR = "DISABLED";
    FD1S3IX baud_counter_i7 (.D(n108[7]), .CK(dac_clk_p_c), .CD(n11549), 
            .Q(baud_counter[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i7.GSR = "DISABLED";
    FD1S3IX baud_counter_i6 (.D(n108[6]), .CK(dac_clk_p_c), .CD(n11549), 
            .Q(baud_counter[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i6.GSR = "DISABLED";
    FD1S3IX baud_counter_i5 (.D(n108[5]), .CK(dac_clk_p_c), .CD(n11549), 
            .Q(baud_counter[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i5.GSR = "DISABLED";
    FD1S3IX baud_counter_i4 (.D(n108[4]), .CK(dac_clk_p_c), .CD(n11549), 
            .Q(baud_counter[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i4.GSR = "DISABLED";
    LUT4 i1_4_lut (.A(n21146), .B(n21154), .C(n21152), .D(n21144), .Z(n20747)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(207[24:43])
    defparam i1_4_lut.init = 16'hfffe;
    FD1S3AX baud_counter_i3 (.D(baud_counter_23__N_482[3]), .CK(dac_clk_p_c), 
            .Q(baud_counter[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i3.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_106 (.A(baud_counter[13]), .B(baud_counter[7]), .C(baud_counter[21]), 
         .D(baud_counter[11]), .Z(n21146)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(207[24:43])
    defparam i1_4_lut_adj_106.init = 16'hfffe;
    LUT4 i1_4_lut_adj_107 (.A(n21130), .B(baud_counter[0]), .C(n21140), 
         .D(baud_counter[1]), .Z(n21154)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(207[24:43])
    defparam i1_4_lut_adj_107.init = 16'hfffb;
    FD1S3AX baud_counter_i2 (.D(baud_counter_23__N_482[2]), .CK(dac_clk_p_c), 
            .Q(baud_counter[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i2.GSR = "DISABLED";
    FD1S3AX baud_counter_i1 (.D(baud_counter_23__N_482[1]), .CK(dac_clk_p_c), 
            .Q(baud_counter[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i1.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_108 (.A(baud_counter[15]), .B(n21142), .C(n21132), 
         .D(baud_counter[12]), .Z(n21152)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(207[24:43])
    defparam i1_4_lut_adj_108.init = 16'hfffe;
    FD1P3IX lcl_data_i7 (.D(n29969), .SP(zero_baud_counter), .CD(n27281), 
            .CK(dac_clk_p_c), .Q(\lcl_data[7] )) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(139[9] 143[40])
    defparam lcl_data_i7.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_109 (.A(baud_counter[18]), .B(baud_counter[4]), .C(baud_counter[22]), 
         .D(baud_counter[20]), .Z(n21144)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(207[24:43])
    defparam i1_4_lut_adj_109.init = 16'hfffe;
    LUT4 i1_2_lut (.A(baud_counter[8]), .B(baud_counter[17]), .Z(n21130)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(207[24:43])
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i1_4_lut_adj_110 (.A(baud_counter[9]), .B(baud_counter[5]), .C(baud_counter[16]), 
         .D(baud_counter[23]), .Z(n21140)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(207[24:43])
    defparam i1_4_lut_adj_110.init = 16'hfffe;
    LUT4 i1_4_lut_adj_111 (.A(baud_counter[19]), .B(baud_counter[2]), .C(baud_counter[3]), 
         .D(baud_counter[14]), .Z(n21142)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(207[24:43])
    defparam i1_4_lut_adj_111.init = 16'hfffe;
    LUT4 i1_2_lut_adj_112 (.A(baud_counter[6]), .B(baud_counter[10]), .Z(n21132)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(207[24:43])
    defparam i1_2_lut_adj_112.init = 16'heeee;
    LUT4 i1_4_lut_adj_113 (.A(state_c[1]), .B(n27261), .C(state_c[2]), 
         .D(zero_baud_counter), .Z(zero_baud_counter_N_527)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_adj_113.init = 16'h0400;
    CCU2D sub_36_add_2_25 (.A0(baud_counter[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n17970), .S0(n108[23]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_25.INIT0 = 16'h5555;
    defparam sub_36_add_2_25.INIT1 = 16'h0000;
    defparam sub_36_add_2_25.INJECT1_0 = "NO";
    defparam sub_36_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_36_add_2_23 (.A0(baud_counter[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17969), .COUT(n17970), .S0(n108[21]), 
          .S1(n108[22]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_23.INIT0 = 16'h5555;
    defparam sub_36_add_2_23.INIT1 = 16'h5555;
    defparam sub_36_add_2_23.INJECT1_0 = "NO";
    defparam sub_36_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_36_add_2_21 (.A0(baud_counter[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17968), .COUT(n17969), .S0(n108[19]), 
          .S1(n108[20]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_21.INIT0 = 16'h5555;
    defparam sub_36_add_2_21.INIT1 = 16'h5555;
    defparam sub_36_add_2_21.INJECT1_0 = "NO";
    defparam sub_36_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_36_add_2_19 (.A0(baud_counter[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17967), .COUT(n17968), .S0(n108[17]), 
          .S1(n108[18]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_19.INIT0 = 16'h5555;
    defparam sub_36_add_2_19.INIT1 = 16'h5555;
    defparam sub_36_add_2_19.INJECT1_0 = "NO";
    defparam sub_36_add_2_19.INJECT1_1 = "NO";
    FD1P3AY lcl_data_i6 (.D(\lcl_data_7__N_510[6] ), .SP(dac_clk_p_c_enable_346), 
            .CK(dac_clk_p_c), .Q(\lcl_data[6] )) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(139[9] 143[40])
    defparam lcl_data_i6.GSR = "DISABLED";
    FD1P3AY lcl_data_i5 (.D(\lcl_data_7__N_510[5] ), .SP(dac_clk_p_c_enable_346), 
            .CK(dac_clk_p_c), .Q(\lcl_data[5] )) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(139[9] 143[40])
    defparam lcl_data_i5.GSR = "DISABLED";
    FD1P3AY lcl_data_i4 (.D(\lcl_data_7__N_510[4] ), .SP(dac_clk_p_c_enable_346), 
            .CK(dac_clk_p_c), .Q(\lcl_data[4] )) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(139[9] 143[40])
    defparam lcl_data_i4.GSR = "DISABLED";
    FD1P3AY lcl_data_i3 (.D(\lcl_data_7__N_510[3] ), .SP(dac_clk_p_c_enable_346), 
            .CK(dac_clk_p_c), .Q(\lcl_data[3] )) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(139[9] 143[40])
    defparam lcl_data_i3.GSR = "DISABLED";
    FD1P3AY lcl_data_i2 (.D(\lcl_data_7__N_510[2] ), .SP(dac_clk_p_c_enable_346), 
            .CK(dac_clk_p_c), .Q(\lcl_data[2] )) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(139[9] 143[40])
    defparam lcl_data_i2.GSR = "DISABLED";
    FD1P3AY lcl_data_i1 (.D(\lcl_data_7__N_510[1] ), .SP(dac_clk_p_c_enable_346), 
            .CK(dac_clk_p_c), .Q(\lcl_data[1] )) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(139[9] 143[40])
    defparam lcl_data_i1.GSR = "DISABLED";
    LUT4 baud_counter_23__I_10_i14_4_lut (.A(n27281), .B(n133[13]), .C(n27142), 
         .D(zero_baud_counter_N_527), .Z(baud_counter_23__N_482[13])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((C+(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(217[12] 224[43])
    defparam baud_counter_23__I_10_i14_4_lut.init = 16'ha0ac;
    LUT4 i11812_2_lut (.A(n108[13]), .B(zero_baud_counter), .Z(n133[13])) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(224[4:43])
    defparam i11812_2_lut.init = 16'heeee;
    LUT4 baud_counter_23__I_10_i11_4_lut (.A(n27281), .B(n133[10]), .C(n27142), 
         .D(zero_baud_counter_N_527), .Z(baud_counter_23__N_482[10])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((C+(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(217[12] 224[43])
    defparam baud_counter_23__I_10_i11_4_lut.init = 16'ha0ac;
    LUT4 i11813_2_lut (.A(n108[10]), .B(zero_baud_counter), .Z(n133[10])) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(224[4:43])
    defparam i11813_2_lut.init = 16'heeee;
    LUT4 baud_counter_23__I_10_i10_4_lut (.A(n27281), .B(n133[9]), .C(n27142), 
         .D(zero_baud_counter_N_527), .Z(baud_counter_23__N_482[9])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((C+(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(217[12] 224[43])
    defparam baud_counter_23__I_10_i10_4_lut.init = 16'ha0ac;
    LUT4 i11814_2_lut (.A(n108[9]), .B(zero_baud_counter), .Z(n133[9])) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(224[4:43])
    defparam i11814_2_lut.init = 16'heeee;
    LUT4 baud_counter_23__I_10_i9_4_lut (.A(n27281), .B(n133[8]), .C(n27142), 
         .D(zero_baud_counter_N_527), .Z(baud_counter_23__N_482[8])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((C+(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(217[12] 224[43])
    defparam baud_counter_23__I_10_i9_4_lut.init = 16'ha0ac;
    LUT4 i11815_2_lut (.A(n108[8]), .B(zero_baud_counter), .Z(n133[8])) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(224[4:43])
    defparam i11815_2_lut.init = 16'heeee;
    CCU2D sub_36_add_2_17 (.A0(baud_counter[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17966), .COUT(n17967), .S0(n108[15]), 
          .S1(n108[16]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_17.INIT0 = 16'h5555;
    defparam sub_36_add_2_17.INIT1 = 16'h5555;
    defparam sub_36_add_2_17.INJECT1_0 = "NO";
    defparam sub_36_add_2_17.INJECT1_1 = "NO";
    LUT4 baud_counter_23__I_10_i4_4_lut (.A(n27281), .B(n133[3]), .C(n27142), 
         .D(zero_baud_counter_N_527), .Z(baud_counter_23__N_482[3])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((C+(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(217[12] 224[43])
    defparam baud_counter_23__I_10_i4_4_lut.init = 16'ha0ac;
    LUT4 i11816_2_lut (.A(n108[3]), .B(zero_baud_counter), .Z(n133[3])) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(224[4:43])
    defparam i11816_2_lut.init = 16'heeee;
    LUT4 baud_counter_23__I_10_i3_4_lut (.A(n27281), .B(n133[2]), .C(n27142), 
         .D(zero_baud_counter_N_527), .Z(baud_counter_23__N_482[2])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((C+(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(217[12] 224[43])
    defparam baud_counter_23__I_10_i3_4_lut.init = 16'ha0ac;
    LUT4 i11817_2_lut (.A(n108[2]), .B(zero_baud_counter), .Z(n133[2])) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(224[4:43])
    defparam i11817_2_lut.init = 16'heeee;
    LUT4 baud_counter_23__I_10_i2_4_lut (.A(n27281), .B(n133[1]), .C(n27142), 
         .D(zero_baud_counter_N_527), .Z(baud_counter_23__N_482[1])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((C+(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(217[12] 224[43])
    defparam baud_counter_23__I_10_i2_4_lut.init = 16'ha0ac;
    LUT4 i11818_2_lut (.A(n108[1]), .B(zero_baud_counter), .Z(n133[1])) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(224[4:43])
    defparam i11818_2_lut.init = 16'heeee;
    LUT4 i23025_2_lut (.A(o_busy_N_535), .B(zero_baud_counter), .Z(n8982)) /* synthesis lut_function=(!(A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(97[8] 113[6])
    defparam i23025_2_lut.init = 16'h7777;
    LUT4 i790_4_lut (.A(state_c[2]), .B(state_c[3]), .C(state_c[1]), .D(state[0]), 
         .Z(o_busy_N_535)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;
    defparam i790_4_lut.init = 16'hccc8;
    CCU2D sub_36_add_2_15 (.A0(baud_counter[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17965), .COUT(n17966), .S0(n108[13]), 
          .S1(n108[14]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_15.INIT0 = 16'h5555;
    defparam sub_36_add_2_15.INIT1 = 16'h5555;
    defparam sub_36_add_2_15.INJECT1_0 = "NO";
    defparam sub_36_add_2_15.INJECT1_1 = "NO";
    LUT4 state_596_mux_6_i2_4_lut (.A(state_c[1]), .B(n27281), .C(o_busy_N_535), 
         .D(state[0]), .Z(n27[1])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(110[14:26])
    defparam state_596_mux_6_i2_4_lut.init = 16'h353a;
    LUT4 i1_2_lut_rep_596 (.A(state[0]), .B(state_c[3]), .Z(n27261)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(110[14:26])
    defparam i1_2_lut_rep_596.init = 16'h8888;
    LUT4 i1_3_lut_rep_477_4_lut (.A(state[0]), .B(state_c[3]), .C(state_c[1]), 
         .D(state_c[2]), .Z(n27142)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(110[14:26])
    defparam i1_3_lut_rep_477_4_lut.init = 16'h8000;
    LUT4 i11316_2_lut (.A(n108[0]), .B(zero_baud_counter), .Z(n133[0])) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(224[4:43])
    defparam i11316_2_lut.init = 16'heeee;
    CCU2D sub_36_add_2_13 (.A0(baud_counter[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17964), .COUT(n17965), .S0(n108[11]), 
          .S1(n108[12]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_13.INIT0 = 16'h5555;
    defparam sub_36_add_2_13.INIT1 = 16'h5555;
    defparam sub_36_add_2_13.INJECT1_0 = "NO";
    defparam sub_36_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_36_add_2_11 (.A0(baud_counter[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17963), .COUT(n17964), .S0(n108[9]), .S1(n108[10]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_11.INIT0 = 16'h5555;
    defparam sub_36_add_2_11.INIT1 = 16'h5555;
    defparam sub_36_add_2_11.INJECT1_0 = "NO";
    defparam sub_36_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_36_add_2_9 (.A0(baud_counter[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17962), .COUT(n17963), .S0(n108[7]), .S1(n108[8]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_9.INIT0 = 16'h5555;
    defparam sub_36_add_2_9.INIT1 = 16'h5555;
    defparam sub_36_add_2_9.INJECT1_0 = "NO";
    defparam sub_36_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_36_add_2_7 (.A0(baud_counter[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17961), .COUT(n17962), .S0(n108[5]), .S1(n108[6]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_7.INIT0 = 16'h5555;
    defparam sub_36_add_2_7.INIT1 = 16'h5555;
    defparam sub_36_add_2_7.INJECT1_0 = "NO";
    defparam sub_36_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_36_add_2_5 (.A0(baud_counter[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17960), .COUT(n17961), .S0(n108[3]), .S1(n108[4]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_5.INIT0 = 16'h5555;
    defparam sub_36_add_2_5.INIT1 = 16'h5555;
    defparam sub_36_add_2_5.INJECT1_0 = "NO";
    defparam sub_36_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_36_add_2_3 (.A0(baud_counter[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17959), .COUT(n17960), .S0(n108[1]), .S1(n108[2]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_3.INIT0 = 16'h5555;
    defparam sub_36_add_2_3.INIT1 = 16'h5555;
    defparam sub_36_add_2_3.INJECT1_0 = "NO";
    defparam sub_36_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_36_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(baud_counter[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n17959), .S1(n108[0]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_1.INIT0 = 16'hF000;
    defparam sub_36_add_2_1.INIT1 = 16'h5555;
    defparam sub_36_add_2_1.INJECT1_0 = "NO";
    defparam sub_36_add_2_1.INJECT1_1 = "NO";
    FD1S3JX r_busy_45 (.D(n8982), .CK(dac_clk_p_c), .PD(n27281), .Q(tx_busy)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(92[9] 114[5])
    defparam r_busy_45.GSR = "DISABLED";
    FD1P3AX state_596__i3 (.D(n27487), .SP(zero_baud_counter), .CK(dac_clk_p_c), 
            .Q(state_c[3]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(110[14:26])
    defparam state_596__i3.GSR = "DISABLED";
    FD1P3AX state_596__i2 (.D(n27484), .SP(zero_baud_counter), .CK(dac_clk_p_c), 
            .Q(state_c[2]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(110[14:26])
    defparam state_596__i2.GSR = "DISABLED";
    FD1P3AX state_596__i1 (.D(n27[1]), .SP(zero_baud_counter), .CK(dac_clk_p_c), 
            .Q(state_c[1]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(110[14:26])
    defparam state_596__i1.GSR = "DISABLED";
    FD1P3AX state_596__i0 (.D(n18134), .SP(zero_baud_counter), .CK(dac_clk_p_c), 
            .Q(state[0]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(110[14:26])
    defparam state_596__i0.GSR = "DISABLED";
    PFUMX i25162 (.BLUT(n27485), .ALUT(n27486), .C0(state_c[3]), .Z(n27487));
    
endmodule
//
// Verilog Description of module TSALL
// module not written out since it is a black-box. 
//

//
// Verilog Description of module efb_inst
//

module efb_inst (dac_clk_p_c, i_sw0_c, wb_cyc, wb_lo_data_7__N_96, wb_we, 
            \wb_addr[7] , \wb_addr[6] , \wb_addr[5] , \wb_addr[4] , 
            \wb_addr[3] , \wb_addr[2] , \wb_addr[1] , \wb_addr[0] , 
            \wb_odata[7] , \wb_odata[6] , \wb_odata[5] , \wb_odata[4] , 
            \wb_odata[3] , \wb_odata[2] , \wb_odata[1] , \wb_odata[0] , 
            pll_data_o, pll_ack, wb_lo_data, wb_lo_ack, pll_clk, pll_rst, 
            pll_stb, pll_we, pll_addr, pll_data_i, GND_net, VCC_net) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;
    input dac_clk_p_c;
    input i_sw0_c;
    input wb_cyc;
    input wb_lo_data_7__N_96;
    input wb_we;
    input \wb_addr[7] ;
    input \wb_addr[6] ;
    input \wb_addr[5] ;
    input \wb_addr[4] ;
    input \wb_addr[3] ;
    input \wb_addr[2] ;
    input \wb_addr[1] ;
    input \wb_addr[0] ;
    input \wb_odata[7] ;
    input \wb_odata[6] ;
    input \wb_odata[5] ;
    input \wb_odata[4] ;
    input \wb_odata[3] ;
    input \wb_odata[2] ;
    input \wb_odata[1] ;
    input \wb_odata[0] ;
    input [7:0]pll_data_o;
    input pll_ack;
    output [7:0]wb_lo_data;
    output wb_lo_ack;
    output pll_clk;
    output pll_rst;
    output pll_stb;
    output pll_we;
    output [4:0]pll_addr;
    output [7:0]pll_data_i;
    input GND_net;
    input VCC_net;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[49:58])
    
    EFB EFBInst_0 (.WBCLKI(dac_clk_p_c), .WBRSTI(i_sw0_c), .WBCYCI(wb_cyc), 
        .WBSTBI(wb_lo_data_7__N_96), .WBWEI(wb_we), .WBADRI0(\wb_addr[0] ), 
        .WBADRI1(\wb_addr[1] ), .WBADRI2(\wb_addr[2] ), .WBADRI3(\wb_addr[3] ), 
        .WBADRI4(\wb_addr[4] ), .WBADRI5(\wb_addr[5] ), .WBADRI6(\wb_addr[6] ), 
        .WBADRI7(\wb_addr[7] ), .WBDATI0(\wb_odata[0] ), .WBDATI1(\wb_odata[1] ), 
        .WBDATI2(\wb_odata[2] ), .WBDATI3(\wb_odata[3] ), .WBDATI4(\wb_odata[4] ), 
        .WBDATI5(\wb_odata[5] ), .WBDATI6(\wb_odata[6] ), .WBDATI7(\wb_odata[7] ), 
        .I2C1SCLI(GND_net), .I2C1SDAI(GND_net), .I2C2SCLI(GND_net), .I2C2SDAI(GND_net), 
        .SPISCKI(GND_net), .SPIMISOI(GND_net), .SPIMOSII(GND_net), .SPISCSN(GND_net), 
        .TCCLKI(GND_net), .TCRSTN(GND_net), .TCIC(GND_net), .UFMSN(VCC_net), 
        .PLL0DATI0(pll_data_o[0]), .PLL0DATI1(pll_data_o[1]), .PLL0DATI2(pll_data_o[2]), 
        .PLL0DATI3(pll_data_o[3]), .PLL0DATI4(pll_data_o[4]), .PLL0DATI5(pll_data_o[5]), 
        .PLL0DATI6(pll_data_o[6]), .PLL0DATI7(pll_data_o[7]), .PLL0ACKI(pll_ack), 
        .PLL1DATI0(GND_net), .PLL1DATI1(GND_net), .PLL1DATI2(GND_net), 
        .PLL1DATI3(GND_net), .PLL1DATI4(GND_net), .PLL1DATI5(GND_net), 
        .PLL1DATI6(GND_net), .PLL1DATI7(GND_net), .PLL1ACKI(GND_net), 
        .WBDATO0(wb_lo_data[0]), .WBDATO1(wb_lo_data[1]), .WBDATO2(wb_lo_data[2]), 
        .WBDATO3(wb_lo_data[3]), .WBDATO4(wb_lo_data[4]), .WBDATO5(wb_lo_data[5]), 
        .WBDATO6(wb_lo_data[6]), .WBDATO7(wb_lo_data[7]), .WBACKO(wb_lo_ack), 
        .PLLCLKO(pll_clk), .PLLRSTO(pll_rst), .PLL0STBO(pll_stb), .PLLWEO(pll_we), 
        .PLLADRO0(pll_addr[0]), .PLLADRO1(pll_addr[1]), .PLLADRO2(pll_addr[2]), 
        .PLLADRO3(pll_addr[3]), .PLLADRO4(pll_addr[4]), .PLLDATO0(pll_data_i[0]), 
        .PLLDATO1(pll_data_i[1]), .PLLDATO2(pll_data_i[2]), .PLLDATO3(pll_data_i[3]), 
        .PLLDATO4(pll_data_i[4]), .PLLDATO5(pll_data_i[5]), .PLLDATO6(pll_data_i[6]), 
        .PLLDATO7(pll_data_i[7])) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=8, LSE_LCOL=11, LSE_RCOL=4, LSE_LLINE=187, LSE_RLINE=199 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(187[11] 199[4])
    defparam EFBInst_0.EFB_I2C1 = "DISABLED";
    defparam EFBInst_0.EFB_I2C2 = "DISABLED";
    defparam EFBInst_0.EFB_SPI = "DISABLED";
    defparam EFBInst_0.EFB_TC = "DISABLED";
    defparam EFBInst_0.EFB_TC_PORTMODE = "WB";
    defparam EFBInst_0.EFB_UFM = "DISABLED";
    defparam EFBInst_0.EFB_WB_CLK_FREQ = "50.0";
    defparam EFBInst_0.DEV_DENSITY = "6900L";
    defparam EFBInst_0.UFM_INIT_PAGES = 0;
    defparam EFBInst_0.UFM_INIT_START_PAGE = 0;
    defparam EFBInst_0.UFM_INIT_ALL_ZEROS = "ENABLED";
    defparam EFBInst_0.UFM_INIT_FILE_NAME = "NONE";
    defparam EFBInst_0.UFM_INIT_FILE_FORMAT = "HEX";
    defparam EFBInst_0.I2C1_ADDRESSING = "7BIT";
    defparam EFBInst_0.I2C2_ADDRESSING = "7BIT";
    defparam EFBInst_0.I2C1_SLAVE_ADDR = "0b1000001";
    defparam EFBInst_0.I2C2_SLAVE_ADDR = "0b1000010";
    defparam EFBInst_0.I2C1_BUS_PERF = "100kHz";
    defparam EFBInst_0.I2C2_BUS_PERF = "100kHz";
    defparam EFBInst_0.I2C1_CLK_DIVIDER = 1;
    defparam EFBInst_0.I2C2_CLK_DIVIDER = 1;
    defparam EFBInst_0.I2C1_GEN_CALL = "DISABLED";
    defparam EFBInst_0.I2C2_GEN_CALL = "DISABLED";
    defparam EFBInst_0.I2C1_WAKEUP = "DISABLED";
    defparam EFBInst_0.I2C2_WAKEUP = "DISABLED";
    defparam EFBInst_0.SPI_MODE = "MASTER";
    defparam EFBInst_0.SPI_CLK_DIVIDER = 1;
    defparam EFBInst_0.SPI_LSB_FIRST = "DISABLED";
    defparam EFBInst_0.SPI_CLK_INV = "DISABLED";
    defparam EFBInst_0.SPI_PHASE_ADJ = "DISABLED";
    defparam EFBInst_0.SPI_SLAVE_HANDSHAKE = "DISABLED";
    defparam EFBInst_0.SPI_INTR_TXRDY = "DISABLED";
    defparam EFBInst_0.SPI_INTR_RXRDY = "DISABLED";
    defparam EFBInst_0.SPI_INTR_TXOVR = "DISABLED";
    defparam EFBInst_0.SPI_INTR_RXOVR = "DISABLED";
    defparam EFBInst_0.SPI_WAKEUP = "DISABLED";
    defparam EFBInst_0.TC_MODE = "CTCM";
    defparam EFBInst_0.TC_SCLK_SEL = "PCLOCK";
    defparam EFBInst_0.TC_CCLK_SEL = 1;
    defparam EFBInst_0.GSR = "ENABLED";
    defparam EFBInst_0.TC_TOP_SET = 65535;
    defparam EFBInst_0.TC_OCR_SET = 32767;
    defparam EFBInst_0.TC_OC_MODE = "TOGGLE";
    defparam EFBInst_0.TC_RESETN = "ENABLED";
    defparam EFBInst_0.TC_TOP_SEL = "OFF";
    defparam EFBInst_0.TC_OV_INT = "OFF";
    defparam EFBInst_0.TC_OCR_INT = "OFF";
    defparam EFBInst_0.TC_ICR_INT = "OFF";
    defparam EFBInst_0.TC_OVERFLOW = "DISABLED";
    defparam EFBInst_0.TC_ICAPTURE = "DISABLED";
    
endmodule
//
// Verilog Description of module clock_phase_shifter
//

module clock_phase_shifter (q_clk_p_c, i_clk_2f_N_2268, q_clk_n_c, i_clk_p_c, 
            lo_pll_out, i_clk_n_c) /* synthesis syn_module_defined=1 */ ;
    output q_clk_p_c;
    input i_clk_2f_N_2268;
    input q_clk_n_c;
    output i_clk_p_c;
    input lo_pll_out;
    input i_clk_n_c;
    
    wire i_clk_2f_N_2268 /* synthesis is_inv_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/clock_phase_shifter.v(11[21:28])
    wire lo_pll_out /* synthesis is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(166[6:16])
    
    FD1S3AX o_clk_q_10 (.D(q_clk_n_c), .CK(i_clk_2f_N_2268), .Q(q_clk_p_c)) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=21, LSE_RCOL=2, LSE_LLINE=167, LSE_RLINE=171 */ ;   // d:/documents/git_local/fm_modulator/rtl/clock_phase_shifter.v(17[8] 19[4])
    defparam o_clk_q_10.GSR = "DISABLED";
    FD1S3AX o_clk_i_9 (.D(i_clk_n_c), .CK(lo_pll_out), .Q(i_clk_p_c)) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=21, LSE_RCOL=2, LSE_LLINE=167, LSE_RLINE=171 */ ;   // d:/documents/git_local/fm_modulator/rtl/clock_phase_shifter.v(13[8] 15[4])
    defparam o_clk_i_9.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module sys_clk
//

module sys_clk (i_ref_clk_c, dac_clk_p_c, GND_net) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;
    input i_ref_clk_c;
    output dac_clk_p_c;
    input GND_net;
    
    wire i_ref_clk_c /* synthesis is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(26[12:21])
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[49:58])
    
    EHXPLLJ PLLInst_0 (.CLKI(i_ref_clk_c), .CLKFB(dac_clk_p_c), .PHASESEL0(GND_net), 
            .PHASESEL1(GND_net), .PHASEDIR(GND_net), .PHASESTEP(GND_net), 
            .LOADREG(GND_net), .STDBY(GND_net), .PLLWAKESYNC(GND_net), 
            .RST(GND_net), .RESETC(GND_net), .RESETD(GND_net), .RESETM(GND_net), 
            .ENCLKOP(GND_net), .ENCLKOS(GND_net), .ENCLKOS2(GND_net), 
            .ENCLKOS3(GND_net), .PLLCLK(GND_net), .PLLRST(GND_net), .PLLSTB(GND_net), 
            .PLLWE(GND_net), .PLLDATI0(GND_net), .PLLDATI1(GND_net), .PLLDATI2(GND_net), 
            .PLLDATI3(GND_net), .PLLDATI4(GND_net), .PLLDATI5(GND_net), 
            .PLLDATI6(GND_net), .PLLDATI7(GND_net), .PLLADDR0(GND_net), 
            .PLLADDR1(GND_net), .PLLADDR2(GND_net), .PLLADDR3(GND_net), 
            .PLLADDR4(GND_net), .CLKOP(dac_clk_p_c)) /* synthesis FREQUENCY_PIN_CLKOP="72.000000", FREQUENCY_PIN_CLKI="12.000000", ICP_CURRENT="9", LPF_RESISTOR="72", syn_instantiated=1, LSE_LINE_FILE_ID=8, LSE_LCOL=10, LSE_RCOL=54, LSE_LLINE=47, LSE_RLINE=47 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(47[10:54])
    defparam PLLInst_0.CLKI_DIV = 1;
    defparam PLLInst_0.CLKFB_DIV = 6;
    defparam PLLInst_0.CLKOP_DIV = 7;
    defparam PLLInst_0.CLKOS_DIV = 1;
    defparam PLLInst_0.CLKOS2_DIV = 1;
    defparam PLLInst_0.CLKOS3_DIV = 1;
    defparam PLLInst_0.CLKOP_ENABLE = "ENABLED";
    defparam PLLInst_0.CLKOS_ENABLE = "DISABLED";
    defparam PLLInst_0.CLKOS2_ENABLE = "DISABLED";
    defparam PLLInst_0.CLKOS3_ENABLE = "DISABLED";
    defparam PLLInst_0.VCO_BYPASS_A0 = "DISABLED";
    defparam PLLInst_0.VCO_BYPASS_B0 = "DISABLED";
    defparam PLLInst_0.VCO_BYPASS_C0 = "DISABLED";
    defparam PLLInst_0.VCO_BYPASS_D0 = "DISABLED";
    defparam PLLInst_0.CLKOP_CPHASE = 6;
    defparam PLLInst_0.CLKOS_CPHASE = 0;
    defparam PLLInst_0.CLKOS2_CPHASE = 0;
    defparam PLLInst_0.CLKOS3_CPHASE = 0;
    defparam PLLInst_0.CLKOP_FPHASE = 0;
    defparam PLLInst_0.CLKOS_FPHASE = 0;
    defparam PLLInst_0.CLKOS2_FPHASE = 0;
    defparam PLLInst_0.CLKOS3_FPHASE = 0;
    defparam PLLInst_0.FEEDBK_PATH = "CLKOP";
    defparam PLLInst_0.FRACN_ENABLE = "DISABLED";
    defparam PLLInst_0.FRACN_DIV = 0;
    defparam PLLInst_0.CLKOP_TRIM_POL = "RISING";
    defparam PLLInst_0.CLKOP_TRIM_DELAY = 0;
    defparam PLLInst_0.CLKOS_TRIM_POL = "FALLING";
    defparam PLLInst_0.CLKOS_TRIM_DELAY = 0;
    defparam PLLInst_0.PLL_USE_WB = "DISABLED";
    defparam PLLInst_0.PREDIVIDER_MUXA1 = 0;
    defparam PLLInst_0.PREDIVIDER_MUXB1 = 0;
    defparam PLLInst_0.PREDIVIDER_MUXC1 = 0;
    defparam PLLInst_0.PREDIVIDER_MUXD1 = 0;
    defparam PLLInst_0.OUTDIVIDER_MUXA2 = "DIVA";
    defparam PLLInst_0.OUTDIVIDER_MUXB2 = "DIVB";
    defparam PLLInst_0.OUTDIVIDER_MUXC2 = "DIVC";
    defparam PLLInst_0.OUTDIVIDER_MUXD2 = "DIVD";
    defparam PLLInst_0.PLL_LOCK_MODE = 0;
    defparam PLLInst_0.STDBY_ENABLE = "DISABLED";
    defparam PLLInst_0.DPHASE_SOURCE = "DISABLED";
    defparam PLLInst_0.PLLRST_ENA = "DISABLED";
    defparam PLLInst_0.MRST_ENA = "DISABLED";
    defparam PLLInst_0.DCRST_ENA = "DISABLED";
    defparam PLLInst_0.DDRST_ENA = "DISABLED";
    defparam PLLInst_0.INTFB_WAKE = "DISABLED";
    
endmodule
//
// Verilog Description of module dynamic_pll
//

module dynamic_pll (i_clk_2f_N_2268, lo_pll_out, i_ref_clk_c, pll_clk, 
            pll_rst, pll_stb, pll_we, pll_data_i, pll_addr, pll_data_o, 
            pll_ack, GND_net) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;
    output i_clk_2f_N_2268;
    output lo_pll_out;
    input i_ref_clk_c;
    input pll_clk;
    input pll_rst;
    input pll_stb;
    input pll_we;
    input [7:0]pll_data_i;
    input [4:0]pll_addr;
    output [7:0]pll_data_o;
    output pll_ack;
    input GND_net;
    
    wire i_clk_2f_N_2268 /* synthesis is_inv_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/clock_phase_shifter.v(11[21:28])
    wire lo_pll_out /* synthesis is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(166[6:16])
    wire i_ref_clk_c /* synthesis is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(26[12:21])
    
    INV i26979 (.A(lo_pll_out), .Z(i_clk_2f_N_2268));
    EHXPLLJ PLLInst_0 (.CLKI(i_ref_clk_c), .CLKFB(lo_pll_out), .PHASESEL0(GND_net), 
            .PHASESEL1(GND_net), .PHASEDIR(GND_net), .PHASESTEP(GND_net), 
            .LOADREG(GND_net), .STDBY(GND_net), .PLLWAKESYNC(GND_net), 
            .RST(GND_net), .RESETC(GND_net), .RESETD(GND_net), .RESETM(GND_net), 
            .ENCLKOP(GND_net), .ENCLKOS(GND_net), .ENCLKOS2(GND_net), 
            .ENCLKOS3(GND_net), .PLLCLK(pll_clk), .PLLRST(pll_rst), .PLLSTB(pll_stb), 
            .PLLWE(pll_we), .PLLDATI0(pll_data_i[0]), .PLLDATI1(pll_data_i[1]), 
            .PLLDATI2(pll_data_i[2]), .PLLDATI3(pll_data_i[3]), .PLLDATI4(pll_data_i[4]), 
            .PLLDATI5(pll_data_i[5]), .PLLDATI6(pll_data_i[6]), .PLLDATI7(pll_data_i[7]), 
            .PLLADDR0(pll_addr[0]), .PLLADDR1(pll_addr[1]), .PLLADDR2(pll_addr[2]), 
            .PLLADDR3(pll_addr[3]), .PLLADDR4(pll_addr[4]), .CLKOP(lo_pll_out), 
            .PLLDATO0(pll_data_o[0]), .PLLDATO1(pll_data_o[1]), .PLLDATO2(pll_data_o[2]), 
            .PLLDATO3(pll_data_o[3]), .PLLDATO4(pll_data_o[4]), .PLLDATO5(pll_data_o[5]), 
            .PLLDATO6(pll_data_o[6]), .PLLDATO7(pll_data_o[7]), .PLLACK(pll_ack)) /* synthesis FREQUENCY_PIN_CLKOP="420.000000", FREQUENCY_PIN_CLKI="12.000000", ICP_CURRENT="6", LPF_RESISTOR="8", syn_instantiated=1, LSE_LINE_FILE_ID=8, LSE_LCOL=14, LSE_RCOL=5, LSE_LLINE=174, LSE_RLINE=185 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(174[14] 185[5])
    defparam PLLInst_0.CLKI_DIV = 1;
    defparam PLLInst_0.CLKFB_DIV = 35;
    defparam PLLInst_0.CLKOP_DIV = 1;
    defparam PLLInst_0.CLKOS_DIV = 1;
    defparam PLLInst_0.CLKOS2_DIV = 1;
    defparam PLLInst_0.CLKOS3_DIV = 1;
    defparam PLLInst_0.CLKOP_ENABLE = "ENABLED";
    defparam PLLInst_0.CLKOS_ENABLE = "DISABLED";
    defparam PLLInst_0.CLKOS2_ENABLE = "DISABLED";
    defparam PLLInst_0.CLKOS3_ENABLE = "DISABLED";
    defparam PLLInst_0.VCO_BYPASS_A0 = "DISABLED";
    defparam PLLInst_0.VCO_BYPASS_B0 = "DISABLED";
    defparam PLLInst_0.VCO_BYPASS_C0 = "DISABLED";
    defparam PLLInst_0.VCO_BYPASS_D0 = "DISABLED";
    defparam PLLInst_0.CLKOP_CPHASE = 0;
    defparam PLLInst_0.CLKOS_CPHASE = 0;
    defparam PLLInst_0.CLKOS2_CPHASE = 0;
    defparam PLLInst_0.CLKOS3_CPHASE = 0;
    defparam PLLInst_0.CLKOP_FPHASE = 0;
    defparam PLLInst_0.CLKOS_FPHASE = 0;
    defparam PLLInst_0.CLKOS2_FPHASE = 0;
    defparam PLLInst_0.CLKOS3_FPHASE = 0;
    defparam PLLInst_0.FEEDBK_PATH = "CLKOP";
    defparam PLLInst_0.FRACN_ENABLE = "ENABLED";
    defparam PLLInst_0.FRACN_DIV = 2731;
    defparam PLLInst_0.CLKOP_TRIM_POL = "RISING";
    defparam PLLInst_0.CLKOP_TRIM_DELAY = 0;
    defparam PLLInst_0.CLKOS_TRIM_POL = "FALLING";
    defparam PLLInst_0.CLKOS_TRIM_DELAY = 0;
    defparam PLLInst_0.PLL_USE_WB = "ENABLED";
    defparam PLLInst_0.PREDIVIDER_MUXA1 = 0;
    defparam PLLInst_0.PREDIVIDER_MUXB1 = 0;
    defparam PLLInst_0.PREDIVIDER_MUXC1 = 0;
    defparam PLLInst_0.PREDIVIDER_MUXD1 = 0;
    defparam PLLInst_0.OUTDIVIDER_MUXA2 = "DIVA";
    defparam PLLInst_0.OUTDIVIDER_MUXB2 = "DIVB";
    defparam PLLInst_0.OUTDIVIDER_MUXC2 = "DIVC";
    defparam PLLInst_0.OUTDIVIDER_MUXD2 = "DIVD";
    defparam PLLInst_0.PLL_LOCK_MODE = 0;
    defparam PLLInst_0.STDBY_ENABLE = "DISABLED";
    defparam PLLInst_0.DPHASE_SOURCE = "DISABLED";
    defparam PLLInst_0.PLLRST_ENA = "DISABLED";
    defparam PLLInst_0.MRST_ENA = "DISABLED";
    defparam PLLInst_0.DCRST_ENA = "DISABLED";
    defparam PLLInst_0.DDRST_ENA = "DISABLED";
    defparam PLLInst_0.INTFB_WAKE = "DISABLED";
    
endmodule
//
// Verilog Description of module fm_generator_wb_slave
//

module fm_generator_wb_slave (dac_clk_p_c, wb_odata, i_sw0_c, wb_fm_data, 
            wb_fm_ack, o_dac_a_9__N_1, \wb_addr[0] , \wb_addr[1] , \power_counter[1] , 
            \smpl_register[1] , n2122, n27114, n27304, n27313, \wb_addr[15] , 
            \wb_addr[8] , \wb_addr[12] , GND_net, o_dac_a_c_7, o_dac_a_c_6, 
            o_dac_a_c_5, o_dac_a_c_4, o_dac_a_c_3, o_dac_a_c_2, o_dac_a_c_1, 
            o_dac_a_c_0, o_dac_b_c_15, o_dac_b_c_9, o_dac_cw_b_c, n27380, 
            o_dac_a_c_9, n21102, n38, n2, \smpl_register[5] , n27049, 
            n2_adj_1, \smpl_register[20] , n27061, n2_adj_2, \smpl_register[18] , 
            n27059, n2_adj_3, \smpl_register[17] , n27058, n2_adj_4, 
            \smpl_register[16] , n27057, n2_adj_5, \smpl_register[29] , 
            n27056, n2_adj_6, \smpl_register[10] , n27051, n2_adj_7, 
            \smpl_register[9] , n27050, n21088, n21078, n21044, n29969, 
            o_dac_b_c_7, n29968, o_dac_b_c_14, o_dac_b_c_13, o_dac_b_c_12, 
            o_dac_b_c_11, o_dac_b_c_10, n3639, o_dac_b_c_8) /* synthesis syn_module_defined=1 */ ;
    input dac_clk_p_c;
    input [31:0]wb_odata;
    input i_sw0_c;
    output [31:0]wb_fm_data;
    output wb_fm_ack;
    input o_dac_a_9__N_1;
    input \wb_addr[0] ;
    input \wb_addr[1] ;
    input \power_counter[1] ;
    input \smpl_register[1] ;
    output n2122;
    input n27114;
    input n27304;
    input n27313;
    input \wb_addr[15] ;
    input \wb_addr[8] ;
    input \wb_addr[12] ;
    input GND_net;
    output o_dac_a_c_7;
    output o_dac_a_c_6;
    output o_dac_a_c_5;
    output o_dac_a_c_4;
    output o_dac_a_c_3;
    output o_dac_a_c_2;
    output o_dac_a_c_1;
    output o_dac_a_c_0;
    output o_dac_b_c_15;
    output o_dac_b_c_9;
    output o_dac_cw_b_c;
    output n27380;
    output o_dac_a_c_9;
    input n21102;
    input n38;
    input n2;
    input \smpl_register[5] ;
    output n27049;
    input n2_adj_1;
    input \smpl_register[20] ;
    output n27061;
    input n2_adj_2;
    input \smpl_register[18] ;
    output n27059;
    input n2_adj_3;
    input \smpl_register[17] ;
    output n27058;
    input n2_adj_4;
    input \smpl_register[16] ;
    output n27057;
    input n2_adj_5;
    input \smpl_register[29] ;
    output n27056;
    input n2_adj_6;
    input \smpl_register[10] ;
    output n27051;
    input n2_adj_7;
    input \smpl_register[9] ;
    output n27050;
    input n21088;
    input n21078;
    input n21044;
    input n29969;
    output o_dac_b_c_7;
    input n29968;
    output o_dac_b_c_14;
    output o_dac_b_c_13;
    output o_dac_b_c_12;
    output o_dac_b_c_11;
    output o_dac_b_c_10;
    output n3639;
    output o_dac_b_c_8;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[49:58])
    wire [15:0]modulation_output /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(73[39:56])
    wire [15:0]o_sample_i /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[39:49])
    wire o_dac_b_c_15 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire o_dac_b_c_7 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire o_dac_b_c_14 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire o_dac_b_c_13 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire o_dac_b_c_12 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire o_dac_b_c_11 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire o_dac_b_c_10 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire n3639 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire o_dac_b_c_8 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire [31:0]\addr_space[3] ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(36[12:22])
    
    wire dac_clk_p_c_enable_149;
    wire [31:0]\addr_space[0] ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(36[12:22])
    
    wire dac_clk_p_c_enable_116;
    wire [31:0]\addr_space[1] ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(36[12:22])
    
    wire dac_clk_p_c_enable_73;
    wire [31:0]\addr_space[2] ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(36[12:22])
    
    wire dac_clk_p_c_enable_105;
    wire [31:0]o_wb_data_31__N_1336;
    wire [30:0]carrier_center_increment_offset_rs;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(63[67:101])
    wire [30:0]carrier_center_increment_offset_rs_30__N_1559;
    wire [30:0]carrier_increment;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(64[31:48])
    wire [30:0]carrier_increment_30__N_1590;
    wire [16:0]sine_lookup_width_minus_modulation_deviation_amount;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(85[27:78])
    wire [31:0]sine_lookup_width_minus_modulation_deviation_amount_16__N_1621;
    wire [16:0]modulation_deviation_amount_minus_sine_lookup_width;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(85[80:131])
    wire [30:0]carrier_center_increment_offset_ls;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(63[31:65])
    
    wire n20732;
    wire [15:0]n1109;
    wire [15:0]n31;
    
    wire n178, n27121, n69, n100, n22746, n25046, cw_mux_dac_a_mux_sel, 
        dac_clk_p_c_enable_218, cw_N_1877, n21208, n63, n94, n22774, 
        n64, n95, n25141, n43, n25039, n21206, n21210, n21196, 
        n178_adj_2995, n25041, n25042, n40, n25044, n36, n44, 
        n25045, n14, n25048, n37, n41, n25049, n22482, n22483, 
        n4, n6, n25040, n27250, n124, dac_clk_p_c_enable_488, n3, 
        n5, n25139, n25140, n73, n17925, n14676, n17924;
    wire [15:0]n61;
    wire [30:0]n62;
    
    wire n20736;
    wire [17:0]modulation_deviation_amount_minus_sine_lookup_width_16__N_1638;
    
    wire n17923, n17922, n17921, n27284, n72, n22468, n17920, 
        n22467, n17919, n17918, n22453, n22452, n22441, n22440, 
        n78, n101, n22438, n79, n102, n22437, n82, n59_adj_3003, 
        n27272, n105, n8, n10, n39_adj_3004, n12, n47_adj_3005, 
        n74, n83, n60_adj_3006, n106, n48_adj_3007, n75, n21276, 
        n21278, n21280, n21266, n22435, n22434, n77, n85, n108, 
        n22429, n22428, n7, n9, n11, n13, n15, n22426, n22425, 
        n9093, n22423, n27105, n22422, n38_adj_3008, n42_adj_3009, 
        n22420, n22419, n22417, n22416, n22414, n22413, n22411, 
        n22410, n22408, n22407, n22405, n22404, n21691, n21690, 
        n21688, n21687, n21685, n25050, n21684, n21682, n21681, 
        n22540, n22539, n32_adj_3010, n71, n1, n33_adj_3011, n45_adj_3012, 
        n72_adj_3013, n2_c, n46_adj_3014, n21068, n21058, n22537, 
        n22536, n22534, n17917, n22533, n22531, n73_adj_3015, n104, 
        n22608, n135, n22530, n103, n134, n22528, n22527, n22522, 
        n22521, n22519, n22518, n17976, n17916, n22516, n22515, 
        n22513, n22512, n22510, n22509, n20994, n21008, n21006, 
        n22507, n17915, n22506, n20992, n20996, n17914, n22501, 
        n17913, n22500, n22492, n22491, n55_adj_3016, n27109, n56_adj_3017, 
        n27110, n27080, n52_adj_3018, n25, n27, n29, n17, n19, 
        n21, n23, n95_adj_3019, n27079, n27154, n49_adj_3020, n53_adj_3021, 
        n80, n57_adj_3022, n30, n88, n26, n28, n18, n20, n22, 
        n24, n17975, n17912, n96, n27078, n27283, n50_adj_3023, 
        n54_adj_3024, n81, n58_adj_3025, n89, n97, n113, n16, 
        n27092, n51_adj_3026, n98, n114, n99, n115, n76, n45_adj_3027, 
        n84, n27282, n100_adj_3028, n116, n17911, n46_adj_3029, 
        n27138, n17974, n17973, n17972, n132, n17971, n133, n136, 
        n137, n107, n123, n139, n17909, n9095, n70, n17908, 
        n17907, n17906, dac_clk_p_c_enable_432, n27082, n117, n118, 
        dac_clk_p_c_enable_486, n17905, n17904, n17903, n17902, cw;
    wire [15:0]quarter_wave_sample_register_q;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(22[56:86])
    
    FD1P3AX \addr_space_3[[30__281  (.D(wb_odata[30]), .SP(dac_clk_p_c_enable_149), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[30__281 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[29__283  (.D(wb_odata[29]), .SP(dac_clk_p_c_enable_149), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[29__283 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[28__285  (.D(wb_odata[28]), .SP(dac_clk_p_c_enable_149), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[28__285 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[27__287  (.D(wb_odata[27]), .SP(dac_clk_p_c_enable_149), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[27__287 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[26__289  (.D(wb_odata[26]), .SP(dac_clk_p_c_enable_149), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[26__289 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[25__291  (.D(wb_odata[25]), .SP(dac_clk_p_c_enable_149), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[25__291 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[30__182  (.D(wb_odata[30]), .SP(dac_clk_p_c_enable_116), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[30__182 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[29__183  (.D(wb_odata[29]), .SP(dac_clk_p_c_enable_116), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[29__183 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[28__184  (.D(wb_odata[28]), .SP(dac_clk_p_c_enable_116), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[28__184 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[27__185  (.D(wb_odata[27]), .SP(dac_clk_p_c_enable_116), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[27__185 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[25__188  (.D(wb_odata[25]), .SP(dac_clk_p_c_enable_116), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[25__188 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[24__189  (.D(wb_odata[24]), .SP(dac_clk_p_c_enable_116), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[24__189 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[23__190  (.D(wb_odata[23]), .SP(dac_clk_p_c_enable_116), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[23__190 .GSR = "DISABLED";
    FD1P3BX \addr_space_0[[22__191  (.D(wb_odata[22]), .SP(dac_clk_p_c_enable_116), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(\addr_space[0] [22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[22__191 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[21__192  (.D(wb_odata[21]), .SP(dac_clk_p_c_enable_116), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[21__192 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[20__193  (.D(wb_odata[20]), .SP(dac_clk_p_c_enable_116), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[20__193 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[19__194  (.D(wb_odata[19]), .SP(dac_clk_p_c_enable_116), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[19__194 .GSR = "DISABLED";
    FD1P3BX \addr_space_0[[18__195  (.D(wb_odata[18]), .SP(dac_clk_p_c_enable_116), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(\addr_space[0] [18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[18__195 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[17__196  (.D(wb_odata[17]), .SP(dac_clk_p_c_enable_116), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[17__196 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[16__197  (.D(wb_odata[16]), .SP(dac_clk_p_c_enable_116), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[16__197 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[15__198  (.D(wb_odata[15]), .SP(dac_clk_p_c_enable_116), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[15__198 .GSR = "DISABLED";
    FD1P3BX \addr_space_0[[14__199  (.D(wb_odata[14]), .SP(dac_clk_p_c_enable_116), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(\addr_space[0] [14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[14__199 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[13__200  (.D(wb_odata[13]), .SP(dac_clk_p_c_enable_116), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[13__200 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[12__201  (.D(wb_odata[12]), .SP(dac_clk_p_c_enable_116), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[12__201 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[11__202  (.D(wb_odata[11]), .SP(dac_clk_p_c_enable_116), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[11__202 .GSR = "DISABLED";
    FD1P3BX \addr_space_0[[10__203  (.D(wb_odata[10]), .SP(dac_clk_p_c_enable_116), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(\addr_space[0] [10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[10__203 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[9__204  (.D(wb_odata[9]), .SP(dac_clk_p_c_enable_116), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[9__204 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[8__205  (.D(wb_odata[8]), .SP(dac_clk_p_c_enable_116), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[8__205 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[7__206  (.D(wb_odata[7]), .SP(dac_clk_p_c_enable_116), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[7__206 .GSR = "DISABLED";
    FD1P3BX \addr_space_0[[6__207  (.D(wb_odata[6]), .SP(dac_clk_p_c_enable_116), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(\addr_space[0] [6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[6__207 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[5__208  (.D(wb_odata[5]), .SP(dac_clk_p_c_enable_116), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[5__208 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[4__209  (.D(wb_odata[4]), .SP(dac_clk_p_c_enable_116), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[4__209 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[3__210  (.D(wb_odata[3]), .SP(dac_clk_p_c_enable_116), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[3__210 .GSR = "DISABLED";
    FD1P3BX \addr_space_0[[2__211  (.D(wb_odata[2]), .SP(dac_clk_p_c_enable_116), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(\addr_space[0] [2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[2__211 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[1__212  (.D(wb_odata[1]), .SP(dac_clk_p_c_enable_116), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[1__212 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[0__213  (.D(wb_odata[0]), .SP(dac_clk_p_c_enable_116), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[0__213 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[31__214  (.D(wb_odata[31]), .SP(dac_clk_p_c_enable_73), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[1] [31])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[31__214 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[30__215  (.D(wb_odata[30]), .SP(dac_clk_p_c_enable_73), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[1] [30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[30__215 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[29__216  (.D(wb_odata[29]), .SP(dac_clk_p_c_enable_73), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[1] [29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[29__216 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[28__217  (.D(wb_odata[28]), .SP(dac_clk_p_c_enable_73), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[1] [28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[28__217 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[27__218  (.D(wb_odata[27]), .SP(dac_clk_p_c_enable_73), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[1] [27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[27__218 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[26__219  (.D(wb_odata[26]), .SP(dac_clk_p_c_enable_73), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[1] [26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[26__219 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[25__220  (.D(wb_odata[25]), .SP(dac_clk_p_c_enable_73), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[1] [25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[25__220 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[24__221  (.D(wb_odata[24]), .SP(dac_clk_p_c_enable_73), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[1] [24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[24__221 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[23__222  (.D(wb_odata[23]), .SP(dac_clk_p_c_enable_73), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[1] [23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[23__222 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[22__223  (.D(wb_odata[22]), .SP(dac_clk_p_c_enable_73), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[1] [22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[22__223 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[21__224  (.D(wb_odata[21]), .SP(dac_clk_p_c_enable_73), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[1] [21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[21__224 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[20__225  (.D(wb_odata[20]), .SP(dac_clk_p_c_enable_73), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[1] [20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[20__225 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[19__226  (.D(wb_odata[19]), .SP(dac_clk_p_c_enable_73), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[1] [19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[19__226 .GSR = "DISABLED";
    FD1P3BX \addr_space_1[[18__227  (.D(wb_odata[18]), .SP(dac_clk_p_c_enable_73), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(\addr_space[1] [18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[18__227 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[17__228  (.D(wb_odata[17]), .SP(dac_clk_p_c_enable_73), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[1] [17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[17__228 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[16__229  (.D(wb_odata[16]), .SP(dac_clk_p_c_enable_73), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[1] [16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[16__229 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[15__230  (.D(wb_odata[15]), .SP(dac_clk_p_c_enable_73), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[1] [15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[15__230 .GSR = "DISABLED";
    FD1P3BX \addr_space_1[[14__231  (.D(wb_odata[14]), .SP(dac_clk_p_c_enable_73), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(\addr_space[1] [14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[14__231 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[13__232  (.D(wb_odata[13]), .SP(dac_clk_p_c_enable_73), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[1] [13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[13__232 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[12__233  (.D(wb_odata[12]), .SP(dac_clk_p_c_enable_73), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[1] [12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[12__233 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[11__234  (.D(wb_odata[11]), .SP(dac_clk_p_c_enable_73), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[1] [11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[11__234 .GSR = "DISABLED";
    FD1P3BX \addr_space_1[[10__235  (.D(wb_odata[10]), .SP(dac_clk_p_c_enable_73), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(\addr_space[1] [10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[10__235 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[9__236  (.D(wb_odata[9]), .SP(dac_clk_p_c_enable_73), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[1] [9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[9__236 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[8__237  (.D(wb_odata[8]), .SP(dac_clk_p_c_enable_73), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[1] [8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[8__237 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[7__238  (.D(wb_odata[7]), .SP(dac_clk_p_c_enable_73), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[1] [7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[7__238 .GSR = "DISABLED";
    FD1P3BX \addr_space_1[[6__239  (.D(wb_odata[6]), .SP(dac_clk_p_c_enable_73), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(\addr_space[1] [6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[6__239 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[5__240  (.D(wb_odata[5]), .SP(dac_clk_p_c_enable_73), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[1] [5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[5__240 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[4__241  (.D(wb_odata[4]), .SP(dac_clk_p_c_enable_73), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[1] [4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[4__241 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[3__242  (.D(wb_odata[3]), .SP(dac_clk_p_c_enable_73), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[1] [3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[3__242 .GSR = "DISABLED";
    FD1P3BX \addr_space_1[[2__243  (.D(wb_odata[2]), .SP(dac_clk_p_c_enable_73), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(\addr_space[1] [2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[2__243 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[1__244  (.D(wb_odata[1]), .SP(dac_clk_p_c_enable_73), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[1] [1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[1__244 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[0__245  (.D(wb_odata[0]), .SP(dac_clk_p_c_enable_73), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[1] [0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[0__245 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[31__246  (.D(wb_odata[31]), .SP(dac_clk_p_c_enable_105), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[2] [31])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[31__246 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[30__247  (.D(wb_odata[30]), .SP(dac_clk_p_c_enable_105), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[2] [30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[30__247 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[29__248  (.D(wb_odata[29]), .SP(dac_clk_p_c_enable_105), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[2] [29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[29__248 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[28__249  (.D(wb_odata[28]), .SP(dac_clk_p_c_enable_105), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[2] [28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[28__249 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[27__250  (.D(wb_odata[27]), .SP(dac_clk_p_c_enable_105), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[2] [27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[27__250 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[26__251  (.D(wb_odata[26]), .SP(dac_clk_p_c_enable_105), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[2] [26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[26__251 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[25__252  (.D(wb_odata[25]), .SP(dac_clk_p_c_enable_105), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[2] [25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[25__252 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[24__253  (.D(wb_odata[24]), .SP(dac_clk_p_c_enable_105), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[2] [24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[24__253 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[23__254  (.D(wb_odata[23]), .SP(dac_clk_p_c_enable_105), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[2] [23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[23__254 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[22__255  (.D(wb_odata[22]), .SP(dac_clk_p_c_enable_105), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[2] [22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[22__255 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[21__256  (.D(wb_odata[21]), .SP(dac_clk_p_c_enable_105), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[2] [21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[21__256 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[20__257  (.D(wb_odata[20]), .SP(dac_clk_p_c_enable_105), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[2] [20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[20__257 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[19__258  (.D(wb_odata[19]), .SP(dac_clk_p_c_enable_105), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[2] [19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[19__258 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[18__259  (.D(wb_odata[18]), .SP(dac_clk_p_c_enable_105), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[2] [18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[18__259 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[17__260  (.D(wb_odata[17]), .SP(dac_clk_p_c_enable_105), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[2] [17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[17__260 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[16__261  (.D(wb_odata[16]), .SP(dac_clk_p_c_enable_105), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[2] [16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[16__261 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[15__262  (.D(wb_odata[15]), .SP(dac_clk_p_c_enable_105), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[2] [15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[15__262 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[14__263  (.D(wb_odata[14]), .SP(dac_clk_p_c_enable_105), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[2] [14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[14__263 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[13__264  (.D(wb_odata[13]), .SP(dac_clk_p_c_enable_105), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[2] [13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[13__264 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[12__265  (.D(wb_odata[12]), .SP(dac_clk_p_c_enable_105), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[2] [12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[12__265 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[11__266  (.D(wb_odata[11]), .SP(dac_clk_p_c_enable_105), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[2] [11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[11__266 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[10__267  (.D(wb_odata[10]), .SP(dac_clk_p_c_enable_105), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[2] [10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[10__267 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[9__268  (.D(wb_odata[9]), .SP(dac_clk_p_c_enable_105), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[2] [9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[9__268 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[8__269  (.D(wb_odata[8]), .SP(dac_clk_p_c_enable_105), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[2] [8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[8__269 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[7__270  (.D(wb_odata[7]), .SP(dac_clk_p_c_enable_105), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[2] [7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[7__270 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[6__271  (.D(wb_odata[6]), .SP(dac_clk_p_c_enable_105), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[2] [6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[6__271 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[5__272  (.D(wb_odata[5]), .SP(dac_clk_p_c_enable_105), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[2] [5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[5__272 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[4__273  (.D(wb_odata[4]), .SP(dac_clk_p_c_enable_105), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[2] [4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[4__273 .GSR = "DISABLED";
    FD1P3BX \addr_space_2[[3__274  (.D(wb_odata[3]), .SP(dac_clk_p_c_enable_105), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(\addr_space[2] [3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[3__274 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[2__275  (.D(wb_odata[2]), .SP(dac_clk_p_c_enable_105), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[2] [2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[2__275 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[1__276  (.D(wb_odata[1]), .SP(dac_clk_p_c_enable_105), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[2] [1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[1__276 .GSR = "DISABLED";
    FD1P3BX \addr_space_2[[0__277  (.D(wb_odata[0]), .SP(dac_clk_p_c_enable_105), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(\addr_space[2] [0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[0__277 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[24__293  (.D(wb_odata[24]), .SP(dac_clk_p_c_enable_149), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[24__293 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[23__295  (.D(wb_odata[23]), .SP(dac_clk_p_c_enable_149), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[23__295 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[22__297  (.D(wb_odata[22]), .SP(dac_clk_p_c_enable_149), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[22__297 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[21__299  (.D(wb_odata[21]), .SP(dac_clk_p_c_enable_149), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[21__299 .GSR = "DISABLED";
    FD1S3AX o_wb_data_i0 (.D(o_wb_data_31__N_1336[0]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i0.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_rs_i1 (.D(carrier_center_increment_offset_rs_30__N_1559[0]), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(carrier_center_increment_offset_rs[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_center_increment_offset_rs_i1.GSR = "DISABLED";
    FD1S3DX carrier_increment_i0 (.D(carrier_increment_30__N_1590[0]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_increment[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_increment_i0.GSR = "DISABLED";
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i0 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1621[0]), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(sine_lookup_width_minus_modulation_deviation_amount[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i0.GSR = "DISABLED";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i0 (.D(\addr_space[2] [0]), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(modulation_deviation_amount_minus_sine_lookup_width[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i0.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i0 (.D(n20732), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_center_increment_offset_ls[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_center_increment_offset_ls__i0.GSR = "DISABLED";
    FD1P3AX \addr_space_3[[20__301  (.D(wb_odata[20]), .SP(dac_clk_p_c_enable_149), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[20__301 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[31__181  (.D(wb_odata[31]), .SP(dac_clk_p_c_enable_116), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [31])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[31__181 .GSR = "DISABLED";
    FD1P3BX \addr_space_0[[26__187  (.D(wb_odata[26]), .SP(dac_clk_p_c_enable_116), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(\addr_space[0] [26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[26__187 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[19__303  (.D(wb_odata[19]), .SP(dac_clk_p_c_enable_149), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[19__303 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[18__305  (.D(wb_odata[18]), .SP(dac_clk_p_c_enable_149), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[18__305 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[17__307  (.D(wb_odata[17]), .SP(dac_clk_p_c_enable_149), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[17__307 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[16__309  (.D(wb_odata[16]), .SP(dac_clk_p_c_enable_149), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[16__309 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[15__311  (.D(wb_odata[15]), .SP(dac_clk_p_c_enable_149), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[15__311 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[14__313  (.D(wb_odata[14]), .SP(dac_clk_p_c_enable_149), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[14__313 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[13__315  (.D(wb_odata[13]), .SP(dac_clk_p_c_enable_149), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[13__315 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[12__317  (.D(wb_odata[12]), .SP(dac_clk_p_c_enable_149), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[12__317 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[11__319  (.D(wb_odata[11]), .SP(dac_clk_p_c_enable_149), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[11__319 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[10__321  (.D(wb_odata[10]), .SP(dac_clk_p_c_enable_149), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[10__321 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[9__323  (.D(wb_odata[9]), .SP(dac_clk_p_c_enable_149), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[9__323 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[8__325  (.D(wb_odata[8]), .SP(dac_clk_p_c_enable_149), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[8__325 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[7__327  (.D(wb_odata[7]), .SP(dac_clk_p_c_enable_149), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[7__327 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[6__329  (.D(wb_odata[6]), .SP(dac_clk_p_c_enable_149), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[6__329 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[5__331  (.D(wb_odata[5]), .SP(dac_clk_p_c_enable_149), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[5__331 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[4__333  (.D(wb_odata[4]), .SP(dac_clk_p_c_enable_149), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[4__333 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[3__335  (.D(wb_odata[3]), .SP(dac_clk_p_c_enable_149), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[3__335 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[2__337  (.D(wb_odata[2]), .SP(dac_clk_p_c_enable_149), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[2__337 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[1__339  (.D(wb_odata[1]), .SP(dac_clk_p_c_enable_149), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[1__339 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[0__341  (.D(wb_odata[0]), .SP(dac_clk_p_c_enable_149), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[0__341 .GSR = "DISABLED";
    LUT4 sub_437_inv_0_i1_1_lut (.A(\addr_space[2] [0]), .Z(sine_lookup_width_minus_modulation_deviation_amount_16__N_1621[0])) /* synthesis lut_function=(!(A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(96[58:109])
    defparam sub_437_inv_0_i1_1_lut.init = 16'h5555;
    FD1S3IX o_wb_ack_343 (.D(o_dac_a_9__N_1), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(wb_fm_ack)) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(54[8] 59[4])
    defparam o_wb_ack_343.GSR = "DISABLED";
    FD1S3BX startup_timer_FSM_i0_i0 (.D(n31[0]), .CK(dac_clk_p_c), .PD(i_sw0_c), 
            .Q(n1109[0]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(143[21:41])
    defparam startup_timer_FSM_i0_i0.GSR = "DISABLED";
    FD1P3AX \addr_space_3[[31__279  (.D(wb_odata[31]), .SP(dac_clk_p_c_enable_149), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [31])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[31__279 .GSR = "DISABLED";
    LUT4 i6715_2_lut_rep_456 (.A(sine_lookup_width_minus_modulation_deviation_amount[4]), 
         .B(n178), .Z(n27121)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(100[41:116])
    defparam i6715_2_lut_rep_456.init = 16'heeee;
    PFUMX i6718 (.BLUT(n69), .ALUT(n100), .C0(n22746), .Z(carrier_center_increment_offset_rs_30__N_1559[6]));
    LUT4 n25046_bdd_3_lut_4_lut (.A(sine_lookup_width_minus_modulation_deviation_amount[4]), 
         .B(n178), .C(modulation_output[15]), .D(n25046), .Z(carrier_center_increment_offset_rs_30__N_1559[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(100[41:116])
    defparam n25046_bdd_3_lut_4_lut.init = 16'hf1e0;
    FD1P3AX cw_mux_dac_a_mux_sel_351 (.D(cw_N_1877), .SP(dac_clk_p_c_enable_218), 
            .CK(dac_clk_p_c), .Q(cw_mux_dac_a_mux_sel)) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(133[11] 145[5])
    defparam cw_mux_dac_a_mux_sel_351.GSR = "DISABLED";
    LUT4 i1_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[6]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[15]), .C(modulation_deviation_amount_minus_sine_lookup_width[12]), 
         .D(modulation_deviation_amount_minus_sine_lookup_width[9]), .Z(n21208)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam i1_4_lut.init = 16'hfffe;
    LUT4 i23078_2_lut_2_lut_3_lut (.A(sine_lookup_width_minus_modulation_deviation_amount[4]), 
         .B(n178), .C(sine_lookup_width_minus_modulation_deviation_amount[3]), 
         .Z(n22746)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(100[41:116])
    defparam i23078_2_lut_2_lut_3_lut.init = 16'hfefe;
    PFUMX i6706 (.BLUT(n63), .ALUT(n94), .C0(n22774), .Z(carrier_center_increment_offset_rs_30__N_1559[0]));
    PFUMX i6708 (.BLUT(n64), .ALUT(n95), .C0(n22774), .Z(carrier_center_increment_offset_rs_30__N_1559[1]));
    LUT4 n25141_bdd_3_lut_4_lut (.A(sine_lookup_width_minus_modulation_deviation_amount[4]), 
         .B(n178), .C(modulation_output[15]), .D(n25141), .Z(carrier_center_increment_offset_rs_30__N_1559[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(100[41:116])
    defparam n25141_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n39_bdd_3_lut_23432 (.A(n43), .B(modulation_output[15]), .C(sine_lookup_width_minus_modulation_deviation_amount[2]), 
         .Z(n25039)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n39_bdd_3_lut_23432.init = 16'hcaca;
    LUT4 i1_4_lut_adj_91 (.A(n21206), .B(n21208), .C(n21210), .D(n21196), 
         .Z(n178_adj_2995)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam i1_4_lut_adj_91.init = 16'hfffe;
    LUT4 n25041_bdd_3_lut (.A(n25041), .B(n25039), .C(sine_lookup_width_minus_modulation_deviation_amount[3]), 
         .Z(n25042)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n25041_bdd_3_lut.init = 16'hcaca;
    LUT4 mux_434_Mux_1_i3_4_lut_4_lut_4_lut (.A(\wb_addr[0] ), .B(\wb_addr[1] ), 
         .C(\power_counter[1] ), .D(\smpl_register[1] ), .Z(n2122)) /* synthesis lut_function=(A (B (C)+!B (D))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(45[4:25])
    defparam mux_434_Mux_1_i3_4_lut_4_lut_4_lut.init = 16'hb391;
    LUT4 n36_bdd_3_lut_23435 (.A(n40), .B(sine_lookup_width_minus_modulation_deviation_amount[3]), 
         .C(modulation_output[15]), .Z(n25044)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n36_bdd_3_lut_23435.init = 16'he2e2;
    LUT4 n36_bdd_3_lut_25492 (.A(n36), .B(n44), .C(sine_lookup_width_minus_modulation_deviation_amount[3]), 
         .Z(n25045)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n36_bdd_3_lut_25492.init = 16'hcaca;
    LUT4 n37_bdd_4_lut_25070 (.A(n14), .B(modulation_output[15]), .C(sine_lookup_width_minus_modulation_deviation_amount[2]), 
         .D(sine_lookup_width_minus_modulation_deviation_amount[1]), .Z(n25048)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;
    defparam n37_bdd_4_lut_25070.init = 16'hccca;
    LUT4 n37_bdd_3_lut_25071 (.A(n37), .B(n41), .C(sine_lookup_width_minus_modulation_deviation_amount[2]), 
         .Z(n25049)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n37_bdd_3_lut_25071.init = 16'hcaca;
    PFUMX i20129 (.BLUT(n22482), .ALUT(n22483), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1336[18]));
    LUT4 i1_4_lut_adj_92 (.A(modulation_deviation_amount_minus_sine_lookup_width[5]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[16]), .C(modulation_deviation_amount_minus_sine_lookup_width[11]), 
         .D(modulation_deviation_amount_minus_sine_lookup_width[8]), .Z(n21210)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam i1_4_lut_adj_92.init = 16'hfffe;
    LUT4 i1_2_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[14]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[13]), .Z(n21206)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam i1_2_lut.init = 16'heeee;
    LUT4 n39_bdd_3_lut_25105 (.A(n4), .B(n6), .C(sine_lookup_width_minus_modulation_deviation_amount[1]), 
         .Z(n25040)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n39_bdd_3_lut_25105.init = 16'hcaca;
    LUT4 i12215_2_lut_3_lut_4_lut (.A(n27250), .B(modulation_deviation_amount_minus_sine_lookup_width[2]), 
         .C(modulation_output[0]), .D(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .Z(n124)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam i12215_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 i615_1_lut (.A(i_sw0_c), .Z(dac_clk_p_c_enable_488)) /* synthesis lut_function=(!(A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(31[12:17])
    defparam i615_1_lut.init = 16'h5555;
    LUT4 n38_bdd_3_lut_25023 (.A(n3), .B(n5), .C(sine_lookup_width_minus_modulation_deviation_amount[1]), 
         .Z(n25139)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n38_bdd_3_lut_25023.init = 16'hcaca;
    LUT4 n25140_bdd_3_lut (.A(n25140), .B(n73), .C(sine_lookup_width_minus_modulation_deviation_amount[3]), 
         .Z(n25141)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n25140_bdd_3_lut.init = 16'hcaca;
    CCU2D add_425_31 (.A0(\addr_space[0] [29]), .B0(n14676), .C0(carrier_center_increment_offset_rs[30]), 
          .D0(carrier_center_increment_offset_ls[29]), .A1(\addr_space[0] [30]), 
          .B1(n14676), .C1(carrier_center_increment_offset_rs[30]), .D1(carrier_center_increment_offset_ls[30]), 
          .CIN(n17925), .S0(carrier_increment_30__N_1590[29]), .S1(carrier_increment_30__N_1590[30]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(105[4:87])
    defparam add_425_31.INIT0 = 16'h569a;
    defparam add_425_31.INIT1 = 16'h569a;
    defparam add_425_31.INJECT1_0 = "NO";
    defparam add_425_31.INJECT1_1 = "NO";
    CCU2D add_425_29 (.A0(\addr_space[0] [27]), .B0(n14676), .C0(carrier_center_increment_offset_rs[30]), 
          .D0(carrier_center_increment_offset_ls[27]), .A1(\addr_space[0] [28]), 
          .B1(n14676), .C1(carrier_center_increment_offset_rs[30]), .D1(carrier_center_increment_offset_ls[28]), 
          .CIN(n17924), .COUT(n17925), .S0(carrier_increment_30__N_1590[27]), 
          .S1(carrier_increment_30__N_1590[28]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(105[4:87])
    defparam add_425_29.INIT0 = 16'h569a;
    defparam add_425_29.INIT1 = 16'h569a;
    defparam add_425_29.INJECT1_0 = "NO";
    defparam add_425_29.INJECT1_1 = "NO";
    LUT4 i1_2_lut_adj_93 (.A(modulation_deviation_amount_minus_sine_lookup_width[7]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[10]), .Z(n21196)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam i1_2_lut_adj_93.init = 16'heeee;
    LUT4 i6482_2_lut (.A(n1109[0]), .B(n61[15]), .Z(n31[0])) /* synthesis lut_function=(A (B)) */ ;
    defparam i6482_2_lut.init = 16'h8888;
    FD1S3DX carrier_center_increment_offset_ls__i30 (.D(n62[30]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_center_increment_offset_ls[30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_center_increment_offset_ls__i30.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i29 (.D(n62[29]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_center_increment_offset_ls[29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_center_increment_offset_ls__i29.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i28 (.D(n62[28]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_center_increment_offset_ls[28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_center_increment_offset_ls__i28.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i27 (.D(n62[27]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_center_increment_offset_ls[27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_center_increment_offset_ls__i27.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i26 (.D(n62[26]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_center_increment_offset_ls[26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_center_increment_offset_ls__i26.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i25 (.D(n62[25]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_center_increment_offset_ls[25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_center_increment_offset_ls__i25.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i24 (.D(n62[24]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_center_increment_offset_ls[24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_center_increment_offset_ls__i24.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i23 (.D(n62[23]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_center_increment_offset_ls[23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_center_increment_offset_ls__i23.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i22 (.D(n62[22]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_center_increment_offset_ls[22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_center_increment_offset_ls__i22.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i21 (.D(n62[21]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_center_increment_offset_ls[21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_center_increment_offset_ls__i21.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i20 (.D(n62[20]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_center_increment_offset_ls[20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_center_increment_offset_ls__i20.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i19 (.D(n62[19]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_center_increment_offset_ls[19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_center_increment_offset_ls__i19.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i18 (.D(n62[18]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_center_increment_offset_ls[18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_center_increment_offset_ls__i18.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i17 (.D(n62[17]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_center_increment_offset_ls[17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_center_increment_offset_ls__i17.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i16 (.D(n62[16]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_center_increment_offset_ls[16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_center_increment_offset_ls__i16.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i15 (.D(n62[15]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_center_increment_offset_ls[15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_center_increment_offset_ls__i15.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i14 (.D(n62[14]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_center_increment_offset_ls[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_center_increment_offset_ls__i14.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i13 (.D(n62[13]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_center_increment_offset_ls[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_center_increment_offset_ls__i13.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i12 (.D(n62[12]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_center_increment_offset_ls[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_center_increment_offset_ls__i12.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i11 (.D(n62[11]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_center_increment_offset_ls[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_center_increment_offset_ls__i11.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i10 (.D(n62[10]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_center_increment_offset_ls[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_center_increment_offset_ls__i10.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i9 (.D(n62[9]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_center_increment_offset_ls[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_center_increment_offset_ls__i9.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i8 (.D(n62[8]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_center_increment_offset_ls[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_center_increment_offset_ls__i8.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i7 (.D(n62[7]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_center_increment_offset_ls[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_center_increment_offset_ls__i7.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i6 (.D(n62[6]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_center_increment_offset_ls[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_center_increment_offset_ls__i6.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i5 (.D(n62[5]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_center_increment_offset_ls[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_center_increment_offset_ls__i5.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i4 (.D(n62[4]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_center_increment_offset_ls[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_center_increment_offset_ls__i4.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i3 (.D(n62[3]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_center_increment_offset_ls[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_center_increment_offset_ls__i3.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i2 (.D(n62[2]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_center_increment_offset_ls[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_center_increment_offset_ls__i2.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i1 (.D(n20736), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_center_increment_offset_ls[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_center_increment_offset_ls__i1.GSR = "DISABLED";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i16 (.D(modulation_deviation_amount_minus_sine_lookup_width_16__N_1638[16]), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(modulation_deviation_amount_minus_sine_lookup_width[16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i16.GSR = "DISABLED";
    CCU2D add_425_27 (.A0(\addr_space[0] [25]), .B0(n14676), .C0(carrier_center_increment_offset_rs[30]), 
          .D0(carrier_center_increment_offset_ls[25]), .A1(\addr_space[0] [26]), 
          .B1(n14676), .C1(carrier_center_increment_offset_rs[30]), .D1(carrier_center_increment_offset_ls[26]), 
          .CIN(n17923), .COUT(n17924), .S0(carrier_increment_30__N_1590[25]), 
          .S1(carrier_increment_30__N_1590[26]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(105[4:87])
    defparam add_425_27.INIT0 = 16'h569a;
    defparam add_425_27.INIT1 = 16'h569a;
    defparam add_425_27.INJECT1_0 = "NO";
    defparam add_425_27.INJECT1_1 = "NO";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i15 (.D(modulation_deviation_amount_minus_sine_lookup_width_16__N_1638[15]), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(modulation_deviation_amount_minus_sine_lookup_width[15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i15.GSR = "DISABLED";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i14 (.D(modulation_deviation_amount_minus_sine_lookup_width_16__N_1638[14]), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(modulation_deviation_amount_minus_sine_lookup_width[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i14.GSR = "DISABLED";
    CCU2D add_425_25 (.A0(\addr_space[0] [23]), .B0(n14676), .C0(carrier_center_increment_offset_rs[30]), 
          .D0(carrier_center_increment_offset_ls[23]), .A1(\addr_space[0] [24]), 
          .B1(n14676), .C1(carrier_center_increment_offset_rs[30]), .D1(carrier_center_increment_offset_ls[24]), 
          .CIN(n17922), .COUT(n17923), .S0(carrier_increment_30__N_1590[23]), 
          .S1(carrier_increment_30__N_1590[24]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(105[4:87])
    defparam add_425_25.INIT0 = 16'h569a;
    defparam add_425_25.INIT1 = 16'h569a;
    defparam add_425_25.INJECT1_0 = "NO";
    defparam add_425_25.INJECT1_1 = "NO";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i13 (.D(modulation_deviation_amount_minus_sine_lookup_width_16__N_1638[13]), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(modulation_deviation_amount_minus_sine_lookup_width[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i13.GSR = "DISABLED";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i12 (.D(modulation_deviation_amount_minus_sine_lookup_width_16__N_1638[12]), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(modulation_deviation_amount_minus_sine_lookup_width[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i12.GSR = "DISABLED";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i11 (.D(modulation_deviation_amount_minus_sine_lookup_width_16__N_1638[11]), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(modulation_deviation_amount_minus_sine_lookup_width[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i11.GSR = "DISABLED";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i10 (.D(modulation_deviation_amount_minus_sine_lookup_width_16__N_1638[10]), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(modulation_deviation_amount_minus_sine_lookup_width[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i10.GSR = "DISABLED";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i9 (.D(modulation_deviation_amount_minus_sine_lookup_width_16__N_1638[9]), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(modulation_deviation_amount_minus_sine_lookup_width[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i9.GSR = "DISABLED";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i8 (.D(modulation_deviation_amount_minus_sine_lookup_width_16__N_1638[8]), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(modulation_deviation_amount_minus_sine_lookup_width[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i8.GSR = "DISABLED";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i7 (.D(modulation_deviation_amount_minus_sine_lookup_width_16__N_1638[7]), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(modulation_deviation_amount_minus_sine_lookup_width[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i7.GSR = "DISABLED";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i6 (.D(modulation_deviation_amount_minus_sine_lookup_width_16__N_1638[6]), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(modulation_deviation_amount_minus_sine_lookup_width[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i6.GSR = "DISABLED";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i5 (.D(modulation_deviation_amount_minus_sine_lookup_width_16__N_1638[5]), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(modulation_deviation_amount_minus_sine_lookup_width[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i5.GSR = "DISABLED";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i4 (.D(modulation_deviation_amount_minus_sine_lookup_width_16__N_1638[4]), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(modulation_deviation_amount_minus_sine_lookup_width[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i4.GSR = "DISABLED";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i3 (.D(\addr_space[2] [3]), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(modulation_deviation_amount_minus_sine_lookup_width[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i3.GSR = "DISABLED";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i2 (.D(\addr_space[2] [2]), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(modulation_deviation_amount_minus_sine_lookup_width[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i2.GSR = "DISABLED";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i1 (.D(\addr_space[2] [1]), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(modulation_deviation_amount_minus_sine_lookup_width[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i1.GSR = "DISABLED";
    CCU2D add_425_23 (.A0(\addr_space[0] [21]), .B0(n14676), .C0(carrier_center_increment_offset_rs[30]), 
          .D0(carrier_center_increment_offset_ls[21]), .A1(\addr_space[0] [22]), 
          .B1(n14676), .C1(carrier_center_increment_offset_rs[30]), .D1(carrier_center_increment_offset_ls[22]), 
          .CIN(n17921), .COUT(n17922), .S0(carrier_increment_30__N_1590[21]), 
          .S1(carrier_increment_30__N_1590[22]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(105[4:87])
    defparam add_425_23.INIT0 = 16'h569a;
    defparam add_425_23.INIT1 = 16'h569a;
    defparam add_425_23.INJECT1_0 = "NO";
    defparam add_425_23.INJECT1_1 = "NO";
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i16 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1621[16]), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(sine_lookup_width_minus_modulation_deviation_amount[16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i16.GSR = "DISABLED";
    LUT4 i6627_3_lut_4_lut (.A(n27284), .B(modulation_deviation_amount_minus_sine_lookup_width[2]), 
         .C(modulation_output[14]), .D(modulation_output[15]), .Z(n72)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam i6627_3_lut_4_lut.init = 16'hf780;
    LUT4 i20113_3_lut (.A(\addr_space[2] [19]), .B(\addr_space[3] [19]), 
         .C(\wb_addr[0] ), .Z(n22468)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20113_3_lut.init = 16'hcaca;
    CCU2D add_425_21 (.A0(\addr_space[0] [19]), .B0(n14676), .C0(carrier_center_increment_offset_rs[30]), 
          .D0(carrier_center_increment_offset_ls[19]), .A1(\addr_space[0] [20]), 
          .B1(n14676), .C1(carrier_center_increment_offset_rs[30]), .D1(carrier_center_increment_offset_ls[20]), 
          .CIN(n17920), .COUT(n17921), .S0(carrier_increment_30__N_1590[19]), 
          .S1(carrier_increment_30__N_1590[20]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(105[4:87])
    defparam add_425_21.INIT0 = 16'h569a;
    defparam add_425_21.INIT1 = 16'h569a;
    defparam add_425_21.INJECT1_0 = "NO";
    defparam add_425_21.INJECT1_1 = "NO";
    LUT4 i20112_3_lut (.A(\addr_space[0] [19]), .B(\addr_space[1] [19]), 
         .C(\wb_addr[0] ), .Z(n22467)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20112_3_lut.init = 16'hcaca;
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i15 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1621[15]), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(sine_lookup_width_minus_modulation_deviation_amount[15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i15.GSR = "DISABLED";
    CCU2D add_425_19 (.A0(\addr_space[0] [17]), .B0(n14676), .C0(carrier_center_increment_offset_rs[30]), 
          .D0(carrier_center_increment_offset_ls[17]), .A1(\addr_space[0] [18]), 
          .B1(n14676), .C1(carrier_center_increment_offset_rs[30]), .D1(carrier_center_increment_offset_ls[18]), 
          .CIN(n17919), .COUT(n17920), .S0(carrier_increment_30__N_1590[17]), 
          .S1(carrier_increment_30__N_1590[18]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(105[4:87])
    defparam add_425_19.INIT0 = 16'h569a;
    defparam add_425_19.INIT1 = 16'h569a;
    defparam add_425_19.INJECT1_0 = "NO";
    defparam add_425_19.INJECT1_1 = "NO";
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i14 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1621[14]), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(sine_lookup_width_minus_modulation_deviation_amount[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i14.GSR = "DISABLED";
    CCU2D add_425_17 (.A0(\addr_space[0] [15]), .B0(n14676), .C0(carrier_center_increment_offset_rs[30]), 
          .D0(carrier_center_increment_offset_ls[15]), .A1(\addr_space[0] [16]), 
          .B1(n14676), .C1(carrier_center_increment_offset_rs[30]), .D1(carrier_center_increment_offset_ls[16]), 
          .CIN(n17918), .COUT(n17919), .S0(carrier_increment_30__N_1590[15]), 
          .S1(carrier_increment_30__N_1590[16]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(105[4:87])
    defparam add_425_17.INIT0 = 16'h569a;
    defparam add_425_17.INIT1 = 16'h569a;
    defparam add_425_17.INJECT1_0 = "NO";
    defparam add_425_17.INJECT1_1 = "NO";
    LUT4 i20098_3_lut (.A(\addr_space[2] [20]), .B(\addr_space[3] [20]), 
         .C(\wb_addr[0] ), .Z(n22453)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20098_3_lut.init = 16'hcaca;
    LUT4 i20097_3_lut (.A(\addr_space[0] [20]), .B(\addr_space[1] [20]), 
         .C(\wb_addr[0] ), .Z(n22452)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20097_3_lut.init = 16'hcaca;
    LUT4 i20086_3_lut (.A(\addr_space[2] [21]), .B(\addr_space[3] [21]), 
         .C(\wb_addr[0] ), .Z(n22441)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20086_3_lut.init = 16'hcaca;
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i13 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1621[13]), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(sine_lookup_width_minus_modulation_deviation_amount[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i13.GSR = "DISABLED";
    LUT4 i20085_3_lut (.A(\addr_space[0] [21]), .B(\addr_space[1] [21]), 
         .C(\wb_addr[0] ), .Z(n22440)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20085_3_lut.init = 16'hcaca;
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i12 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1621[12]), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(sine_lookup_width_minus_modulation_deviation_amount[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i12.GSR = "DISABLED";
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i11 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1621[11]), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(sine_lookup_width_minus_modulation_deviation_amount[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i11.GSR = "DISABLED";
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i10 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1621[10]), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(sine_lookup_width_minus_modulation_deviation_amount[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i10.GSR = "DISABLED";
    LUT4 modulation_output_15__I_0_355_i101_3_lut (.A(modulation_output[15]), 
         .B(n78), .C(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .Z(n101)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_355_i101_3_lut.init = 16'hcaca;
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i9 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1621[9]), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(sine_lookup_width_minus_modulation_deviation_amount[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i9.GSR = "DISABLED";
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i8 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1621[8]), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(sine_lookup_width_minus_modulation_deviation_amount[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i8.GSR = "DISABLED";
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i7 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1621[7]), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(sine_lookup_width_minus_modulation_deviation_amount[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i7.GSR = "DISABLED";
    LUT4 i20083_3_lut (.A(\addr_space[2] [22]), .B(\addr_space[3] [22]), 
         .C(\wb_addr[0] ), .Z(n22438)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20083_3_lut.init = 16'hcaca;
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i6 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1621[6]), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(sine_lookup_width_minus_modulation_deviation_amount[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i6.GSR = "DISABLED";
    LUT4 modulation_output_15__I_0_i4_3_lut (.A(modulation_output[3]), .B(modulation_output[4]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[0]), .Z(n4)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(100[41:116])
    defparam modulation_output_15__I_0_i4_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i6_3_lut (.A(modulation_output[5]), .B(modulation_output[6]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[0]), .Z(n6)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(100[41:116])
    defparam modulation_output_15__I_0_i6_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_355_i102_3_lut (.A(modulation_output[15]), 
         .B(n79), .C(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .Z(n102)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_355_i102_3_lut.init = 16'hcaca;
    LUT4 i20082_3_lut (.A(\addr_space[0] [22]), .B(\addr_space[1] [22]), 
         .C(\wb_addr[0] ), .Z(n22437)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20082_3_lut.init = 16'hcaca;
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i5 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1621[5]), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(sine_lookup_width_minus_modulation_deviation_amount[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i5.GSR = "DISABLED";
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i4 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1621[4]), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(sine_lookup_width_minus_modulation_deviation_amount[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i4.GSR = "DISABLED";
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i3 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1621[3]), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(sine_lookup_width_minus_modulation_deviation_amount[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i3.GSR = "DISABLED";
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i2 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1621[2]), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(sine_lookup_width_minus_modulation_deviation_amount[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i2.GSR = "DISABLED";
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i1 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1621[1]), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(sine_lookup_width_minus_modulation_deviation_amount[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i1.GSR = "DISABLED";
    LUT4 modulation_output_15__I_0_355_i105_4_lut (.A(n82), .B(n59_adj_3003), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[4]), .D(n27272), 
         .Z(n105)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_355_i105_4_lut.init = 16'hca0a;
    FD1S3DX carrier_increment_i30 (.D(carrier_increment_30__N_1590[30]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_increment[30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_increment_i30.GSR = "DISABLED";
    FD1S3DX carrier_increment_i29 (.D(carrier_increment_30__N_1590[29]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_increment[29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_increment_i29.GSR = "DISABLED";
    LUT4 modulation_output_15__I_0_i39_3_lut (.A(n8), .B(n10), .C(sine_lookup_width_minus_modulation_deviation_amount[1]), 
         .Z(n39_adj_3004)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(100[41:116])
    defparam modulation_output_15__I_0_i39_3_lut.init = 16'hcaca;
    FD1S3DX carrier_increment_i28 (.D(carrier_increment_30__N_1590[28]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_increment[28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_increment_i28.GSR = "DISABLED";
    LUT4 modulation_output_15__I_0_i43_3_lut (.A(n12), .B(n14), .C(sine_lookup_width_minus_modulation_deviation_amount[1]), 
         .Z(n43)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(100[41:116])
    defparam modulation_output_15__I_0_i43_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_355_i74_3_lut (.A(modulation_output[15]), 
         .B(n47_adj_3005), .C(modulation_deviation_amount_minus_sine_lookup_width[2]), 
         .Z(n74)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_355_i74_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i8_3_lut (.A(modulation_output[7]), .B(modulation_output[8]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[0]), .Z(n8)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(100[41:116])
    defparam modulation_output_15__I_0_i8_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i10_3_lut (.A(modulation_output[9]), .B(modulation_output[10]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[0]), .Z(n10)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(100[41:116])
    defparam modulation_output_15__I_0_i10_3_lut.init = 16'hcaca;
    FD1S3DX carrier_increment_i27 (.D(carrier_increment_30__N_1590[27]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_increment[27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_increment_i27.GSR = "DISABLED";
    FD1S3DX carrier_increment_i26 (.D(carrier_increment_30__N_1590[26]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_increment[26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_increment_i26.GSR = "DISABLED";
    FD1S3DX carrier_increment_i25 (.D(carrier_increment_30__N_1590[25]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_increment[25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_increment_i25.GSR = "DISABLED";
    LUT4 modulation_output_15__I_0_355_i106_4_lut (.A(n83), .B(n60_adj_3006), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[4]), .D(n27272), 
         .Z(n106)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_355_i106_4_lut.init = 16'hca0a;
    FD1S3DX carrier_increment_i24 (.D(carrier_increment_30__N_1590[24]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_increment[24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_increment_i24.GSR = "DISABLED";
    FD1S3DX carrier_increment_i23 (.D(carrier_increment_30__N_1590[23]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_increment[23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_increment_i23.GSR = "DISABLED";
    FD1S3DX carrier_increment_i22 (.D(carrier_increment_30__N_1590[22]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_increment[22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_increment_i22.GSR = "DISABLED";
    FD1S3DX carrier_increment_i21 (.D(carrier_increment_30__N_1590[21]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_increment[21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_increment_i21.GSR = "DISABLED";
    FD1S3DX carrier_increment_i20 (.D(carrier_increment_30__N_1590[20]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_increment[20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_increment_i20.GSR = "DISABLED";
    FD1S3DX carrier_increment_i19 (.D(carrier_increment_30__N_1590[19]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_increment[19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_increment_i19.GSR = "DISABLED";
    FD1S3DX carrier_increment_i18 (.D(carrier_increment_30__N_1590[18]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_increment[18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_increment_i18.GSR = "DISABLED";
    FD1S3DX carrier_increment_i17 (.D(carrier_increment_30__N_1590[17]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_increment[17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_increment_i17.GSR = "DISABLED";
    FD1S3DX carrier_increment_i16 (.D(carrier_increment_30__N_1590[16]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_increment[16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_increment_i16.GSR = "DISABLED";
    LUT4 modulation_output_15__I_0_i12_3_lut (.A(modulation_output[11]), .B(modulation_output[12]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[0]), .Z(n12)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(100[41:116])
    defparam modulation_output_15__I_0_i12_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i14_3_lut (.A(modulation_output[13]), .B(modulation_output[14]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[0]), .Z(n14)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(100[41:116])
    defparam modulation_output_15__I_0_i14_3_lut.init = 16'hcaca;
    FD1S3DX carrier_increment_i15 (.D(carrier_increment_30__N_1590[15]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_increment[15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_increment_i15.GSR = "DISABLED";
    FD1S3DX carrier_increment_i14 (.D(carrier_increment_30__N_1590[14]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_increment[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_increment_i14.GSR = "DISABLED";
    FD1S3DX carrier_increment_i13 (.D(carrier_increment_30__N_1590[13]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_increment[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_increment_i13.GSR = "DISABLED";
    FD1S3DX carrier_increment_i12 (.D(carrier_increment_30__N_1590[12]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_increment[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_increment_i12.GSR = "DISABLED";
    FD1S3DX carrier_increment_i11 (.D(carrier_increment_30__N_1590[11]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_increment[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_increment_i11.GSR = "DISABLED";
    LUT4 modulation_output_15__I_0_355_i75_3_lut (.A(modulation_output[15]), 
         .B(n48_adj_3007), .C(modulation_deviation_amount_minus_sine_lookup_width[2]), 
         .Z(n75)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_355_i75_3_lut.init = 16'hcaca;
    FD1S3DX carrier_increment_i10 (.D(carrier_increment_30__N_1590[10]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_increment[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_increment_i10.GSR = "DISABLED";
    FD1S3DX carrier_increment_i9 (.D(carrier_increment_30__N_1590[9]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_increment[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_increment_i9.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_94 (.A(n21276), .B(n21278), .C(n21280), .D(n21266), 
         .Z(n178)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(100[41:116])
    defparam i1_4_lut_adj_94.init = 16'hfffe;
    LUT4 i1_2_lut_adj_95 (.A(sine_lookup_width_minus_modulation_deviation_amount[14]), 
         .B(sine_lookup_width_minus_modulation_deviation_amount[5]), .Z(n21276)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(100[41:116])
    defparam i1_2_lut_adj_95.init = 16'heeee;
    FD1S3DX carrier_increment_i8 (.D(carrier_increment_30__N_1590[8]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_increment[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_increment_i8.GSR = "DISABLED";
    FD1S3DX carrier_increment_i7 (.D(carrier_increment_30__N_1590[7]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_increment[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_increment_i7.GSR = "DISABLED";
    LUT4 i20080_3_lut (.A(\addr_space[2] [23]), .B(\addr_space[3] [23]), 
         .C(\wb_addr[0] ), .Z(n22435)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20080_3_lut.init = 16'hcaca;
    LUT4 i20079_3_lut (.A(\addr_space[0] [23]), .B(\addr_space[1] [23]), 
         .C(\wb_addr[0] ), .Z(n22434)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20079_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_96 (.A(sine_lookup_width_minus_modulation_deviation_amount[6]), 
         .B(sine_lookup_width_minus_modulation_deviation_amount[15]), .C(sine_lookup_width_minus_modulation_deviation_amount[16]), 
         .D(sine_lookup_width_minus_modulation_deviation_amount[9]), .Z(n21278)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(100[41:116])
    defparam i1_4_lut_adj_96.init = 16'hfffe;
    LUT4 i1_4_lut_adj_97 (.A(sine_lookup_width_minus_modulation_deviation_amount[12]), 
         .B(sine_lookup_width_minus_modulation_deviation_amount[8]), .C(sine_lookup_width_minus_modulation_deviation_amount[11]), 
         .D(sine_lookup_width_minus_modulation_deviation_amount[13]), .Z(n21280)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(100[41:116])
    defparam i1_4_lut_adj_97.init = 16'hfffe;
    FD1S3DX carrier_increment_i6 (.D(carrier_increment_30__N_1590[6]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_increment[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_increment_i6.GSR = "DISABLED";
    LUT4 i1_2_lut_adj_98 (.A(sine_lookup_width_minus_modulation_deviation_amount[7]), 
         .B(sine_lookup_width_minus_modulation_deviation_amount[10]), .Z(n21266)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(100[41:116])
    defparam i1_2_lut_adj_98.init = 16'heeee;
    LUT4 modulation_output_15__I_0_355_i108_3_lut (.A(n77), .B(n85), .C(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .Z(n108)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_355_i108_3_lut.init = 16'hcaca;
    FD1S3DX carrier_increment_i5 (.D(carrier_increment_30__N_1590[5]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_increment[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_increment_i5.GSR = "DISABLED";
    FD1S3DX carrier_increment_i4 (.D(carrier_increment_30__N_1590[4]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_increment[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_increment_i4.GSR = "DISABLED";
    LUT4 i20074_3_lut (.A(\addr_space[2] [24]), .B(\addr_space[3] [24]), 
         .C(\wb_addr[0] ), .Z(n22429)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20074_3_lut.init = 16'hcaca;
    LUT4 i20073_3_lut (.A(\addr_space[0] [24]), .B(\addr_space[1] [24]), 
         .C(\wb_addr[0] ), .Z(n22428)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20073_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i36_3_lut (.A(n5), .B(n7), .C(sine_lookup_width_minus_modulation_deviation_amount[1]), 
         .Z(n36)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(100[41:116])
    defparam modulation_output_15__I_0_i36_3_lut.init = 16'hcaca;
    FD1S3DX carrier_increment_i3 (.D(carrier_increment_30__N_1590[3]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_increment[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_increment_i3.GSR = "DISABLED";
    FD1S3DX carrier_increment_i2 (.D(carrier_increment_30__N_1590[2]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_increment[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_increment_i2.GSR = "DISABLED";
    LUT4 modulation_output_15__I_0_i40_3_lut (.A(n9), .B(n11), .C(sine_lookup_width_minus_modulation_deviation_amount[1]), 
         .Z(n40)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(100[41:116])
    defparam modulation_output_15__I_0_i40_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i9_3_lut (.A(modulation_output[8]), .B(modulation_output[9]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[0]), .Z(n9)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(100[41:116])
    defparam modulation_output_15__I_0_i9_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i11_3_lut (.A(modulation_output[10]), .B(modulation_output[11]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[0]), .Z(n11)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(100[41:116])
    defparam modulation_output_15__I_0_i11_3_lut.init = 16'hcaca;
    FD1S3DX carrier_increment_i1 (.D(carrier_increment_30__N_1590[1]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_increment[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_increment_i1.GSR = "DISABLED";
    LUT4 modulation_output_15__I_0_i5_3_lut (.A(modulation_output[4]), .B(modulation_output[5]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[0]), .Z(n5)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(100[41:116])
    defparam modulation_output_15__I_0_i5_3_lut.init = 16'hcaca;
    FD1S3DX carrier_center_increment_offset_rs_i16 (.D(modulation_output[15]), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(carrier_center_increment_offset_rs[30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_center_increment_offset_rs_i16.GSR = "DISABLED";
    LUT4 modulation_output_15__I_0_i7_3_lut (.A(modulation_output[6]), .B(modulation_output[7]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[0]), .Z(n7)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(100[41:116])
    defparam modulation_output_15__I_0_i7_3_lut.init = 16'hcaca;
    FD1S3DX carrier_center_increment_offset_rs_i15 (.D(carrier_center_increment_offset_rs_30__N_1559[14]), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(carrier_center_increment_offset_rs[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_center_increment_offset_rs_i15.GSR = "DISABLED";
    LUT4 modulation_output_15__I_0_i44_3_lut (.A(n13), .B(n15), .C(sine_lookup_width_minus_modulation_deviation_amount[1]), 
         .Z(n44)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(100[41:116])
    defparam modulation_output_15__I_0_i44_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i15_3_lut (.A(modulation_output[14]), .B(modulation_output[15]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[0]), .Z(n15)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(100[41:116])
    defparam modulation_output_15__I_0_i15_3_lut.init = 16'hcaca;
    FD1S3DX carrier_center_increment_offset_rs_i14 (.D(carrier_center_increment_offset_rs_30__N_1559[13]), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(carrier_center_increment_offset_rs[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_center_increment_offset_rs_i14.GSR = "DISABLED";
    LUT4 modulation_output_15__I_0_i13_3_lut (.A(modulation_output[12]), .B(modulation_output[13]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[0]), .Z(n13)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(100[41:116])
    defparam modulation_output_15__I_0_i13_3_lut.init = 16'hcaca;
    LUT4 i20071_3_lut (.A(\addr_space[2] [25]), .B(\addr_space[3] [25]), 
         .C(\wb_addr[0] ), .Z(n22426)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20071_3_lut.init = 16'hcaca;
    FD1S3DX carrier_center_increment_offset_rs_i13 (.D(carrier_center_increment_offset_rs_30__N_1559[12]), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(carrier_center_increment_offset_rs[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_center_increment_offset_rs_i13.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_rs_i12 (.D(carrier_center_increment_offset_rs_30__N_1559[11]), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(carrier_center_increment_offset_rs[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_center_increment_offset_rs_i12.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_rs_i11 (.D(carrier_center_increment_offset_rs_30__N_1559[10]), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(carrier_center_increment_offset_rs[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_center_increment_offset_rs_i11.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_rs_i10 (.D(carrier_center_increment_offset_rs_30__N_1559[9]), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(carrier_center_increment_offset_rs[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_center_increment_offset_rs_i10.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_rs_i9 (.D(carrier_center_increment_offset_rs_30__N_1559[8]), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(carrier_center_increment_offset_rs[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_center_increment_offset_rs_i9.GSR = "DISABLED";
    LUT4 i20070_3_lut (.A(\addr_space[0] [25]), .B(\addr_space[1] [25]), 
         .C(\wb_addr[0] ), .Z(n22425)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20070_3_lut.init = 16'hcaca;
    FD1S3DX carrier_center_increment_offset_rs_i8 (.D(carrier_center_increment_offset_rs_30__N_1559[7]), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(carrier_center_increment_offset_rs[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_center_increment_offset_rs_i8.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_rs_i7 (.D(carrier_center_increment_offset_rs_30__N_1559[6]), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(carrier_center_increment_offset_rs[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_center_increment_offset_rs_i7.GSR = "DISABLED";
    LUT4 modulation_output_15__I_0_i37_3_lut (.A(n6), .B(n8), .C(sine_lookup_width_minus_modulation_deviation_amount[1]), 
         .Z(n37)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(100[41:116])
    defparam modulation_output_15__I_0_i37_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i41_3_lut (.A(n10), .B(n12), .C(sine_lookup_width_minus_modulation_deviation_amount[1]), 
         .Z(n41)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(100[41:116])
    defparam modulation_output_15__I_0_i41_3_lut.init = 16'hcaca;
    FD1S3DX carrier_center_increment_offset_rs_i6 (.D(carrier_center_increment_offset_rs_30__N_1559[5]), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(carrier_center_increment_offset_rs[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_center_increment_offset_rs_i6.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_rs_i5 (.D(carrier_center_increment_offset_rs_30__N_1559[4]), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(carrier_center_increment_offset_rs[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_center_increment_offset_rs_i5.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_rs_i4 (.D(carrier_center_increment_offset_rs_30__N_1559[3]), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(carrier_center_increment_offset_rs[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_center_increment_offset_rs_i4.GSR = "DISABLED";
    LUT4 i6672_2_lut (.A(sine_lookup_width_minus_modulation_deviation_amount[1]), 
         .B(sine_lookup_width_minus_modulation_deviation_amount[2]), .Z(n9093)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(100[41:116])
    defparam i6672_2_lut.init = 16'heeee;
    FD1S3DX carrier_center_increment_offset_rs_i3 (.D(carrier_center_increment_offset_rs_30__N_1559[2]), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(carrier_center_increment_offset_rs[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_center_increment_offset_rs_i3.GSR = "DISABLED";
    LUT4 i20068_3_lut (.A(\addr_space[2] [26]), .B(\addr_space[3] [26]), 
         .C(\wb_addr[0] ), .Z(n22423)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20068_3_lut.init = 16'hcaca;
    FD1S3DX carrier_center_increment_offset_rs_i2 (.D(carrier_center_increment_offset_rs_30__N_1559[1]), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(carrier_center_increment_offset_rs[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam carrier_center_increment_offset_rs_i2.GSR = "DISABLED";
    LUT4 i1_3_lut_rep_440 (.A(sine_lookup_width_minus_modulation_deviation_amount[3]), 
         .B(n178), .C(sine_lookup_width_minus_modulation_deviation_amount[4]), 
         .Z(n27105)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(100[41:116])
    defparam i1_3_lut_rep_440.init = 16'hfefe;
    LUT4 i20067_3_lut (.A(\addr_space[0] [26]), .B(\addr_space[1] [26]), 
         .C(\wb_addr[0] ), .Z(n22422)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20067_3_lut.init = 16'hcaca;
    FD1S3AX o_wb_data_i31 (.D(o_wb_data_31__N_1336[31]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[31])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i31.GSR = "DISABLED";
    LUT4 modulation_output_15__I_0_i38_3_lut (.A(n7), .B(n9), .C(sine_lookup_width_minus_modulation_deviation_amount[1]), 
         .Z(n38_adj_3008)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(100[41:116])
    defparam modulation_output_15__I_0_i38_3_lut.init = 16'hcaca;
    FD1S3AX o_wb_data_i30 (.D(o_wb_data_31__N_1336[30]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i30.GSR = "DISABLED";
    FD1S3AX o_wb_data_i29 (.D(o_wb_data_31__N_1336[29]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i29.GSR = "DISABLED";
    FD1S3AX o_wb_data_i28 (.D(o_wb_data_31__N_1336[28]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i28.GSR = "DISABLED";
    LUT4 modulation_output_15__I_0_i42_3_lut (.A(n11), .B(n13), .C(sine_lookup_width_minus_modulation_deviation_amount[1]), 
         .Z(n42_adj_3009)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(100[41:116])
    defparam modulation_output_15__I_0_i42_3_lut.init = 16'hcaca;
    FD1S3AX o_wb_data_i27 (.D(o_wb_data_31__N_1336[27]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i27.GSR = "DISABLED";
    LUT4 i20065_3_lut (.A(\addr_space[2] [27]), .B(\addr_space[3] [27]), 
         .C(\wb_addr[0] ), .Z(n22420)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20065_3_lut.init = 16'hcaca;
    FD1S3AX o_wb_data_i26 (.D(o_wb_data_31__N_1336[26]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i26.GSR = "DISABLED";
    FD1S3AX o_wb_data_i25 (.D(o_wb_data_31__N_1336[25]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i25.GSR = "DISABLED";
    FD1S3AX o_wb_data_i24 (.D(o_wb_data_31__N_1336[24]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i24.GSR = "DISABLED";
    FD1S3AX o_wb_data_i23 (.D(o_wb_data_31__N_1336[23]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i23.GSR = "DISABLED";
    FD1S3AX o_wb_data_i22 (.D(o_wb_data_31__N_1336[22]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i22.GSR = "DISABLED";
    FD1S3AX o_wb_data_i21 (.D(o_wb_data_31__N_1336[21]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i21.GSR = "DISABLED";
    FD1S3AX o_wb_data_i20 (.D(o_wb_data_31__N_1336[20]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i20.GSR = "DISABLED";
    FD1S3AX o_wb_data_i19 (.D(o_wb_data_31__N_1336[19]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i19.GSR = "DISABLED";
    FD1S3AX o_wb_data_i18 (.D(o_wb_data_31__N_1336[18]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i18.GSR = "DISABLED";
    FD1S3AX o_wb_data_i17 (.D(o_wb_data_31__N_1336[17]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i17.GSR = "DISABLED";
    FD1S3AX o_wb_data_i16 (.D(o_wb_data_31__N_1336[16]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i16.GSR = "DISABLED";
    FD1S3AX o_wb_data_i15 (.D(o_wb_data_31__N_1336[15]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i15.GSR = "DISABLED";
    LUT4 i20064_3_lut (.A(\addr_space[0] [27]), .B(\addr_space[1] [27]), 
         .C(\wb_addr[0] ), .Z(n22419)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20064_3_lut.init = 16'hcaca;
    FD1S3AX o_wb_data_i14 (.D(o_wb_data_31__N_1336[14]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i14.GSR = "DISABLED";
    FD1S3AX o_wb_data_i13 (.D(o_wb_data_31__N_1336[13]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i13.GSR = "DISABLED";
    FD1S3AX o_wb_data_i12 (.D(o_wb_data_31__N_1336[12]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i12.GSR = "DISABLED";
    FD1S3AX o_wb_data_i11 (.D(o_wb_data_31__N_1336[11]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i11.GSR = "DISABLED";
    LUT4 i20062_3_lut (.A(\addr_space[2] [28]), .B(\addr_space[3] [28]), 
         .C(\wb_addr[0] ), .Z(n22417)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20062_3_lut.init = 16'hcaca;
    LUT4 i20061_3_lut (.A(\addr_space[0] [28]), .B(\addr_space[1] [28]), 
         .C(\wb_addr[0] ), .Z(n22416)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20061_3_lut.init = 16'hcaca;
    LUT4 i20059_3_lut (.A(\addr_space[2] [29]), .B(\addr_space[3] [29]), 
         .C(\wb_addr[0] ), .Z(n22414)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20059_3_lut.init = 16'hcaca;
    LUT4 i20058_3_lut (.A(\addr_space[0] [29]), .B(\addr_space[1] [29]), 
         .C(\wb_addr[0] ), .Z(n22413)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20058_3_lut.init = 16'hcaca;
    LUT4 i20056_3_lut (.A(\addr_space[2] [30]), .B(\addr_space[3] [30]), 
         .C(\wb_addr[0] ), .Z(n22411)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20056_3_lut.init = 16'hcaca;
    LUT4 i20055_3_lut (.A(\addr_space[0] [30]), .B(\addr_space[1] [30]), 
         .C(\wb_addr[0] ), .Z(n22410)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20055_3_lut.init = 16'hcaca;
    FD1S3AX o_wb_data_i10 (.D(o_wb_data_31__N_1336[10]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i10.GSR = "DISABLED";
    LUT4 i20053_3_lut (.A(\addr_space[2] [31]), .B(\addr_space[3] [31]), 
         .C(\wb_addr[0] ), .Z(n22408)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20053_3_lut.init = 16'hcaca;
    LUT4 i20052_3_lut (.A(\addr_space[0] [31]), .B(\addr_space[1] [31]), 
         .C(\wb_addr[0] ), .Z(n22407)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20052_3_lut.init = 16'hcaca;
    FD1S3AX o_wb_data_i9 (.D(o_wb_data_31__N_1336[9]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i9.GSR = "DISABLED";
    FD1S3AX o_wb_data_i8 (.D(o_wb_data_31__N_1336[8]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i8.GSR = "DISABLED";
    FD1S3AX o_wb_data_i7 (.D(o_wb_data_31__N_1336[7]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i7.GSR = "DISABLED";
    FD1S3AX o_wb_data_i6 (.D(o_wb_data_31__N_1336[6]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i6.GSR = "DISABLED";
    LUT4 i20050_3_lut (.A(\addr_space[2] [0]), .B(\addr_space[3] [0]), .C(\wb_addr[0] ), 
         .Z(n22405)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20050_3_lut.init = 16'hcaca;
    FD1S3AX o_wb_data_i5 (.D(o_wb_data_31__N_1336[5]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i5.GSR = "DISABLED";
    LUT4 i20049_3_lut (.A(\addr_space[0] [0]), .B(\addr_space[1] [0]), .C(\wb_addr[0] ), 
         .Z(n22404)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20049_3_lut.init = 16'hcaca;
    FD1S3AX o_wb_data_i4 (.D(o_wb_data_31__N_1336[4]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i4.GSR = "DISABLED";
    FD1S3AX o_wb_data_i3 (.D(o_wb_data_31__N_1336[3]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i3.GSR = "DISABLED";
    FD1S3AX o_wb_data_i2 (.D(o_wb_data_31__N_1336[2]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i2.GSR = "DISABLED";
    LUT4 i19336_3_lut (.A(\addr_space[2] [1]), .B(\addr_space[3] [1]), .C(\wb_addr[0] ), 
         .Z(n21691)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19336_3_lut.init = 16'hcaca;
    FD1S3AX o_wb_data_i1 (.D(o_wb_data_31__N_1336[1]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i1.GSR = "DISABLED";
    LUT4 i19335_3_lut (.A(\addr_space[0] [1]), .B(\addr_space[1] [1]), .C(\wb_addr[0] ), 
         .Z(n21690)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19335_3_lut.init = 16'hcaca;
    LUT4 i19333_3_lut (.A(\addr_space[2] [2]), .B(\addr_space[3] [2]), .C(\wb_addr[0] ), 
         .Z(n21688)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19333_3_lut.init = 16'hcaca;
    LUT4 i23050_4_lut (.A(n61[15]), .B(i_sw0_c), .C(cw_N_1877), .D(n61[10]), 
         .Z(dac_clk_p_c_enable_218)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C)))) */ ;
    defparam i23050_4_lut.init = 16'h3032;
    LUT4 i19332_3_lut (.A(\addr_space[0] [2]), .B(\addr_space[1] [2]), .C(\wb_addr[0] ), 
         .Z(n21687)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19332_3_lut.init = 16'hcaca;
    LUT4 i19330_3_lut (.A(\addr_space[2] [3]), .B(\addr_space[3] [3]), .C(\wb_addr[0] ), 
         .Z(n21685)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19330_3_lut.init = 16'hcaca;
    LUT4 n25050_bdd_3_lut_4_lut (.A(sine_lookup_width_minus_modulation_deviation_amount[4]), 
         .B(n178), .C(modulation_output[15]), .D(n25050), .Z(carrier_center_increment_offset_rs_30__N_1559[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(100[41:116])
    defparam n25050_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i19329_3_lut (.A(\addr_space[0] [3]), .B(\addr_space[1] [3]), .C(\wb_addr[0] ), 
         .Z(n21684)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19329_3_lut.init = 16'hcaca;
    LUT4 i19327_3_lut (.A(\addr_space[2] [4]), .B(\addr_space[3] [4]), .C(\wb_addr[0] ), 
         .Z(n21682)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19327_3_lut.init = 16'hcaca;
    LUT4 i19326_3_lut (.A(\addr_space[0] [4]), .B(\addr_space[1] [4]), .C(\wb_addr[0] ), 
         .Z(n21681)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19326_3_lut.init = 16'hcaca;
    LUT4 i20185_3_lut (.A(\addr_space[2] [5]), .B(\addr_space[3] [5]), .C(\wb_addr[0] ), 
         .Z(n22540)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20185_3_lut.init = 16'hcaca;
    LUT4 i20184_3_lut (.A(\addr_space[0] [5]), .B(\addr_space[1] [5]), .C(\wb_addr[0] ), 
         .Z(n22539)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20184_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i32_3_lut (.A(n3), .B(n36), .C(sine_lookup_width_minus_modulation_deviation_amount[2]), 
         .Z(n32_adj_3010)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(100[41:116])
    defparam modulation_output_15__I_0_i32_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i71_3_lut (.A(n40), .B(n44), .C(sine_lookup_width_minus_modulation_deviation_amount[2]), 
         .Z(n71)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(100[41:116])
    defparam modulation_output_15__I_0_i71_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i3_3_lut (.A(modulation_output[2]), .B(modulation_output[3]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[0]), .Z(n3)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(100[41:116])
    defparam modulation_output_15__I_0_i3_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i1_3_lut (.A(modulation_output[0]), .B(modulation_output[1]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[0]), .Z(n1)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(100[41:116])
    defparam modulation_output_15__I_0_i1_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i33_3_lut (.A(n4), .B(n37), .C(sine_lookup_width_minus_modulation_deviation_amount[2]), 
         .Z(n33_adj_3011)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(100[41:116])
    defparam modulation_output_15__I_0_i33_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i72_3_lut (.A(n41), .B(n45_adj_3012), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[2]), .Z(n72_adj_3013)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(100[41:116])
    defparam modulation_output_15__I_0_i72_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i45_3_lut (.A(n14), .B(modulation_output[15]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[1]), .Z(n45_adj_3012)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(100[41:116])
    defparam modulation_output_15__I_0_i45_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i2_3_lut (.A(modulation_output[1]), .B(modulation_output[2]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[0]), .Z(n2_c)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(100[41:116])
    defparam modulation_output_15__I_0_i2_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i73_3_lut (.A(n42_adj_3009), .B(n46_adj_3014), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[2]), .Z(n73)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(100[41:116])
    defparam modulation_output_15__I_0_i73_3_lut.init = 16'hcaca;
    LUT4 i23171_4_lut (.A(n21068), .B(n27114), .C(n27304), .D(\wb_addr[0] ), 
         .Z(dac_clk_p_c_enable_149)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i23171_4_lut.init = 16'h1000;
    LUT4 i1_4_lut_adj_99 (.A(n27313), .B(\wb_addr[1] ), .C(\wb_addr[15] ), 
         .D(n21058), .Z(n21068)) /* synthesis lut_function=(A+(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_99.init = 16'hffbf;
    LUT4 i1_3_lut (.A(\wb_addr[8] ), .B(\wb_addr[12] ), .C(i_sw0_c), .Z(n21058)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_3_lut.init = 16'hfefe;
    LUT4 i20182_3_lut (.A(\addr_space[2] [6]), .B(\addr_space[3] [6]), .C(\wb_addr[0] ), 
         .Z(n22537)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20182_3_lut.init = 16'hcaca;
    LUT4 i20181_3_lut (.A(\addr_space[0] [6]), .B(\addr_space[1] [6]), .C(\wb_addr[0] ), 
         .Z(n22536)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20181_3_lut.init = 16'hcaca;
    LUT4 i20179_3_lut (.A(\addr_space[2] [7]), .B(\addr_space[3] [7]), .C(\wb_addr[0] ), 
         .Z(n22534)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20179_3_lut.init = 16'hcaca;
    CCU2D add_425_15 (.A0(\addr_space[0] [13]), .B0(n14676), .C0(carrier_center_increment_offset_rs[13]), 
          .D0(carrier_center_increment_offset_ls[13]), .A1(\addr_space[0] [14]), 
          .B1(n14676), .C1(carrier_center_increment_offset_rs[14]), .D1(carrier_center_increment_offset_ls[14]), 
          .CIN(n17917), .COUT(n17918), .S0(carrier_increment_30__N_1590[13]), 
          .S1(carrier_increment_30__N_1590[14]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(105[4:87])
    defparam add_425_15.INIT0 = 16'h569a;
    defparam add_425_15.INIT1 = 16'h569a;
    defparam add_425_15.INJECT1_0 = "NO";
    defparam add_425_15.INJECT1_1 = "NO";
    LUT4 i20178_3_lut (.A(\addr_space[0] [7]), .B(\addr_space[1] [7]), .C(\wb_addr[0] ), 
         .Z(n22533)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20178_3_lut.init = 16'hcaca;
    LUT4 i20176_3_lut (.A(\addr_space[2] [8]), .B(\addr_space[3] [8]), .C(\wb_addr[0] ), 
         .Z(n22531)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20176_3_lut.init = 16'hcaca;
    LUT4 i6730_3_lut_4_lut (.A(sine_lookup_width_minus_modulation_deviation_amount[2]), 
         .B(n27105), .C(modulation_output[15]), .D(n44), .Z(carrier_center_increment_offset_rs_30__N_1559[12])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(100[41:116])
    defparam i6730_3_lut_4_lut.init = 16'hf1e0;
    PFUMX modulation_output_15__I_0_355_i135 (.BLUT(n73_adj_3015), .ALUT(n104), 
          .C0(n22608), .Z(n135)) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;
    LUT4 i20175_3_lut (.A(\addr_space[0] [8]), .B(\addr_space[1] [8]), .C(\wb_addr[0] ), 
         .Z(n22530)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20175_3_lut.init = 16'hcaca;
    PFUMX modulation_output_15__I_0_355_i134 (.BLUT(n72), .ALUT(n103), .C0(n22608), 
          .Z(n134)) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;
    LUT4 i20173_3_lut (.A(\addr_space[2] [9]), .B(\addr_space[3] [9]), .C(\wb_addr[0] ), 
         .Z(n22528)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20173_3_lut.init = 16'hcaca;
    LUT4 n25042_bdd_3_lut_4_lut (.A(sine_lookup_width_minus_modulation_deviation_amount[4]), 
         .B(n178), .C(modulation_output[15]), .D(n25042), .Z(carrier_center_increment_offset_rs_30__N_1559[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(100[41:116])
    defparam n25042_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i6728_3_lut_4_lut (.A(sine_lookup_width_minus_modulation_deviation_amount[2]), 
         .B(n27105), .C(modulation_output[15]), .D(n43), .Z(carrier_center_increment_offset_rs_30__N_1559[11])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(100[41:116])
    defparam i6728_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i20172_3_lut (.A(\addr_space[0] [9]), .B(\addr_space[1] [9]), .C(\wb_addr[0] ), 
         .Z(n22527)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20172_3_lut.init = 16'hcaca;
    LUT4 i20167_3_lut (.A(\addr_space[2] [10]), .B(\addr_space[3] [10]), 
         .C(\wb_addr[0] ), .Z(n22522)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20167_3_lut.init = 16'hcaca;
    LUT4 i20166_3_lut (.A(\addr_space[0] [10]), .B(\addr_space[1] [10]), 
         .C(\wb_addr[0] ), .Z(n22521)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20166_3_lut.init = 16'hcaca;
    LUT4 i20164_3_lut (.A(\addr_space[2] [11]), .B(\addr_space[3] [11]), 
         .C(\wb_addr[0] ), .Z(n22519)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20164_3_lut.init = 16'hcaca;
    LUT4 i20163_3_lut (.A(\addr_space[0] [11]), .B(\addr_space[1] [11]), 
         .C(\wb_addr[0] ), .Z(n22518)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20163_3_lut.init = 16'hcaca;
    CCU2D sub_106_add_2_13 (.A0(\addr_space[2] [15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\addr_space[2] [16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17976), .S0(modulation_deviation_amount_minus_sine_lookup_width_16__N_1638[15]), 
          .S1(modulation_deviation_amount_minus_sine_lookup_width_16__N_1638[16]));
    defparam sub_106_add_2_13.INIT0 = 16'h5555;
    defparam sub_106_add_2_13.INIT1 = 16'h5555;
    defparam sub_106_add_2_13.INJECT1_0 = "NO";
    defparam sub_106_add_2_13.INJECT1_1 = "NO";
    CCU2D add_425_13 (.A0(\addr_space[0] [11]), .B0(n14676), .C0(carrier_center_increment_offset_rs[11]), 
          .D0(carrier_center_increment_offset_ls[11]), .A1(\addr_space[0] [12]), 
          .B1(n14676), .C1(carrier_center_increment_offset_rs[12]), .D1(carrier_center_increment_offset_ls[12]), 
          .CIN(n17916), .COUT(n17917), .S0(carrier_increment_30__N_1590[11]), 
          .S1(carrier_increment_30__N_1590[12]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(105[4:87])
    defparam add_425_13.INIT0 = 16'h569a;
    defparam add_425_13.INIT1 = 16'h569a;
    defparam add_425_13.INJECT1_0 = "NO";
    defparam add_425_13.INJECT1_1 = "NO";
    LUT4 i20161_3_lut (.A(\addr_space[2] [12]), .B(\addr_space[3] [12]), 
         .C(\wb_addr[0] ), .Z(n22516)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20161_3_lut.init = 16'hcaca;
    LUT4 i20160_3_lut (.A(\addr_space[0] [12]), .B(\addr_space[1] [12]), 
         .C(\wb_addr[0] ), .Z(n22515)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20160_3_lut.init = 16'hcaca;
    LUT4 i20158_3_lut (.A(\addr_space[2] [13]), .B(\addr_space[3] [13]), 
         .C(\wb_addr[0] ), .Z(n22513)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20158_3_lut.init = 16'hcaca;
    LUT4 i20157_3_lut (.A(\addr_space[0] [13]), .B(\addr_space[1] [13]), 
         .C(\wb_addr[0] ), .Z(n22512)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20157_3_lut.init = 16'hcaca;
    LUT4 i20155_3_lut (.A(\addr_space[2] [14]), .B(\addr_space[3] [14]), 
         .C(\wb_addr[0] ), .Z(n22510)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20155_3_lut.init = 16'hcaca;
    LUT4 i20154_3_lut (.A(\addr_space[0] [14]), .B(\addr_space[1] [14]), 
         .C(\wb_addr[0] ), .Z(n22509)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20154_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_100 (.A(n20994), .B(n21008), .C(n21006), .D(\addr_space[2] [4]), 
         .Z(n14676)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_100.init = 16'hfffe;
    LUT4 i20152_3_lut (.A(\addr_space[2] [15]), .B(\addr_space[3] [15]), 
         .C(\wb_addr[0] ), .Z(n22507)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20152_3_lut.init = 16'hcaca;
    CCU2D add_425_11 (.A0(\addr_space[0] [9]), .B0(n14676), .C0(carrier_center_increment_offset_rs[9]), 
          .D0(carrier_center_increment_offset_ls[9]), .A1(\addr_space[0] [10]), 
          .B1(n14676), .C1(carrier_center_increment_offset_rs[10]), .D1(carrier_center_increment_offset_ls[10]), 
          .CIN(n17915), .COUT(n17916), .S0(carrier_increment_30__N_1590[9]), 
          .S1(carrier_increment_30__N_1590[10]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(105[4:87])
    defparam add_425_11.INIT0 = 16'h569a;
    defparam add_425_11.INIT1 = 16'h569a;
    defparam add_425_11.INJECT1_0 = "NO";
    defparam add_425_11.INJECT1_1 = "NO";
    LUT4 i20151_3_lut (.A(\addr_space[0] [15]), .B(\addr_space[1] [15]), 
         .C(\wb_addr[0] ), .Z(n22506)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20151_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_101 (.A(\addr_space[2] [11]), .B(\addr_space[2] [14]), 
         .Z(n20994)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_101.init = 16'heeee;
    LUT4 i1_4_lut_adj_102 (.A(\addr_space[2] [12]), .B(n20992), .C(n20996), 
         .D(\addr_space[2] [13]), .Z(n21008)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_102.init = 16'hfffe;
    LUT4 i1_4_lut_adj_103 (.A(\addr_space[2] [15]), .B(\addr_space[2] [8]), 
         .C(\addr_space[2] [6]), .D(\addr_space[2] [7]), .Z(n21006)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_103.init = 16'hfffe;
    LUT4 i1_2_lut_adj_104 (.A(\addr_space[2] [5]), .B(\addr_space[2] [10]), 
         .Z(n20992)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_104.init = 16'heeee;
    LUT4 i1_2_lut_adj_105 (.A(\addr_space[2] [9]), .B(\addr_space[2] [16]), 
         .Z(n20996)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_105.init = 16'heeee;
    CCU2D add_425_9 (.A0(\addr_space[0] [7]), .B0(n14676), .C0(carrier_center_increment_offset_rs[7]), 
          .D0(carrier_center_increment_offset_ls[7]), .A1(\addr_space[0] [8]), 
          .B1(n14676), .C1(carrier_center_increment_offset_rs[8]), .D1(carrier_center_increment_offset_ls[8]), 
          .CIN(n17914), .COUT(n17915), .S0(carrier_increment_30__N_1590[7]), 
          .S1(carrier_increment_30__N_1590[8]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(105[4:87])
    defparam add_425_9.INIT0 = 16'h569a;
    defparam add_425_9.INIT1 = 16'h569a;
    defparam add_425_9.INJECT1_0 = "NO";
    defparam add_425_9.INJECT1_1 = "NO";
    LUT4 i20146_3_lut (.A(\addr_space[2] [16]), .B(\addr_space[3] [16]), 
         .C(\wb_addr[0] ), .Z(n22501)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20146_3_lut.init = 16'hcaca;
    CCU2D add_425_7 (.A0(\addr_space[0] [5]), .B0(n14676), .C0(carrier_center_increment_offset_rs[5]), 
          .D0(carrier_center_increment_offset_ls[5]), .A1(\addr_space[0] [6]), 
          .B1(n14676), .C1(carrier_center_increment_offset_rs[6]), .D1(carrier_center_increment_offset_ls[6]), 
          .CIN(n17913), .COUT(n17914), .S0(carrier_increment_30__N_1590[5]), 
          .S1(carrier_increment_30__N_1590[6]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(105[4:87])
    defparam add_425_7.INIT0 = 16'h569a;
    defparam add_425_7.INIT1 = 16'h569a;
    defparam add_425_7.INJECT1_0 = "NO";
    defparam add_425_7.INJECT1_1 = "NO";
    LUT4 i20145_3_lut (.A(\addr_space[0] [16]), .B(\addr_space[1] [16]), 
         .C(\wb_addr[0] ), .Z(n22500)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20145_3_lut.init = 16'hcaca;
    LUT4 i20137_3_lut (.A(\addr_space[2] [17]), .B(\addr_space[3] [17]), 
         .C(\wb_addr[0] ), .Z(n22492)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20137_3_lut.init = 16'hcaca;
    LUT4 i20136_3_lut (.A(\addr_space[0] [17]), .B(\addr_space[1] [17]), 
         .C(\wb_addr[0] ), .Z(n22491)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20136_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_355_i86_3_lut_rep_444 (.A(n55_adj_3016), 
         .B(n59_adj_3003), .C(modulation_deviation_amount_minus_sine_lookup_width[2]), 
         .Z(n27109)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_355_i86_3_lut_rep_444.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_355_i87_3_lut_rep_445 (.A(n56_adj_3017), 
         .B(n60_adj_3006), .C(modulation_deviation_amount_minus_sine_lookup_width[2]), 
         .Z(n27110)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_355_i87_3_lut_rep_445.init = 16'hcaca;
    LUT4 i11326_4_lut (.A(modulation_output[15]), .B(n178_adj_2995), .C(n27080), 
         .D(modulation_deviation_amount_minus_sine_lookup_width[4]), .Z(n62[30])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam i11326_4_lut.init = 16'h3022;
    LUT4 modulation_output_15__I_0_355_i79_3_lut (.A(n48_adj_3007), .B(n52_adj_3018), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[2]), .Z(n79)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_355_i79_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_355_i56_3_lut (.A(n25), .B(n27), .C(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .Z(n56_adj_3017)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_355_i56_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_355_i60_4_lut (.A(n29), .B(modulation_output[0]), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[1]), .D(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .Z(n60_adj_3006)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_355_i60_4_lut.init = 16'h0aca;
    LUT4 modulation_output_15__I_0_355_i29_3_lut (.A(modulation_output[2]), 
         .B(modulation_output[1]), .C(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .Z(n29)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_355_i29_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_355_i48_3_lut (.A(n17), .B(n19), .C(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .Z(n48_adj_3007)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_355_i48_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_355_i52_3_lut (.A(n21), .B(n23), .C(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .Z(n52_adj_3018)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_355_i52_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_355_i21_3_lut (.A(modulation_output[10]), 
         .B(modulation_output[9]), .C(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .Z(n21)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_355_i21_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_355_i23_3_lut (.A(modulation_output[8]), 
         .B(modulation_output[7]), .C(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .Z(n23)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_355_i23_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_355_i17_3_lut (.A(modulation_output[14]), 
         .B(modulation_output[13]), .C(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .Z(n17)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_355_i17_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_355_i19_3_lut (.A(modulation_output[12]), 
         .B(modulation_output[11]), .C(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .Z(n19)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_355_i19_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_355_i25_3_lut (.A(modulation_output[6]), 
         .B(modulation_output[5]), .C(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .Z(n25)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_355_i25_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_355_i27_3_lut (.A(modulation_output[4]), 
         .B(modulation_output[3]), .C(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .Z(n27)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_355_i27_3_lut.init = 16'hcaca;
    LUT4 i11328_4_lut (.A(n95_adj_3019), .B(n178_adj_2995), .C(n27079), 
         .D(modulation_deviation_amount_minus_sine_lookup_width[4]), .Z(n62[29])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam i11328_4_lut.init = 16'h3022;
    LUT4 i6635_4_lut (.A(modulation_output[15]), .B(modulation_output[14]), 
         .C(n27154), .D(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .Z(n95_adj_3019)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C (D)))) */ ;
    defparam i6635_4_lut.init = 16'hcaaa;
    LUT4 modulation_output_15__I_0_355_i80_3_lut (.A(n49_adj_3020), .B(n53_adj_3021), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[2]), .Z(n80)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_355_i80_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_355_i88_4_lut (.A(n57_adj_3022), .B(n30), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[2]), .D(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .Z(n88)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_355_i88_4_lut.init = 16'h0aca;
    LUT4 modulation_output_15__I_0_355_i57_3_lut (.A(n26), .B(n28), .C(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .Z(n57_adj_3022)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_355_i57_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_355_i30_3_lut (.A(modulation_output[1]), 
         .B(modulation_output[0]), .C(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .Z(n30)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_355_i30_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_355_i26_3_lut (.A(modulation_output[5]), 
         .B(modulation_output[4]), .C(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .Z(n26)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_355_i26_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_355_i28_3_lut (.A(modulation_output[3]), 
         .B(modulation_output[2]), .C(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .Z(n28)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_355_i28_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_355_i49_3_lut (.A(n18), .B(n20), .C(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .Z(n49_adj_3020)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_355_i49_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_355_i53_3_lut (.A(n22), .B(n24), .C(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .Z(n53_adj_3021)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_355_i53_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_355_i22_3_lut (.A(modulation_output[9]), 
         .B(modulation_output[8]), .C(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .Z(n22)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_355_i22_3_lut.init = 16'hcaca;
    LUT4 i11794_2_lut (.A(o_sample_i[14]), .B(cw_mux_dac_a_mux_sel), .Z(o_dac_a_c_7)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(29[18:140])
    defparam i11794_2_lut.init = 16'h2222;
    LUT4 modulation_output_15__I_0_355_i24_3_lut (.A(modulation_output[7]), 
         .B(modulation_output[6]), .C(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .Z(n24)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_355_i24_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_355_i18_3_lut (.A(modulation_output[13]), 
         .B(modulation_output[12]), .C(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .Z(n18)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_355_i18_3_lut.init = 16'hcaca;
    CCU2D sub_106_add_2_11 (.A0(\addr_space[2] [13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\addr_space[2] [14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17975), .COUT(n17976), .S0(modulation_deviation_amount_minus_sine_lookup_width_16__N_1638[13]), 
          .S1(modulation_deviation_amount_minus_sine_lookup_width_16__N_1638[14]));
    defparam sub_106_add_2_11.INIT0 = 16'h5555;
    defparam sub_106_add_2_11.INIT1 = 16'h5555;
    defparam sub_106_add_2_11.INJECT1_0 = "NO";
    defparam sub_106_add_2_11.INJECT1_1 = "NO";
    CCU2D add_425_5 (.A0(\addr_space[0] [3]), .B0(n14676), .C0(carrier_center_increment_offset_rs[3]), 
          .D0(carrier_center_increment_offset_ls[3]), .A1(\addr_space[0] [4]), 
          .B1(n14676), .C1(carrier_center_increment_offset_rs[4]), .D1(carrier_center_increment_offset_ls[4]), 
          .CIN(n17912), .COUT(n17913), .S0(carrier_increment_30__N_1590[3]), 
          .S1(carrier_increment_30__N_1590[4]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(105[4:87])
    defparam add_425_5.INIT0 = 16'h569a;
    defparam add_425_5.INIT1 = 16'h569a;
    defparam add_425_5.INJECT1_0 = "NO";
    defparam add_425_5.INJECT1_1 = "NO";
    LUT4 modulation_output_15__I_0_355_i20_3_lut (.A(modulation_output[11]), 
         .B(modulation_output[10]), .C(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .Z(n20)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_355_i20_3_lut.init = 16'hcaca;
    LUT4 i11346_4_lut (.A(n96), .B(n178_adj_2995), .C(n27078), .D(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .Z(n62[28])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam i11346_4_lut.init = 16'h3022;
    LUT4 i6637_4_lut (.A(modulation_output[15]), .B(n17), .C(n27283), 
         .D(modulation_deviation_amount_minus_sine_lookup_width[3]), .Z(n96)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C (D)))) */ ;
    defparam i6637_4_lut.init = 16'hcaaa;
    LUT4 modulation_output_15__I_0_355_i81_3_lut (.A(n50_adj_3023), .B(n54_adj_3024), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[2]), .Z(n81)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_355_i81_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_355_i89_4_lut (.A(n58_adj_3025), .B(modulation_output[0]), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[2]), .D(n27250), 
         .Z(n89)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_355_i89_4_lut.init = 16'h0aca;
    LUT4 modulation_output_15__I_0_355_i50_3_lut (.A(n19), .B(n21), .C(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .Z(n50_adj_3023)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_355_i50_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_355_i54_3_lut (.A(n23), .B(n25), .C(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .Z(n54_adj_3024)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_355_i54_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_355_i58_3_lut (.A(n27), .B(n29), .C(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .Z(n58_adj_3025)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_355_i58_3_lut.init = 16'hcaca;
    LUT4 i11352_4_lut (.A(n97), .B(n178_adj_2995), .C(n113), .D(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .Z(n62[27])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam i11352_4_lut.init = 16'h3022;
    LUT4 modulation_output_15__I_0_355_i47_3_lut (.A(n16), .B(n18), .C(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .Z(n47_adj_3005)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_355_i47_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_355_i16_3_lut (.A(modulation_output[15]), 
         .B(modulation_output[14]), .C(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .Z(n16)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_355_i16_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_355_i112_3_lut_rep_413 (.A(n81), .B(n89), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[3]), .Z(n27078)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_355_i112_3_lut_rep_413.init = 16'hcaca;
    LUT4 i11385_2_lut_4_lut (.A(n81), .B(n89), .C(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .D(n27092), .Z(n62[12])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam i11385_2_lut_4_lut.init = 16'h00ca;
    LUT4 modulation_output_15__I_0_355_i111_3_lut_rep_414 (.A(n80), .B(n88), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[3]), .Z(n27079)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_355_i111_3_lut_rep_414.init = 16'hcaca;
    LUT4 i11386_2_lut_4_lut (.A(n80), .B(n88), .C(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .D(n27092), .Z(n62[13])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam i11386_2_lut_4_lut.init = 16'h00ca;
    LUT4 modulation_output_15__I_0_355_i113_4_lut (.A(n82), .B(n59_adj_3003), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[3]), .D(modulation_deviation_amount_minus_sine_lookup_width[2]), 
         .Z(n113)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_355_i113_4_lut.init = 16'h0aca;
    LUT4 modulation_output_15__I_0_355_i82_3_lut (.A(n51_adj_3026), .B(n55_adj_3016), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[2]), .Z(n82)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_355_i82_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_355_i59_3_lut (.A(n28), .B(n30), .C(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .Z(n59_adj_3003)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_355_i59_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_355_i51_3_lut (.A(n20), .B(n22), .C(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .Z(n51_adj_3026)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_355_i51_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_355_i55_3_lut (.A(n24), .B(n26), .C(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .Z(n55_adj_3016)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_355_i55_3_lut.init = 16'hcaca;
    LUT4 i11369_4_lut (.A(n98), .B(n178_adj_2995), .C(n114), .D(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .Z(n62[26])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam i11369_4_lut.init = 16'h3022;
    LUT4 modulation_output_15__I_0_355_i114_4_lut (.A(n83), .B(n60_adj_3006), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[3]), .D(modulation_deviation_amount_minus_sine_lookup_width[2]), 
         .Z(n114)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_355_i114_4_lut.init = 16'h0aca;
    LUT4 modulation_output_15__I_0_355_i83_3_lut (.A(n52_adj_3018), .B(n56_adj_3017), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[2]), .Z(n83)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_355_i83_3_lut.init = 16'hcaca;
    LUT4 i11373_4_lut (.A(n99), .B(n178_adj_2995), .C(n115), .D(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .Z(n62[25])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam i11373_4_lut.init = 16'h3022;
    LUT4 modulation_output_15__I_0_355_i99_3_lut (.A(modulation_output[15]), 
         .B(n76), .C(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .Z(n99)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_355_i99_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_355_i76_3_lut (.A(n45_adj_3027), .B(n49_adj_3020), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[2]), .Z(n76)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_355_i76_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_355_i115_4_lut (.A(n84), .B(n30), .C(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .D(n27282), .Z(n115)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_355_i115_4_lut.init = 16'h0aca;
    LUT4 modulation_output_15__I_0_355_i84_3_lut (.A(n53_adj_3021), .B(n57_adj_3022), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[2]), .Z(n84)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_355_i84_3_lut.init = 16'hcaca;
    LUT4 i11380_4_lut (.A(n100_adj_3028), .B(n178_adj_2995), .C(n116), 
         .D(modulation_deviation_amount_minus_sine_lookup_width[4]), .Z(n62[24])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam i11380_4_lut.init = 16'h3022;
    CCU2D add_425_3 (.A0(\addr_space[0] [1]), .B0(n14676), .C0(carrier_center_increment_offset_rs[1]), 
          .D0(carrier_center_increment_offset_ls[1]), .A1(\addr_space[0] [2]), 
          .B1(n14676), .C1(carrier_center_increment_offset_rs[2]), .D1(carrier_center_increment_offset_ls[2]), 
          .CIN(n17911), .COUT(n17912), .S0(carrier_increment_30__N_1590[1]), 
          .S1(carrier_increment_30__N_1590[2]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(105[4:87])
    defparam add_425_3.INIT0 = 16'h569a;
    defparam add_425_3.INIT1 = 16'h569a;
    defparam add_425_3.INJECT1_0 = "NO";
    defparam add_425_3.INJECT1_1 = "NO";
    LUT4 modulation_output_15__I_0_355_i100_3_lut (.A(modulation_output[15]), 
         .B(n77), .C(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .Z(n100_adj_3028)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_355_i100_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_355_i77_3_lut (.A(n46_adj_3029), .B(n50_adj_3023), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[2]), .Z(n77)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_355_i77_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_355_i46_3_lut (.A(modulation_output[15]), 
         .B(n17), .C(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .Z(n46_adj_3029)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_355_i46_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_355_i116_4_lut (.A(n85), .B(modulation_output[0]), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[3]), .D(n27138), 
         .Z(n116)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_355_i116_4_lut.init = 16'h0aca;
    CCU2D sub_106_add_2_9 (.A0(\addr_space[2] [11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\addr_space[2] [12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17974), .COUT(n17975), .S0(modulation_deviation_amount_minus_sine_lookup_width_16__N_1638[11]), 
          .S1(modulation_deviation_amount_minus_sine_lookup_width_16__N_1638[12]));
    defparam sub_106_add_2_9.INIT0 = 16'h5555;
    defparam sub_106_add_2_9.INIT1 = 16'h5555;
    defparam sub_106_add_2_9.INJECT1_0 = "NO";
    defparam sub_106_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_106_add_2_7 (.A0(\addr_space[2] [9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\addr_space[2] [10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17973), .COUT(n17974), .S0(modulation_deviation_amount_minus_sine_lookup_width_16__N_1638[9]), 
          .S1(modulation_deviation_amount_minus_sine_lookup_width_16__N_1638[10]));
    defparam sub_106_add_2_7.INIT0 = 16'h5555;
    defparam sub_106_add_2_7.INIT1 = 16'h5555;
    defparam sub_106_add_2_7.INJECT1_0 = "NO";
    defparam sub_106_add_2_7.INJECT1_1 = "NO";
    LUT4 modulation_output_15__I_0_355_i85_3_lut (.A(n54_adj_3024), .B(n58_adj_3025), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[2]), .Z(n85)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_355_i85_3_lut.init = 16'hcaca;
    CCU2D add_425_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\addr_space[0] [0]), .B1(n14676), .C1(carrier_center_increment_offset_rs[0]), 
          .D1(carrier_center_increment_offset_ls[0]), .COUT(n17911), .S1(carrier_increment_30__N_1590[0]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(105[4:87])
    defparam add_425_1.INIT0 = 16'hF000;
    defparam add_425_1.INIT1 = 16'h569a;
    defparam add_425_1.INJECT1_0 = "NO";
    defparam add_425_1.INJECT1_1 = "NO";
    CCU2D sub_106_add_2_5 (.A0(\addr_space[2] [7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\addr_space[2] [8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17972), .COUT(n17973), .S0(modulation_deviation_amount_minus_sine_lookup_width_16__N_1638[7]), 
          .S1(modulation_deviation_amount_minus_sine_lookup_width_16__N_1638[8]));
    defparam sub_106_add_2_5.INIT0 = 16'h5555;
    defparam sub_106_add_2_5.INIT1 = 16'h5555;
    defparam sub_106_add_2_5.INJECT1_0 = "NO";
    defparam sub_106_add_2_5.INJECT1_1 = "NO";
    LUT4 i11381_2_lut (.A(n132), .B(n178_adj_2995), .Z(n62[23])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam i11381_2_lut.init = 16'h2222;
    CCU2D sub_106_add_2_3 (.A0(\addr_space[2] [5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\addr_space[2] [6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17971), .COUT(n17972), .S0(modulation_deviation_amount_minus_sine_lookup_width_16__N_1638[5]), 
          .S1(modulation_deviation_amount_minus_sine_lookup_width_16__N_1638[6]));
    defparam sub_106_add_2_3.INIT0 = 16'h5555;
    defparam sub_106_add_2_3.INIT1 = 16'h5555;
    defparam sub_106_add_2_3.INJECT1_0 = "NO";
    defparam sub_106_add_2_3.INJECT1_1 = "NO";
    LUT4 i11382_2_lut (.A(n133), .B(n178_adj_2995), .Z(n62[22])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam i11382_2_lut.init = 16'h2222;
    LUT4 i11388_2_lut (.A(n134), .B(n178_adj_2995), .Z(n62[21])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam i11388_2_lut.init = 16'h2222;
    LUT4 i11389_2_lut (.A(n135), .B(n178_adj_2995), .Z(n62[20])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam i11389_2_lut.init = 16'h2222;
    LUT4 i11390_2_lut (.A(n136), .B(n178_adj_2995), .Z(n62[19])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam i11390_2_lut.init = 16'h2222;
    LUT4 i11399_2_lut (.A(n137), .B(n178_adj_2995), .Z(n62[18])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam i11399_2_lut.init = 16'h2222;
    LUT4 modulation_output_15__I_0_355_i110_3_lut_rep_415 (.A(n79), .B(n27110), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[3]), .Z(n27080)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_355_i110_3_lut_rep_415.init = 16'hcaca;
    LUT4 i11387_2_lut_4_lut (.A(n79), .B(n27110), .C(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .D(n27092), .Z(n62[14])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam i11387_2_lut_4_lut.init = 16'h00ca;
    LUT4 i11310_4_lut (.A(n107), .B(n178_adj_2995), .C(n123), .D(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .Z(n62[17])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam i11310_4_lut.init = 16'h3022;
    LUT4 modulation_output_15__I_0_355_i107_3_lut (.A(n76), .B(n84), .C(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .Z(n107)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_355_i107_3_lut.init = 16'hcaca;
    LUT4 i11311_2_lut (.A(n139), .B(n178_adj_2995), .Z(n62[16])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam i11311_2_lut.init = 16'h2222;
    LUT4 i11392_4_lut (.A(n78), .B(n27092), .C(n27109), .D(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .Z(n62[15])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam i11392_4_lut.init = 16'h3022;
    LUT4 modulation_output_15__I_0_355_i78_3_lut (.A(n47_adj_3005), .B(n51_adj_3026), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[2]), .Z(n78)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_355_i78_3_lut.init = 16'hcaca;
    CCU2D sub_437_add_2_17 (.A0(\addr_space[2] [15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\addr_space[2] [16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17909), .S0(sine_lookup_width_minus_modulation_deviation_amount_16__N_1621[15]), 
          .S1(sine_lookup_width_minus_modulation_deviation_amount_16__N_1621[16]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(96[58:109])
    defparam sub_437_add_2_17.INIT0 = 16'hf555;
    defparam sub_437_add_2_17.INIT1 = 16'hf555;
    defparam sub_437_add_2_17.INJECT1_0 = "NO";
    defparam sub_437_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_106_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\addr_space[2] [4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n17971), .S1(modulation_deviation_amount_minus_sine_lookup_width_16__N_1638[4]));
    defparam sub_106_add_2_1.INIT0 = 16'hF000;
    defparam sub_106_add_2_1.INIT1 = 16'h5555;
    defparam sub_106_add_2_1.INJECT1_0 = "NO";
    defparam sub_106_add_2_1.INJECT1_1 = "NO";
    LUT4 i6734_4_lut (.A(modulation_output[14]), .B(modulation_output[15]), 
         .C(n9095), .D(n27105), .Z(carrier_center_increment_offset_rs_30__N_1559[14])) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(100[41:116])
    defparam i6734_4_lut.init = 16'hccca;
    LUT4 i6732_4_lut (.A(n14), .B(modulation_output[15]), .C(n9093), .D(n27105), 
         .Z(carrier_center_increment_offset_rs_30__N_1559[13])) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(100[41:116])
    defparam i6732_4_lut.init = 16'hccca;
    LUT4 i6726_3_lut (.A(n73), .B(modulation_output[15]), .C(n27105), 
         .Z(carrier_center_increment_offset_rs_30__N_1559[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(100[41:116])
    defparam i6726_3_lut.init = 16'hcaca;
    LUT4 i6724_3_lut (.A(n72_adj_3013), .B(modulation_output[15]), .C(n27105), 
         .Z(carrier_center_increment_offset_rs_30__N_1559[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(100[41:116])
    defparam i6724_3_lut.init = 16'hcaca;
    LUT4 i6722_3_lut (.A(n71), .B(modulation_output[15]), .C(n27105), 
         .Z(carrier_center_increment_offset_rs_30__N_1559[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(100[41:116])
    defparam i6722_3_lut.init = 16'hcaca;
    LUT4 i6720_3_lut (.A(n70), .B(modulation_output[15]), .C(n27105), 
         .Z(carrier_center_increment_offset_rs_30__N_1559[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(100[41:116])
    defparam i6720_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i70_3_lut (.A(n39_adj_3004), .B(n43), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[2]), .Z(n70)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(100[41:116])
    defparam modulation_output_15__I_0_i70_3_lut.init = 16'hcaca;
    CCU2D sub_437_add_2_15 (.A0(\addr_space[2] [13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\addr_space[2] [14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17908), .COUT(n17909), .S0(sine_lookup_width_minus_modulation_deviation_amount_16__N_1621[13]), 
          .S1(sine_lookup_width_minus_modulation_deviation_amount_16__N_1621[14]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(96[58:109])
    defparam sub_437_add_2_15.INIT0 = 16'hf555;
    defparam sub_437_add_2_15.INIT1 = 16'hf555;
    defparam sub_437_add_2_15.INJECT1_0 = "NO";
    defparam sub_437_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_437_add_2_13 (.A0(\addr_space[2] [11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\addr_space[2] [12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17907), .COUT(n17908), .S0(sine_lookup_width_minus_modulation_deviation_amount_16__N_1621[11]), 
          .S1(sine_lookup_width_minus_modulation_deviation_amount_16__N_1621[12]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(96[58:109])
    defparam sub_437_add_2_13.INIT0 = 16'hf555;
    defparam sub_437_add_2_13.INIT1 = 16'hf555;
    defparam sub_437_add_2_13.INJECT1_0 = "NO";
    defparam sub_437_add_2_13.INJECT1_1 = "NO";
    LUT4 i23143_2_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[3]), .Z(n22608)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam i23143_2_lut.init = 16'heeee;
    LUT4 i1_3_lut_4_lut (.A(n27138), .B(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .C(modulation_output[0]), .D(n27092), .Z(n20732)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam i1_3_lut_4_lut.init = 16'h0010;
    LUT4 i6557_2_lut_rep_427 (.A(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .B(n178_adj_2995), .Z(n27092)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam i6557_2_lut_rep_427.init = 16'heeee;
    LUT4 i11945_2_lut_3_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .B(n178_adj_2995), .C(n27110), .D(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .Z(n62[6])) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam i11945_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 i12208_2_lut_3_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .B(n178_adj_2995), .C(n60_adj_3006), .D(n27272), .Z(n62[2])) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam i12208_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 i11946_2_lut_3_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .B(n178_adj_2995), .C(n88), .D(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .Z(n62[5])) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam i11946_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 i11944_2_lut_3_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .B(n178_adj_2995), .C(n27109), .D(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .Z(n62[7])) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam i11944_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 i12211_2_lut_3_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .B(n178_adj_2995), .C(n59_adj_3003), .D(n27272), .Z(n62[3])) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam i12211_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 i11947_2_lut_3_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .B(n178_adj_2995), .C(n89), .D(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .Z(n62[4])) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam i11947_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 i11377_2_lut_3_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .B(n178_adj_2995), .C(n115), .Z(n62[9])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam i11377_2_lut_3_lut.init = 16'h1010;
    LUT4 i11383_2_lut_3_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .B(n178_adj_2995), .C(n114), .Z(n62[10])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam i11383_2_lut_3_lut.init = 16'h1010;
    LUT4 i11384_2_lut_3_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .B(n178_adj_2995), .C(n113), .Z(n62[11])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam i11384_2_lut_3_lut.init = 16'h1010;
    LUT4 i11682_2_lut_3_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .B(n178_adj_2995), .C(n116), .Z(n62[8])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam i11682_2_lut_3_lut.init = 16'h1010;
    LUT4 i1_2_lut_3_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .B(n178_adj_2995), .C(n123), .Z(n20736)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam i1_2_lut_3_lut.init = 16'h1010;
    LUT4 modulation_output_15__I_0_i94_3_lut_4_lut (.A(sine_lookup_width_minus_modulation_deviation_amount[4]), 
         .B(n178), .C(modulation_output[15]), .D(n1), .Z(n94)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(100[41:116])
    defparam modulation_output_15__I_0_i94_3_lut_4_lut.init = 16'hf1e0;
    CCU2D sub_437_add_2_11 (.A0(\addr_space[2] [9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\addr_space[2] [10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17906), .COUT(n17907), .S0(sine_lookup_width_minus_modulation_deviation_amount_16__N_1621[9]), 
          .S1(sine_lookup_width_minus_modulation_deviation_amount_16__N_1621[10]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(96[58:109])
    defparam sub_437_add_2_11.INIT0 = 16'hf555;
    defparam sub_437_add_2_11.INIT1 = 16'hf555;
    defparam sub_437_add_2_11.INJECT1_0 = "NO";
    defparam sub_437_add_2_11.INJECT1_1 = "NO";
    LUT4 i23027_3_lut (.A(n61[10]), .B(i_sw0_c), .C(cw_N_1877), .Z(dac_clk_p_c_enable_432)) /* synthesis lut_function=(!(A (B)+!A (B+!(C)))) */ ;
    defparam i23027_3_lut.init = 16'h3232;
    LUT4 i10107_3_lut_rep_417_4_lut (.A(sine_lookup_width_minus_modulation_deviation_amount[4]), 
         .B(n178), .C(sine_lookup_width_minus_modulation_deviation_amount[3]), 
         .D(n9095), .Z(n27082)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(100[41:116])
    defparam i10107_3_lut_rep_417_4_lut.init = 16'hfeee;
    LUT4 modulation_output_15__I_0_i95_3_lut_4_lut (.A(sine_lookup_width_minus_modulation_deviation_amount[4]), 
         .B(n178), .C(modulation_output[15]), .D(n2_c), .Z(n95)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(100[41:116])
    defparam modulation_output_15__I_0_i95_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i11795_2_lut (.A(o_sample_i[13]), .B(cw_mux_dac_a_mux_sel), .Z(o_dac_a_c_6)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(29[18:140])
    defparam i11795_2_lut.init = 16'h2222;
    LUT4 modulation_output_15__I_0_355_i104_4_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[4]), .C(n89), 
         .D(n81), .Z(n104)) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C)+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam modulation_output_15__I_0_355_i104_4_lut_4_lut.init = 16'h7340;
    LUT4 i11354_2_lut_4_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[2]), .C(n59_adj_3003), 
         .D(n55_adj_3016), .Z(n117)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam i11354_2_lut_4_lut_4_lut.init = 16'h5140;
    LUT4 i11355_2_lut_4_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[2]), .C(n60_adj_3006), 
         .D(n56_adj_3017), .Z(n118)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam i11355_2_lut_4_lut_4_lut.init = 16'h5140;
    LUT4 modulation_output_15__I_0_355_i103_4_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[4]), .C(n88), 
         .D(n80), .Z(n103)) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C)+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam modulation_output_15__I_0_355_i103_4_lut_4_lut.init = 16'h7340;
    LUT4 i10017_1_lut (.A(n61[15]), .Z(dac_clk_p_c_enable_486)) /* synthesis lut_function=(!(A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(143[21:41])
    defparam i10017_1_lut.init = 16'h5555;
    CCU2D sub_437_add_2_9 (.A0(\addr_space[2] [7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\addr_space[2] [8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17905), .COUT(n17906), .S0(sine_lookup_width_minus_modulation_deviation_amount_16__N_1621[7]), 
          .S1(sine_lookup_width_minus_modulation_deviation_amount_16__N_1621[8]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(96[58:109])
    defparam sub_437_add_2_9.INIT0 = 16'hf555;
    defparam sub_437_add_2_9.INIT1 = 16'hf555;
    defparam sub_437_add_2_9.INJECT1_0 = "NO";
    defparam sub_437_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_437_add_2_7 (.A0(\addr_space[2] [5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\addr_space[2] [6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17904), .COUT(n17905), .S0(sine_lookup_width_minus_modulation_deviation_amount_16__N_1621[5]), 
          .S1(sine_lookup_width_minus_modulation_deviation_amount_16__N_1621[6]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(96[58:109])
    defparam sub_437_add_2_7.INIT0 = 16'hf555;
    defparam sub_437_add_2_7.INIT1 = 16'hf555;
    defparam sub_437_add_2_7.INJECT1_0 = "NO";
    defparam sub_437_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_437_add_2_5 (.A0(\addr_space[2] [3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\addr_space[2] [4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17903), .COUT(n17904), .S0(sine_lookup_width_minus_modulation_deviation_amount_16__N_1621[3]), 
          .S1(sine_lookup_width_minus_modulation_deviation_amount_16__N_1621[4]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(96[58:109])
    defparam sub_437_add_2_5.INIT0 = 16'hf555;
    defparam sub_437_add_2_5.INIT1 = 16'h0aaa;
    defparam sub_437_add_2_5.INJECT1_0 = "NO";
    defparam sub_437_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_437_add_2_3 (.A0(\addr_space[2] [1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\addr_space[2] [2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17902), .COUT(n17903), .S0(sine_lookup_width_minus_modulation_deviation_amount_16__N_1621[1]), 
          .S1(sine_lookup_width_minus_modulation_deviation_amount_16__N_1621[2]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(96[58:109])
    defparam sub_437_add_2_3.INIT0 = 16'hf555;
    defparam sub_437_add_2_3.INIT1 = 16'hf555;
    defparam sub_437_add_2_3.INJECT1_0 = "NO";
    defparam sub_437_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_437_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\addr_space[2] [0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n17902));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(96[58:109])
    defparam sub_437_add_2_1.INIT0 = 16'h0000;
    defparam sub_437_add_2_1.INIT1 = 16'h0aaa;
    defparam sub_437_add_2_1.INJECT1_0 = "NO";
    defparam sub_437_add_2_1.INJECT1_1 = "NO";
    LUT4 i11796_2_lut (.A(o_sample_i[12]), .B(cw_mux_dac_a_mux_sel), .Z(o_dac_a_c_5)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(29[18:140])
    defparam i11796_2_lut.init = 16'heeee;
    LUT4 i11797_2_lut (.A(o_sample_i[11]), .B(cw_mux_dac_a_mux_sel), .Z(o_dac_a_c_4)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(29[18:140])
    defparam i11797_2_lut.init = 16'h2222;
    LUT4 i11798_2_lut (.A(o_sample_i[10]), .B(cw_mux_dac_a_mux_sel), .Z(o_dac_a_c_3)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(29[18:140])
    defparam i11798_2_lut.init = 16'h2222;
    LUT4 i11799_2_lut (.A(o_sample_i[9]), .B(cw_mux_dac_a_mux_sel), .Z(o_dac_a_c_2)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(29[18:140])
    defparam i11799_2_lut.init = 16'h2222;
    LUT4 i11800_2_lut (.A(o_sample_i[8]), .B(cw_mux_dac_a_mux_sel), .Z(o_dac_a_c_1)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(29[18:140])
    defparam i11800_2_lut.init = 16'h2222;
    LUT4 i11321_2_lut (.A(o_sample_i[7]), .B(cw_mux_dac_a_mux_sel), .Z(o_dac_a_c_0)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(29[18:140])
    defparam i11321_2_lut.init = 16'h2222;
    PFUMX i20138 (.BLUT(n22491), .ALUT(n22492), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1336[17]));
    LUT4 i849_1_lut (.A(o_dac_b_c_15), .Z(o_dac_b_c_9)) /* synthesis lut_function=(!(A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(28[31:66])
    defparam i849_1_lut.init = 16'h5555;
    LUT4 cw_I_0_1_lut (.A(cw), .Z(o_dac_cw_b_c)) /* synthesis lut_function=(!(A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(111[17:20])
    defparam cw_I_0_1_lut.init = 16'h5555;
    PFUMX i20147 (.BLUT(n22500), .ALUT(n22501), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1336[16]));
    LUT4 i23164_2_lut_rep_607 (.A(modulation_deviation_amount_minus_sine_lookup_width[2]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[3]), .Z(n27272)) /* synthesis lut_function=(!(A+(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam i23164_2_lut_rep_607.init = 16'h1111;
    PFUMX i20153 (.BLUT(n22506), .ALUT(n22507), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1336[15]));
    PFUMX i20156 (.BLUT(n22509), .ALUT(n22510), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1336[14]));
    PFUMX i20159 (.BLUT(n22512), .ALUT(n22513), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1336[13]));
    PFUMX i20162 (.BLUT(n22515), .ALUT(n22516), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1336[12]));
    LUT4 i6630_2_lut_rep_617 (.A(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[2]), .Z(n27282)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam i6630_2_lut_rep_617.init = 16'heeee;
    LUT4 i12217_3_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[2]), .C(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .D(n30), .Z(n123)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam i12217_3_lut_4_lut.init = 16'h0100;
    LUT4 i6639_3_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[2]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[3]), .C(n47_adj_3005), 
         .D(modulation_output[15]), .Z(n97)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam i6639_3_lut_4_lut.init = 16'hf780;
    LUT4 i6641_3_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[2]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[3]), .C(n48_adj_3007), 
         .D(modulation_output[15]), .Z(n98)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam i6641_3_lut_4_lut.init = 16'hf780;
    LUT4 i6628_2_lut_rep_618 (.A(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[2]), .Z(n27283)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam i6628_2_lut_rep_618.init = 16'h8888;
    LUT4 i6629_3_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[2]), .C(n17), 
         .D(modulation_output[15]), .Z(n73_adj_3015)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam i6629_3_lut_4_lut.init = 16'hf780;
    LUT4 i6622_2_lut_rep_619 (.A(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[1]), .Z(n27284)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam i6622_2_lut_rep_619.init = 16'h8888;
    LUT4 i6626_2_lut_rep_489_3_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[1]), .C(modulation_deviation_amount_minus_sine_lookup_width[2]), 
         .Z(n27154)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam i6626_2_lut_rep_489_3_lut.init = 16'h8080;
    LUT4 i6623_3_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[1]), .C(modulation_output[14]), 
         .D(modulation_output[15]), .Z(n45_adj_3027)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam i6623_3_lut_4_lut.init = 16'hf780;
    PFUMX i20165 (.BLUT(n22518), .ALUT(n22519), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1336[11]));
    PFUMX i20168 (.BLUT(n22521), .ALUT(n22522), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1336[10]));
    PFUMX i20174 (.BLUT(n22527), .ALUT(n22528), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1336[9]));
    PFUMX i20177 (.BLUT(n22530), .ALUT(n22531), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1336[8]));
    PFUMX i20180 (.BLUT(n22533), .ALUT(n22534), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1336[7]));
    PFUMX i20183 (.BLUT(n22536), .ALUT(n22537), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1336[6]));
    LUT4 i20128_3_lut (.A(\addr_space[2] [18]), .B(\addr_space[3] [18]), 
         .C(\wb_addr[0] ), .Z(n22483)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20128_3_lut.init = 16'hcaca;
    LUT4 i20127_3_lut (.A(\addr_space[0] [18]), .B(\addr_space[1] [18]), 
         .C(\wb_addr[0] ), .Z(n22482)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20127_3_lut.init = 16'hcaca;
    PFUMX i20186 (.BLUT(n22539), .ALUT(n22540), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1336[5]));
    PFUMX i19328 (.BLUT(n21681), .ALUT(n21682), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1336[4]));
    PFUMX i19331 (.BLUT(n21684), .ALUT(n21685), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1336[3]));
    PFUMX i19334 (.BLUT(n21687), .ALUT(n21688), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1336[2]));
    LUT4 i12507_2_lut_rep_715 (.A(o_sample_i[15]), .B(cw_mux_dac_a_mux_sel), 
         .Z(n27380)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i12507_2_lut_rep_715.init = 16'heeee;
    LUT4 i12508_1_lut_2_lut (.A(o_sample_i[15]), .B(cw_mux_dac_a_mux_sel), 
         .Z(o_dac_a_c_9)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i12508_1_lut_2_lut.init = 16'h1111;
    PFUMX i19337 (.BLUT(n21690), .ALUT(n21691), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1336[1]));
    PFUMX i20051 (.BLUT(n22404), .ALUT(n22405), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1336[0]));
    PFUMX i20054 (.BLUT(n22407), .ALUT(n22408), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1336[31]));
    PFUMX i20057 (.BLUT(n22410), .ALUT(n22411), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1336[30]));
    PFUMX i20060 (.BLUT(n22413), .ALUT(n22414), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1336[29]));
    LUT4 i23142_4_lut (.A(n21102), .B(n27304), .C(n38), .D(\wb_addr[15] ), 
         .Z(dac_clk_p_c_enable_116)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(44[3] 46[6])
    defparam i23142_4_lut.init = 16'h0400;
    PFUMX i20063 (.BLUT(n22416), .ALUT(n22417), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1336[28]));
    PFUMX i20066 (.BLUT(n22419), .ALUT(n22420), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1336[27]));
    LUT4 smpl_register_5__bdd_4_lut_4_lut (.A(\wb_addr[0] ), .B(\wb_addr[1] ), 
         .C(n2), .D(\smpl_register[5] ), .Z(n27049)) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(45[4:25])
    defparam smpl_register_5__bdd_4_lut_4_lut.init = 16'hf3d1;
    LUT4 smpl_register_20__bdd_4_lut_4_lut (.A(\wb_addr[0] ), .B(\wb_addr[1] ), 
         .C(n2_adj_1), .D(\smpl_register[20] ), .Z(n27061)) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(45[4:25])
    defparam smpl_register_20__bdd_4_lut_4_lut.init = 16'hf3d1;
    LUT4 modulation_output_15__I_0_i64_3_lut (.A(n33_adj_3011), .B(n72_adj_3013), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[3]), .Z(n64)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(100[41:116])
    defparam modulation_output_15__I_0_i64_3_lut.init = 16'hcaca;
    LUT4 smpl_register_18__bdd_4_lut_4_lut (.A(\wb_addr[0] ), .B(\wb_addr[1] ), 
         .C(n2_adj_2), .D(\smpl_register[18] ), .Z(n27059)) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(45[4:25])
    defparam smpl_register_18__bdd_4_lut_4_lut.init = 16'hf3d1;
    LUT4 smpl_register_17__bdd_4_lut_4_lut (.A(\wb_addr[0] ), .B(\wb_addr[1] ), 
         .C(n2_adj_3), .D(\smpl_register[17] ), .Z(n27058)) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(45[4:25])
    defparam smpl_register_17__bdd_4_lut_4_lut.init = 16'hf3d1;
    LUT4 modulation_output_15__I_0_i63_3_lut (.A(n32_adj_3010), .B(n71), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[3]), .Z(n63)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(100[41:116])
    defparam modulation_output_15__I_0_i63_3_lut.init = 16'hcaca;
    LUT4 smpl_register_16__bdd_4_lut_4_lut (.A(\wb_addr[0] ), .B(\wb_addr[1] ), 
         .C(n2_adj_4), .D(\smpl_register[16] ), .Z(n27057)) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(45[4:25])
    defparam smpl_register_16__bdd_4_lut_4_lut.init = 16'hf3d1;
    LUT4 smpl_register_29__bdd_4_lut_4_lut (.A(\wb_addr[0] ), .B(\wb_addr[1] ), 
         .C(n2_adj_5), .D(\smpl_register[29] ), .Z(n27056)) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(45[4:25])
    defparam smpl_register_29__bdd_4_lut_4_lut.init = 16'hf3d1;
    LUT4 smpl_register_10__bdd_4_lut_4_lut (.A(\wb_addr[0] ), .B(\wb_addr[1] ), 
         .C(n2_adj_6), .D(\smpl_register[10] ), .Z(n27051)) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(45[4:25])
    defparam smpl_register_10__bdd_4_lut_4_lut.init = 16'hf3d1;
    LUT4 smpl_register_9__bdd_4_lut_4_lut (.A(\wb_addr[0] ), .B(\wb_addr[1] ), 
         .C(n2_adj_7), .D(\smpl_register[9] ), .Z(n27050)) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(45[4:25])
    defparam smpl_register_9__bdd_4_lut_4_lut.init = 16'hf3d1;
    PFUMX i20069 (.BLUT(n22422), .ALUT(n22423), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1336[26]));
    PFUMX i20072 (.BLUT(n22425), .ALUT(n22426), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1336[25]));
    PFUMX i20075 (.BLUT(n22428), .ALUT(n22429), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1336[24]));
    PFUMX modulation_output_15__I_0_355_i139 (.BLUT(n108), .ALUT(n124), 
          .C0(modulation_deviation_amount_minus_sine_lookup_width[4]), .Z(n139)) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;
    PFUMX i20081 (.BLUT(n22434), .ALUT(n22435), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1336[23]));
    PFUMX modulation_output_15__I_0_355_i137 (.BLUT(n75), .ALUT(n106), .C0(n22608), 
          .Z(n137)) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;
    PFUMX modulation_output_15__I_0_355_i136 (.BLUT(n74), .ALUT(n105), .C0(n22608), 
          .Z(n136)) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;
    PFUMX modulation_output_15__I_0_355_i133 (.BLUT(n102), .ALUT(n118), 
          .C0(modulation_deviation_amount_minus_sine_lookup_width[4]), .Z(n133)) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;
    PFUMX i20084 (.BLUT(n22437), .ALUT(n22438), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1336[22]));
    PFUMX modulation_output_15__I_0_355_i132 (.BLUT(n101), .ALUT(n117), 
          .C0(modulation_deviation_amount_minus_sine_lookup_width[4]), .Z(n132)) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;
    PFUMX i20087 (.BLUT(n22440), .ALUT(n22441), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1336[21]));
    PFUMX i20099 (.BLUT(n22452), .ALUT(n22453), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1336[20]));
    PFUMX i20114 (.BLUT(n22467), .ALUT(n22468), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1336[19]));
    LUT4 i23138_4_lut (.A(n21088), .B(\wb_addr[0] ), .C(n21078), .D(\wb_addr[15] ), 
         .Z(dac_clk_p_c_enable_73)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(44[3] 46[6])
    defparam i23138_4_lut.init = 16'h0400;
    FD1P3AX cw_350 (.D(cw_N_1877), .SP(dac_clk_p_c_enable_432), .CK(dac_clk_p_c), 
            .Q(cw)) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=129, LSE_RLINE=141 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(133[11] 145[5])
    defparam cw_350.GSR = "DISABLED";
    PFUMX i23489 (.BLUT(n25139), .ALUT(n38_adj_3008), .C0(sine_lookup_width_minus_modulation_deviation_amount[2]), 
          .Z(n25140));
    LUT4 i23133_4_lut (.A(n21088), .B(n21044), .C(\wb_addr[1] ), .D(\wb_addr[15] ), 
         .Z(dac_clk_p_c_enable_105)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(44[3] 46[6])
    defparam i23133_4_lut.init = 16'h1000;
    LUT4 i6674_2_lut_3_lut (.A(sine_lookup_width_minus_modulation_deviation_amount[0]), 
         .B(sine_lookup_width_minus_modulation_deviation_amount[1]), .C(sine_lookup_width_minus_modulation_deviation_amount[2]), 
         .Z(n9095)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(100[41:116])
    defparam i6674_2_lut_3_lut.init = 16'hfefe;
    LUT4 modulation_output_15__I_0_i100_4_lut (.A(modulation_output[14]), 
         .B(modulation_output[15]), .C(n27082), .D(n9095), .Z(n100)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(100[41:116])
    defparam modulation_output_15__I_0_i100_4_lut.init = 16'hc0ca;
    LUT4 modulation_output_15__I_0_i69_3_lut (.A(n38_adj_3008), .B(n42_adj_3009), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[2]), .Z(n69)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(100[41:116])
    defparam modulation_output_15__I_0_i69_3_lut.init = 16'hcaca;
    LUT4 i6671_3_lut_4_lut (.A(sine_lookup_width_minus_modulation_deviation_amount[0]), 
         .B(sine_lookup_width_minus_modulation_deviation_amount[1]), .C(modulation_output[15]), 
         .D(modulation_output[14]), .Z(n46_adj_3014)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(100[41:116])
    defparam i6671_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i23071_4_lut_4_lut (.A(sine_lookup_width_minus_modulation_deviation_amount[2]), 
         .B(sine_lookup_width_minus_modulation_deviation_amount[1]), .C(sine_lookup_width_minus_modulation_deviation_amount[3]), 
         .D(n27121), .Z(n22774)) /* synthesis lut_function=(A (D)+!A (B (D)+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 107[5])
    defparam i23071_4_lut_4_lut.init = 16'hff01;
    LUT4 i6624_2_lut_rep_585 (.A(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[1]), .Z(n27250)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam i6624_2_lut_rep_585.init = 16'heeee;
    LUT4 i6632_2_lut_rep_473_3_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[1]), .C(modulation_deviation_amount_minus_sine_lookup_width[2]), 
         .Z(n27138)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam i6632_2_lut_rep_473_3_lut.init = 16'hfefe;
    PFUMX i23438 (.BLUT(n25049), .ALUT(n25048), .C0(sine_lookup_width_minus_modulation_deviation_amount[3]), 
          .Z(n25050));
    PFUMX i23436 (.BLUT(n25045), .ALUT(n25044), .C0(sine_lookup_width_minus_modulation_deviation_amount[2]), 
          .Z(n25046));
    FD1P3DX startup_timer_FSM_i0_i15 (.D(n29969), .SP(n1109[14]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(n61[15]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(143[21:41])
    defparam startup_timer_FSM_i0_i15.GSR = "DISABLED";
    FD1P3DX startup_timer_FSM_i0_i14 (.D(n1109[13]), .SP(dac_clk_p_c_enable_486), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(n1109[14]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(143[21:41])
    defparam startup_timer_FSM_i0_i14.GSR = "DISABLED";
    FD1P3DX startup_timer_FSM_i0_i13 (.D(n1109[12]), .SP(dac_clk_p_c_enable_486), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(n1109[13]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(143[21:41])
    defparam startup_timer_FSM_i0_i13.GSR = "DISABLED";
    FD1P3DX startup_timer_FSM_i0_i12 (.D(n1109[11]), .SP(dac_clk_p_c_enable_486), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(n1109[12]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(143[21:41])
    defparam startup_timer_FSM_i0_i12.GSR = "DISABLED";
    FD1P3DX startup_timer_FSM_i0_i11 (.D(n61[10]), .SP(dac_clk_p_c_enable_486), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(n1109[11]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(143[21:41])
    defparam startup_timer_FSM_i0_i11.GSR = "DISABLED";
    FD1P3DX startup_timer_FSM_i0_i10 (.D(n1109[9]), .SP(dac_clk_p_c_enable_486), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(n61[10]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(143[21:41])
    defparam startup_timer_FSM_i0_i10.GSR = "DISABLED";
    FD1P3DX startup_timer_FSM_i0_i9 (.D(n1109[8]), .SP(dac_clk_p_c_enable_486), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(n1109[9]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(143[21:41])
    defparam startup_timer_FSM_i0_i9.GSR = "DISABLED";
    FD1P3DX startup_timer_FSM_i0_i8 (.D(n1109[7]), .SP(dac_clk_p_c_enable_486), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(n1109[8]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(143[21:41])
    defparam startup_timer_FSM_i0_i8.GSR = "DISABLED";
    FD1P3DX startup_timer_FSM_i0_i7 (.D(n1109[6]), .SP(dac_clk_p_c_enable_486), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(n1109[7]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(143[21:41])
    defparam startup_timer_FSM_i0_i7.GSR = "DISABLED";
    FD1P3DX startup_timer_FSM_i0_i6 (.D(n1109[5]), .SP(dac_clk_p_c_enable_486), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(n1109[6]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(143[21:41])
    defparam startup_timer_FSM_i0_i6.GSR = "DISABLED";
    FD1P3DX startup_timer_FSM_i0_i5 (.D(n1109[4]), .SP(dac_clk_p_c_enable_486), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(n1109[5]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(143[21:41])
    defparam startup_timer_FSM_i0_i5.GSR = "DISABLED";
    FD1P3DX startup_timer_FSM_i0_i4 (.D(cw_N_1877), .SP(dac_clk_p_c_enable_486), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(n1109[4]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(143[21:41])
    defparam startup_timer_FSM_i0_i4.GSR = "DISABLED";
    FD1P3DX startup_timer_FSM_i0_i3 (.D(n1109[2]), .SP(dac_clk_p_c_enable_486), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(cw_N_1877));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(143[21:41])
    defparam startup_timer_FSM_i0_i3.GSR = "DISABLED";
    FD1P3DX startup_timer_FSM_i0_i2 (.D(n1109[1]), .SP(dac_clk_p_c_enable_486), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(n1109[2]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(143[21:41])
    defparam startup_timer_FSM_i0_i2.GSR = "DISABLED";
    FD1P3DX startup_timer_FSM_i0_i1 (.D(n1109[0]), .SP(dac_clk_p_c_enable_486), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(n1109[1]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(143[21:41])
    defparam startup_timer_FSM_i0_i1.GSR = "DISABLED";
    PFUMX i23433 (.BLUT(n25040), .ALUT(n39_adj_3004), .C0(sine_lookup_width_minus_modulation_deviation_amount[2]), 
          .Z(n25041));
    dds modulation (.dac_clk_p_c(dac_clk_p_c), .i_sw0_c(i_sw0_c), .\addr_space[1][0] (\addr_space[1] [0]), 
        .\addr_space[1][30] (\addr_space[1] [30]), .\addr_space[1][29] (\addr_space[1] [29]), 
        .\addr_space[1][28] (\addr_space[1] [28]), .\addr_space[1][27] (\addr_space[1] [27]), 
        .\addr_space[1][26] (\addr_space[1] [26]), .\addr_space[1][25] (\addr_space[1] [25]), 
        .\addr_space[1][24] (\addr_space[1] [24]), .\addr_space[1][23] (\addr_space[1] [23]), 
        .\addr_space[1][22] (\addr_space[1] [22]), .\addr_space[1][21] (\addr_space[1] [21]), 
        .\addr_space[1][20] (\addr_space[1] [20]), .\addr_space[1][19] (\addr_space[1] [19]), 
        .\addr_space[1][18] (\addr_space[1] [18]), .\addr_space[1][17] (\addr_space[1] [17]), 
        .\addr_space[1][16] (\addr_space[1] [16]), .\addr_space[1][15] (\addr_space[1] [15]), 
        .\addr_space[1][14] (\addr_space[1] [14]), .\addr_space[1][13] (\addr_space[1] [13]), 
        .\addr_space[1][12] (\addr_space[1] [12]), .\addr_space[1][11] (\addr_space[1] [11]), 
        .\addr_space[1][10] (\addr_space[1] [10]), .\addr_space[1][9] (\addr_space[1] [9]), 
        .\addr_space[1][8] (\addr_space[1] [8]), .\addr_space[1][7] (\addr_space[1] [7]), 
        .\addr_space[1][6] (\addr_space[1] [6]), .\addr_space[1][5] (\addr_space[1] [5]), 
        .\addr_space[1][4] (\addr_space[1] [4]), .\addr_space[1][3] (\addr_space[1] [3]), 
        .\addr_space[1][2] (\addr_space[1] [2]), .\addr_space[1][1] (\addr_space[1] [1]), 
        .dac_clk_p_c_enable_488(dac_clk_p_c_enable_488), .modulation_output({modulation_output}), 
        .\quarter_wave_sample_register_q[15] (quarter_wave_sample_register_q[15]), 
        .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(83[4:161])
    dds_U2 carrier (.dac_clk_p_c(dac_clk_p_c), .i_sw0_c(i_sw0_c), .carrier_increment({carrier_increment}), 
           .dac_clk_p_c_enable_488(dac_clk_p_c_enable_488), .o_dac_b_c_7(o_dac_b_c_7), 
           .\o_sample_i[7] (o_sample_i[7]), .\o_sample_i[15] (o_sample_i[15]), 
           .\o_sample_i[14] (o_sample_i[14]), .\o_sample_i[13] (o_sample_i[13]), 
           .\o_sample_i[12] (o_sample_i[12]), .\o_sample_i[11] (o_sample_i[11]), 
           .\o_sample_i[10] (o_sample_i[10]), .\o_sample_i[9] (o_sample_i[9]), 
           .\o_sample_i[8] (o_sample_i[8]), .GND_net(GND_net), .\quarter_wave_sample_register_q[15] (quarter_wave_sample_register_q[15]), 
           .n29968(n29968), .o_dac_b_c_15(o_dac_b_c_15), .o_dac_b_c_14(o_dac_b_c_14), 
           .o_dac_b_c_13(o_dac_b_c_13), .o_dac_b_c_12(o_dac_b_c_12), .o_dac_b_c_11(o_dac_b_c_11), 
           .o_dac_b_c_10(o_dac_b_c_10), .n3639(n3639), .o_dac_b_c_8(o_dac_b_c_8)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(78[4:158])
    
endmodule
//
// Verilog Description of module dds
//

module dds (dac_clk_p_c, i_sw0_c, \addr_space[1][0] , \addr_space[1][30] , 
            \addr_space[1][29] , \addr_space[1][28] , \addr_space[1][27] , 
            \addr_space[1][26] , \addr_space[1][25] , \addr_space[1][24] , 
            \addr_space[1][23] , \addr_space[1][22] , \addr_space[1][21] , 
            \addr_space[1][20] , \addr_space[1][19] , \addr_space[1][18] , 
            \addr_space[1][17] , \addr_space[1][16] , \addr_space[1][15] , 
            \addr_space[1][14] , \addr_space[1][13] , \addr_space[1][12] , 
            \addr_space[1][11] , \addr_space[1][10] , \addr_space[1][9] , 
            \addr_space[1][8] , \addr_space[1][7] , \addr_space[1][6] , 
            \addr_space[1][5] , \addr_space[1][4] , \addr_space[1][3] , 
            \addr_space[1][2] , \addr_space[1][1] , dac_clk_p_c_enable_488, 
            modulation_output, \quarter_wave_sample_register_q[15] , GND_net) /* synthesis syn_module_defined=1 */ ;
    input dac_clk_p_c;
    input i_sw0_c;
    input \addr_space[1][0] ;
    input \addr_space[1][30] ;
    input \addr_space[1][29] ;
    input \addr_space[1][28] ;
    input \addr_space[1][27] ;
    input \addr_space[1][26] ;
    input \addr_space[1][25] ;
    input \addr_space[1][24] ;
    input \addr_space[1][23] ;
    input \addr_space[1][22] ;
    input \addr_space[1][21] ;
    input \addr_space[1][20] ;
    input \addr_space[1][19] ;
    input \addr_space[1][18] ;
    input \addr_space[1][17] ;
    input \addr_space[1][16] ;
    input \addr_space[1][15] ;
    input \addr_space[1][14] ;
    input \addr_space[1][13] ;
    input \addr_space[1][12] ;
    input \addr_space[1][11] ;
    input \addr_space[1][10] ;
    input \addr_space[1][9] ;
    input \addr_space[1][8] ;
    input \addr_space[1][7] ;
    input \addr_space[1][6] ;
    input \addr_space[1][5] ;
    input \addr_space[1][4] ;
    input \addr_space[1][3] ;
    input \addr_space[1][2] ;
    input \addr_space[1][1] ;
    input dac_clk_p_c_enable_488;
    output [15:0]modulation_output;
    input \quarter_wave_sample_register_q[15] ;
    input GND_net;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[49:58])
    wire [15:0]modulation_output_c /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(73[39:56])
    wire [30:0]increment;   // d:/documents/git_local/fm_modulator/rtl/dds.v(14[31:40])
    wire [11:0]o_phase;   // d:/documents/git_local/fm_modulator/rtl/dds.v(18[26:33])
    
    FD1S3DX increment_i0 (.D(\addr_space[1][0] ), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[0])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=83, LSE_RLINE=83 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i0.GSR = "DISABLED";
    FD1S3DX increment_i30 (.D(\addr_space[1][30] ), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[30])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=83, LSE_RLINE=83 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i30.GSR = "DISABLED";
    FD1S3DX increment_i29 (.D(\addr_space[1][29] ), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[29])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=83, LSE_RLINE=83 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i29.GSR = "DISABLED";
    FD1S3DX increment_i28 (.D(\addr_space[1][28] ), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[28])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=83, LSE_RLINE=83 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i28.GSR = "DISABLED";
    FD1S3DX increment_i27 (.D(\addr_space[1][27] ), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[27])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=83, LSE_RLINE=83 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i27.GSR = "DISABLED";
    FD1S3DX increment_i26 (.D(\addr_space[1][26] ), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[26])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=83, LSE_RLINE=83 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i26.GSR = "DISABLED";
    FD1S3DX increment_i25 (.D(\addr_space[1][25] ), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[25])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=83, LSE_RLINE=83 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i25.GSR = "DISABLED";
    FD1S3DX increment_i24 (.D(\addr_space[1][24] ), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[24])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=83, LSE_RLINE=83 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i24.GSR = "DISABLED";
    FD1S3DX increment_i23 (.D(\addr_space[1][23] ), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[23])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=83, LSE_RLINE=83 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i23.GSR = "DISABLED";
    FD1S3DX increment_i22 (.D(\addr_space[1][22] ), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[22])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=83, LSE_RLINE=83 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i22.GSR = "DISABLED";
    FD1S3DX increment_i21 (.D(\addr_space[1][21] ), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[21])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=83, LSE_RLINE=83 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i21.GSR = "DISABLED";
    FD1S3DX increment_i20 (.D(\addr_space[1][20] ), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[20])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=83, LSE_RLINE=83 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i20.GSR = "DISABLED";
    FD1S3DX increment_i19 (.D(\addr_space[1][19] ), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[19])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=83, LSE_RLINE=83 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i19.GSR = "DISABLED";
    FD1S3DX increment_i18 (.D(\addr_space[1][18] ), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[18])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=83, LSE_RLINE=83 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i18.GSR = "DISABLED";
    FD1S3DX increment_i17 (.D(\addr_space[1][17] ), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[17])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=83, LSE_RLINE=83 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i17.GSR = "DISABLED";
    FD1S3DX increment_i16 (.D(\addr_space[1][16] ), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[16])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=83, LSE_RLINE=83 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i16.GSR = "DISABLED";
    FD1S3DX increment_i15 (.D(\addr_space[1][15] ), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[15])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=83, LSE_RLINE=83 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i15.GSR = "DISABLED";
    FD1S3DX increment_i14 (.D(\addr_space[1][14] ), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[14])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=83, LSE_RLINE=83 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i14.GSR = "DISABLED";
    FD1S3DX increment_i13 (.D(\addr_space[1][13] ), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[13])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=83, LSE_RLINE=83 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i13.GSR = "DISABLED";
    FD1S3DX increment_i12 (.D(\addr_space[1][12] ), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[12])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=83, LSE_RLINE=83 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i12.GSR = "DISABLED";
    FD1S3DX increment_i11 (.D(\addr_space[1][11] ), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[11])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=83, LSE_RLINE=83 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i11.GSR = "DISABLED";
    FD1S3DX increment_i10 (.D(\addr_space[1][10] ), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[10])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=83, LSE_RLINE=83 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i10.GSR = "DISABLED";
    FD1S3DX increment_i9 (.D(\addr_space[1][9] ), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[9])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=83, LSE_RLINE=83 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i9.GSR = "DISABLED";
    FD1S3DX increment_i8 (.D(\addr_space[1][8] ), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[8])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=83, LSE_RLINE=83 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i8.GSR = "DISABLED";
    FD1S3DX increment_i7 (.D(\addr_space[1][7] ), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[7])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=83, LSE_RLINE=83 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i7.GSR = "DISABLED";
    FD1S3DX increment_i6 (.D(\addr_space[1][6] ), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[6])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=83, LSE_RLINE=83 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i6.GSR = "DISABLED";
    FD1S3DX increment_i5 (.D(\addr_space[1][5] ), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[5])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=83, LSE_RLINE=83 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i5.GSR = "DISABLED";
    FD1S3DX increment_i4 (.D(\addr_space[1][4] ), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[4])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=83, LSE_RLINE=83 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i4.GSR = "DISABLED";
    FD1S3DX increment_i3 (.D(\addr_space[1][3] ), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[3])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=83, LSE_RLINE=83 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i3.GSR = "DISABLED";
    FD1S3DX increment_i2 (.D(\addr_space[1][2] ), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[2])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=83, LSE_RLINE=83 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i2.GSR = "DISABLED";
    FD1S3DX increment_i1 (.D(\addr_space[1][1] ), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[1])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=83, LSE_RLINE=83 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i1.GSR = "DISABLED";
    quarter_wave_sine_lookup qtr_inst (.dac_clk_p_c(dac_clk_p_c), .dac_clk_p_c_enable_488(dac_clk_p_c_enable_488), 
            .o_phase({o_phase}), .i_sw0_c(i_sw0_c), .modulation_output({modulation_output}), 
            .\quarter_wave_sample_register_q[15] (\quarter_wave_sample_register_q[15] ), 
            .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(21[70:134])
    \nco(OW=12)  nco_inst (.dac_clk_p_c(dac_clk_p_c), .i_sw0_c(i_sw0_c), 
            .increment({increment}), .o_phase({o_phase}), .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(20[49:100])
    
endmodule
//
// Verilog Description of module quarter_wave_sine_lookup
//

module quarter_wave_sine_lookup (dac_clk_p_c, dac_clk_p_c_enable_488, o_phase, 
            i_sw0_c, modulation_output, \quarter_wave_sample_register_q[15] , 
            GND_net) /* synthesis syn_module_defined=1 */ ;
    input dac_clk_p_c;
    input dac_clk_p_c_enable_488;
    input [11:0]o_phase;
    input i_sw0_c;
    output [15:0]modulation_output;
    input \quarter_wave_sample_register_q[15] ;
    input GND_net;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[49:58])
    wire [15:0]modulation_output_c /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(73[39:56])
    wire [15:0]\o_val_pipeline_i[0]  /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(15[24:40])
    
    wire n23640, n23641;
    wire [9:0]index_i;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(31[17:24])
    wire [14:0]quarter_wave_sample_register_i_15__N_2145;
    
    wire n25804, n25801, n22816, n25803, n25802, n25800, n25799, 
        n23249, n23250, n23733, n23734, n723, n27404, n22254, 
        n22378, n27205, n348, n349, n27143, n27318, n14735, n204, 
        n27399, n23351, n124, n25280, n635, n14736, n636, n27408, 
        n14, n589, n526, n25282, n93, n27336, n908, n908_adj_2793, 
        n27489, n22252, n22253, n23048, n23049;
    wire [11:0]phase_i;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(11[17:24])
    
    wire n23337, n23338, n23341, n21753, n21754;
    wire [1:0]phase_negation_i;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(23[12:28])
    wire [9:0]index_i_9__N_2125;
    wire [15:0]quarter_wave_sample_register_i;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(22[24:54])
    
    wire n23339, n23340, n23342, n25743, n25742, n25744, n620, 
        n635_adj_2794, n636_adj_2795, n23344, n23345, n23348, n23346, 
        n23347, n23349, n27122, n27160, n20708, n27324, n892, 
        n20171, n23775, n23776, n23779, n22802, n22803, n23430, 
        n23461, n23368, n27326, n924, n955, n23765, n27578, n27579, 
        n62, n511, n20537, n23352, n23355, n23353, n23354, n23356, 
        n22464, n22465, n22466, n27169, n23570, n23571, n23574, 
        n23572, n23573, n23575, n23243, n23244, n23248, n22470, 
        n22471, n22472, n23753, n26283, n23768, n23358, n23359, 
        n23362, n23727, n23728, n23732, n27416, n333, n23767, 
        n23769, n23770, n23360, n23361, n23363, n27417, n348_adj_2796, 
        n397, n21912, n21913, n21914, n27571, n27572, n27573, 
        n23428, n23429, n574, n637, n21777, n23459, n23460, n23038, 
        n23039, n23045, n23040, n23041, n23046, n27395, n29957, 
        n605, n23042, n23043, n23047, n844, n12122, n23441, n23566, 
        n23567, n23568, n23569, n844_adj_2797, n23725, n23726, n23731, 
        n23715, n23716, n604, n142, n23628, n23629, n23636, n428, 
        n23630, n23631, n23637, n27329, n812, n443, n22270, n18102, 
        n21879, n23231, n23232, n23242, n23233, n23234, n23239, 
        n23240, n23246, n762, n27552, n27553, n27554, n21774, 
        n21775, n21776, n27222, n860, n25183, n27073, n15342, 
        n252, n27100, n46, n21826, n890, n27144, n189, n12018, 
        n27221, n317, n9462, n765, n404, n27370, n21993, n25683, 
        n25680, n25684, n21994, n21995, n21847, n29939, n21988, 
        n890_adj_2798, n891, n25658, n25682, n25681, n142_adj_2799, 
        n157, n158, n21984, n21985, n21986, n27421, n21982, n21981, 
        n21983, n316, n23275, n12119, n23717, n23718, n23721, 
        n23722, n23729, n23723, n23724, n23730, n844_adj_2800, n860_adj_2801, 
        n27225, n27146, n23283, n413, n412, n23281, n23771, n23772, 
        n23777, n22640, n381, n22794, n22795, n22800, n29920, 
        n252_adj_2802, n27067, n701, n24866, n21978, n21979, n21980, 
        n251, n460, n109, n22796, n22797, n22801, n93_adj_2803, 
        n23402, n21910, n22817, n24869, n22811, n24870, n15, n22809, 
        n22810, n379, n443_adj_2804, n684, n23277, n25679, n25678, 
        n716, n699, n27546, n27547, n27548, n412_adj_2805, n22359, 
        n445, n890_adj_2806, n252_adj_2807, n46_adj_2808, n23401, 
        n25661, n25659, n21800, n27196, n221, n22808, n28001, 
        n28002, n25660, n28003, n27413, n28004, n23022, n23023, 
        n23037, n23024, n23025, n28000, n23026, n23027, n27325, 
        n526_adj_2809, n542, n635_adj_2810, n21844, n25657, n23028, 
        n23029, n27999, n28005, n28006, n27543, n27544, n27545, 
        n23030, n23031, n892_adj_2811, n23350, n23357, n23562, n27337, 
        n29076, n29908, n23247, n27262, n700, n21860, n21863, 
        n23565, n21929, n21935, n684_adj_2812, n29927, n27407, n29930, 
        n22351, n27490, n27360, n26045, n731, n27376, n26054, 
        n27492, n24889, n77, n475, n25286, n23044, n27377, n22261, 
        n24890, n24895, n21938, n21941, n26056, n21944, n892_adj_2813, 
        n508, n173, n189_adj_2814, n27491, n22498, n22497, n22499, 
        n22494, n22495, n22496, n22360, n15328, n25642, n25639, 
        n25643, n23622, n23623, n23633, n25641, n27364, n27401, 
        n251_adj_2815, n444, n25638, n22489, n29933, n747, n25636, 
        n25634, n25637, n25635, n285, n620_adj_2816, n14250, n21934, 
        n25633, n25632, n325, n21931, n124_adj_2817, n21930, n21932, 
        n29917, n27402, n21925, n22323, n173_adj_2818, n27412, n25168, 
        n301, n25180, n27266, n475_adj_2819, n27398, n491, n27065, 
        n142_adj_2820, n157_adj_2821, n23404, n27369, n22486, n21928, 
        n27406, n22485, n684_adj_2822, n653, n21921, n21922, n21923, 
        n475_adj_2823, n21933, n173_adj_2824, n188, n23405, n23612, 
        n23613, n23614, n23615, n23616, n23617, n23618, n23619, 
        n23620, n23621, n23632, n23624, n23625, n23634, n21022, 
        n23643, n23644, n23659, n254, n732, n763, n22480, n22361, 
        n891_adj_2825, n38, n23645, n23646, n23660, n23647, n23648, 
        n23661, n23221, n23222, n23237, n23225, n23226, n23651, 
        n23652, n23663, n23227, n23228, n23653, n23654, n23664, 
        n23655, n23656, n23665, n23657, n23658, n23666, n23235, 
        n23236, n27331, n22479, n333_adj_2826, n348_adj_2827, n23410, 
        n364, n23411, n397_adj_2828, n23412, n23278, n23279, n23280, 
        n20104, n23285, n23286, n23287, n23413, n23414, n491_adj_2829, 
        n11349, n23415, n797, n828, n27400, n26189, n23705, n23706, 
        n23707, n23708, n23709, n23710, n23711, n23712, n23713, 
        n23714, n23719, n23720, n23759, n23760, n286, n23761, 
        n23762, n23763, n23764, n23773, n653_adj_2830, n23766, n23774, 
        n27403, n26205, n21827, n21830, n22790, n11982, n21833, 
        n22791, n190, n26581, n23563, n23364, n21857, n23564, 
        n21839, n21842, n22793, n557, n572, n23432, n574_adj_2831, 
        n21845, n21848, n764, n23433, n27534, n27535, n27536, 
        n22255, n22256, n22257, n22258, n22259, n29942, n22805, 
        n22806, n22807, n12158, n22814, n22815, n29943, n796, 
        n620_adj_2832, n635_adj_2833, n23434, n12113, n27397, n12114, 
        n26436, n23343, n22792, n653_adj_2834, n668, n23435, n699_adj_2835, 
        n23436, n716_adj_2836, n23437, n20184, n1018, n700_adj_2837, 
        n747_adj_2838, n762_adj_2839, n23438, n11192, n26281, n23416, 
        n23417, n23424, n23422, n23423, n23427, n732_adj_2840, n476, 
        n25281, n22455, n22456, n22457, n22278, n22279, n22280, 
        n28834, n28835, n23447, n23448, n23455, n875, n891_adj_2841, 
        n23449, n23450, n23456, n781, n23439, n23418, n29079, 
        n23425, n23451, n23452, n23457, n26501, n23421, n23426, 
        n25285, n859, n860_adj_2842, n21861, n23453, n23454, n23458, 
        n443_adj_2843, n21859, n412_adj_2844, n21858, n364_adj_2845, 
        n379_adj_2846, n21856, n21855, n812_adj_2847, n23440, n318, 
        n526_adj_2848, n541, n23431, n124_adj_2849, n875_adj_2850, 
        n23442, n29074, n27531, n27532, n27533, n923, n23443, 
        n25579, n27054, n23294, n25578, n25577, n939, n954, n23444, 
        n29073, n27128, n25574, n22287, n22288, n22289, n732_adj_2851, 
        n27452, n27453, n27454, n22296, n22297, n22298, n684_adj_2852, 
        n700_adj_2853, n747_adj_2854, n763_adj_2855, n541_adj_2856, 
        n23400, n24972, n24969, n158_adj_2857, n22305, n22306, n22307, 
        n221_adj_2858, n971, n986, n23445, n1002, n1017, n23446, 
        n27130, n286_adj_2859, n317_adj_2860, n349_adj_2861, n413_adj_2862, 
        n21989, n507, n21849, n21850, n21851, n21992, n573, n21877, 
        n23662, n24941, n21927, n491_adj_2863, n541_adj_2864, n21841, 
        n397_adj_2865, n475_adj_2866, n21840, n605_adj_2867, n669, 
        n21838, n732_adj_2868, n763_adj_2869, n15042, n21837, n23033, 
        n18130, n18131, n18132, n78, n93_adj_2870, n21828, n27359, 
        n24939, n22324, n22325, n21871, n27379, n460_adj_2871, n30, 
        n21825, n27396, n24942, n731_adj_2872, n732_adj_2873, n27422, 
        n26498, n21936, n21937, n24971, n24970, n27373, n61, n62_adj_2874, 
        n15_adj_2875, n31, n22341, n22342, n22343, n22350, n22352, 
        n781_adj_2876, n30_adj_2877, n31_adj_2878, n21939, n21940, 
        n21864, n21865, n21866, n27362, n890_adj_2879, n27367, n956, 
        n20737, n668_adj_2880, n763_adj_2881, n23245, n21867, n21868, 
        n21869, n11986, n30_adj_2882, n23276, n27519, n27520, n27521, 
        n27372, n573_adj_2883, n27419, n26577, n124_adj_2884, n285_adj_2885, 
        n23274, n573_adj_2886, n557_adj_2887, n890_adj_2888, n891_adj_2889, 
        n812_adj_2890, n14276, n828_adj_2891, n27511, n27076, n797_adj_2892, 
        n653_adj_2893, n668_adj_2894, n669_adj_2895, n541_adj_2896, 
        n542_adj_2897, n27112, n27119, n27510, n21972, n27564, n21974, 
        n908_adj_2898, n924_adj_2899, n891_adj_2900, n669_adj_2901, 
        n12030, n21918, n21919, n21920, n476_adj_2902, n21870, n21872, 
        n397_adj_2903, n413_adj_2904, n93_adj_2905, n15081, n286_adj_2906, 
        n21904, n21903, n21905, n142_adj_2907, n27132, n158_adj_2908, 
        n15075, n125, n21900, n27374, n21876, n21878, n25478, 
        n25479, n24968, n21898, n444_adj_2909, n25482, n27514, n908_adj_2910, 
        n924_adj_2911, n22332, n22333, n22334, n21911, n1002_adj_2912, 
        n506, n860_adj_2913, n21901, n21902, n22736, n21897, n21899, 
        n348_adj_2914, n349_adj_2915, n22260, n22262, n684_adj_2916, 
        n700_adj_2917, n21891, n668_adj_2918, n669_adj_2919, n542_adj_2920, 
        n15304, n27207, n27512, n27103, n93_adj_2921, n94, n270, 
        n286_adj_2922, n27330, n94_adj_2923, n27513, n27516, n27517, 
        n27518, n21886, n21885, n875_adj_2924, n891_adj_2925, n15_adj_2926, 
        n859_adj_2927, n860_adj_2928, n21887, n27366, n21883, n21882, 
        n21884, n21873, n21874, n21875, n27206, n636_adj_2929, n21880, 
        n21881, n18103, n18104, n491_adj_2930, n507_adj_2931, n460_adj_2932, 
        n475_adj_2933, n476_adj_2934, n397_adj_2935, n413_adj_2936, 
        n18120, n18121, n18122, n109_adj_2937, n125_adj_2938, n94_adj_2939, 
        n30_adj_2940, n31_adj_2941, n27405, n270_adj_2942, n316_adj_2943, 
        n397_adj_2944, n573_adj_2945, n605_adj_2946, n25166, n700_adj_2947, 
        n797_adj_2948, n828_adj_2949, n11985, n27515, n27171, n21843, 
        n27089, n27375, n22377, n22379, n491_adj_2950, n859_adj_2951, 
        n860_adj_2952, n221_adj_2953, n252_adj_2954, n22368, n22369, 
        n22370, n349_adj_2955, n21806, n23223, n21892, n747_adj_2956, 
        n762_adj_2957, n491_adj_2958, n506_adj_2959, n21862, n716_adj_2960, 
        n317_adj_2961, n22271, n27415, n828_adj_2962, n250, n27333, 
        n348_adj_2963, n108, n27204, n766, n27083, n986_adj_2964, 
        n1021, n23230, n716_adj_2965, n731_adj_2966, n653_adj_2967, 
        n604_adj_2968, n954_adj_2969, n526_adj_2970, n27577, n21991, 
        n21987, n987, n985, n14323, n20892, n254_adj_2971, n27418, 
        n125_adj_2972, n27063, n23282, n22269, n27378, n23284, n94_adj_2973, 
        n924_adj_2974, n27129, n21917, n444_adj_2975, n507_adj_2976, 
        n700_adj_2977, n21926, n101, n26053, n22798, n22799, n25741, 
        n23752, n22481, n23756, n22487, n11994, n23757, n573_adj_2978, 
        n27265, n21909, n26580, n26578, n796_adj_2979, n26579, n882, 
        n890_adj_2980, n21943, n11987, n22459, n27368, n23780, n23778;
    wire [15:0]o_val_pipeline_i_0__15__N_2176;
    wire [15:0]n1087;
    
    wire n27481, n23403, n62_adj_2981, n684_adj_2982, n638, n17958, 
        n26500, n26497, n26499, n24943, n24940, n26082, n205, 
        n26282, n26496, n17957, n21829, n24867, n24868, n23034, 
        n26058, n26435, n26432, n23670, n26434, n26433, n205_adj_2983, 
        n157_adj_2984, n26431, n348_adj_2985, n173_adj_2986, n29075, 
        n12034, n21916, n21915, n25170, n23639, n572_adj_2987, n23638, 
        n21846, n716_adj_2988, n26080, n12157, n221_adj_2989, n26192, 
        n23238, n491_adj_2990, n27493, n17956, n17955, n26194, n1022, 
        n62_adj_2991, n17954, n23241, n26207, n17953, n26047, n17952, 
        n26206, n26203, n26204, n17951, n26202, n27101, n26193, 
        n26191, n572_adj_2992, n26190, n189_adj_2993, n25185, n25184, 
        n21924, n26044, n25169, n25167, n924_adj_2994, n26081, n26057, 
        n26055, n22735, n26042, n26046, n26043, n27077;
    
    PFUMX i21268 (.BLUT(n23640), .ALUT(n23641), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2145[5]));
    L6MUX21 i24092 (.D0(n25804), .D1(n25801), .SD(index_i[6]), .Z(n22816));
    PFUMX i24090 (.BLUT(n25803), .ALUT(n25802), .C0(index_i[5]), .Z(n25804));
    PFUMX i24088 (.BLUT(n25800), .ALUT(n25799), .C0(index_i[5]), .Z(n25801));
    LUT4 n428_bdd_2_lut_24094_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[4]), .D(index_i[1]), .Z(n25800)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n428_bdd_2_lut_24094_3_lut_4_lut.init = 16'h0f1f;
    LUT4 n557_bdd_2_lut_24268_3_lut (.A(index_i[2]), .B(index_i[3]), .C(index_i[4]), 
         .Z(n25803)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n557_bdd_2_lut_24268_3_lut.init = 16'he0e0;
    PFUMX i20877 (.BLUT(n23249), .ALUT(n23250), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2145[1]));
    PFUMX i21361 (.BLUT(n23733), .ALUT(n23734), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2145[3]));
    LUT4 i19899_3_lut (.A(n723), .B(n27404), .C(index_i[3]), .Z(n22254)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19899_3_lut.init = 16'hcaca;
    LUT4 i20023_3_lut_4_lut_3_lut (.A(index_i[1]), .B(index_i[3]), .C(index_i[2]), 
         .Z(n22378)) /* synthesis lut_function=(A (B)+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20023_3_lut_4_lut_3_lut.init = 16'hd9d9;
    LUT4 i11558_2_lut_rep_540_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[3]), 
         .Z(n27205)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11558_2_lut_rep_540_3_lut.init = 16'he0e0;
    LUT4 mux_231_Mux_3_i349_3_lut_3_lut (.A(index_i[1]), .B(index_i[4]), 
         .C(n348), .Z(n349)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_3_i349_3_lut_3_lut.init = 16'hd1d1;
    LUT4 i11991_2_lut_rep_478_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[0]), 
         .Z(n27143)) /* synthesis lut_function=(A (C)+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11991_2_lut_rep_478_3_lut.init = 16'hf1f1;
    LUT4 i12137_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(n27318), .C(index_i[4]), 
         .D(index_i[0]), .Z(n14735)) /* synthesis lut_function=(!(A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12137_3_lut_4_lut_4_lut_4_lut.init = 16'h55d5;
    LUT4 i20977_3_lut (.A(n204), .B(n27399), .C(index_i[3]), .Z(n23351)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20977_3_lut.init = 16'hcaca;
    LUT4 n476_bdd_3_lut_23767_3_lut (.A(index_i[1]), .B(index_i[4]), .C(n124), 
         .Z(n25280)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n476_bdd_3_lut_23767_3_lut.init = 16'hd1d1;
    LUT4 mux_231_Mux_6_i636_4_lut_4_lut (.A(index_i[1]), .B(index_i[4]), 
         .C(n635), .D(n14736), .Z(n636)) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_6_i636_4_lut_4_lut.init = 16'hf3d1;
    LUT4 mux_231_Mux_0_i589_3_lut (.A(n27408), .B(n14), .C(index_i[3]), 
         .Z(n589)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_0_i589_3_lut.init = 16'hcaca;
    LUT4 n21976_bdd_3_lut_3_lut (.A(index_i[1]), .B(n526), .C(index_i[4]), 
         .Z(n25282)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n21976_bdd_3_lut_3_lut.init = 16'h5c5c;
    LUT4 mux_231_Mux_9_i93_3_lut_3_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .Z(n93)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_9_i93_3_lut_3_lut_3_lut.init = 16'hc1c1;
    LUT4 i11577_2_lut_rep_671 (.A(index_i[2]), .B(index_i[3]), .Z(n27336)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11577_2_lut_rep_671.init = 16'heeee;
    LUT4 mux_231_Mux_2_i908_3_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .D(index_i[3]), .Z(n908)) /* synthesis lut_function=(!(A (B+!(D))+!A !(B+!(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_2_i908_3_lut_4_lut_4_lut.init = 16'h6645;
    LUT4 mux_231_Mux_0_i908_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n908_adj_2793)) /* synthesis lut_function=(!(A (B (C (D))+!B !(D))+!A (B+((D)+!C)))) */ ;
    defparam mux_231_Mux_0_i908_3_lut_4_lut_4_lut.init = 16'h2a98;
    LUT4 i22293_3_lut (.A(n27489), .B(n22252), .C(index_i[4]), .Z(n22253)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22293_3_lut.init = 16'hcaca;
    PFUMX i20676 (.BLUT(n23048), .ALUT(n23049), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2145[2]));
    FD1P3AX phase_i_i0_i0 (.D(o_phase[0]), .SP(dac_clk_p_c_enable_488), 
            .CK(dac_clk_p_c), .Q(phase_i[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam phase_i_i0_i0.GSR = "DISABLED";
    PFUMX i20967 (.BLUT(n23337), .ALUT(n23338), .C0(index_i[4]), .Z(n23341));
    PFUMX i19400 (.BLUT(n21753), .ALUT(n21754), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2145[11]));
    FD1S3DX phase_negation_i_i0 (.D(phase_i[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(phase_negation_i[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam phase_negation_i_i0.GSR = "DISABLED";
    FD1S3DX index_i_i0 (.D(index_i_9__N_2125[0]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(index_i[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam index_i_i0.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i1 (.D(\o_val_pipeline_i[0] [0]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(modulation_output[0])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i1.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i0 (.D(quarter_wave_sample_register_i_15__N_2145[0]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_i[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_i_i0.GSR = "DISABLED";
    PFUMX i20968 (.BLUT(n23339), .ALUT(n23340), .C0(index_i[4]), .Z(n23342));
    PFUMX i24031 (.BLUT(n25743), .ALUT(n25742), .C0(index_i[5]), .Z(n25744));
    PFUMX mux_231_Mux_1_i636 (.BLUT(n620), .ALUT(n635_adj_2794), .C0(index_i[4]), 
          .Z(n636_adj_2795)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    PFUMX i20974 (.BLUT(n23344), .ALUT(n23345), .C0(index_i[4]), .Z(n23348));
    PFUMX i20975 (.BLUT(n23346), .ALUT(n23347), .C0(index_i[4]), .Z(n23349));
    LUT4 i11559_2_lut_rep_457_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[4]), .D(index_i[3]), .Z(n27122)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11559_2_lut_rep_457_3_lut_4_lut.init = 16'hfef0;
    LUT4 i1_4_lut (.A(index_i[6]), .B(n27160), .C(index_i[5]), .D(index_i[4]), 
         .Z(n20708)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_4_lut.init = 16'hfffe;
    LUT4 i17961_4_lut (.A(n27324), .B(n892), .C(index_i[6]), .D(index_i[5]), 
         .Z(n20171)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D))))) */ ;
    defparam i17961_4_lut.init = 16'h3a35;
    FD1P3AX phase_i_i0_i11 (.D(o_phase[11]), .SP(dac_clk_p_c_enable_488), 
            .CK(dac_clk_p_c), .Q(phase_i[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam phase_i_i0_i11.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i10 (.D(o_phase[10]), .SP(dac_clk_p_c_enable_488), 
            .CK(dac_clk_p_c), .Q(phase_i[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam phase_i_i0_i10.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i9 (.D(o_phase[9]), .SP(dac_clk_p_c_enable_488), 
            .CK(dac_clk_p_c), .Q(phase_i[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam phase_i_i0_i9.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i8 (.D(o_phase[8]), .SP(dac_clk_p_c_enable_488), 
            .CK(dac_clk_p_c), .Q(phase_i[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam phase_i_i0_i8.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i7 (.D(o_phase[7]), .SP(dac_clk_p_c_enable_488), 
            .CK(dac_clk_p_c), .Q(phase_i[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam phase_i_i0_i7.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i6 (.D(o_phase[6]), .SP(dac_clk_p_c_enable_488), 
            .CK(dac_clk_p_c), .Q(phase_i[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam phase_i_i0_i6.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i5 (.D(o_phase[5]), .SP(dac_clk_p_c_enable_488), 
            .CK(dac_clk_p_c), .Q(phase_i[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam phase_i_i0_i5.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i4 (.D(o_phase[4]), .SP(dac_clk_p_c_enable_488), 
            .CK(dac_clk_p_c), .Q(phase_i[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam phase_i_i0_i4.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i3 (.D(o_phase[3]), .SP(dac_clk_p_c_enable_488), 
            .CK(dac_clk_p_c), .Q(phase_i[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam phase_i_i0_i3.GSR = "DISABLED";
    L6MUX21 i21405 (.D0(n23775), .D1(n23776), .SD(index_i[8]), .Z(n23779));
    PFUMX i20430 (.BLUT(n22802), .ALUT(n22803), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2145[8]));
    FD1P3AX phase_i_i0_i2 (.D(o_phase[2]), .SP(dac_clk_p_c_enable_488), 
            .CK(dac_clk_p_c), .Q(phase_i[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam phase_i_i0_i2.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i1 (.D(o_phase[1]), .SP(dac_clk_p_c_enable_488), 
            .CK(dac_clk_p_c), .Q(phase_i[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam phase_i_i0_i1.GSR = "DISABLED";
    L6MUX21 i13238356_i1 (.D0(n23430), .D1(n23461), .SD(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2145[0]));
    LUT4 i22841_3_lut (.A(n20171), .B(n20708), .C(index_i[7]), .Z(n23368)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22841_3_lut.init = 16'hcaca;
    LUT4 i7076_2_lut_rep_661 (.A(index_i[3]), .B(index_i[4]), .Z(n27326)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i7076_2_lut_rep_661.init = 16'heeee;
    LUT4 i22594_3_lut (.A(n924), .B(n955), .C(index_i[5]), .Z(n23765)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22594_3_lut.init = 16'hcaca;
    PFUMX i25224 (.BLUT(n27578), .ALUT(n27579), .C0(index_i[3]), .Z(n62));
    PFUMX mux_231_Mux_13_i1023 (.BLUT(n511), .ALUT(n20537), .C0(index_i[9]), 
          .Z(quarter_wave_sample_register_i_15__N_2145[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    PFUMX i20981 (.BLUT(n23351), .ALUT(n23352), .C0(index_i[4]), .Z(n23355));
    PFUMX i20982 (.BLUT(n23353), .ALUT(n23354), .C0(index_i[4]), .Z(n23356));
    PFUMX i20111 (.BLUT(n22464), .ALUT(n22465), .C0(index_i[4]), .Z(n22466));
    LUT4 i12048_2_lut_rep_504_3_lut (.A(index_i[2]), .B(index_i[3]), .C(index_i[1]), 
         .Z(n27169)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12048_2_lut_rep_504_3_lut.init = 16'hfefe;
    PFUMX i21200 (.BLUT(n23570), .ALUT(n23571), .C0(index_i[8]), .Z(n23574));
    L6MUX21 i21201 (.D0(n23572), .D1(n23573), .SD(index_i[8]), .Z(n23575));
    L6MUX21 i20874 (.D0(n23243), .D1(n23244), .SD(index_i[7]), .Z(n23248));
    PFUMX i20117 (.BLUT(n22470), .ALUT(n22471), .C0(index_i[4]), .Z(n22472));
    LUT4 i22844_3_lut (.A(n23753), .B(n26283), .C(index_i[6]), .Z(n23768)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22844_3_lut.init = 16'hcaca;
    PFUMX i20988 (.BLUT(n23358), .ALUT(n23359), .C0(index_i[4]), .Z(n23362));
    L6MUX21 i21358 (.D0(n23727), .D1(n23728), .SD(index_i[7]), .Z(n23732));
    LUT4 mux_231_Mux_7_i333_3_lut (.A(n27416), .B(n204), .C(index_i[3]), 
         .Z(n333)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_7_i333_3_lut.init = 16'hcaca;
    PFUMX i21401 (.BLUT(n23767), .ALUT(n23768), .C0(index_i[7]), .Z(n23775));
    PFUMX i21402 (.BLUT(n23769), .ALUT(n23770), .C0(index_i[7]), .Z(n23776));
    PFUMX i20989 (.BLUT(n23360), .ALUT(n23361), .C0(index_i[4]), .Z(n23363));
    LUT4 mux_231_Mux_7_i348_3_lut (.A(n27417), .B(n27408), .C(index_i[3]), 
         .Z(n348_adj_2796)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_7_i348_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_7_i397_3_lut (.A(n27417), .B(n27416), .C(index_i[3]), 
         .Z(n397)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_7_i397_3_lut.init = 16'hcaca;
    LUT4 i22238_3_lut (.A(n21912), .B(n21913), .C(index_i[4]), .Z(n21914)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22238_3_lut.init = 16'hcaca;
    PFUMX i25219 (.BLUT(n27571), .ALUT(n27572), .C0(index_i[0]), .Z(n27573));
    PFUMX i21056 (.BLUT(n23428), .ALUT(n23429), .C0(index_i[8]), .Z(n23430));
    LUT4 i22923_3_lut (.A(n574), .B(n637), .C(index_i[6]), .Z(n21777)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22923_3_lut.init = 16'hcaca;
    PFUMX i21087 (.BLUT(n23459), .ALUT(n23460), .C0(index_i[8]), .Z(n23461));
    L6MUX21 i20671 (.D0(n23038), .D1(n23039), .SD(index_i[7]), .Z(n23045));
    L6MUX21 i20672 (.D0(n23040), .D1(n23041), .SD(index_i[7]), .Z(n23046));
    LUT4 i9514_3_lut_4_lut (.A(index_i[3]), .B(index_i[4]), .C(n27395), 
         .D(n29957), .Z(n605)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9514_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i20673 (.BLUT(n23042), .ALUT(n23043), .C0(index_i[7]), .Z(n23047));
    PFUMX i21067 (.BLUT(n844), .ALUT(n12122), .C0(index_i[4]), .Z(n23441));
    L6MUX21 i21198 (.D0(n23566), .D1(n23567), .SD(index_i[7]), .Z(n23572));
    L6MUX21 i21199 (.D0(n23568), .D1(n23569), .SD(index_i[7]), .Z(n23573));
    LUT4 i9551_3_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[3]), .C(index_i[0]), 
         .D(index_i[1]), .Z(n844_adj_2797)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9551_3_lut_4_lut_4_lut.init = 16'hf00e;
    LUT4 i21357_3_lut (.A(n23725), .B(n23726), .C(index_i[7]), .Z(n23731)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21357_3_lut.init = 16'hcaca;
    LUT4 i21352_3_lut (.A(n23715), .B(n23716), .C(index_i[6]), .Z(n23726)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21352_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_0_i604_3_lut_4_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[1]), .D(index_i[3]), .Z(n604)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A !(B (D)+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_0_i604_3_lut_4_lut_4_lut_4_lut.init = 16'h5439;
    LUT4 mux_231_Mux_2_i142_3_lut_4_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n142)) /* synthesis lut_function=(!(A (B+(C))+!A !(B+(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_2_i142_3_lut_4_lut_4_lut_4_lut.init = 16'h5646;
    L6MUX21 i21262 (.D0(n23628), .D1(n23629), .SD(index_i[7]), .Z(n23636));
    LUT4 mux_231_Mux_0_i428_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[2]), 
         .B(index_i[0]), .C(index_i[1]), .D(index_i[3]), .Z(n428)) /* synthesis lut_function=(A (B (C+!(D))+!B !((D)+!C))+!A (B (D)+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_0_i428_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hd5a9;
    L6MUX21 i21263 (.D0(n23630), .D1(n23631), .SD(index_i[7]), .Z(n23637));
    LUT4 mux_231_Mux_4_i236_3_lut_4_lut_3_lut_rep_664_4_lut (.A(index_i[0]), 
         .B(index_i[3]), .C(index_i[1]), .D(index_i[2]), .Z(n27329)) /* synthesis lut_function=(A (B)+!A !(B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_4_i236_3_lut_4_lut_3_lut_rep_664_4_lut.init = 16'h999d;
    LUT4 mux_231_Mux_4_i812_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[4]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n812)) /* synthesis lut_function=(A (B (C+(D)))+!A !(B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_4_i812_3_lut_3_lut_4_lut.init = 16'h9995;
    LUT4 mux_231_Mux_0_i443_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n443)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (D))+!A !(B (D)+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_0_i443_3_lut_4_lut_4_lut_4_lut.init = 16'h54b3;
    LUT4 i19915_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n22270)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(D))+!A (B (D)+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19915_3_lut_4_lut_4_lut_4_lut.init = 16'hd52b;
    LUT4 i15916_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[1]), .Z(n18102)) /* synthesis lut_function=(A (B (C (D))+!B !(C))+!A (B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i15916_3_lut_4_lut_4_lut_4_lut.init = 16'hd656;
    LUT4 i19524_3_lut_4_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[3]), 
         .C(index_i[1]), .D(index_i[2]), .Z(n21879)) /* synthesis lut_function=(!(A (B)+!A !(B (C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19524_3_lut_4_lut_3_lut_4_lut.init = 16'h6662;
    L6MUX21 i20868 (.D0(n23231), .D1(n23232), .SD(index_i[6]), .Z(n23242));
    L6MUX21 i20869 (.D0(n23233), .D1(n23234), .SD(index_i[6]), .Z(n23243));
    L6MUX21 i20872 (.D0(n23239), .D1(n23240), .SD(index_i[7]), .Z(n23246));
    LUT4 i9546_3_lut_3_lut_4_lut_4_lut (.A(index_i[3]), .B(index_i[2]), 
         .C(index_i[0]), .D(index_i[1]), .Z(n762)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C (D)+!C !(D)))+!A !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9546_3_lut_3_lut_4_lut_4_lut.init = 16'h700f;
    PFUMX i25206 (.BLUT(n27552), .ALUT(n27553), .C0(index_i[8]), .Z(n27554));
    L6MUX21 i19421 (.D0(n21774), .D1(n21775), .SD(index_i[7]), .Z(n21776));
    LUT4 mux_231_Mux_8_i860_3_lut_4_lut (.A(n27222), .B(index_i[3]), .C(index_i[4]), 
         .D(n27160), .Z(n860)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_8_i860_3_lut_4_lut.init = 16'h08f8;
    LUT4 index_i_4__bdd_3_lut_23531_4_lut (.A(n27222), .B(index_i[3]), .C(index_i[5]), 
         .D(index_i[4]), .Z(n25183)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam index_i_4__bdd_3_lut_23531_4_lut.init = 16'hf080;
    LUT4 n557_bdd_3_lut_24267_4_lut (.A(n27222), .B(index_i[3]), .C(index_i[4]), 
         .D(n27160), .Z(n25802)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n557_bdd_3_lut_24267_4_lut.init = 16'hf707;
    LUT4 mux_231_Mux_6_i955_3_lut_4_lut (.A(n27222), .B(index_i[3]), .C(index_i[4]), 
         .D(n27073), .Z(n955)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_6_i955_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_231_Mux_3_i252_3_lut_4_lut (.A(n27222), .B(index_i[3]), .C(index_i[4]), 
         .D(n15342), .Z(n252)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_3_i252_3_lut_4_lut.init = 16'h08f8;
    LUT4 i19471_3_lut_3_lut (.A(n27100), .B(index_i[4]), .C(n46), .Z(n21826)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam i19471_3_lut_3_lut.init = 16'h7474;
    LUT4 mux_231_Mux_2_i890_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n890)) /* synthesis lut_function=(A (B (C)+!B !(C+!(D)))+!A !(B (C+(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_2_i890_3_lut_4_lut_4_lut.init = 16'h9394;
    LUT4 mux_231_Mux_3_i189_3_lut_3_lut_4_lut (.A(n27222), .B(index_i[3]), 
         .C(index_i[4]), .D(n27144), .Z(n189)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_3_i189_3_lut_3_lut_4_lut.init = 16'h08f8;
    LUT4 i9532_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n12018)) /* synthesis lut_function=(!(A (B (C)+!B ((D)+!C))+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9532_3_lut_4_lut_4_lut.init = 16'h4969;
    LUT4 mux_231_Mux_10_i317_3_lut_3_lut_4_lut (.A(n27221), .B(index_i[3]), 
         .C(n27144), .D(index_i[4]), .Z(n317)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_10_i317_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 i11543_3_lut_4_lut (.A(n27221), .B(index_i[3]), .C(n9462), .D(index_i[6]), 
         .Z(n765)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11543_3_lut_4_lut.init = 16'hffe0;
    LUT4 i19638_3_lut (.A(n404), .B(n27370), .C(index_i[3]), .Z(n21993)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19638_3_lut.init = 16'hcaca;
    L6MUX21 i23972 (.D0(n25683), .D1(n25680), .SD(index_i[5]), .Z(n25684));
    LUT4 i22453_3_lut (.A(n21993), .B(n21994), .C(index_i[4]), .Z(n21995)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22453_3_lut.init = 16'hcaca;
    LUT4 i19492_3_lut_3_lut_4_lut (.A(n27221), .B(index_i[3]), .C(n93), 
         .D(index_i[4]), .Z(n21847)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19492_3_lut_3_lut_4_lut.init = 16'h11f0;
    LUT4 i19633_3_lut (.A(n404), .B(n29939), .C(index_i[3]), .Z(n21988)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19633_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_7_i891_3_lut_4_lut (.A(n27221), .B(index_i[3]), .C(index_i[4]), 
         .D(n890_adj_2798), .Z(n891)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_7_i891_3_lut_4_lut.init = 16'hfe0e;
    LUT4 n124_bdd_3_lut_4_lut (.A(n27221), .B(index_i[3]), .C(index_i[4]), 
         .D(n93), .Z(n25658)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n124_bdd_3_lut_4_lut.init = 16'hfe0e;
    PFUMX i23970 (.BLUT(n25682), .ALUT(n25681), .C0(index_i[4]), .Z(n25683));
    LUT4 mux_231_Mux_4_i158_3_lut (.A(n142_adj_2799), .B(n157), .C(index_i[4]), 
         .Z(n158)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_4_i158_3_lut.init = 16'hcaca;
    LUT4 i22460_3_lut (.A(n21984), .B(n21985), .C(index_i[4]), .Z(n21986)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22460_3_lut.init = 16'hcaca;
    LUT4 i19627_3_lut (.A(n29939), .B(n27421), .C(index_i[3]), .Z(n21982)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19627_3_lut.init = 16'hcaca;
    LUT4 i22462_3_lut (.A(n21981), .B(n21982), .C(index_i[4]), .Z(n21983)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22462_3_lut.init = 16'hcaca;
    LUT4 i20901_3_lut_3_lut_4_lut (.A(n27221), .B(index_i[3]), .C(n316), 
         .D(index_i[4]), .Z(n23275)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20901_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 i9633_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n12119)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))+!A !(B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9633_3_lut_4_lut_4_lut.init = 16'hb5b3;
    LUT4 i9636_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n12122)) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B ((D)+!C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9636_3_lut_4_lut_4_lut.init = 16'hcdad;
    L6MUX21 i21353 (.D0(n23717), .D1(n23718), .SD(index_i[6]), .Z(n23727));
    L6MUX21 i21355 (.D0(n23721), .D1(n23722), .SD(index_i[7]), .Z(n23729));
    L6MUX21 i21356 (.D0(n23723), .D1(n23724), .SD(index_i[7]), .Z(n23730));
    LUT4 mux_231_Mux_6_i860_3_lut_3_lut (.A(n27100), .B(index_i[4]), .C(n844_adj_2800), 
         .Z(n860_adj_2801)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam mux_231_Mux_6_i860_3_lut_3_lut.init = 16'h7474;
    LUT4 i20909_3_lut_4_lut (.A(n27225), .B(index_i[3]), .C(index_i[4]), 
         .D(n27146), .Z(n23283)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20909_3_lut_4_lut.init = 16'hfe0e;
    LUT4 mux_231_Mux_10_i413_3_lut_3_lut_4_lut (.A(n27225), .B(index_i[3]), 
         .C(n27144), .D(index_i[4]), .Z(n413)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_10_i413_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 i20907_3_lut_3_lut_4_lut (.A(n27225), .B(index_i[3]), .C(n412), 
         .D(index_i[4]), .Z(n23281)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20907_3_lut_3_lut_4_lut.init = 16'hf011;
    L6MUX21 i21403 (.D0(n23771), .D1(n23772), .SD(index_i[7]), .Z(n23777));
    LUT4 i23127_2_lut (.A(index_i[5]), .B(index_i[4]), .Z(n22640)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i23127_2_lut.init = 16'heeee;
    LUT4 i12794_1_lut_2_lut_3_lut_4_lut (.A(n27225), .B(index_i[3]), .C(index_i[5]), 
         .D(index_i[4]), .Z(n381)) /* synthesis lut_function=(!(A (C+(D))+!A (B (C+(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12794_1_lut_2_lut_3_lut_4_lut.init = 16'h010f;
    L6MUX21 i20426 (.D0(n22794), .D1(n22795), .SD(index_i[7]), .Z(n22800));
    LUT4 mux_231_Mux_10_i252_3_lut_4_lut_4_lut (.A(n27225), .B(index_i[3]), 
         .C(index_i[4]), .D(n29920), .Z(n252_adj_2802)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B (C (D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_10_i252_3_lut_4_lut_4_lut.init = 16'h3efe;
    LUT4 n21777_bdd_3_lut_25067 (.A(n27067), .B(n701), .C(index_i[6]), 
         .Z(n24866)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n21777_bdd_3_lut_25067.init = 16'hacac;
    LUT4 i22465_3_lut (.A(n21978), .B(n21979), .C(index_i[4]), .Z(n21980)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22465_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_8_i251_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[2]), .D(index_i[3]), .Z(n251)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_8_i251_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h07e0;
    LUT4 mux_231_Mux_8_i61_3_lut_rep_435_4_lut_4_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[2]), .D(index_i[3]), .Z(n27100)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A (B (C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_8_i61_3_lut_rep_435_4_lut_4_lut_4_lut.init = 16'he0f8;
    LUT4 mux_231_Mux_0_i460_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n460)) /* synthesis lut_function=(A (B+(C (D)+!C !(D)))+!A (B (C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_0_i460_3_lut_4_lut_4_lut.init = 16'hf8cb;
    LUT4 mux_231_Mux_8_i109_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n109)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C+!(D)))+!A (B (C (D)+!C !(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_8_i109_3_lut_4_lut_4_lut.init = 16'hf83e;
    LUT4 i20966_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n23340)) /* synthesis lut_function=(A (B (C+!(D))+!B !((D)+!C))+!A !(B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20966_3_lut_4_lut_4_lut.init = 16'h81f8;
    LUT4 i20964_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n23338)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20964_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hf81f;
    PFUMX i20427 (.BLUT(n22796), .ALUT(n22797), .C0(index_i[7]), .Z(n22801));
    LUT4 i21028_3_lut_3_lut_4_lut (.A(n29920), .B(index_i[3]), .C(n93_adj_2803), 
         .D(index_i[4]), .Z(n23402)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21028_3_lut_3_lut_4_lut.init = 16'hf077;
    LUT4 i19555_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n21910)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C))+!A (B (C)+!B !((D)+!C))) */ ;
    defparam i19555_3_lut_4_lut_4_lut_4_lut.init = 16'he078;
    LUT4 i20965_3_lut_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n23339)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C+!(D))+!B !((D)+!C)))) */ ;
    defparam i20965_3_lut_3_lut_4_lut_4_lut.init = 16'h1f81;
    LUT4 n22811_bdd_3_lut (.A(n22816), .B(n22817), .C(index_i[7]), .Z(n24869)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n22811_bdd_3_lut.init = 16'hcaca;
    LUT4 n24869_bdd_3_lut (.A(n24869), .B(n22811), .C(index_i[8]), .Z(n24870)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n24869_bdd_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_8_i15_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n15)) /* synthesis lut_function=(A (B (C)+!B !(C (D)+!C !(D)))+!A !(B ((D)+!C)+!B (C+!(D)))) */ ;
    defparam mux_231_Mux_8_i15_3_lut_4_lut_4_lut.init = 16'h83e0;
    L6MUX21 i20437 (.D0(n22809), .D1(n22810), .SD(index_i[7]), .Z(n22811));
    LUT4 mux_231_Mux_0_i379_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n379)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !((D)+!C))+!A !(B ((D)+!C)+!B (D))) */ ;
    defparam mux_231_Mux_0_i379_3_lut_4_lut_4_lut.init = 16'h8079;
    LUT4 mux_231_Mux_8_i443_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n443_adj_2804)) /* synthesis lut_function=(A (B (C+!(D))+!B !((D)+!C))+!A !(B (D)+!B ((D)+!C))) */ ;
    defparam mux_231_Mux_8_i443_3_lut_4_lut_4_lut.init = 16'h80fc;
    LUT4 i20116_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n22471)) /* synthesis lut_function=(A (C)+!A !(B (C)+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20116_3_lut_4_lut_4_lut.init = 16'hb4b5;
    LUT4 mux_231_Mux_1_i684_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n684)) /* synthesis lut_function=(A (B ((D)+!C)+!B !((D)+!C))+!A !(B (C+(D))+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_1_i684_3_lut_4_lut_4_lut.init = 16'h992d;
    LUT4 i20903_3_lut_4_lut_4_lut (.A(n27225), .B(index_i[3]), .C(n27222), 
         .D(index_i[4]), .Z(n23277)) /* synthesis lut_function=(A (B (C (D))+!B !((D)+!C))+!A (B (C+!(D))+!B !((D)+!C))) */ ;
    defparam i20903_3_lut_4_lut_4_lut.init = 16'hc074;
    PFUMX i23967 (.BLUT(n25679), .ALUT(n25678), .C0(index_i[4]), .Z(n25680));
    LUT4 mux_231_Mux_1_i716_3_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[1]), .D(index_i[3]), .Z(n716)) /* synthesis lut_function=(!(A (B (D)+!B !(C))+!A !(B (C (D))+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_1_i716_3_lut_4_lut_4_lut.init = 16'h70a9;
    LUT4 mux_231_Mux_7_i699_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n699)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C+!(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_7_i699_3_lut_4_lut_4_lut.init = 16'hf07e;
    PFUMX i25202 (.BLUT(n27546), .ALUT(n27547), .C0(index_i[1]), .Z(n27548));
    LUT4 mux_231_Mux_0_i412_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n412_adj_2805)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(D))+!A (B (D)+!B !(C+!(D)))) */ ;
    defparam mux_231_Mux_0_i412_3_lut_4_lut_4_lut.init = 16'hcd2a;
    LUT4 i20004_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n22359)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B+(C+(D))))) */ ;
    defparam i20004_3_lut_4_lut_4_lut_4_lut.init = 16'h2aab;
    LUT4 mux_231_Mux_11_i445_3_lut_4_lut_4_lut_4_lut (.A(index_i[3]), .B(index_i[4]), 
         .C(index_i[5]), .D(n27225), .Z(n445)) /* synthesis lut_function=(!(A (B (C))+!A !(B+(C+(D))))) */ ;
    defparam mux_231_Mux_11_i445_3_lut_4_lut_4_lut_4_lut.init = 16'h7f7e;
    LUT4 mux_231_Mux_0_i890_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n890_adj_2806)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)+!C !(D)))+!A !(B (C)+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_0_i890_3_lut_4_lut_4_lut.init = 16'h70ca;
    LUT4 mux_231_Mux_5_i252_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[4]), .Z(n252_adj_2807)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+(D)))+!A (B (C (D))+!B !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_5_i252_3_lut_4_lut.init = 16'hc993;
    LUT4 i21027_3_lut_4_lut (.A(n29920), .B(index_i[3]), .C(index_i[4]), 
         .D(n46_adj_2808), .Z(n23401)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21027_3_lut_4_lut.init = 16'h8f80;
    L6MUX21 i23952 (.D0(n25661), .D1(n25659), .SD(index_i[6]), .Z(n21800));
    LUT4 mux_231_Mux_3_i221_3_lut_4_lut (.A(n29920), .B(index_i[3]), .C(index_i[4]), 
         .D(n27196), .Z(n221)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_3_i221_3_lut_4_lut.init = 16'h08f8;
    LUT4 i20434_3_lut_4_lut_4_lut (.A(n27146), .B(index_i[4]), .C(index_i[5]), 
         .D(n27144), .Z(n22808)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C)+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20434_3_lut_4_lut_4_lut.init = 16'h0434;
    LUT4 index_i_5__bdd_3_lut_25666 (.A(index_i[5]), .B(n28001), .C(index_i[3]), 
         .Z(n28002)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam index_i_5__bdd_3_lut_25666.init = 16'hcaca;
    PFUMX i23950 (.BLUT(n25660), .ALUT(n62), .C0(index_i[5]), .Z(n25661));
    LUT4 n27413_bdd_3_lut_25605 (.A(n27221), .B(index_i[6]), .C(index_i[5]), 
         .Z(n28003)) /* synthesis lut_function=(!(A (B)+!A (C))) */ ;
    defparam n27413_bdd_3_lut_25605.init = 16'h2727;
    LUT4 n27413_bdd_4_lut_25519 (.A(n27413), .B(index_i[6]), .C(index_i[2]), 
         .D(index_i[5]), .Z(n28004)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A !(B (C+(D))+!B (D)))) */ ;
    defparam n27413_bdd_4_lut_25519.init = 16'h5fe0;
    L6MUX21 i20663 (.D0(n23022), .D1(n23023), .SD(index_i[6]), .Z(n23037));
    L6MUX21 i20664 (.D0(n23024), .D1(n23025), .SD(index_i[6]), .Z(n23038));
    LUT4 index_i_6__bdd_4_lut_25566 (.A(index_i[6]), .B(index_i[5]), .C(index_i[1]), 
         .D(index_i[0]), .Z(n28000)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C))+!A (B (C)+!B !(C)))) */ ;
    defparam index_i_6__bdd_4_lut_25566.init = 16'h3cbc;
    L6MUX21 i20665 (.D0(n23026), .D1(n23027), .SD(index_i[6]), .Z(n23039));
    LUT4 mux_231_Mux_8_i542_3_lut_4_lut (.A(n27325), .B(index_i[3]), .C(index_i[4]), 
         .D(n526_adj_2809), .Z(n542)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_8_i542_3_lut_4_lut.init = 16'h6f60;
    LUT4 i19489_3_lut_4_lut (.A(n27325), .B(index_i[3]), .C(index_i[4]), 
         .D(n635_adj_2810), .Z(n21844)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19489_3_lut_4_lut.init = 16'hf606;
    PFUMX i23948 (.BLUT(n25658), .ALUT(n25657), .C0(index_i[5]), .Z(n25659));
    L6MUX21 i20666 (.D0(n23028), .D1(n23029), .SD(index_i[6]), .Z(n23040));
    LUT4 index_i_6__bdd_1_lut_25663 (.A(index_i[5]), .Z(n27999)) /* synthesis lut_function=(!(A)) */ ;
    defparam index_i_6__bdd_1_lut_25663.init = 16'h5555;
    LUT4 n28005_bdd_3_lut (.A(n28005), .B(n28002), .C(index_i[4]), .Z(n28006)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n28005_bdd_3_lut.init = 16'hcaca;
    PFUMX i25200 (.BLUT(n27543), .ALUT(n27544), .C0(index_i[1]), .Z(n27545));
    L6MUX21 i20667 (.D0(n23030), .D1(n23031), .SD(index_i[6]), .Z(n23041));
    LUT4 mux_231_Mux_8_i892_3_lut_4_lut (.A(n27146), .B(index_i[4]), .C(index_i[5]), 
         .D(n860), .Z(n892_adj_2811)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_8_i892_3_lut_4_lut.init = 16'h4f40;
    L6MUX21 i21188 (.D0(n23350), .D1(n23357), .SD(index_i[6]), .Z(n23562));
    LUT4 n27337_bdd_4_lut (.A(n27337), .B(index_i[4]), .C(n29076), .D(index_i[5]), 
         .Z(n29908)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C (D))) */ ;
    defparam n27337_bdd_4_lut.init = 16'hf088;
    LUT4 i20876_3_lut (.A(n23247), .B(n23248), .C(index_i[8]), .Z(n23250)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20876_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_1_i700_3_lut_4_lut (.A(n27262), .B(index_i[3]), .C(index_i[4]), 
         .D(n684), .Z(n700)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_1_i700_3_lut_4_lut.init = 16'hefe0;
    L6MUX21 i21191 (.D0(n21860), .D1(n21863), .SD(index_i[6]), .Z(n23565));
    LUT4 index_i_1__bdd_4_lut_25164 (.A(index_i[1]), .B(index_i[0]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n27489)) /* synthesis lut_function=(!(A (B (D)+!B (C+!(D)))+!A !(B (C (D)+!C !(D))+!B !((D)+!C)))) */ ;
    defparam index_i_1__bdd_4_lut_25164.init = 16'h429c;
    L6MUX21 i21192 (.D0(n21929), .D1(n21935), .SD(index_i[6]), .Z(n23566));
    LUT4 i21360_3_lut (.A(n23731), .B(n23732), .C(index_i[8]), .Z(n23734)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21360_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_0_i684_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n684_adj_2812)) /* synthesis lut_function=(!(A ((D)+!B)+!A !(B (D)+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_0_i684_3_lut_4_lut_4_lut_4_lut.init = 16'h5498;
    LUT4 mux_231_Mux_6_i467_3_lut_3_lut_rep_800 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29927)) /* synthesis lut_function=(!(A (B)+!A (B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_6_i467_3_lut_3_lut_rep_800.init = 16'h3636;
    LUT4 i19996_3_lut_4_lut (.A(n27407), .B(index_i[2]), .C(index_i[3]), 
         .D(n29930), .Z(n22351)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19996_3_lut_4_lut.init = 16'hf404;
    LUT4 index_i_1__bdd_4_lut_26126 (.A(index_i[1]), .B(index_i[0]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n27490)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A !(B ((D)+!C)+!B (D))) */ ;
    defparam index_i_1__bdd_4_lut_26126.init = 16'h8a51;
    LUT4 n300_bdd_3_lut_24326 (.A(n27360), .B(n29927), .C(index_i[3]), 
         .Z(n26045)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n300_bdd_3_lut_24326.init = 16'hcaca;
    LUT4 mux_231_Mux_0_i731_3_lut_4_lut (.A(n27407), .B(index_i[2]), .C(index_i[3]), 
         .D(n27417), .Z(n731)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_0_i731_3_lut_4_lut.init = 16'h4f40;
    LUT4 n442_bdd_3_lut_24332 (.A(n27376), .B(n29957), .C(index_i[3]), 
         .Z(n26054)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n442_bdd_3_lut_24332.init = 16'hcaca;
    LUT4 mux_231_Mux_2_i955_then_4_lut (.A(index_i[4]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n27492)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B (C+!(D))+!B !(C (D)))) */ ;
    defparam mux_231_Mux_2_i955_then_4_lut.init = 16'he95d;
    LUT4 n254_bdd_4_lut_25020 (.A(index_i[5]), .B(index_i[3]), .C(index_i[6]), 
         .D(index_i[4]), .Z(n24889)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;
    defparam n254_bdd_4_lut_25020.init = 16'hf8f0;
    LUT4 i11648_3_lut (.A(index_i[2]), .B(index_i[1]), .C(index_i[0]), 
         .Z(n77)) /* synthesis lut_function=(!(A (B (C))+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11648_3_lut.init = 16'h3b3b;
    LUT4 mux_231_Mux_6_i475_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n475)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A !(B (C+(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_6_i475_3_lut_4_lut_4_lut.init = 16'h9936;
    LUT4 i20670_3_lut (.A(n25286), .B(n23037), .C(index_i[7]), .Z(n23044)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20670_3_lut.init = 16'hcaca;
    LUT4 i19906_3_lut_4_lut (.A(index_i[0]), .B(n27325), .C(index_i[3]), 
         .D(n27377), .Z(n22261)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19906_3_lut_4_lut.init = 16'hfb0b;
    LUT4 n24894_bdd_3_lut (.A(n27554), .B(n24890), .C(index_i[7]), .Z(n24895)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n24894_bdd_3_lut.init = 16'hcaca;
    L6MUX21 i21193 (.D0(n21938), .D1(n21941), .SD(index_i[6]), .Z(n23567));
    LUT4 n300_bdd_3_lut_24514 (.A(n27360), .B(n14), .C(index_i[3]), .Z(n26056)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n300_bdd_3_lut_24514.init = 16'hacac;
    PFUMX i21194 (.BLUT(n21944), .ALUT(n892_adj_2813), .C0(index_i[6]), 
          .Z(n23568));
    LUT4 i11557_2_lut_3_lut_4_lut (.A(index_i[1]), .B(n27318), .C(index_i[5]), 
         .D(index_i[4]), .Z(n508)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;
    defparam i11557_2_lut_3_lut_4_lut.init = 16'hf080;
    LUT4 mux_231_Mux_2_i189_3_lut_3_lut_4_lut (.A(index_i[1]), .B(n27318), 
         .C(n173), .D(index_i[4]), .Z(n189_adj_2814)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(C+(D)))) */ ;
    defparam mux_231_Mux_2_i189_3_lut_3_lut_4_lut.init = 16'h77f0;
    LUT4 mux_231_Mux_2_i955_else_4_lut (.A(index_i[4]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n27491)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+(D)))+!A !(B (C+!(D))+!B !(C+!(D))))) */ ;
    defparam mux_231_Mux_2_i955_else_4_lut.init = 16'h49c6;
    LUT4 i20143_3_lut (.A(n27421), .B(n29957), .C(index_i[3]), .Z(n22498)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20143_3_lut.init = 16'hcaca;
    LUT4 i22339_3_lut (.A(n22497), .B(n22498), .C(index_i[4]), .Z(n22499)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22339_3_lut.init = 16'hcaca;
    LUT4 i22202_3_lut (.A(n22494), .B(n22495), .C(index_i[4]), .Z(n22496)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22202_3_lut.init = 16'hcaca;
    LUT4 i20005_3_lut_4_lut (.A(n27413), .B(index_i[2]), .C(index_i[3]), 
         .D(n27404), .Z(n22360)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20005_3_lut_4_lut.init = 16'hdfd0;
    LUT4 i6481_2_lut (.A(phase_i[0]), .B(phase_i[10]), .Z(index_i_9__N_2125[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(60[14] 63[8])
    defparam i6481_2_lut.init = 16'h6666;
    LUT4 i7041_2_lut (.A(index_i[4]), .B(index_i[5]), .Z(n9462)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i7041_2_lut.init = 16'h8888;
    LUT4 mux_231_Mux_8_i763_3_lut_4_lut (.A(n27407), .B(n27336), .C(index_i[4]), 
         .D(n27160), .Z(n15328)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam mux_231_Mux_8_i763_3_lut_4_lut.init = 16'hfe0e;
    L6MUX21 i23932 (.D0(n25642), .D1(n25639), .SD(index_i[5]), .Z(n25643));
    LUT4 i21259_3_lut (.A(n23622), .B(n23623), .C(index_i[6]), .Z(n23633)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21259_3_lut.init = 16'hcaca;
    PFUMX i23930 (.BLUT(n25641), .ALUT(n475), .C0(index_i[4]), .Z(n25642));
    LUT4 mux_231_Mux_6_i251_3_lut_4_lut (.A(n27364), .B(index_i[2]), .C(index_i[3]), 
         .D(n27401), .Z(n251_adj_2815)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_6_i251_3_lut_4_lut.init = 16'hf606;
    LUT4 i9526_3_lut_4_lut (.A(n27364), .B(index_i[2]), .C(n27324), .D(n27401), 
         .Z(n444)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9526_3_lut_4_lut.init = 16'h6f60;
    PFUMX i23927 (.BLUT(n25638), .ALUT(n22489), .C0(index_i[4]), .Z(n25639));
    LUT4 mux_231_Mux_4_i747_3_lut_4_lut (.A(n27364), .B(index_i[2]), .C(index_i[3]), 
         .D(n29933), .Z(n747)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_4_i747_3_lut_4_lut.init = 16'hf606;
    L6MUX21 i23925 (.D0(n25636), .D1(n25634), .SD(index_i[5]), .Z(n25637));
    PFUMX i23923 (.BLUT(n25635), .ALUT(n285), .C0(index_i[4]), .Z(n25636));
    LUT4 i22441_3_lut (.A(n620_adj_2816), .B(n14250), .C(index_i[4]), 
         .Z(n21934)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22441_3_lut.init = 16'hcaca;
    PFUMX i23921 (.BLUT(n25633), .ALUT(n25632), .C0(index_i[4]), .Z(n25634));
    LUT4 mux_231_Mux_6_i518_3_lut_3_lut_rep_803 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29930)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_6_i518_3_lut_3_lut_rep_803.init = 16'h6c6c;
    LUT4 i19576_3_lut (.A(n325), .B(n27404), .C(index_i[3]), .Z(n21931)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19576_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_0_i124_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n124_adj_2817)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A !(B (D)+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_0_i124_3_lut_4_lut_4_lut.init = 16'h6c99;
    LUT4 i22223_3_lut (.A(n21930), .B(n21931), .C(index_i[4]), .Z(n21932)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22223_3_lut.init = 16'hcaca;
    LUT4 i11646_3_lut_3_lut_3_lut_rep_790 (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .Z(n29917)) /* synthesis lut_function=(!(A+!(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11646_3_lut_3_lut_3_lut_rep_790.init = 16'h4545;
    LUT4 i19570_3_lut (.A(n27402), .B(n29933), .C(index_i[3]), .Z(n21925)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19570_3_lut.init = 16'hcaca;
    LUT4 i19968_3_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[0]), 
         .D(index_i[3]), .Z(n22323)) /* synthesis lut_function=(!(A ((D)+!B)+!A !(B (D)+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19968_3_lut_4_lut_4_lut.init = 16'h4588;
    LUT4 mux_231_Mux_5_i371_3_lut_4_lut_3_lut_rep_806 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29933)) /* synthesis lut_function=(A ((C)+!B)+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_5_i371_3_lut_4_lut_3_lut_rep_806.init = 16'hb6b6;
    LUT4 n173_bdd_4_lut (.A(n173_adj_2818), .B(n27412), .C(index_i[4]), 
         .D(index_i[3]), .Z(n25168)) /* synthesis lut_function=(A (B+(C+!(D)))+!A !((C+!(D))+!B)) */ ;
    defparam n173_bdd_4_lut.init = 16'hacaa;
    LUT4 mux_231_Mux_1_i301_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n301)) /* synthesis lut_function=(A (B (C+(D))+!B !(D))+!A !(B (C+(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_1_i301_3_lut_4_lut_4_lut.init = 16'h99b6;
    LUT4 i20134_3_lut (.A(n404), .B(n27404), .C(index_i[3]), .Z(n22489)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20134_3_lut.init = 16'hcaca;
    LUT4 index_i_4__bdd_4_lut_24167 (.A(index_i[4]), .B(n27196), .C(index_i[7]), 
         .D(n27169), .Z(n25180)) /* synthesis lut_function=(A (C+!(D))+!A (B+!(C))) */ ;
    defparam index_i_4__bdd_4_lut_24167.init = 16'he5ef;
    LUT4 mux_231_Mux_0_i475_3_lut_4_lut (.A(n27266), .B(index_i[1]), .C(index_i[3]), 
         .D(n29920), .Z(n475_adj_2819)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_0_i475_3_lut_4_lut.init = 16'h4f40;
    LUT4 mux_231_Mux_3_i491_3_lut_4_lut (.A(n27266), .B(index_i[1]), .C(index_i[3]), 
         .D(n27398), .Z(n491)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_3_i491_3_lut_4_lut.init = 16'h4f40;
    LUT4 i11517_3_lut_4_lut (.A(n27065), .B(index_i[7]), .C(index_i[8]), 
         .D(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2145[14])) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11517_3_lut_4_lut.init = 16'hffe0;
    PFUMX i21030 (.BLUT(n142_adj_2820), .ALUT(n157_adj_2821), .C0(index_i[4]), 
          .Z(n23404));
    LUT4 i20131_3_lut (.A(n404), .B(n27369), .C(index_i[3]), .Z(n22486)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20131_3_lut.init = 16'hcaca;
    LUT4 i19573_3_lut_4_lut_4_lut_4_lut (.A(n27413), .B(index_i[2]), .C(index_i[3]), 
         .D(index_i[4]), .Z(n21928)) /* synthesis lut_function=(A (B)+!A (B (C (D))+!B !(C (D)))) */ ;
    defparam i19573_3_lut_4_lut_4_lut_4_lut.init = 16'hc999;
    LUT4 i20140_3_lut_4_lut (.A(n27413), .B(index_i[2]), .C(index_i[3]), 
         .D(n27337), .Z(n22495)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;
    defparam i20140_3_lut_4_lut.init = 16'h6f60;
    LUT4 i20130_3_lut (.A(n27406), .B(n325), .C(index_i[3]), .Z(n22485)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20130_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_2_i684_3_lut_4_lut (.A(n27413), .B(index_i[2]), .C(index_i[3]), 
         .D(n29917), .Z(n684_adj_2822)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;
    defparam mux_231_Mux_2_i684_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_231_Mux_7_i653_3_lut_4_lut (.A(n27413), .B(index_i[2]), .C(index_i[3]), 
         .D(n27412), .Z(n653)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam mux_231_Mux_7_i653_3_lut_4_lut.init = 16'hf606;
    LUT4 i22228_3_lut (.A(n21921), .B(n21922), .C(index_i[4]), .Z(n21923)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22228_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_7_i475_3_lut_3_lut_4_lut (.A(n27413), .B(index_i[2]), 
         .C(n27408), .D(index_i[3]), .Z(n475_adj_2823)) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))+!A !(B ((D)+!C)+!B !(C+(D)))) */ ;
    defparam mux_231_Mux_7_i475_3_lut_3_lut_4_lut.init = 16'h99f0;
    LUT4 i19578_4_lut_4_lut_4_lut (.A(n27413), .B(index_i[2]), .C(index_i[4]), 
         .D(index_i[3]), .Z(n21933)) /* synthesis lut_function=(A (B)+!A !(B (C+(D))+!B !(C+(D)))) */ ;
    defparam i19578_4_lut_4_lut_4_lut.init = 16'h999c;
    PFUMX i21031 (.BLUT(n173_adj_2824), .ALUT(n188), .C0(index_i[4]), 
          .Z(n23405));
    L6MUX21 i21254 (.D0(n23612), .D1(n23613), .SD(index_i[6]), .Z(n23628));
    L6MUX21 i21255 (.D0(n23614), .D1(n23615), .SD(index_i[6]), .Z(n23629));
    L6MUX21 i21256 (.D0(n23616), .D1(n23617), .SD(index_i[6]), .Z(n23630));
    L6MUX21 i21257 (.D0(n23618), .D1(n23619), .SD(index_i[6]), .Z(n23631));
    L6MUX21 i21258 (.D0(n23620), .D1(n23621), .SD(index_i[6]), .Z(n23632));
    L6MUX21 i21260 (.D0(n23624), .D1(n23625), .SD(index_i[6]), .Z(n23634));
    LUT4 i1_3_lut (.A(index_i[0]), .B(index_i[4]), .C(index_i[2]), .Z(n21022)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_3_lut.init = 16'hfefe;
    L6MUX21 i21285 (.D0(n23643), .D1(n23644), .SD(index_i[6]), .Z(n23659));
    LUT4 mux_231_Mux_13_i511_4_lut_4_lut (.A(n27065), .B(index_i[7]), .C(index_i[8]), 
         .D(n254), .Z(n511)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (B (C+!(D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_13_i511_4_lut_4_lut.init = 16'h1c10;
    PFUMX i20858 (.BLUT(n732), .ALUT(n763), .C0(index_i[5]), .Z(n23232));
    LUT4 i20125_3_lut (.A(n27406), .B(n27369), .C(index_i[3]), .Z(n22480)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20125_3_lut.init = 16'hcaca;
    L6MUX21 i20860 (.D0(n22361), .D1(n891_adj_2825), .SD(index_i[5]), 
            .Z(n23234));
    LUT4 i12449_3_lut (.A(index_i[2]), .B(index_i[1]), .C(index_i[0]), 
         .Z(n38)) /* synthesis lut_function=(A (B)+!A (B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12449_3_lut.init = 16'hdcdc;
    L6MUX21 i21286 (.D0(n23645), .D1(n23646), .SD(index_i[6]), .Z(n23660));
    L6MUX21 i21287 (.D0(n23647), .D1(n23648), .SD(index_i[6]), .Z(n23661));
    L6MUX21 i20863 (.D0(n23221), .D1(n23222), .SD(index_i[6]), .Z(n23237));
    L6MUX21 i20865 (.D0(n23225), .D1(n23226), .SD(index_i[6]), .Z(n23239));
    PFUMX i21289 (.BLUT(n23651), .ALUT(n23652), .C0(index_i[6]), .Z(n23663));
    L6MUX21 i20866 (.D0(n23227), .D1(n23228), .SD(index_i[6]), .Z(n23240));
    L6MUX21 i21290 (.D0(n23653), .D1(n23654), .SD(index_i[6]), .Z(n23664));
    L6MUX21 i21291 (.D0(n23655), .D1(n23656), .SD(index_i[6]), .Z(n23665));
    PFUMX i21292 (.BLUT(n23657), .ALUT(n23658), .C0(index_i[6]), .Z(n23666));
    L6MUX21 i20870 (.D0(n23235), .D1(n23236), .SD(index_i[6]), .Z(n23244));
    LUT4 i20124_3_lut (.A(n325), .B(n27331), .C(index_i[3]), .Z(n22479)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20124_3_lut.init = 16'hcaca;
    PFUMX i21036 (.BLUT(n333_adj_2826), .ALUT(n348_adj_2827), .C0(index_i[4]), 
          .Z(n23410));
    PFUMX i21037 (.BLUT(n364), .ALUT(n379), .C0(index_i[4]), .Z(n23411));
    PFUMX i21038 (.BLUT(n397_adj_2828), .ALUT(n412_adj_2805), .C0(index_i[4]), 
          .Z(n23412));
    L6MUX21 i20906 (.D0(n23278), .D1(n23279), .SD(index_i[6]), .Z(n23280));
    LUT4 i1_2_lut (.A(index_i[6]), .B(index_i[7]), .Z(n20104)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_2_lut.init = 16'heeee;
    L6MUX21 i20913 (.D0(n23285), .D1(n23286), .SD(index_i[6]), .Z(n23287));
    PFUMX i21039 (.BLUT(n428), .ALUT(n443), .C0(index_i[4]), .Z(n23413));
    PFUMX i21040 (.BLUT(n460), .ALUT(n475_adj_2819), .C0(index_i[4]), 
          .Z(n23414));
    PFUMX i21041 (.BLUT(n491_adj_2829), .ALUT(n11349), .C0(index_i[4]), 
          .Z(n23415));
    PFUMX i21343 (.BLUT(n797), .ALUT(n828), .C0(index_i[5]), .Z(n23717));
    LUT4 n308_bdd_3_lut_24465 (.A(n27400), .B(n29927), .C(index_i[3]), 
         .Z(n26189)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n308_bdd_3_lut_24465.init = 16'hacac;
    L6MUX21 i21347 (.D0(n23705), .D1(n23706), .SD(index_i[6]), .Z(n23721));
    L6MUX21 i21348 (.D0(n23707), .D1(n23708), .SD(index_i[6]), .Z(n23722));
    L6MUX21 i21349 (.D0(n23709), .D1(n23710), .SD(index_i[6]), .Z(n23723));
    L6MUX21 i21350 (.D0(n23711), .D1(n23712), .SD(index_i[6]), .Z(n23724));
    L6MUX21 i21351 (.D0(n23713), .D1(n23714), .SD(index_i[6]), .Z(n23725));
    L6MUX21 i21354 (.D0(n23719), .D1(n23720), .SD(index_i[6]), .Z(n23728));
    L6MUX21 i21397 (.D0(n23759), .D1(n23760), .SD(index_i[6]), .Z(n23771));
    LUT4 i15954_4_lut (.A(index_i[0]), .B(index_i[4]), .C(index_i[1]), 
         .D(n27336), .Z(n286)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i15954_4_lut.init = 16'hccc8;
    L6MUX21 i21398 (.D0(n23761), .D1(n23762), .SD(index_i[6]), .Z(n23772));
    L6MUX21 i21399 (.D0(n23763), .D1(n23764), .SD(index_i[6]), .Z(n23773));
    LUT4 mux_231_Mux_3_i652_rep_812 (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .Z(n29939)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_3_i652_rep_812.init = 16'h4d4d;
    LUT4 mux_231_Mux_3_i653_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n653_adj_2830)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A !(B (D)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_3_i653_3_lut_4_lut_4_lut.init = 16'h4d99;
    PFUMX i21400 (.BLUT(n23765), .ALUT(n23766), .C0(index_i[6]), .Z(n23774));
    LUT4 n715_bdd_3_lut_24516 (.A(n27416), .B(n27403), .C(index_i[3]), 
         .Z(n26205)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n715_bdd_3_lut_24516.init = 16'hcaca;
    L6MUX21 i20416 (.D0(n21827), .D1(n21830), .SD(index_i[6]), .Z(n22790));
    PFUMX i20417 (.BLUT(n11982), .ALUT(n21833), .C0(index_i[6]), .Z(n22791));
    LUT4 i21189_3_lut (.A(n190), .B(n26581), .C(index_i[6]), .Z(n23563)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21189_3_lut.init = 16'hcaca;
    LUT4 i21190_3_lut (.A(n23364), .B(n21857), .C(index_i[6]), .Z(n23564)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21190_3_lut.init = 16'hcaca;
    L6MUX21 i20419 (.D0(n21839), .D1(n21842), .SD(index_i[6]), .Z(n22793));
    PFUMX i21058 (.BLUT(n557), .ALUT(n572), .C0(index_i[4]), .Z(n23432));
    L6MUX21 i20420 (.D0(n574_adj_2831), .D1(n21845), .SD(index_i[6]), 
            .Z(n22794));
    L6MUX21 i20421 (.D0(n21848), .D1(n764), .SD(index_i[6]), .Z(n22795));
    PFUMX i21059 (.BLUT(n589), .ALUT(n604), .C0(index_i[4]), .Z(n23433));
    PFUMX i25194 (.BLUT(n27534), .ALUT(n27535), .C0(index_i[0]), .Z(n27536));
    PFUMX i19901 (.BLUT(n22254), .ALUT(n22255), .C0(index_i[4]), .Z(n22256));
    PFUMX i19904 (.BLUT(n22257), .ALUT(n22258), .C0(index_i[4]), .Z(n22259));
    LUT4 mux_231_Mux_6_i435_3_lut_4_lut_3_lut_rep_815 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29942)) /* synthesis lut_function=(A (B+!(C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_6_i435_3_lut_4_lut_3_lut_rep_815.init = 16'hdbdb;
    PFUMX i20435 (.BLUT(n22805), .ALUT(n22806), .C0(index_i[6]), .Z(n22809));
    PFUMX i20436 (.BLUT(n22807), .ALUT(n22808), .C0(index_i[6]), .Z(n22810));
    LUT4 i9669_3_lut_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n12158)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A !(B (C+(D))+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9669_3_lut_3_lut_4_lut_4_lut.init = 16'h44db;
    PFUMX i20443 (.BLUT(n22814), .ALUT(n22815), .C0(index_i[6]), .Z(n22817));
    LUT4 mux_231_Mux_5_i505_3_lut_3_lut_rep_816 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29943)) /* synthesis lut_function=(A (B+(C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_5_i505_3_lut_3_lut_rep_816.init = 16'hadad;
    LUT4 mux_231_Mux_0_i796_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n796)) /* synthesis lut_function=(A (B (C+(D))+!B (C (D)))+!A !(B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_0_i796_3_lut_4_lut_4_lut.init = 16'hadc0;
    LUT4 i11606_2_lut_rep_793 (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .Z(n29920)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11606_2_lut_rep_793.init = 16'hf8f8;
    PFUMX i21060 (.BLUT(n620_adj_2832), .ALUT(n635_adj_2833), .C0(index_i[4]), 
          .Z(n23434));
    LUT4 i9628_3_lut (.A(n12113), .B(n27397), .C(index_i[3]), .Z(n12114)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9628_3_lut.init = 16'hcaca;
    LUT4 i20418_3_lut (.A(n26436), .B(n23343), .C(index_i[6]), .Z(n22792)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20418_3_lut.init = 16'hcaca;
    PFUMX i21061 (.BLUT(n653_adj_2834), .ALUT(n668), .C0(index_i[4]), 
          .Z(n23435));
    PFUMX i21062 (.BLUT(n684_adj_2812), .ALUT(n699_adj_2835), .C0(index_i[4]), 
          .Z(n23436));
    PFUMX i21063 (.BLUT(n716_adj_2836), .ALUT(n731), .C0(index_i[4]), 
          .Z(n23437));
    LUT4 i11597_3_lut_4_lut (.A(n27318), .B(index_i[4]), .C(index_i[5]), 
         .D(n27413), .Z(n892)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11597_3_lut_4_lut.init = 16'hf8f0;
    LUT4 mux_231_Mux_3_i1018_3_lut_4_lut (.A(index_i[1]), .B(n27336), .C(index_i[4]), 
         .D(n20184), .Z(n1018)) /* synthesis lut_function=(A (C+!(D))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_3_i1018_3_lut_4_lut.init = 16'he0ef;
    LUT4 mux_231_Mux_2_i700_3_lut_4_lut (.A(index_i[1]), .B(n27336), .C(index_i[4]), 
         .D(n684_adj_2822), .Z(n700_adj_2837)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_2_i700_3_lut_4_lut.init = 16'hefe0;
    PFUMX i21064 (.BLUT(n747_adj_2838), .ALUT(n762_adj_2839), .C0(index_i[4]), 
          .Z(n23438));
    LUT4 n251_bdd_4_lut_26381 (.A(n251_adj_2815), .B(n11192), .C(index_i[2]), 
         .D(index_i[4]), .Z(n26281)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C+(D)))+!A !(B (C+(D))+!B ((D)+!C))) */ ;
    defparam n251_bdd_4_lut_26381.init = 16'haa3c;
    L6MUX21 i21050 (.D0(n23416), .D1(n23417), .SD(index_i[6]), .Z(n23424));
    L6MUX21 i21053 (.D0(n23422), .D1(n23423), .SD(index_i[6]), .Z(n23427));
    LUT4 mux_231_Mux_8_i732_3_lut (.A(index_i[3]), .B(n15328), .C(index_i[5]), 
         .Z(n732_adj_2840)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_8_i732_3_lut.init = 16'h3a3a;
    LUT4 n25280_bdd_3_lut (.A(n25280), .B(n476), .C(index_i[5]), .Z(n25281)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n25280_bdd_3_lut.init = 16'hcaca;
    LUT4 i22044_3_lut (.A(n22455), .B(n22456), .C(index_i[4]), .Z(n22457)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i22044_3_lut.init = 16'hcaca;
    PFUMX i19925 (.BLUT(n22278), .ALUT(n22279), .C0(index_i[4]), .Z(n22280));
    LUT4 n28834_bdd_3_lut (.A(n28834), .B(index_i[1]), .C(index_i[4]), 
         .Z(n28835)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n28834_bdd_3_lut.init = 16'hcaca;
    LUT4 index_i_1__bdd_4_lut_26738 (.A(index_i[1]), .B(index_i[3]), .C(index_i[0]), 
         .D(index_i[2]), .Z(n28834)) /* synthesis lut_function=(A (B (C+(D))+!B (C (D)))+!A !(B (C)+!B !(C+(D)))) */ ;
    defparam index_i_1__bdd_4_lut_26738.init = 16'hbd94;
    L6MUX21 i21081 (.D0(n23447), .D1(n23448), .SD(index_i[6]), .Z(n23455));
    PFUMX mux_231_Mux_2_i891 (.BLUT(n875), .ALUT(n890), .C0(index_i[4]), 
          .Z(n891_adj_2841)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    L6MUX21 i21082 (.D0(n23449), .D1(n23450), .SD(index_i[6]), .Z(n23456));
    PFUMX i21065 (.BLUT(n781), .ALUT(n796), .C0(index_i[4]), .Z(n23439));
    LUT4 i21051_3_lut (.A(n23418), .B(n29079), .C(index_i[6]), .Z(n23425)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21051_3_lut.init = 16'hcaca;
    L6MUX21 i21083 (.D0(n23451), .D1(n23452), .SD(index_i[6]), .Z(n23457));
    LUT4 i21052_3_lut (.A(n26501), .B(n23421), .C(index_i[6]), .Z(n23426)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21052_3_lut.init = 16'hcaca;
    LUT4 n25284_bdd_3_lut_25033 (.A(n27545), .B(n25282), .C(index_i[5]), 
         .Z(n25285)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n25284_bdd_3_lut_25033.init = 16'hcaca;
    PFUMX mux_231_Mux_2_i860 (.BLUT(n844_adj_2797), .ALUT(n859), .C0(index_i[4]), 
          .Z(n860_adj_2842)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 i19506_3_lut (.A(n397), .B(n475_adj_2823), .C(index_i[4]), .Z(n21861)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19506_3_lut.init = 16'hcaca;
    L6MUX21 i21084 (.D0(n23453), .D1(n23454), .SD(index_i[6]), .Z(n23458));
    LUT4 i19504_3_lut (.A(n348_adj_2796), .B(n443_adj_2843), .C(index_i[4]), 
         .Z(n21859)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19504_3_lut.init = 16'hcaca;
    LUT4 i19503_3_lut (.A(n397), .B(n412_adj_2844), .C(index_i[4]), .Z(n21858)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19503_3_lut.init = 16'hcaca;
    LUT4 i19501_3_lut (.A(n364_adj_2845), .B(n379_adj_2846), .C(index_i[4]), 
         .Z(n21856)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19501_3_lut.init = 16'hcaca;
    LUT4 i19500_3_lut (.A(n333), .B(n348_adj_2796), .C(index_i[4]), .Z(n21855)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19500_3_lut.init = 16'hcaca;
    PFUMX i21066 (.BLUT(n812_adj_2847), .ALUT(n12119), .C0(index_i[4]), 
          .Z(n23440));
    PFUMX i19419 (.BLUT(n318), .ALUT(n381), .C0(index_i[6]), .Z(n21774));
    PFUMX i21057 (.BLUT(n526_adj_2848), .ALUT(n541), .C0(index_i[4]), 
          .Z(n23431));
    LUT4 mux_231_Mux_8_i124_3_lut_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n124_adj_2849)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C+!(D)))+!A (B (C (D)+!C !(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_8_i124_3_lut_3_lut_4_lut_4_lut.init = 16'h07c1;
    PFUMX i21068 (.BLUT(n875_adj_2850), .ALUT(n890_adj_2806), .C0(index_i[4]), 
          .Z(n23442));
    LUT4 n27226_bdd_3_lut_26276_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[5]), .Z(n29074)) /* synthesis lut_function=(A (B+(C+(D)))+!A !((D)+!C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n27226_bdd_3_lut_26276_4_lut.init = 16'haaf8;
    PFUMX i25192 (.BLUT(n27531), .ALUT(n27532), .C0(index_i[0]), .Z(n27533));
    PFUMX i21069 (.BLUT(n908_adj_2793), .ALUT(n923), .C0(index_i[4]), 
          .Z(n23443));
    L6MUX21 i23867 (.D0(n25579), .D1(n27054), .SD(index_i[6]), .Z(n23294));
    PFUMX i23865 (.BLUT(n25578), .ALUT(n25577), .C0(index_i[5]), .Z(n25579));
    PFUMX i21070 (.BLUT(n939), .ALUT(n954), .C0(index_i[4]), .Z(n23444));
    LUT4 n27226_bdd_4_lut_26275 (.A(index_i[5]), .B(index_i[2]), .C(index_i[0]), 
         .D(index_i[1]), .Z(n29073)) /* synthesis lut_function=(!(A (B (D)+!B ((D)+!C))+!A !(B (C (D)+!C !(D))+!B !(D)))) */ ;
    defparam n27226_bdd_4_lut_26275.init = 16'h40bd;
    LUT4 n557_bdd_4_lut (.A(n27128), .B(index_i[4]), .C(n25574), .D(index_i[5]), 
         .Z(n27054)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (B (C (D))+!B (C+!(D)))) */ ;
    defparam n557_bdd_4_lut.init = 16'hf099;
    PFUMX i19934 (.BLUT(n22287), .ALUT(n22288), .C0(index_i[4]), .Z(n22289));
    LUT4 mux_231_Mux_6_i844_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n844_adj_2800)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (B (C)+!B !(C+!(D)))) */ ;
    defparam mux_231_Mux_6_i844_3_lut_4_lut_4_lut.init = 16'hc1e0;
    LUT4 n27337_bdd_3_lut_26279 (.A(index_i[2]), .B(index_i[0]), .C(index_i[4]), 
         .Z(n29076)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B (C)+!B !(C)))) */ ;
    defparam n27337_bdd_3_lut_26279.init = 16'h6969;
    LUT4 mux_231_Mux_6_i732_3_lut_4_lut (.A(n27416), .B(index_i[3]), .C(index_i[4]), 
         .D(n412_adj_2844), .Z(n732_adj_2851)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_6_i732_3_lut_4_lut.init = 16'hf909;
    PFUMX i25142 (.BLUT(n27452), .ALUT(n27453), .C0(index_i[1]), .Z(n27454));
    PFUMX i19943 (.BLUT(n22296), .ALUT(n22297), .C0(index_i[4]), .Z(n22298));
    LUT4 mux_231_Mux_6_i700_3_lut_4_lut (.A(n27416), .B(index_i[3]), .C(index_i[4]), 
         .D(n684_adj_2852), .Z(n700_adj_2853)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_6_i700_3_lut_4_lut.init = 16'h9f90;
    PFUMX mux_231_Mux_3_i763 (.BLUT(n747_adj_2854), .ALUT(n762), .C0(index_i[4]), 
          .Z(n763_adj_2855)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 i21026_3_lut (.A(n541_adj_2856), .B(n27490), .C(index_i[4]), 
         .Z(n23400)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21026_3_lut.init = 16'hcaca;
    L6MUX21 i23372 (.D0(n24972), .D1(n24969), .SD(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2145[9]));
    PFUMX i20648 (.BLUT(n158_adj_2857), .ALUT(n189_adj_2814), .C0(index_i[5]), 
          .Z(n23022));
    PFUMX i19952 (.BLUT(n22305), .ALUT(n22306), .C0(index_i[4]), .Z(n22307));
    PFUMX i20649 (.BLUT(n221_adj_2858), .ALUT(n21980), .C0(index_i[5]), 
          .Z(n23023));
    PFUMX i21071 (.BLUT(n971), .ALUT(n986), .C0(index_i[4]), .Z(n23445));
    PFUMX i21072 (.BLUT(n1002), .ALUT(n1017), .C0(index_i[4]), .Z(n23446));
    LUT4 i20440_4_lut_4_lut (.A(n27130), .B(n27205), .C(index_i[5]), .D(index_i[4]), 
         .Z(n22814)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C+(D))+!B !(C (D)+!C !(D)))) */ ;
    defparam i20440_4_lut_4_lut.init = 16'hcf50;
    PFUMX i20650 (.BLUT(n286_adj_2859), .ALUT(n317_adj_2860), .C0(index_i[5]), 
          .Z(n23024));
    PFUMX i20651 (.BLUT(n349_adj_2861), .ALUT(n21983), .C0(index_i[5]), 
          .Z(n23025));
    PFUMX i20652 (.BLUT(n413_adj_2862), .ALUT(n21986), .C0(index_i[5]), 
          .Z(n23026));
    PFUMX i20653 (.BLUT(n21989), .ALUT(n507), .C0(index_i[5]), .Z(n23027));
    PFUMX i19496 (.BLUT(n21849), .ALUT(n21850), .C0(index_i[4]), .Z(n21851));
    PFUMX i20654 (.BLUT(n21992), .ALUT(n573), .C0(index_i[5]), .Z(n23028));
    LUT4 i19522_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21877)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A (B (C (D)+!C !(D))+!B (D))) */ ;
    defparam i19522_3_lut_4_lut.init = 16'hd926;
    LUT4 n23662_bdd_3_lut_23342 (.A(n23662), .B(n23661), .C(index_i[7]), 
         .Z(n24941)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n23662_bdd_3_lut_23342.init = 16'hacac;
    LUT4 mux_231_Mux_5_i124_3_lut (.A(n204), .B(n27421), .C(index_i[3]), 
         .Z(n124)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_5_i124_3_lut.init = 16'hcaca;
    PFUMX i19574 (.BLUT(n21927), .ALUT(n21928), .C0(index_i[5]), .Z(n21929));
    LUT4 i19486_3_lut (.A(n491_adj_2863), .B(n541_adj_2864), .C(index_i[4]), 
         .Z(n21841)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19486_3_lut.init = 16'hcaca;
    LUT4 i19485_3_lut (.A(n397_adj_2865), .B(n475_adj_2866), .C(index_i[4]), 
         .Z(n21840)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19485_3_lut.init = 16'hcaca;
    PFUMX i20655 (.BLUT(n605_adj_2867), .ALUT(n21995), .C0(index_i[5]), 
          .Z(n23029));
    PFUMX i20656 (.BLUT(n669), .ALUT(n700_adj_2837), .C0(index_i[5]), 
          .Z(n23030));
    LUT4 i19483_3_lut (.A(n251), .B(n443_adj_2804), .C(index_i[4]), .Z(n21838)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19483_3_lut.init = 16'hcaca;
    PFUMX i20657 (.BLUT(n732_adj_2868), .ALUT(n763_adj_2869), .C0(index_i[5]), 
          .Z(n23031));
    LUT4 i19482_3_lut (.A(n397_adj_2865), .B(n15042), .C(index_i[4]), 
         .Z(n21837)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;
    defparam i19482_3_lut.init = 16'h3a3a;
    LUT4 i22578_3_lut (.A(n27533), .B(n27536), .C(index_i[5]), .Z(n21833)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22578_3_lut.init = 16'hcaca;
    L6MUX21 i20659 (.D0(n860_adj_2842), .D1(n891_adj_2841), .SD(index_i[5]), 
            .Z(n23033));
    PFUMX i15946 (.BLUT(n18130), .ALUT(n18131), .C0(index_i[4]), .Z(n18132));
    LUT4 i19473_3_lut (.A(n78), .B(n93_adj_2870), .C(index_i[4]), .Z(n21828)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19473_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_6_i285_3_lut_4_lut (.A(n27359), .B(index_i[2]), .C(index_i[3]), 
         .D(n27400), .Z(n285)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_6_i285_3_lut_4_lut.init = 16'hf606;
    LUT4 n23670_bdd_3_lut (.A(n23663), .B(n23664), .C(index_i[7]), .Z(n24939)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n23670_bdd_3_lut.init = 16'hcaca;
    PFUMX i19970 (.BLUT(n22323), .ALUT(n22324), .C0(index_i[4]), .Z(n22325));
    LUT4 i19516_3_lut_4_lut (.A(n27359), .B(index_i[2]), .C(index_i[3]), 
         .D(n29933), .Z(n21871)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19516_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_231_Mux_3_i460_3_lut_4_lut (.A(n27359), .B(index_i[2]), .C(index_i[3]), 
         .D(n27379), .Z(n460_adj_2871)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_3_i460_3_lut_4_lut.init = 16'h6f60;
    LUT4 i19470_3_lut (.A(n15), .B(n30), .C(index_i[4]), .Z(n21825)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19470_3_lut.init = 16'hcaca;
    LUT4 i19897_3_lut_4_lut (.A(n27359), .B(index_i[2]), .C(index_i[3]), 
         .D(n27396), .Z(n22252)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19897_3_lut_4_lut.init = 16'hf606;
    LUT4 n23662_bdd_3_lut_24594 (.A(n23659), .B(n23660), .C(index_i[7]), 
         .Z(n24942)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n23662_bdd_3_lut_24594.init = 16'hcaca;
    PFUMX i19580 (.BLUT(n21933), .ALUT(n21934), .C0(index_i[5]), .Z(n21935));
    PFUMX mux_231_Mux_5_i732 (.BLUT(n12018), .ALUT(n731_adj_2872), .C0(index_i[4]), 
          .Z(n732_adj_2873)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 n123_bdd_3_lut_24699 (.A(n27422), .B(n29957), .C(index_i[3]), 
         .Z(n26498)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n123_bdd_3_lut_24699.init = 16'hcaca;
    PFUMX i19583 (.BLUT(n21936), .ALUT(n21937), .C0(index_i[5]), .Z(n21938));
    LUT4 i21359_3_lut (.A(n23729), .B(n23730), .C(index_i[8]), .Z(n23733)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21359_3_lut.init = 16'hcaca;
    PFUMX i23370 (.BLUT(n24971), .ALUT(n24970), .C0(index_i[8]), .Z(n24972));
    LUT4 mux_231_Mux_4_i62_4_lut (.A(n27373), .B(n61), .C(index_i[4]), 
         .D(index_i[3]), .Z(n62_adj_2874)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_4_i62_4_lut.init = 16'hc5ca;
    LUT4 mux_231_Mux_4_i31_4_lut (.A(n15_adj_2875), .B(n27143), .C(index_i[4]), 
         .D(index_i[3]), .Z(n31)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_4_i31_4_lut.init = 16'h3aca;
    PFUMX i19988 (.BLUT(n22341), .ALUT(n22342), .C0(index_i[4]), .Z(n22343));
    PFUMX i19997 (.BLUT(n22350), .ALUT(n22351), .C0(index_i[4]), .Z(n22352));
    LUT4 mux_231_Mux_3_i31_3_lut (.A(n781_adj_2876), .B(n30_adj_2877), .C(index_i[4]), 
         .Z(n31_adj_2878)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_3_i31_3_lut.init = 16'hcaca;
    PFUMX i19586 (.BLUT(n21939), .ALUT(n21940), .C0(index_i[5]), .Z(n21941));
    PFUMX i19511 (.BLUT(n21864), .ALUT(n21865), .C0(index_i[4]), .Z(n21866));
    LUT4 n269_bdd_3_lut_24318_4_lut (.A(n27362), .B(index_i[2]), .C(index_i[3]), 
         .D(n27360), .Z(n25633)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n269_bdd_3_lut_24318_4_lut.init = 16'hf606;
    LUT4 mux_231_Mux_3_i890_3_lut_4_lut (.A(n27362), .B(index_i[2]), .C(index_i[3]), 
         .D(n325), .Z(n890_adj_2879)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_3_i890_3_lut_4_lut.init = 16'h6f60;
    LUT4 i20110_3_lut_4_lut (.A(n27362), .B(index_i[2]), .C(index_i[3]), 
         .D(n27400), .Z(n22465)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20110_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_231_Mux_0_i348_3_lut_4_lut (.A(n27362), .B(index_i[2]), .C(index_i[3]), 
         .D(n29917), .Z(n348_adj_2827)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_0_i348_3_lut_4_lut.init = 16'h6f60;
    LUT4 n53_bdd_3_lut_23966_4_lut (.A(n27367), .B(index_i[2]), .C(n27377), 
         .D(index_i[3]), .Z(n25678)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n53_bdd_3_lut_23966_4_lut.init = 16'hf066;
    PFUMX i21195 (.BLUT(n956), .ALUT(n20737), .C0(index_i[6]), .Z(n23569));
    LUT4 mux_231_Mux_3_i668_3_lut_4_lut (.A(n27367), .B(index_i[2]), .C(index_i[3]), 
         .D(n27406), .Z(n668_adj_2880)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_3_i668_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_231_Mux_4_i763_3_lut_4_lut (.A(n27367), .B(index_i[2]), .C(index_i[4]), 
         .D(n747), .Z(n763_adj_2881)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_4_i763_3_lut_4_lut.init = 16'h6f60;
    LUT4 i20875_3_lut (.A(n23245), .B(n23246), .C(index_i[8]), .Z(n23249)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20875_3_lut.init = 16'hcaca;
    PFUMX i19514 (.BLUT(n21867), .ALUT(n21868), .C0(index_i[4]), .Z(n21869));
    LUT4 i9500_3_lut_4_lut_4_lut (.A(n27325), .B(index_i[3]), .C(index_i[5]), 
         .D(n27221), .Z(n11986)) /* synthesis lut_function=(A (B+(C (D)))+!A (B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9500_3_lut_4_lut_4_lut.init = 16'hf8c8;
    PFUMX i20006 (.BLUT(n22359), .ALUT(n22360), .C0(index_i[4]), .Z(n22361));
    LUT4 n62_bdd_3_lut_4_lut (.A(n27325), .B(index_i[3]), .C(index_i[4]), 
         .D(n30_adj_2882), .Z(n25660)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n62_bdd_3_lut_4_lut.init = 16'hf808;
    LUT4 i20902_3_lut_3_lut_4_lut_4_lut (.A(n27325), .B(index_i[3]), .C(index_i[4]), 
         .D(n27225), .Z(n23276)) /* synthesis lut_function=(!(A (B (C)+!B ((D)+!C))+!A (B+((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20902_3_lut_3_lut_4_lut_4_lut.init = 16'h0838;
    LUT4 n557_bdd_3_lut_24043_4_lut_4_lut (.A(n27325), .B(index_i[3]), .C(index_i[4]), 
         .D(n29920), .Z(n25578)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C))+!A !(B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n557_bdd_3_lut_24043_4_lut_4_lut.init = 16'h838f;
    PFUMX i25184 (.BLUT(n27519), .ALUT(n27520), .C0(index_i[2]), .Z(n27521));
    LUT4 mux_231_Mux_4_i573_3_lut_3_lut_4_lut_4_lut (.A(n27372), .B(index_i[3]), 
         .C(index_i[4]), .D(n27225), .Z(n573_adj_2883)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_4_i573_3_lut_3_lut_4_lut_4_lut.init = 16'h1f1c;
    LUT4 n22459_bdd_3_lut (.A(n27399), .B(n27419), .C(index_i[3]), .Z(n26577)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n22459_bdd_3_lut.init = 16'hcaca;
    LUT4 n124_bdd_3_lut_23947_4_lut (.A(n27372), .B(index_i[3]), .C(index_i[4]), 
         .D(n124_adj_2884), .Z(n25657)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n124_bdd_3_lut_23947_4_lut.init = 16'hf101;
    LUT4 i20900_3_lut_4_lut (.A(n27372), .B(index_i[3]), .C(index_i[4]), 
         .D(n285_adj_2885), .Z(n23274)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20900_3_lut_4_lut.init = 16'hfe0e;
    LUT4 n428_bdd_3_lut_24095_4_lut_4_lut (.A(n27372), .B(index_i[3]), .C(index_i[4]), 
         .D(n29920), .Z(n25799)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B (C (D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n428_bdd_3_lut_24095_4_lut_4_lut.init = 16'h3efe;
    LUT4 mux_231_Mux_3_i573_3_lut_3_lut_4_lut (.A(n27372), .B(index_i[3]), 
         .C(n397_adj_2865), .D(index_i[4]), .Z(n573_adj_2886)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_3_i573_3_lut_3_lut_4_lut.init = 16'h11f0;
    LUT4 mux_231_Mux_2_i573_3_lut_3_lut_4_lut (.A(n27372), .B(index_i[3]), 
         .C(n557_adj_2887), .D(index_i[4]), .Z(n573)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_2_i573_3_lut_3_lut_4_lut.init = 16'h11f0;
    LUT4 mux_231_Mux_6_i891_3_lut (.A(n78), .B(n890_adj_2888), .C(index_i[4]), 
         .Z(n891_adj_2889)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_6_i891_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_6_i828_4_lut (.A(n812_adj_2890), .B(n14276), .C(index_i[4]), 
         .D(index_i[2]), .Z(n828_adj_2891)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_6_i828_4_lut.init = 16'hfaca;
    LUT4 i19541_then_4_lut (.A(index_i[2]), .B(index_i[1]), .C(index_i[4]), 
         .D(index_i[3]), .Z(n27511)) /* synthesis lut_function=(A (B (C+(D))+!B !(C))+!A !(B (C+(D))+!B !(C+!(D)))) */ ;
    defparam i19541_then_4_lut.init = 16'h9a97;
    LUT4 mux_231_Mux_6_i797_3_lut (.A(n781_adj_2876), .B(n27076), .C(index_i[4]), 
         .Z(n797_adj_2892)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_6_i797_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_6_i669_3_lut (.A(n653_adj_2893), .B(n668_adj_2894), 
         .C(index_i[4]), .Z(n669_adj_2895)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_6_i669_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_6_i542_3_lut (.A(n526), .B(n541_adj_2896), .C(index_i[4]), 
         .Z(n542_adj_2897)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_6_i542_3_lut.init = 16'hcaca;
    LUT4 i20423_3_lut_4_lut (.A(n27112), .B(n27119), .C(index_i[5]), .D(index_i[6]), 
         .Z(n22797)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (B+((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20423_3_lut_4_lut.init = 16'hffc5;
    LUT4 i20432_3_lut_4_lut_4_lut (.A(n27160), .B(index_i[4]), .C(index_i[5]), 
         .D(n27130), .Z(n22806)) /* synthesis lut_function=(A ((C+!(D))+!B)+!A (B (C+!(D))+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20432_3_lut_4_lut_4_lut.init = 16'he3ef;
    LUT4 i19541_else_4_lut (.A(index_i[2]), .B(index_i[1]), .C(index_i[4]), 
         .D(index_i[3]), .Z(n27510)) /* synthesis lut_function=(!(A (B (C)+!B (C+(D)))+!A !(B (C (D)+!C !(D))+!B (C+!(D))))) */ ;
    defparam i19541_else_4_lut.init = 16'h581f;
    LUT4 i22219_3_lut (.A(n21972), .B(n27564), .C(index_i[4]), .Z(n21974)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22219_3_lut.init = 16'hcaca;
    LUT4 i12451_3_lut_rep_830 (.A(index_i[2]), .B(index_i[1]), .C(index_i[0]), 
         .Z(n29957)) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12451_3_lut_rep_830.init = 16'hc4c4;
    LUT4 mux_231_Mux_3_i924_3_lut (.A(n908_adj_2898), .B(index_i[0]), .C(index_i[4]), 
         .Z(n924_adj_2899)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_3_i924_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_3_i891_3_lut (.A(n541_adj_2896), .B(n890_adj_2879), 
         .C(index_i[4]), .Z(n891_adj_2900)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_3_i891_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_3_i669_3_lut (.A(n653_adj_2830), .B(n668_adj_2880), 
         .C(index_i[4]), .Z(n669_adj_2901)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_3_i669_3_lut.init = 16'hcaca;
    LUT4 i9544_4_lut (.A(n27372), .B(n29920), .C(index_i[3]), .D(index_i[4]), 
         .Z(n12030)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B ((D)+!C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9544_4_lut.init = 16'h3afa;
    LUT4 i22230_3_lut (.A(n21918), .B(n21919), .C(index_i[4]), .Z(n21920)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22230_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_3_i476_3_lut (.A(n460_adj_2871), .B(n285), .C(index_i[4]), 
         .Z(n476_adj_2902)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_3_i476_3_lut.init = 16'hcaca;
    PFUMX i19517 (.BLUT(n21870), .ALUT(n21871), .C0(index_i[4]), .Z(n21872));
    LUT4 mux_231_Mux_3_i413_3_lut (.A(n397_adj_2903), .B(n27329), .C(index_i[4]), 
         .Z(n413_adj_2904)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_3_i413_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_3_i286_4_lut (.A(n93_adj_2905), .B(index_i[2]), .C(index_i[4]), 
         .D(n15081), .Z(n286_adj_2906)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_3_i286_4_lut.init = 16'h3aca;
    LUT4 i19549_3_lut (.A(n29933), .B(n325), .C(index_i[3]), .Z(n21904)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19549_3_lut.init = 16'hcaca;
    LUT4 i22278_3_lut (.A(n21903), .B(n21904), .C(index_i[4]), .Z(n21905)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22278_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_3_i158_3_lut (.A(n142_adj_2907), .B(n27132), .C(index_i[4]), 
         .Z(n158_adj_2908)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_3_i158_3_lut.init = 16'hcaca;
    LUT4 i12473_3_lut (.A(index_i[3]), .B(index_i[1]), .C(index_i[0]), 
         .Z(n15075)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12473_3_lut.init = 16'hecec;
    LUT4 mux_231_Mux_3_i125_3_lut (.A(n46), .B(n30), .C(index_i[4]), .Z(n125)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_3_i125_3_lut.init = 16'hcaca;
    LUT4 i19545_3_lut (.A(n14), .B(n27379), .C(index_i[3]), .Z(n21900)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19545_3_lut.init = 16'hcaca;
    LUT4 i19495_3_lut_4_lut (.A(n27374), .B(index_i[1]), .C(index_i[3]), 
         .D(n404), .Z(n21850)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19495_3_lut_4_lut.init = 16'hdfd0;
    PFUMX i19523 (.BLUT(n21876), .ALUT(n21877), .C0(index_i[4]), .Z(n21878));
    LUT4 mux_231_Mux_0_i173_3_lut_4_lut (.A(n27374), .B(index_i[1]), .C(index_i[3]), 
         .D(n27406), .Z(n173_adj_2824)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_0_i173_3_lut_4_lut.init = 16'hdfd0;
    LUT4 mux_231_Mux_1_i620_3_lut_4_lut (.A(n27374), .B(index_i[1]), .C(index_i[3]), 
         .D(n27397), .Z(n620)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_1_i620_3_lut_4_lut.init = 16'hdfd0;
    LUT4 n476_bdd_3_lut_24509 (.A(n476), .B(n25478), .C(index_i[5]), .Z(n25479)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n476_bdd_3_lut_24509.init = 16'hcaca;
    PFUMX i23367 (.BLUT(n24968), .ALUT(n23368), .C0(index_i[8]), .Z(n24969));
    LUT4 i19543_3_lut (.A(n723), .B(n325), .C(index_i[3]), .Z(n21898)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19543_3_lut.init = 16'hcaca;
    LUT4 n25481_bdd_3_lut (.A(n27521), .B(n444_adj_2909), .C(index_i[5]), 
         .Z(n25482)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n25481_bdd_3_lut.init = 16'hcaca;
    LUT4 i9653_3_lut_then_4_lut (.A(index_i[4]), .B(index_i[0]), .C(index_i[1]), 
         .D(index_i[2]), .Z(n27514)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C+(D)))+!A (B (C+(D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9653_3_lut_then_4_lut.init = 16'hd54a;
    LUT4 mux_231_Mux_5_i781_3_lut_4_lut_4_lut_then_4_lut (.A(index_i[3]), 
         .B(index_i[0]), .C(index_i[4]), .D(index_i[2]), .Z(n27453)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_5_i781_3_lut_4_lut_4_lut_then_4_lut.init = 16'hece0;
    LUT4 mux_231_Mux_7_i412_3_lut (.A(n27419), .B(n27337), .C(index_i[3]), 
         .Z(n412_adj_2844)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_7_i412_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_1_i924_3_lut (.A(n908_adj_2910), .B(n412), .C(index_i[4]), 
         .Z(n924_adj_2911)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_1_i924_3_lut.init = 16'hcaca;
    LUT4 i22269_3_lut (.A(n22332), .B(n22333), .C(index_i[4]), .Z(n22334)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22269_3_lut.init = 16'hcaca;
    LUT4 i21284_4_lut (.A(n21911), .B(n1002_adj_2912), .C(index_i[5]), 
         .D(index_i[4]), .Z(n23658)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;
    defparam i21284_4_lut.init = 16'hfaca;
    LUT4 mux_231_Mux_4_i860_3_lut (.A(n506), .B(n25682), .C(index_i[4]), 
         .Z(n860_adj_2913)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_4_i860_3_lut.init = 16'hcaca;
    LUT4 i22280_3_lut (.A(n21900), .B(n21901), .C(index_i[4]), .Z(n21902)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22280_3_lut.init = 16'hcaca;
    LUT4 i20362_2_lut (.A(index_i[3]), .B(index_i[5]), .Z(n22736)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20362_2_lut.init = 16'h8888;
    LUT4 i22282_3_lut (.A(n21897), .B(n21898), .C(index_i[4]), .Z(n21899)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22282_3_lut.init = 16'hcaca;
    LUT4 n21800_bdd_3_lut (.A(n21800), .B(n28006), .C(index_i[7]), .Z(n24971)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n21800_bdd_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_1_i349_3_lut (.A(n541_adj_2864), .B(n348_adj_2914), 
         .C(index_i[4]), .Z(n349_adj_2915)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_1_i349_3_lut.init = 16'hcaca;
    LUT4 i22286_3_lut (.A(n22260), .B(n22261), .C(index_i[4]), .Z(n22262)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22286_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_4_i700_3_lut (.A(n684_adj_2916), .B(index_i[1]), .C(index_i[4]), 
         .Z(n700_adj_2917)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_4_i700_3_lut.init = 16'hcaca;
    LUT4 i19536_3_lut (.A(n29957), .B(n29917), .C(index_i[3]), .Z(n21891)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19536_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_4_i669_3_lut (.A(n781_adj_2876), .B(n668_adj_2918), 
         .C(index_i[4]), .Z(n669_adj_2919)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_4_i669_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_4_i542_3_lut (.A(n30), .B(n541_adj_2864), .C(index_i[4]), 
         .Z(n542_adj_2920)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_4_i542_3_lut.init = 16'hcaca;
    LUT4 i12688_2_lut_3_lut_4_lut (.A(n27128), .B(index_i[4]), .C(index_i[6]), 
         .D(index_i[5]), .Z(n15304)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12688_2_lut_3_lut_4_lut.init = 16'hfef0;
    LUT4 i21278_4_lut (.A(n27207), .B(n27512), .C(index_i[5]), .D(index_i[4]), 
         .Z(n23652)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam i21278_4_lut.init = 16'hc5ca;
    LUT4 mux_231_Mux_10_i574_4_lut_4_lut (.A(n27128), .B(index_i[4]), .C(index_i[5]), 
         .D(n27103), .Z(n574)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_10_i574_4_lut_4_lut.init = 16'h1f1c;
    LUT4 mux_231_Mux_1_i94_3_lut (.A(index_i[0]), .B(n93_adj_2921), .C(index_i[4]), 
         .Z(n94)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_1_i94_3_lut.init = 16'hcaca;
    LUT4 n21800_bdd_3_lut_23369 (.A(n23280), .B(n23287), .C(index_i[7]), 
         .Z(n24970)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n21800_bdd_3_lut_23369.init = 16'hcaca;
    LUT4 mux_231_Mux_4_i286_3_lut (.A(n270), .B(n15_adj_2875), .C(index_i[4]), 
         .Z(n286_adj_2922)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_4_i286_3_lut.init = 16'hcaca;
    LUT4 i11514_2_lut_rep_400_3_lut_4_lut (.A(n27130), .B(index_i[4]), .C(index_i[6]), 
         .D(index_i[5]), .Z(n27065)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11514_2_lut_rep_400_3_lut_4_lut.init = 16'hf080;
    LUT4 mux_231_Mux_4_i94_3_lut (.A(n61), .B(n27330), .C(index_i[4]), 
         .Z(n94_adj_2923)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_4_i94_3_lut.init = 16'hcaca;
    LUT4 i9653_3_lut_else_4_lut (.A(index_i[4]), .B(index_i[0]), .C(index_i[1]), 
         .D(index_i[2]), .Z(n27513)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A !(B (D)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9653_3_lut_else_4_lut.init = 16'ha955;
    PFUMX i25182 (.BLUT(n27516), .ALUT(n27517), .C0(index_i[0]), .Z(n27518));
    LUT4 i19531_3_lut (.A(n27406), .B(n27376), .C(index_i[3]), .Z(n21886)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19531_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_6_i158_3_lut_then_4_lut (.A(index_i[4]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n27517)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (D))+!A !(B (D)+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_6_i158_3_lut_then_4_lut.init = 16'h4c33;
    LUT4 i19530_3_lut (.A(n27370), .B(n325), .C(index_i[3]), .Z(n21885)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19530_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_5_i891_3_lut (.A(n875_adj_2924), .B(n379_adj_2846), 
         .C(index_i[4]), .Z(n891_adj_2925)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_5_i891_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_5_i860_3_lut (.A(n15_adj_2926), .B(n859_adj_2927), 
         .C(index_i[4]), .Z(n860_adj_2928)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_5_i860_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_6_i158_3_lut_else_4_lut (.A(index_i[4]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n27516)) /* synthesis lut_function=(A (D)+!A (B (C+!(D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_6_i158_3_lut_else_4_lut.init = 16'hfb44;
    LUT4 i22297_3_lut (.A(n21885), .B(n21886), .C(index_i[4]), .Z(n21887)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22297_3_lut.init = 16'hcaca;
    LUT4 i19528_3_lut (.A(n27377), .B(n27366), .C(index_i[3]), .Z(n21883)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19528_3_lut.init = 16'hcaca;
    LUT4 i22299_3_lut (.A(n21882), .B(n21883), .C(index_i[4]), .Z(n21884)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22299_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_5_i781_3_lut_4_lut_4_lut_else_4_lut (.A(index_i[3]), 
         .B(index_i[0]), .C(index_i[4]), .Z(n27452)) /* synthesis lut_function=(!(A (C)+!A (B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_5_i781_3_lut_4_lut_4_lut_else_4_lut.init = 16'h1f1f;
    LUT4 i22328_3_lut (.A(n21873), .B(n21874), .C(index_i[4]), .Z(n21875)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22328_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_5_i636_4_lut (.A(n157), .B(n27206), .C(index_i[4]), 
         .D(index_i[3]), .Z(n636_adj_2929)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_5_i636_4_lut.init = 16'h3aca;
    LUT4 i22302_3_lut (.A(n21879), .B(n21880), .C(index_i[4]), .Z(n21881)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22302_3_lut.init = 16'hcaca;
    LUT4 i22331_3_lut (.A(n18102), .B(n18103), .C(index_i[4]), .Z(n18104)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22331_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_5_i507_3_lut (.A(n491_adj_2930), .B(n506), .C(index_i[4]), 
         .Z(n507_adj_2931)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_5_i507_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_5_i476_3_lut (.A(n460_adj_2932), .B(n475_adj_2933), 
         .C(index_i[4]), .Z(n476_adj_2934)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_5_i476_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_5_i413_3_lut (.A(n397_adj_2935), .B(n251_adj_2815), 
         .C(index_i[4]), .Z(n413_adj_2936)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_5_i413_3_lut.init = 16'hcaca;
    LUT4 i15936_3_lut (.A(n18120), .B(n18121), .C(index_i[4]), .Z(n18122)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15936_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_5_i125_3_lut (.A(n109_adj_2937), .B(n124), .C(index_i[4]), 
         .Z(n125_adj_2938)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_5_i125_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_5_i94_3_lut (.A(n653_adj_2893), .B(n635), .C(index_i[4]), 
         .Z(n94_adj_2939)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_5_i94_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_5_i31_3_lut (.A(n15_adj_2926), .B(n30_adj_2940), .C(index_i[4]), 
         .Z(n31_adj_2941)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_5_i31_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_2_i270_3_lut (.A(n27399), .B(n27405), .C(index_i[3]), 
         .Z(n270_adj_2942)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_2_i270_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_2_i316_3_lut (.A(n27402), .B(n27379), .C(index_i[3]), 
         .Z(n316_adj_2943)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_2_i316_3_lut.init = 16'hcaca;
    PFUMX i21238 (.BLUT(n31_adj_2941), .ALUT(n22499), .C0(index_i[5]), 
          .Z(n23612));
    LUT4 mux_231_Mux_2_i397_3_lut (.A(n29957), .B(n27419), .C(index_i[3]), 
         .Z(n397_adj_2944)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_2_i397_3_lut.init = 16'hcaca;
    PFUMX i21239 (.BLUT(n94_adj_2939), .ALUT(n125_adj_2938), .C0(index_i[5]), 
          .Z(n23613));
    PFUMX i21240 (.BLUT(n18122), .ALUT(n14735), .C0(index_i[5]), .Z(n23614));
    L6MUX21 i21242 (.D0(n21851), .D1(n21866), .SD(index_i[5]), .Z(n23616));
    L6MUX21 i21243 (.D0(n21869), .D1(n21872), .SD(index_i[5]), .Z(n23617));
    PFUMX i21244 (.BLUT(n413_adj_2936), .ALUT(n444), .C0(index_i[5]), 
          .Z(n23618));
    PFUMX i21245 (.BLUT(n476_adj_2934), .ALUT(n507_adj_2931), .C0(index_i[5]), 
          .Z(n23619));
    PFUMX i21246 (.BLUT(n18104), .ALUT(n573_adj_2945), .C0(index_i[5]), 
          .Z(n23620));
    PFUMX i21247 (.BLUT(n605_adj_2946), .ALUT(n636_adj_2929), .C0(index_i[5]), 
          .Z(n23621));
    LUT4 n699_bdd_4_lut_24029_4_lut_4_lut (.A(index_i[0]), .B(n27372), .C(index_i[4]), 
         .D(index_i[3]), .Z(n25166)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (D))+!A (B (C (D)+!C !(D))+!B (D)))) */ ;
    defparam n699_bdd_4_lut_24029_4_lut_4_lut.init = 16'h0c73;
    PFUMX i21248 (.BLUT(n21875), .ALUT(n700_adj_2947), .C0(index_i[5]), 
          .Z(n23622));
    L6MUX21 i21249 (.D0(n732_adj_2873), .D1(n21878), .SD(index_i[5]), 
            .Z(n23623));
    LUT4 mux_231_Mux_8_i653_3_lut_rep_408_3_lut_4_lut (.A(index_i[0]), .B(n27372), 
         .C(n27225), .D(index_i[3]), .Z(n27073)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(C+(D)))) */ ;
    defparam mux_231_Mux_8_i653_3_lut_rep_408_3_lut_4_lut.init = 16'h77f0;
    PFUMX i21250 (.BLUT(n797_adj_2948), .ALUT(n828_adj_2949), .C0(index_i[5]), 
          .Z(n23624));
    LUT4 i23769_then_4_lut (.A(index_i[0]), .B(index_i[4]), .C(index_i[1]), 
         .D(index_i[3]), .Z(n27520)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam i23769_then_4_lut.init = 16'h3c69;
    LUT4 mux_231_Mux_7_i890_3_lut_3_lut_4_lut (.A(index_i[0]), .B(n27372), 
         .C(index_i[3]), .D(n29920), .Z(n890_adj_2798)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A !(C+(D))) */ ;
    defparam mux_231_Mux_7_i890_3_lut_3_lut_4_lut.init = 16'h808f;
    LUT4 i19932_3_lut_3_lut_4_lut (.A(index_i[0]), .B(n27372), .C(index_i[3]), 
         .D(n27222), .Z(n22287)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A !(C+(D))) */ ;
    defparam i19932_3_lut_3_lut_4_lut.init = 16'h808f;
    LUT4 i11554_3_lut_4_lut (.A(index_i[0]), .B(n27372), .C(n27326), .D(index_i[5]), 
         .Z(n318)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (C (D))) */ ;
    defparam i11554_3_lut_4_lut.init = 16'hf800;
    LUT4 i19629_3_lut_3_lut_4_lut (.A(index_i[0]), .B(n27372), .C(n27222), 
         .D(index_i[3]), .Z(n21984)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(C+(D)))) */ ;
    defparam i19629_3_lut_3_lut_4_lut.init = 16'h77f0;
    LUT4 mux_231_Mux_3_i251_3_lut_4_lut (.A(n27374), .B(index_i[1]), .C(index_i[3]), 
         .D(n27225), .Z(n15342)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_3_i251_3_lut_4_lut.init = 16'hfe0e;
    LUT4 mux_231_Mux_9_i124_3_lut_3_lut_4_lut (.A(n27374), .B(index_i[1]), 
         .C(index_i[3]), .D(n29920), .Z(n124_adj_2884)) /* synthesis lut_function=(!(A (C (D))+!A (B (C (D))+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_9_i124_3_lut_3_lut_4_lut.init = 16'h0efe;
    LUT4 i9499_4_lut_4_lut (.A(n27374), .B(index_i[1]), .C(index_i[3]), 
         .D(n21022), .Z(n11985)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A (B (C)+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9499_4_lut_4_lut.init = 16'h0e3e;
    LUT4 n557_bdd_3_lut_23864_3_lut_4_lut (.A(n27374), .B(index_i[1]), .C(index_i[4]), 
         .D(index_i[3]), .Z(n25577)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n557_bdd_3_lut_23864_3_lut_4_lut.init = 16'hf10f;
    LUT4 i19521_3_lut (.A(n27376), .B(n29942), .C(index_i[3]), .Z(n21876)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19521_3_lut.init = 16'hcaca;
    PFUMX i21251 (.BLUT(n860_adj_2928), .ALUT(n891_adj_2925), .C0(index_i[5]), 
          .Z(n23625));
    LUT4 mux_231_Mux_5_i700_3_lut (.A(n460_adj_2932), .B(n27400), .C(index_i[4]), 
         .Z(n700_adj_2947)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_5_i700_3_lut.init = 16'hcaca;
    LUT4 i19567_3_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[1]), .C(index_i[0]), 
         .D(index_i[3]), .Z(n21922)) /* synthesis lut_function=(A (B (C)+!B !(C+!(D)))+!A (B (C+!(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19567_3_lut_4_lut_4_lut.init = 16'hc3c4;
    LUT4 mux_231_Mux_0_i572_3_lut_4_lut (.A(n27374), .B(index_i[1]), .C(index_i[3]), 
         .D(n29927), .Z(n572)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_0_i572_3_lut_4_lut.init = 16'hefe0;
    PFUMX i25180 (.BLUT(n27513), .ALUT(n27514), .C0(index_i[3]), .Z(n27515));
    LUT4 mux_231_Mux_8_i475_3_lut_3_lut_4_lut (.A(n27374), .B(index_i[1]), 
         .C(index_i[3]), .D(n29920), .Z(n475_adj_2866)) /* synthesis lut_function=(A (C+!(D))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_8_i475_3_lut_3_lut_4_lut.init = 16'he0ef;
    LUT4 i19515_3_lut (.A(n325), .B(n29942), .C(index_i[3]), .Z(n21870)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19515_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_rep_506_4_lut (.A(index_i[3]), .B(index_i[4]), .C(index_i[2]), 
         .D(n27407), .Z(n27171)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_3_lut_rep_506_4_lut.init = 16'hfffe;
    LUT4 i19488_4_lut_4_lut_3_lut_4_lut (.A(n27374), .B(index_i[1]), .C(index_i[4]), 
         .D(index_i[3]), .Z(n21843)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19488_4_lut_4_lut_3_lut_4_lut.init = 16'h11ef;
    LUT4 i11530_2_lut_rep_424_3_lut_4_lut (.A(n27374), .B(index_i[1]), .C(index_i[4]), 
         .D(index_i[3]), .Z(n27089)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11530_2_lut_rep_424_3_lut_4_lut.init = 16'hfef0;
    LUT4 i20022_3_lut (.A(n27366), .B(n27375), .C(index_i[3]), .Z(n22377)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20022_3_lut.init = 16'hcaca;
    LUT4 i22264_3_lut (.A(n22377), .B(n22378), .C(index_i[4]), .Z(n22379)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22264_3_lut.init = 16'hcaca;
    LUT4 n476_bdd_3_lut_23768_4_lut (.A(index_i[2]), .B(n27407), .C(index_i[4]), 
         .D(n491_adj_2950), .Z(n25478)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+(D)))) */ ;
    defparam n476_bdd_3_lut_23768_4_lut.init = 16'h9f90;
    LUT4 i20139_3_lut_3_lut_4_lut (.A(index_i[2]), .B(n27407), .C(n27419), 
         .D(index_i[3]), .Z(n22494)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (B (C (D))+!B (C+!(D)))) */ ;
    defparam i20139_3_lut_3_lut_4_lut.init = 16'hf099;
    PFUMX i21270 (.BLUT(n94_adj_2923), .ALUT(n21881), .C0(index_i[5]), 
          .Z(n23644));
    LUT4 mux_231_Mux_3_i860_3_lut_4_lut (.A(index_i[2]), .B(n27407), .C(index_i[4]), 
         .D(n859_adj_2951), .Z(n860_adj_2952)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam mux_231_Mux_3_i860_3_lut_4_lut.init = 16'hf606;
    LUT4 i19566_3_lut_3_lut_4_lut (.A(index_i[2]), .B(n27407), .C(n204), 
         .D(index_i[3]), .Z(n21921)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (B (C (D))+!B (C+!(D)))) */ ;
    defparam i19566_3_lut_3_lut_4_lut.init = 16'hf099;
    PFUMX i21272 (.BLUT(n221_adj_2953), .ALUT(n252_adj_2954), .C0(index_i[5]), 
          .Z(n23646));
    LUT4 mux_231_Mux_7_i443_3_lut_4_lut (.A(index_i[2]), .B(n27407), .C(index_i[3]), 
         .D(n27419), .Z(n443_adj_2843)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;
    defparam mux_231_Mux_7_i443_3_lut_4_lut.init = 16'h6f60;
    PFUMX i21273 (.BLUT(n286_adj_2922), .ALUT(n21884), .C0(index_i[5]), 
          .Z(n23647));
    LUT4 i20013_3_lut (.A(n38), .B(n14), .C(index_i[3]), .Z(n22368)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20013_3_lut.init = 16'hcaca;
    LUT4 i22266_3_lut (.A(n22368), .B(n22369), .C(index_i[4]), .Z(n22370)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22266_3_lut.init = 16'hcaca;
    PFUMX i21274 (.BLUT(n349_adj_2955), .ALUT(n21887), .C0(index_i[5]), 
          .Z(n23648));
    LUT4 i23769_else_4_lut (.A(index_i[0]), .B(index_i[4]), .C(index_i[1]), 
         .D(index_i[3]), .Z(n27519)) /* synthesis lut_function=(!(A (B (C)+!B !(C (D)+!C !(D)))+!A (B ((D)+!C)+!B !((D)+!C)))) */ ;
    defparam i23769_else_4_lut.init = 16'h394b;
    PFUMX i20848 (.BLUT(n94), .ALUT(n22253), .C0(index_i[5]), .Z(n23222));
    LUT4 i19513_3_lut (.A(n27396), .B(n29933), .C(index_i[3]), .Z(n21868)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19513_3_lut.init = 16'hcaca;
    LUT4 n23294_bdd_3_lut_24305 (.A(n23294), .B(n21806), .C(index_i[7]), 
         .Z(n24968)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n23294_bdd_3_lut_24305.init = 16'hcaca;
    LUT4 i19512_3_lut (.A(n27404), .B(n29927), .C(index_i[3]), .Z(n21867)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19512_3_lut.init = 16'hcaca;
    L6MUX21 i20849 (.D0(n22256), .D1(n22259), .SD(index_i[5]), .Z(n23223));
    PFUMX i21279 (.BLUT(n669_adj_2919), .ALUT(n700_adj_2917), .C0(index_i[5]), 
          .Z(n23653));
    PFUMX i19538 (.BLUT(n21891), .ALUT(n21892), .C0(index_i[4]), .Z(n476));
    LUT4 mux_231_Mux_7_i892_3_lut (.A(n62), .B(n891), .C(index_i[5]), 
         .Z(n892_adj_2813)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_7_i892_3_lut.init = 16'hcaca;
    LUT4 i19510_3_lut (.A(n29939), .B(n29927), .C(index_i[3]), .Z(n21865)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19510_3_lut.init = 16'hcaca;
    LUT4 i19585_3_lut (.A(n747_adj_2956), .B(n762_adj_2957), .C(index_i[4]), 
         .Z(n21940)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19585_3_lut.init = 16'hcaca;
    LUT4 i22053_3_lut (.A(n491_adj_2958), .B(n506_adj_2959), .C(index_i[4]), 
         .Z(n21862)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22053_3_lut.init = 16'hcaca;
    LUT4 i19584_3_lut (.A(n716_adj_2960), .B(n15042), .C(index_i[4]), 
         .Z(n21939)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19584_3_lut.init = 16'hcaca;
    PFUMX i20851 (.BLUT(n22262), .ALUT(n317_adj_2961), .C0(index_i[5]), 
          .Z(n23225));
    PFUMX i20852 (.BLUT(n349_adj_2915), .ALUT(n22271), .C0(index_i[5]), 
          .Z(n23226));
    LUT4 mux_231_Mux_5_i15_3_lut (.A(n27399), .B(n29917), .C(index_i[3]), 
         .Z(n15_adj_2926)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_5_i15_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_6_i653_3_lut (.A(n27415), .B(n77), .C(index_i[3]), 
         .Z(n653_adj_2893)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_6_i653_3_lut.init = 16'hcaca;
    LUT4 i19987_3_lut (.A(n27379), .B(n27404), .C(index_i[3]), .Z(n22342)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19987_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_5_i397_3_lut (.A(n27396), .B(n27331), .C(index_i[3]), 
         .Z(n397_adj_2935)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_5_i397_3_lut.init = 16'hcaca;
    PFUMX i21280 (.BLUT(n21899), .ALUT(n763_adj_2881), .C0(index_i[5]), 
          .Z(n23654));
    LUT4 mux_231_Mux_5_i506_3_lut (.A(n27366), .B(n29943), .C(index_i[3]), 
         .Z(n506)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_5_i506_3_lut.init = 16'hcaca;
    PFUMX i21281 (.BLUT(n21902), .ALUT(n828_adj_2962), .C0(index_i[5]), 
          .Z(n23655));
    LUT4 mux_231_Mux_5_i859_3_lut (.A(n250), .B(n27399), .C(index_i[3]), 
         .Z(n859_adj_2927)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_5_i859_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_5_i875_3_lut (.A(n204), .B(n27417), .C(index_i[3]), 
         .Z(n875_adj_2924)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_5_i875_3_lut.init = 16'hcaca;
    PFUMX i21282 (.BLUT(n860_adj_2913), .ALUT(n21905), .C0(index_i[5]), 
          .Z(n23656));
    LUT4 i19582_3_lut (.A(n93_adj_2870), .B(n699), .C(index_i[4]), .Z(n21937)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19582_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_5_i731_3_lut (.A(n29942), .B(n29933), .C(index_i[3]), 
         .Z(n731_adj_2872)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_5_i731_3_lut.init = 16'hcaca;
    LUT4 i19581_3_lut (.A(n653), .B(n27100), .C(index_i[4]), .Z(n21936)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19581_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_4_i61_3_lut (.A(n27379), .B(n27333), .C(index_i[3]), 
         .Z(n61)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_4_i61_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_4_i270_3_lut (.A(n27397), .B(n27366), .C(index_i[3]), 
         .Z(n270)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_4_i270_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_4_i15_3_lut (.A(n29943), .B(n14), .C(index_i[3]), 
         .Z(n15_adj_2875)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_4_i15_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_4_i348_3_lut (.A(n27360), .B(n27406), .C(index_i[3]), 
         .Z(n348_adj_2963)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_4_i348_3_lut.init = 16'hcaca;
    L6MUX21 i20853 (.D0(n22280), .D1(n22289), .SD(index_i[5]), .Z(n23227));
    LUT4 mux_231_Mux_4_i684_3_lut (.A(n77), .B(n108), .C(index_i[3]), 
         .Z(n684_adj_2916)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_4_i684_3_lut.init = 16'hcaca;
    LUT4 i22917_3_lut_4_lut (.A(n27204), .B(n20104), .C(index_i[8]), .D(n766), 
         .Z(n21754)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i22917_3_lut_4_lut.init = 16'hefe0;
    LUT4 i15945_3_lut (.A(n27369), .B(n27396), .C(index_i[3]), .Z(n18131)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15945_3_lut.init = 16'hcaca;
    LUT4 i15944_3_lut (.A(n27396), .B(n27406), .C(index_i[3]), .Z(n18130)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15944_3_lut.init = 16'hcaca;
    LUT4 i23058_2_lut_rep_418_3_lut_4_lut (.A(n27413), .B(index_i[2]), .C(index_i[5]), 
         .D(n27326), .Z(n27083)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A (C (D)))) */ ;
    defparam i23058_2_lut_rep_418_3_lut_4_lut.init = 16'h0f7f;
    L6MUX21 i20854 (.D0(n22298), .D1(n22307), .SD(index_i[5]), .Z(n23228));
    LUT4 mux_231_Mux_8_i78_3_lut_4_lut (.A(n27413), .B(index_i[2]), .C(index_i[3]), 
         .D(n27412), .Z(n78)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam mux_231_Mux_8_i78_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_231_Mux_1_i986_3_lut (.A(n27417), .B(n27398), .C(index_i[3]), 
         .Z(n986_adj_2964)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_1_i986_3_lut.init = 16'hcaca;
    LUT4 i22857_3_lut_rep_402_4_lut (.A(n27171), .B(index_i[5]), .C(index_i[8]), 
         .D(n1021), .Z(n27067)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i22857_3_lut_rep_402_4_lut.init = 16'hf808;
    L6MUX21 i20856 (.D0(n22325), .D1(n636_adj_2795), .SD(index_i[5]), 
            .Z(n23230));
    PFUMX i20857 (.BLUT(n22334), .ALUT(n700), .C0(index_i[5]), .Z(n23231));
    LUT4 i22450_3_lut (.A(n716_adj_2965), .B(n731_adj_2966), .C(index_i[4]), 
         .Z(n732_adj_2868)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22450_3_lut.init = 16'hcaca;
    L6MUX21 i20859 (.D0(n22343), .D1(n22352), .SD(index_i[5]), .Z(n23233));
    LUT4 mux_231_Mux_2_i669_3_lut (.A(n653_adj_2967), .B(n475), .C(index_i[4]), 
         .Z(n669)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_2_i669_3_lut.init = 16'hcaca;
    PFUMX i20861 (.BLUT(n924_adj_2911), .ALUT(n22370), .C0(index_i[5]), 
          .Z(n23235));
    LUT4 mux_231_Mux_2_i605_3_lut (.A(n142_adj_2907), .B(n604_adj_2968), 
         .C(index_i[4]), .Z(n605_adj_2867)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_2_i605_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_8_i173_3_lut_3_lut_4_lut (.A(n27413), .B(index_i[2]), 
         .C(n954_adj_2969), .D(index_i[4]), .Z(n173_adj_2818)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C+!(D))) */ ;
    defparam mux_231_Mux_8_i173_3_lut_3_lut_4_lut.init = 16'hf077;
    LUT4 i19572_3_lut (.A(n526_adj_2970), .B(n541_adj_2856), .C(index_i[4]), 
         .Z(n21927)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19572_3_lut.init = 16'hcaca;
    LUT4 i12479_3_lut (.A(index_i[3]), .B(index_i[1]), .C(index_i[0]), 
         .Z(n15081)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12479_3_lut.init = 16'hc8c8;
    LUT4 mux_231_Mux_3_i348_3_lut (.A(n27398), .B(n27404), .C(index_i[3]), 
         .Z(n348)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_3_i348_3_lut.init = 16'hcaca;
    LUT4 i22456_3_lut (.A(n27577), .B(n21991), .C(index_i[4]), .Z(n21992)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22456_3_lut.init = 16'hcaca;
    LUT4 i19494_3_lut (.A(n27376), .B(n29927), .C(index_i[3]), .Z(n21849)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19494_3_lut.init = 16'hcaca;
    LUT4 i22458_3_lut (.A(n21987), .B(n21988), .C(index_i[4]), .Z(n21989)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22458_3_lut.init = 16'hcaca;
    PFUMX i20862 (.BLUT(n987), .ALUT(n22379), .C0(index_i[5]), .Z(n23236));
    LUT4 mux_231_Mux_2_i413_3_lut (.A(n397_adj_2944), .B(n954_adj_2969), 
         .C(index_i[4]), .Z(n413_adj_2862)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_2_i413_3_lut.init = 16'hcaca;
    LUT4 i19977_3_lut_3_lut_4_lut (.A(n27413), .B(index_i[2]), .C(n38), 
         .D(index_i[3]), .Z(n22332)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C+!(D))) */ ;
    defparam i19977_3_lut_3_lut_4_lut.init = 16'hf077;
    LUT4 mux_231_Mux_2_i317_3_lut (.A(n668_adj_2880), .B(n316_adj_2943), 
         .C(index_i[4]), .Z(n317_adj_2860)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_2_i317_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_2_i286_3_lut (.A(n270_adj_2942), .B(n653_adj_2830), 
         .C(index_i[4]), .Z(n286_adj_2859)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_2_i286_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_3_i828_3_lut_3_lut_4_lut_4_lut_4_lut (.A(n27413), .B(index_i[2]), 
         .C(index_i[4]), .D(index_i[3]), .Z(n828)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C (D)+!C !(D)))+!A !(B (C+!(D))+!B (C (D)+!C !(D))))) */ ;
    defparam mux_231_Mux_3_i828_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h70c7;
    LUT4 mux_231_Mux_0_i986_3_lut (.A(n29930), .B(n985), .C(index_i[3]), 
         .Z(n986)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_0_i986_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_0_i971_3_lut (.A(n29927), .B(n27422), .C(index_i[3]), 
         .Z(n971)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_0_i971_3_lut.init = 16'hcaca;
    PFUMX i19420 (.BLUT(n445), .ALUT(n508), .C0(index_i[6]), .Z(n21775));
    LUT4 mux_231_Mux_3_i908_3_lut (.A(n27375), .B(n27333), .C(index_i[3]), 
         .Z(n908_adj_2898)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_3_i908_3_lut.init = 16'hcaca;
    LUT4 i22467_3_lut (.A(n142), .B(n14323), .C(index_i[4]), .Z(n158_adj_2857)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22467_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_3_i93_3_lut_4_lut (.A(n27407), .B(index_i[2]), .C(index_i[3]), 
         .D(n27412), .Z(n93_adj_2905)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_3_i93_3_lut_4_lut.init = 16'hefe0;
    LUT4 mux_231_Mux_3_i747_3_lut (.A(n27376), .B(n404), .C(index_i[3]), 
         .Z(n747_adj_2854)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_3_i747_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_6_i890_3_lut_3_lut_4_lut (.A(n27407), .B(index_i[2]), 
         .C(n27422), .D(index_i[3]), .Z(n890_adj_2888)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_6_i890_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 mux_231_Mux_0_i1002_3_lut_3_lut_4_lut (.A(n27407), .B(index_i[2]), 
         .C(n38), .D(index_i[3]), .Z(n1002)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_0_i1002_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 i19942_3_lut (.A(n29943), .B(n27401), .C(index_i[3]), .Z(n22297)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19942_3_lut.init = 16'hcaca;
    PFUMX i23771 (.BLUT(n25482), .ALUT(n25479), .C0(index_i[6]), .Z(n23662));
    PFUMX i25178 (.BLUT(n27510), .ALUT(n27511), .C0(index_i[0]), .Z(n27512));
    LUT4 i11931_3_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .Z(n11192)) /* synthesis lut_function=(!((B (C))+!A)) */ ;
    defparam i11931_3_lut.init = 16'h2a2a;
    LUT4 i19476_3_lut_then_4_lut (.A(index_i[4]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n27532)) /* synthesis lut_function=(A (B (C)+!B !(C (D)+!C !(D)))+!A !(B (C)+!B !(C (D)+!C !(D)))) */ ;
    defparam i19476_3_lut_then_4_lut.init = 16'h96a5;
    LUT4 mux_231_Mux_0_i939_4_lut (.A(n14), .B(n27364), .C(index_i[3]), 
         .D(index_i[2]), .Z(n939)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_0_i939_4_lut.init = 16'hfaca;
    LUT4 i19476_3_lut_else_4_lut (.A(index_i[4]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n27531)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C+!(D)))+!A !(B ((D)+!C)+!B (C (D)+!C !(D))))) */ ;
    defparam i19476_3_lut_else_4_lut.init = 16'h5685;
    LUT4 mux_231_Mux_0_i923_3_lut (.A(n27419), .B(n27408), .C(index_i[3]), 
         .Z(n923)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_0_i923_3_lut.init = 16'hcaca;
    LUT4 i19477_3_lut_then_4_lut (.A(index_i[4]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n27535)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)+!C !(D)))+!A !(B (C+!(D))+!B (C (D)+!C !(D))))) */ ;
    defparam i19477_3_lut_then_4_lut.init = 16'h5a65;
    LUT4 mux_231_Mux_12_i254_4_lut (.A(n27083), .B(n20892), .C(index_i[6]), 
         .D(n29920), .Z(n254_adj_2971)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_12_i254_4_lut.init = 16'hca0a;
    LUT4 i12579_2_lut (.A(index_i[1]), .B(index_i[3]), .Z(n541)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i12579_2_lut.init = 16'h1111;
    LUT4 mux_231_Mux_0_i526_3_lut (.A(n27406), .B(n27379), .C(index_i[3]), 
         .Z(n526_adj_2848)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_0_i526_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_6_i668_3_lut (.A(n108), .B(n27418), .C(index_i[3]), 
         .Z(n668_adj_2894)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_6_i668_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_6_i684_3_lut (.A(n204), .B(n29957), .C(index_i[3]), 
         .Z(n684_adj_2852)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_6_i684_3_lut.init = 16'hcaca;
    LUT4 i19477_3_lut_else_4_lut (.A(index_i[4]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n27534)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A !(B (C+!(D))+!B ((D)+!C)))) */ ;
    defparam i19477_3_lut_else_4_lut.init = 16'h59e5;
    LUT4 index_i_7__bdd_4_lut_25550 (.A(index_i[7]), .B(n125_adj_2972), 
         .C(n25180), .D(index_i[5]), .Z(n27063)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(B (C+(D))+!B !((D)+!C)))) */ ;
    defparam index_i_7__bdd_4_lut_25550.init = 16'h66f0;
    LUT4 i19923_3_lut (.A(n27379), .B(n29942), .C(index_i[3]), .Z(n22278)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19923_3_lut.init = 16'hcaca;
    PFUMX i20904 (.BLUT(n23274), .ALUT(n23275), .C0(index_i[5]), .Z(n23278));
    PFUMX i20905 (.BLUT(n23276), .ALUT(n23277), .C0(index_i[5]), .Z(n23279));
    PFUMX i20911 (.BLUT(n23281), .ALUT(n23282), .C0(index_i[5]), .Z(n23285));
    LUT4 i22284_3_lut (.A(n22269), .B(n22270), .C(index_i[4]), .Z(n22271)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22284_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_0_i716_3_lut (.A(n27378), .B(n27333), .C(index_i[3]), 
         .Z(n716_adj_2836)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_0_i716_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_0_i653_3_lut (.A(n204), .B(n27366), .C(index_i[3]), 
         .Z(n653_adj_2834)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_0_i653_3_lut.init = 16'hcaca;
    PFUMX i20912 (.BLUT(n23283), .ALUT(n23284), .C0(index_i[5]), .Z(n23286));
    LUT4 mux_231_Mux_0_i620_3_lut (.A(n27417), .B(n27397), .C(index_i[3]), 
         .Z(n620_adj_2832)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_0_i620_3_lut.init = 16'hcaca;
    PFUMX i21332 (.BLUT(n94_adj_2973), .ALUT(n125), .C0(index_i[5]), .Z(n23706));
    LUT4 mux_231_Mux_0_i397_3_lut (.A(n27408), .B(n29933), .C(index_i[3]), 
         .Z(n397_adj_2828)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_0_i397_3_lut.init = 16'hcaca;
    PFUMX i21333 (.BLUT(n158_adj_2908), .ALUT(n189), .C0(index_i[5]), 
          .Z(n23707));
    PFUMX i21334 (.BLUT(n221), .ALUT(n252), .C0(index_i[5]), .Z(n23708));
    LUT4 mux_231_Mux_7_i956_3_lut_3_lut_4_lut (.A(n27196), .B(index_i[4]), 
         .C(n924_adj_2974), .D(index_i[5]), .Z(n956)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_7_i956_3_lut_3_lut_4_lut.init = 16'h11f0;
    LUT4 i20441_3_lut_3_lut_4_lut (.A(n27196), .B(index_i[4]), .C(n252_adj_2802), 
         .D(index_i[5]), .Z(n22815)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20441_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 mux_231_Mux_10_i701_4_lut_4_lut (.A(n27196), .B(index_i[4]), .C(index_i[5]), 
         .D(n27129), .Z(n701)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B (C (D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_10_i701_4_lut_4_lut.init = 16'h3efe;
    PFUMX i21335 (.BLUT(n286_adj_2906), .ALUT(n21914), .C0(index_i[5]), 
          .Z(n23709));
    PFUMX i21336 (.BLUT(n349), .ALUT(n21917), .C0(index_i[5]), .Z(n23710));
    LUT4 i22563_3_lut (.A(n286), .B(n317), .C(index_i[5]), .Z(n22805)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22563_3_lut.init = 16'hcaca;
    PFUMX i21337 (.BLUT(n413_adj_2904), .ALUT(n444_adj_2975), .C0(index_i[5]), 
          .Z(n23711));
    LUT4 mux_231_Mux_1_i317_3_lut (.A(n301), .B(n908), .C(index_i[4]), 
         .Z(n317_adj_2961)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_1_i317_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_4_lut (.A(index_i[3]), .B(index_i[4]), .C(index_i[5]), 
         .D(n27372), .Z(n20737)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_3_lut_4_lut.init = 16'hfffe;
    PFUMX i21338 (.BLUT(n476_adj_2902), .ALUT(n507_adj_2976), .C0(index_i[5]), 
          .Z(n23712));
    PFUMX i21339 (.BLUT(n21920), .ALUT(n573_adj_2886), .C0(index_i[5]), 
          .Z(n23713));
    PFUMX i21340 (.BLUT(n12030), .ALUT(n21923), .C0(index_i[5]), .Z(n23714));
    LUT4 i22648_3_lut (.A(n28835), .B(n27548), .C(index_i[5]), .Z(n23657)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22648_3_lut.init = 16'hcaca;
    LUT4 i22653_3_lut (.A(n542_adj_2920), .B(n573_adj_2883), .C(index_i[5]), 
         .Z(n23651)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22653_3_lut.init = 16'hcaca;
    PFUMX i21341 (.BLUT(n669_adj_2901), .ALUT(n700_adj_2977), .C0(index_i[5]), 
          .Z(n23715));
    L6MUX21 i21342 (.D0(n21926), .D1(n763_adj_2855), .SD(index_i[5]), 
            .Z(n23716));
    PFUMX i21344 (.BLUT(n860_adj_2952), .ALUT(n891_adj_2900), .C0(index_i[5]), 
          .Z(n23718));
    PFUMX i21345 (.BLUT(n924_adj_2899), .ALUT(n21932), .C0(index_i[5]), 
          .Z(n23719));
    LUT4 mux_231_Mux_1_i732_3_lut (.A(n716), .B(n491_adj_2930), .C(index_i[4]), 
         .Z(n732)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_1_i732_3_lut.init = 16'hcaca;
    LUT4 i22967_2_lut_rep_597 (.A(index_i[1]), .B(index_i[2]), .Z(n27262)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i22967_2_lut_rep_597.init = 16'h9999;
    LUT4 mux_231_Mux_0_i93_3_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .Z(n93_adj_2803)) /* synthesis lut_function=(A (B)+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_0_i93_3_lut_3_lut.init = 16'h9c9c;
    LUT4 mux_231_Mux_10_i637_3_lut_4_lut_4_lut (.A(n27205), .B(index_i[4]), 
         .C(index_i[5]), .D(n27128), .Z(n637)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_10_i637_3_lut_4_lut_4_lut.init = 16'h1f1c;
    LUT4 mux_231_Mux_0_i188_3_lut (.A(n27418), .B(n101), .C(index_i[3]), 
         .Z(n188)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_0_i188_3_lut.init = 16'hcaca;
    PFUMX i21346 (.BLUT(n21974), .ALUT(n1018), .C0(index_i[5]), .Z(n23720));
    LUT4 n442_bdd_2_lut_24331_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[3]), 
         .Z(n26053)) /* synthesis lut_function=(A (B+(C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n442_bdd_2_lut_24331_3_lut.init = 16'hf9f9;
    LUT4 i22892_3_lut (.A(n22798), .B(n22799), .C(index_i[8]), .Z(n22802)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22892_3_lut.init = 16'hcaca;
    LUT4 n699_bdd_4_lut (.A(n27129), .B(index_i[6]), .C(n27160), .D(index_i[5]), 
         .Z(n25741)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C+!(D))+!B (D))) */ ;
    defparam n699_bdd_4_lut.init = 16'hd1cc;
    L6MUX21 i21378 (.D0(n22466), .D1(n22472), .SD(index_i[5]), .Z(n23752));
    L6MUX21 i21382 (.D0(n22481), .D1(n18132), .SD(index_i[5]), .Z(n23756));
    L6MUX21 i21383 (.D0(n22487), .D1(n11994), .SD(index_i[5]), .Z(n23757));
    PFUMX i21385 (.BLUT(n542_adj_2897), .ALUT(n573_adj_2978), .C0(index_i[5]), 
          .Z(n23759));
    PFUMX i21386 (.BLUT(n605), .ALUT(n636), .C0(index_i[5]), .Z(n23760));
    LUT4 i23116_2_lut_rep_600 (.A(index_i[4]), .B(index_i[3]), .Z(n27265)) /* synthesis lut_function=((B)+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i23116_2_lut_rep_600.init = 16'hdddd;
    PFUMX i19556 (.BLUT(n21909), .ALUT(n21910), .C0(index_i[4]), .Z(n21911));
    PFUMX i21387 (.BLUT(n669_adj_2895), .ALUT(n700_adj_2853), .C0(index_i[5]), 
          .Z(n23761));
    PFUMX i21388 (.BLUT(n732_adj_2851), .ALUT(n22496), .C0(index_i[5]), 
          .Z(n23762));
    L6MUX21 i24771 (.D0(n26580), .D1(n26578), .SD(index_i[5]), .Z(n26581));
    PFUMX i21389 (.BLUT(n797_adj_2892), .ALUT(n828_adj_2891), .C0(index_i[5]), 
          .Z(n23763));
    LUT4 mux_231_Mux_3_i797_3_lut_4_lut (.A(index_i[4]), .B(index_i[3]), 
         .C(n796_adj_2979), .D(n27412), .Z(n797)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_3_i797_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i8904_4_lut_4_lut (.A(index_i[3]), .B(index_i[0]), .C(index_i[1]), 
         .D(index_i[2]), .Z(n11349)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (D)+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i8904_4_lut_4_lut.init = 16'h0bf4;
    PFUMX i21390 (.BLUT(n860_adj_2801), .ALUT(n891_adj_2889), .C0(index_i[5]), 
          .Z(n23764));
    PFUMX i24769 (.BLUT(n26579), .ALUT(n204), .C0(index_i[3]), .Z(n26580));
    PFUMX mux_231_Mux_1_i891 (.BLUT(n882), .ALUT(n890_adj_2980), .C0(n27265), 
          .Z(n891_adj_2825)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    L6MUX21 i20969 (.D0(n23341), .D1(n23342), .SD(index_i[5]), .Z(n23343));
    LUT4 i20908_3_lut_4_lut_3_lut (.A(index_i[3]), .B(index_i[4]), .C(n29920), 
         .Z(n23282)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20908_3_lut_4_lut_3_lut.init = 16'h6464;
    LUT4 mux_231_Mux_1_i987_3_lut_4_lut_4_lut (.A(index_i[3]), .B(n986_adj_2964), 
         .C(index_i[4]), .D(n27337), .Z(n987)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_1_i987_3_lut_4_lut_4_lut.init = 16'hc5c0;
    LUT4 i12022_4_lut_4_lut (.A(index_i[3]), .B(index_i[2]), .C(index_i[0]), 
         .D(index_i[1]), .Z(n875_adj_2850)) /* synthesis lut_function=((B (C)+!B (D))+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12022_4_lut_4_lut.init = 16'hf7d5;
    LUT4 i19588_4_lut_3_lut (.A(index_i[3]), .B(index_i[4]), .C(n27221), 
         .Z(n21943)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19588_4_lut_3_lut.init = 16'h6565;
    LUT4 mux_231_Mux_2_i221_4_lut_4_lut (.A(index_i[3]), .B(index_i[4]), 
         .C(n27221), .D(n27103), .Z(n221_adj_2858)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (B+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_2_i221_4_lut_4_lut.init = 16'hf7c4;
    LUT4 mux_231_Mux_4_i349_3_lut_4_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[4]), .D(n348_adj_2963), .Z(n349_adj_2955)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_4_i349_3_lut_4_lut.init = 16'hf606;
    LUT4 i9501_3_lut_3_lut (.A(index_i[3]), .B(index_i[4]), .C(n11986), 
         .Z(n11987)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9501_3_lut_3_lut.init = 16'h7474;
    L6MUX21 i20976 (.D0(n23348), .D1(n23349), .SD(index_i[5]), .Z(n23350));
    PFUMX i24767 (.BLUT(n26577), .ALUT(n22459), .C0(index_i[4]), .Z(n26578));
    L6MUX21 i20983 (.D0(n23355), .D1(n23356), .SD(index_i[5]), .Z(n23357));
    LUT4 mux_231_Mux_4_i828_3_lut_4_lut (.A(index_i[4]), .B(index_i[3]), 
         .C(n812), .D(n27368), .Z(n828_adj_2962)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_4_i828_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i21202_3_lut (.A(n23574), .B(n23575), .C(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2145[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21202_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_5_i797_3_lut_4_lut (.A(index_i[4]), .B(index_i[3]), 
         .C(n27454), .D(n27376), .Z(n797_adj_2948)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_5_i797_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i21407_3_lut (.A(n23779), .B(n23780), .C(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2145[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21407_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_1_i763_3_lut_4_lut (.A(index_i[4]), .B(index_i[3]), 
         .C(n27573), .D(n27376), .Z(n763)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_1_i763_3_lut_4_lut.init = 16'hf1e0;
    L6MUX21 i20990 (.D0(n23362), .D1(n23363), .SD(index_i[5]), .Z(n23364));
    LUT4 i21406_3_lut (.A(n23777), .B(n23778), .C(index_i[8]), .Z(n23780)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21406_3_lut.init = 16'hcaca;
    LUT4 mux_188_i16_3_lut (.A(\quarter_wave_sample_register_q[15] ), .B(o_val_pipeline_i_0__15__N_2176[15]), 
         .C(phase_negation_i[1]), .Z(n1087[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam mux_188_i16_3_lut.init = 16'hcaca;
    LUT4 i22123_3_lut (.A(n27481), .B(n124_adj_2817), .C(index_i[4]), 
         .Z(n23403)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22123_3_lut.init = 16'hcaca;
    LUT4 i12476_2_lut_rep_601 (.A(index_i[2]), .B(index_i[0]), .Z(n27266)) /* synthesis lut_function=(A (B)) */ ;
    defparam i12476_2_lut_rep_601.init = 16'h8888;
    LUT4 mux_188_i15_3_lut (.A(quarter_wave_sample_register_i[14]), .B(o_val_pipeline_i_0__15__N_2176[14]), 
         .C(phase_negation_i[1]), .Z(n1087[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam mux_188_i15_3_lut.init = 16'hcaca;
    LUT4 mux_188_i14_3_lut (.A(quarter_wave_sample_register_i[13]), .B(o_val_pipeline_i_0__15__N_2176[13]), 
         .C(phase_negation_i[1]), .Z(n1087[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam mux_188_i14_3_lut.init = 16'hcaca;
    LUT4 mux_188_i13_3_lut (.A(quarter_wave_sample_register_i[12]), .B(o_val_pipeline_i_0__15__N_2176[12]), 
         .C(phase_negation_i[1]), .Z(n1087[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam mux_188_i13_3_lut.init = 16'hcaca;
    PFUMX i21331 (.BLUT(n31_adj_2878), .ALUT(n62_adj_2981), .C0(index_i[5]), 
          .Z(n23705));
    LUT4 mux_188_i12_3_lut (.A(quarter_wave_sample_register_i[11]), .B(o_val_pipeline_i_0__15__N_2176[11]), 
         .C(phase_negation_i[1]), .Z(n1087[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam mux_188_i12_3_lut.init = 16'hcaca;
    LUT4 mux_188_i11_3_lut (.A(quarter_wave_sample_register_i[10]), .B(o_val_pipeline_i_0__15__N_2176[10]), 
         .C(phase_negation_i[1]), .Z(n1087[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam mux_188_i11_3_lut.init = 16'hcaca;
    LUT4 mux_188_i10_3_lut (.A(quarter_wave_sample_register_i[9]), .B(o_val_pipeline_i_0__15__N_2176[9]), 
         .C(phase_negation_i[1]), .Z(n1087[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam mux_188_i10_3_lut.init = 16'hcaca;
    LUT4 mux_188_i9_3_lut (.A(quarter_wave_sample_register_i[8]), .B(o_val_pipeline_i_0__15__N_2176[8]), 
         .C(phase_negation_i[1]), .Z(n1087[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam mux_188_i9_3_lut.init = 16'hcaca;
    LUT4 mux_188_i8_3_lut (.A(quarter_wave_sample_register_i[7]), .B(o_val_pipeline_i_0__15__N_2176[7]), 
         .C(phase_negation_i[1]), .Z(n1087[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam mux_188_i8_3_lut.init = 16'hcaca;
    LUT4 n269_bdd_3_lut_23920 (.A(n27370), .B(index_i[3]), .C(n27401), 
         .Z(n25632)) /* synthesis lut_function=(A (B+(C))+!A !(B+!(C))) */ ;
    defparam n269_bdd_3_lut_23920.init = 16'hb8b8;
    LUT4 n285_bdd_3_lut (.A(n27370), .B(n29933), .C(index_i[3]), .Z(n25635)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n285_bdd_3_lut.init = 16'hacac;
    LUT4 mux_188_i7_3_lut (.A(quarter_wave_sample_register_i[6]), .B(o_val_pipeline_i_0__15__N_2176[6]), 
         .C(phase_negation_i[1]), .Z(n1087[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam mux_188_i7_3_lut.init = 16'hcaca;
    LUT4 n22489_bdd_3_lut (.A(n29930), .B(n29927), .C(index_i[3]), .Z(n25638)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n22489_bdd_3_lut.init = 16'hcaca;
    LUT4 mux_188_i6_3_lut (.A(quarter_wave_sample_register_i[5]), .B(o_val_pipeline_i_0__15__N_2176[5]), 
         .C(phase_negation_i[1]), .Z(n1087[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam mux_188_i6_3_lut.init = 16'hcaca;
    LUT4 mux_188_i5_3_lut (.A(quarter_wave_sample_register_i[4]), .B(o_val_pipeline_i_0__15__N_2176[4]), 
         .C(phase_negation_i[1]), .Z(n1087[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam mux_188_i5_3_lut.init = 16'hcaca;
    PFUMX i21269 (.BLUT(n31), .ALUT(n62_adj_2874), .C0(index_i[5]), .Z(n23643));
    LUT4 mux_231_Mux_3_i700_3_lut_4_lut (.A(index_i[4]), .B(index_i[3]), 
         .C(n684_adj_2982), .D(n27368), .Z(n700_adj_2977)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_3_i700_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_188_i4_3_lut (.A(quarter_wave_sample_register_i[3]), .B(o_val_pipeline_i_0__15__N_2176[3]), 
         .C(phase_negation_i[1]), .Z(n1087[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam mux_188_i4_3_lut.init = 16'hcaca;
    LUT4 mux_188_i3_3_lut (.A(quarter_wave_sample_register_i[2]), .B(o_val_pipeline_i_0__15__N_2176[2]), 
         .C(phase_negation_i[1]), .Z(n1087[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam mux_188_i3_3_lut.init = 16'hcaca;
    LUT4 n652_bdd_3_lut (.A(n29939), .B(n27398), .C(index_i[3]), .Z(n25641)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n652_bdd_3_lut.init = 16'hacac;
    LUT4 mux_188_i2_3_lut (.A(quarter_wave_sample_register_i[1]), .B(o_val_pipeline_i_0__15__N_2176[1]), 
         .C(phase_negation_i[1]), .Z(n1087[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam mux_188_i2_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_11_i638_4_lut_4_lut (.A(n27089), .B(index_i[5]), .C(index_i[6]), 
         .D(n27122), .Z(n638)) /* synthesis lut_function=(A (B (C (D))+!B !(C))+!A (B ((D)+!C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_11_i638_4_lut_4_lut.init = 16'hc707;
    LUT4 mux_188_i1_3_lut (.A(quarter_wave_sample_register_i[0]), .B(o_val_pipeline_i_0__15__N_2176[0]), 
         .C(phase_negation_i[1]), .Z(n1087[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam mux_188_i1_3_lut.init = 16'hcaca;
    LUT4 i6483_2_lut (.A(phase_i[9]), .B(phase_i[10]), .Z(index_i_9__N_2125[9])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(60[14] 63[8])
    defparam i6483_2_lut.init = 16'h6666;
    LUT4 i6484_2_lut (.A(phase_i[8]), .B(phase_i[10]), .Z(index_i_9__N_2125[8])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(60[14] 63[8])
    defparam i6484_2_lut.init = 16'h6666;
    LUT4 i6485_2_lut (.A(phase_i[7]), .B(phase_i[10]), .Z(index_i_9__N_2125[7])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(60[14] 63[8])
    defparam i6485_2_lut.init = 16'h6666;
    LUT4 i6486_2_lut (.A(phase_i[6]), .B(phase_i[10]), .Z(index_i_9__N_2125[6])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(60[14] 63[8])
    defparam i6486_2_lut.init = 16'h6666;
    LUT4 i6487_2_lut (.A(phase_i[5]), .B(phase_i[10]), .Z(index_i_9__N_2125[5])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(60[14] 63[8])
    defparam i6487_2_lut.init = 16'h6666;
    LUT4 i6488_2_lut (.A(phase_i[4]), .B(phase_i[10]), .Z(index_i_9__N_2125[4])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(60[14] 63[8])
    defparam i6488_2_lut.init = 16'h6666;
    CCU2D unary_minus_10_add_3_17 (.A0(\quarter_wave_sample_register_q[15] ), 
          .B0(GND_net), .C0(GND_net), .D0(GND_net), .A1(GND_net), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n17958), .S0(o_val_pipeline_i_0__15__N_2176[15]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam unary_minus_10_add_3_17.INIT0 = 16'hf555;
    defparam unary_minus_10_add_3_17.INIT1 = 16'h0000;
    defparam unary_minus_10_add_3_17.INJECT1_0 = "NO";
    defparam unary_minus_10_add_3_17.INJECT1_1 = "NO";
    L6MUX21 i24702 (.D0(n26500), .D1(n26497), .SD(index_i[5]), .Z(n26501));
    LUT4 i6489_2_lut (.A(phase_i[3]), .B(phase_i[10]), .Z(index_i_9__N_2125[3])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(60[14] 63[8])
    defparam i6489_2_lut.init = 16'h6666;
    LUT4 i6490_2_lut (.A(phase_i[2]), .B(phase_i[10]), .Z(index_i_9__N_2125[2])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(60[14] 63[8])
    defparam i6490_2_lut.init = 16'h6666;
    PFUMX i24700 (.BLUT(n26499), .ALUT(n26498), .C0(index_i[4]), .Z(n26500));
    L6MUX21 i23345 (.D0(n24943), .D1(n24940), .SD(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2145[4]));
    LUT4 i6491_2_lut (.A(phase_i[1]), .B(phase_i[10]), .Z(index_i_9__N_2125[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(60[14] 63[8])
    defparam i6491_2_lut.init = 16'h6666;
    LUT4 i22716_3_lut (.A(n26082), .B(n21943), .C(index_i[5]), .Z(n21944)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22716_3_lut.init = 16'hcaca;
    PFUMX i23343 (.BLUT(n24942), .ALUT(n24941), .C0(index_i[8]), .Z(n24943));
    LUT4 i11519_2_lut_3_lut_4_lut (.A(n27225), .B(n27326), .C(index_i[6]), 
         .D(index_i[5]), .Z(n254)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11519_2_lut_3_lut_4_lut.init = 16'hfef0;
    LUT4 n251_bdd_3_lut_4_lut (.A(index_i[0]), .B(index_i[2]), .C(index_i[4]), 
         .D(n205), .Z(n26282)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n251_bdd_3_lut_4_lut.init = 16'h6f60;
    PFUMX i24697 (.BLUT(n26496), .ALUT(n908_adj_2910), .C0(index_i[4]), 
          .Z(n26497));
    LUT4 i23602_then_3_lut (.A(index_i[0]), .B(index_i[4]), .C(index_i[3]), 
         .Z(n27544)) /* synthesis lut_function=(A (B)+!A (B (C)+!B !(C))) */ ;
    defparam i23602_then_3_lut.init = 16'hc9c9;
    LUT4 i23602_else_3_lut (.A(index_i[2]), .B(index_i[0]), .C(index_i[4]), 
         .D(index_i[3]), .Z(n27543)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)+!C !(D)))+!A (B (C+!(D))+!B !(C)))) */ ;
    defparam i23602_else_3_lut.init = 16'h1e38;
    PFUMX i19472 (.BLUT(n21825), .ALUT(n21826), .C0(index_i[5]), .Z(n21827));
    CCU2D unary_minus_10_add_3_15 (.A0(quarter_wave_sample_register_i[13]), 
          .B0(GND_net), .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[14]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17957), .COUT(n17958), 
          .S0(o_val_pipeline_i_0__15__N_2176[13]), .S1(o_val_pipeline_i_0__15__N_2176[14]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam unary_minus_10_add_3_15.INIT0 = 16'hf555;
    defparam unary_minus_10_add_3_15.INIT1 = 16'hf555;
    defparam unary_minus_10_add_3_15.INJECT1_0 = "NO";
    defparam unary_minus_10_add_3_15.INJECT1_1 = "NO";
    PFUMX i19475 (.BLUT(n21828), .ALUT(n21829), .C0(index_i[5]), .Z(n21830));
    LUT4 i21379_3_lut_4_lut (.A(index_i[0]), .B(index_i[2]), .C(index_i[5]), 
         .D(n27518), .Z(n23753)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21379_3_lut_4_lut.init = 16'h6f60;
    PFUMX i19484 (.BLUT(n21837), .ALUT(n21838), .C0(index_i[5]), .Z(n21839));
    LUT4 n24867_bdd_3_lut_3_lut (.A(n1021), .B(index_i[8]), .C(n24867), 
         .Z(n24868)) /* synthesis lut_function=(A (B+(C))+!A !(B+!(C))) */ ;
    defparam n24867_bdd_3_lut_3_lut.init = 16'hb8b8;
    LUT4 i1_3_lut_4_lut_adj_90 (.A(n27089), .B(index_i[5]), .C(index_i[8]), 
         .D(n20104), .Z(n20537)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_3_lut_4_lut_adj_90.init = 16'hfff8;
    PFUMX i19487 (.BLUT(n21840), .ALUT(n21841), .C0(index_i[5]), .Z(n21842));
    LUT4 i15917_3_lut_3_lut (.A(index_i[0]), .B(index_i[2]), .C(index_i[3]), 
         .Z(n18103)) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i15917_3_lut_3_lut.init = 16'h6a6a;
    LUT4 i11675_2_lut_rep_694 (.A(index_i[0]), .B(index_i[1]), .Z(n27359)) /* synthesis lut_function=((B)+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11675_2_lut_rep_694.init = 16'hdddd;
    LUT4 mux_231_Mux_0_i635_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n635_adj_2833)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_0_i635_3_lut_4_lut_4_lut.init = 16'hfd0a;
    LUT4 i21266_3_lut (.A(n23636), .B(n23637), .C(index_i[8]), .Z(n23640)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21266_3_lut.init = 16'hcaca;
    LUT4 i20104_3_lut (.A(n27417), .B(n250), .C(index_i[3]), .Z(n22459)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20104_3_lut.init = 16'hcaca;
    LUT4 i20115_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n22470)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (D))+!A !(D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20115_3_lut_4_lut_4_lut_4_lut.init = 16'ha25d;
    LUT4 i22817_3_lut (.A(n23034), .B(n26058), .C(index_i[6]), .Z(n23043)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22817_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_1_i908_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n908_adj_2910)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+(D)))+!A (B (C+(D))+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_1_i908_3_lut_4_lut_4_lut_4_lut.init = 16'h332d;
    L6MUX21 i24643 (.D0(n26435), .D1(n26432), .SD(index_i[5]), .Z(n26436));
    PFUMX i23340 (.BLUT(n24939), .ALUT(n23670), .C0(index_i[8]), .Z(n24940));
    LUT4 mux_231_Mux_4_i340_3_lut_rep_695 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27360)) /* synthesis lut_function=(A (B+!(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_4_i340_3_lut_rep_695.init = 16'hdada;
    LUT4 i19905_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n22260)) /* synthesis lut_function=(!(A (B (C (D))+!B (C (D)+!C !(D)))+!A !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19905_3_lut_4_lut_4_lut.init = 16'h5aad;
    LUT4 n53_bdd_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n25679)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n53_bdd_3_lut_4_lut_4_lut.init = 16'ha5ad;
    PFUMX i24641 (.BLUT(n26434), .ALUT(n26433), .C0(index_i[4]), .Z(n26435));
    LUT4 i19548_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21903)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19548_3_lut_4_lut_4_lut.init = 16'hda5a;
    LUT4 i19969_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n22324)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C))+!A !(B (C)+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19969_3_lut_4_lut_4_lut.init = 16'h5ad3;
    LUT4 i11761_2_lut_rep_697 (.A(index_i[0]), .B(index_i[1]), .Z(n27362)) /* synthesis lut_function=(A+!(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11761_2_lut_rep_697.init = 16'hbbbb;
    LUT4 i9553_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n875)) /* synthesis lut_function=(A (C (D))+!A !(B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9553_3_lut_4_lut_4_lut_4_lut.init = 16'hb555;
    LUT4 mux_231_Mux_6_i204_3_lut_3_lut_rep_666_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27331)) /* synthesis lut_function=(!(A (C)+!A !((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_6_i204_3_lut_3_lut_rep_666_3_lut.init = 16'h5b5b;
    LUT4 mux_231_Mux_6_i205_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n205)) /* synthesis lut_function=(!(A (D)+!A !(B (D)+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_6_i205_3_lut_4_lut_4_lut_4_lut.init = 16'h54bb;
    LUT4 i19639_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n21994)) /* synthesis lut_function=(A (C+(D))+!A !(B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19639_3_lut_4_lut_4_lut.init = 16'haba5;
    LUT4 i24518_then_4_lut (.A(index_i[0]), .B(index_i[4]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n27547)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)+!C !(D))+!B (C (D)))) */ ;
    defparam i24518_then_4_lut.init = 16'hda0e;
    LUT4 i24518_else_4_lut (.A(index_i[0]), .B(index_i[4]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n27546)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C))+!A (B (C)+!B (C+(D)))) */ ;
    defparam i24518_else_4_lut.init = 16'hf178;
    LUT4 i19636_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21991)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D))+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19636_3_lut_4_lut.init = 16'hccdb;
    LUT4 mux_231_Mux_0_i364_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n364)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A ((C+!(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_0_i364_3_lut_3_lut_4_lut.init = 16'hdb55;
    LUT4 i11727_2_lut_rep_699 (.A(index_i[0]), .B(index_i[1]), .Z(n27364)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11727_2_lut_rep_699.init = 16'h2222;
    LUT4 mux_231_Mux_4_i723_3_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n723)) /* synthesis lut_function=(A ((C)+!B)+!A !(B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_4_i723_3_lut_4_lut_3_lut.init = 16'hb2b2;
    LUT4 mux_231_Mux_4_i205_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n205_adj_2983)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_4_i205_3_lut_4_lut_4_lut.init = 16'h5a2a;
    LUT4 mux_231_Mux_0_i985_3_lut_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n985)) /* synthesis lut_function=(!(A (B+!(C))+!A (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_0_i985_3_lut_3_lut_3_lut.init = 16'h2525;
    LUT4 mux_231_Mux_6_i157_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n157_adj_2984)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (D))+!A !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_6_i157_3_lut_4_lut_4_lut_4_lut.init = 16'h5d22;
    LUT4 mux_231_Mux_4_i204_3_lut_rep_701 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27366)) /* synthesis lut_function=(!(A (B+(C))+!A !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_4_i204_3_lut_rep_701.init = 16'h5252;
    LUT4 n908_bdd_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n26496)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A !(B ((D)+!C)+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n908_bdd_3_lut_3_lut_4_lut.init = 16'h552c;
    PFUMX i24637 (.BLUT(n78), .ALUT(n26431), .C0(index_i[4]), .Z(n26432));
    LUT4 i20109_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n22464)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C))+!A !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20109_3_lut_4_lut_4_lut.init = 16'h5a52;
    LUT4 i20973_3_lut (.A(n27408), .B(n27418), .C(index_i[3]), .Z(n23347)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20973_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_2_i348_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n348_adj_2985)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_2_i348_3_lut_4_lut_4_lut.init = 16'h52a5;
    PFUMX i21042 (.BLUT(n23400), .ALUT(n23401), .C0(index_i[5]), .Z(n23416));
    LUT4 i19527_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21882)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A !(B (C+!(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19527_3_lut_4_lut_4_lut.init = 16'ha52b;
    LUT4 i11676_2_lut_rep_702 (.A(index_i[0]), .B(index_i[1]), .Z(n27367)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11676_2_lut_rep_702.init = 16'h4444;
    LUT4 i7483_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n157)) /* synthesis lut_function=(!(A (C (D))+!A !(B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i7483_3_lut_4_lut_4_lut.init = 16'h4aaa;
    PFUMX i21043 (.BLUT(n23402), .ALUT(n23403), .C0(index_i[5]), .Z(n23417));
    LUT4 mux_231_Mux_0_i954_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n954)) /* synthesis lut_function=(A (D)+!A !(B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_0_i954_3_lut_4_lut_4_lut.init = 16'haf40;
    LUT4 i20972_3_lut (.A(n38), .B(n27405), .C(index_i[3]), .Z(n23346)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20972_3_lut.init = 16'hcaca;
    L6MUX21 i21044 (.D0(n23404), .D1(n23405), .SD(index_i[5]), .Z(n23418));
    LUT4 mux_231_Mux_5_i483_rep_703 (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .Z(n27368)) /* synthesis lut_function=(!(A (C)+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_5_i483_rep_703.init = 16'h4a4a;
    LUT4 i21392_3_lut_4_lut_4_lut (.A(n27207), .B(index_i[5]), .C(index_i[4]), 
         .D(n27129), .Z(n23766)) /* synthesis lut_function=(A (B+(C (D)))+!A (B+((D)+!C))) */ ;
    defparam i21392_3_lut_4_lut_4_lut.init = 16'hfdcd;
    LUT4 mux_231_Mux_6_i347_3_lut_4_lut_3_lut_rep_704 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27369)) /* synthesis lut_function=(!(A (B+!(C))+!A ((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_6_i347_3_lut_4_lut_3_lut_rep_704.init = 16'h2424;
    LUT4 i20970_3_lut (.A(n27418), .B(n204), .C(index_i[3]), .Z(n23344)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20970_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_6_i315_rep_705 (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .Z(n27370)) /* synthesis lut_function=(A (C)+!A !((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_6_i315_rep_705.init = 16'ha4a4;
    LUT4 i19978_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n22333)) /* synthesis lut_function=(!(A ((D)+!C)+!A !(B ((D)+!C)+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19978_3_lut_3_lut_4_lut.init = 16'h55a4;
    LUT4 mux_231_Mux_0_i491_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n491_adj_2829)) /* synthesis lut_function=(!(A (B (D)+!B !(C+!(D)))+!A ((C+!(D))+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_0_i491_3_lut_4_lut.init = 16'h24aa;
    LUT4 mux_231_Mux_5_i491_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n491_adj_2930)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A !(B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_5_i491_3_lut_4_lut_4_lut.init = 16'ha54a;
    LUT4 mux_231_Mux_5_i475_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n475_adj_2933)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_5_i475_3_lut_4_lut_4_lut.init = 16'hd4a5;
    LUT4 mux_231_Mux_0_i157_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n157_adj_2821)) /* synthesis lut_function=(A (B (C+!(D))+!B !(D))+!A (B (D)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_0_i157_3_lut_4_lut.init = 16'hd4aa;
    L6MUX21 i21047 (.D0(n23410), .D1(n23411), .SD(index_i[5]), .Z(n23421));
    LUT4 i20101_3_lut (.A(n27417), .B(n204), .C(index_i[3]), .Z(n22456)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20101_3_lut.init = 16'hcaca;
    LUT4 i20100_3_lut (.A(n27418), .B(n250), .C(index_i[3]), .Z(n22455)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20100_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_0_i781_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n781)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A (B (C)+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_0_i781_4_lut_4_lut_4_lut.init = 16'h0cb4;
    L6MUX21 i21048 (.D0(n23412), .D1(n23413), .SD(index_i[5]), .Z(n23422));
    LUT4 mux_231_Mux_7_i173_3_lut (.A(n27399), .B(n204), .C(index_i[3]), 
         .Z(n173_adj_2986)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_7_i173_3_lut.init = 16'hcaca;
    L6MUX21 i21049 (.D0(n23414), .D1(n23415), .SD(index_i[5]), .Z(n23423));
    LUT4 index_i_8__bdd_3_lut_then_4_lut (.A(index_i[4]), .B(index_i[6]), 
         .C(index_i[5]), .D(n27130), .Z(n27553)) /* synthesis lut_function=(!(A (B (C+(D)))+!A (B (C)))) */ ;
    defparam index_i_8__bdd_3_lut_then_4_lut.init = 16'h373f;
    LUT4 index_i_8__bdd_3_lut_else_4_lut (.A(n27169), .B(index_i[4]), .C(index_i[6]), 
         .D(index_i[5]), .Z(n27552)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;
    defparam index_i_8__bdd_3_lut_else_4_lut.init = 16'hf080;
    L6MUX21 i26270 (.D0(n29908), .D1(n29075), .SD(index_i[3]), .Z(n29079));
    PFUMX i26266 (.BLUT(n29074), .ALUT(n29073), .C0(index_i[4]), .Z(n29075));
    LUT4 i22758_3_lut (.A(n11987), .B(n892_adj_2811), .C(index_i[6]), 
         .Z(n22796)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22758_3_lut.init = 16'hcaca;
    LUT4 i11853_2_lut_rep_707 (.A(index_i[1]), .B(index_i[2]), .Z(n27372)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11853_2_lut_rep_707.init = 16'h8888;
    LUT4 i9548_2_lut_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[3]), 
         .Z(n12034)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9548_2_lut_3_lut.init = 16'h8080;
    LUT4 i19561_3_lut (.A(n29942), .B(n27366), .C(index_i[3]), .Z(n21916)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19561_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_8_i412_3_lut_4_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .Z(n15042)) /* synthesis lut_function=(A (B+!(C))+!A !((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_8_i412_3_lut_4_lut_3_lut.init = 16'h8e8e;
    LUT4 mux_231_Mux_4_i93_3_lut_4_lut_3_lut_rep_665_4_lut (.A(index_i[1]), 
         .B(index_i[2]), .C(index_i[3]), .D(index_i[0]), .Z(n27330)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_4_i93_3_lut_4_lut_3_lut_rep_665_4_lut.init = 16'h07f0;
    LUT4 i12135_2_lut_rep_541_2_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .Z(n27206)) /* synthesis lut_function=(A (B+!(C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12135_2_lut_rep_541_2_lut_3_lut.init = 16'h8f8f;
    LUT4 i11579_2_lut_rep_542_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[3]), 
         .Z(n27207)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11579_2_lut_rep_542_3_lut.init = 16'hf8f8;
    LUT4 i19560_3_lut (.A(n29927), .B(n27396), .C(index_i[3]), .Z(n21915)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19560_3_lut.init = 16'hcaca;
    LUT4 i19546_3_lut_4_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n21901)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19546_3_lut_4_lut_3_lut_4_lut.init = 16'hf80f;
    LUT4 i21265_3_lut (.A(n23634), .B(n25170), .C(index_i[7]), .Z(n23639)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21265_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_9_i412_3_lut_3_lut_4_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .Z(n412)) /* synthesis lut_function=(!(A (B (C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_9_i412_3_lut_3_lut_4_lut_3_lut.init = 16'h7e7e;
    LUT4 i19630_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .D(index_i[3]), .Z(n21985)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(D))+!A (B+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19630_3_lut_4_lut_4_lut_4_lut.init = 16'h3380;
    LUT4 i19525_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n21880)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C (D)+!C !(D)))+!A !(B (D)+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19525_3_lut_4_lut_4_lut_4_lut.init = 16'h7c03;
    LUT4 mux_231_Mux_5_i573_3_lut_3_lut (.A(index_i[0]), .B(index_i[4]), 
         .C(n572_adj_2987), .Z(n573_adj_2945)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_5_i573_3_lut_3_lut.init = 16'hd1d1;
    PFUMX i19490 (.BLUT(n21843), .ALUT(n21844), .C0(index_i[5]), .Z(n21845));
    LUT4 i21264_3_lut (.A(n23632), .B(n23633), .C(index_i[7]), .Z(n23638)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21264_3_lut.init = 16'hcaca;
    LUT4 i11998_2_lut_rep_556_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[0]), 
         .Z(n27221)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11998_2_lut_rep_556_3_lut.init = 16'h8080;
    LUT4 mux_231_Mux_9_i30_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .D(index_i[3]), .Z(n30_adj_2882)) /* synthesis lut_function=(A (B (C (D))+!B !(D))+!A !(B+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_9_i30_3_lut_4_lut_4_lut_4_lut.init = 16'h8033;
    LUT4 i11542_2_lut_rep_464_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n27129)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11542_2_lut_rep_464_3_lut_4_lut.init = 16'hf8f0;
    LUT4 mux_231_Mux_8_i491_3_lut_3_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n491_adj_2863)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_8_i491_3_lut_3_lut_3_lut_4_lut.init = 16'h7870;
    LUT4 mux_231_Mux_3_i142_3_lut_3_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .Z(n142_adj_2907)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_3_i142_3_lut_3_lut_3_lut.init = 16'h3838;
    LUT4 i11957_2_lut_rep_708 (.A(index_i[1]), .B(index_i[2]), .C(index_i[0]), 
         .Z(n27373)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11957_2_lut_rep_708.init = 16'h7070;
    PFUMX i19493 (.BLUT(n21846), .ALUT(n21847), .C0(index_i[5]), .Z(n21848));
    LUT4 i22933_3_lut (.A(n23638), .B(n23639), .C(index_i[8]), .Z(n23641)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22933_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_0_i1017_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .D(index_i[3]), .Z(n1017)) /* synthesis lut_function=(A (B (D)+!B !((D)+!C))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_0_i1017_4_lut_4_lut_4_lut.init = 16'hdd70;
    LUT4 i12474_2_lut_rep_709 (.A(index_i[2]), .B(index_i[0]), .Z(n27374)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12474_2_lut_rep_709.init = 16'heeee;
    LUT4 i1_2_lut_rep_557_3_lut (.A(index_i[2]), .B(index_i[0]), .C(index_i[1]), 
         .Z(n27222)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_2_lut_rep_557_3_lut.init = 16'hfefe;
    LUT4 mux_231_Mux_2_i173_3_lut_4_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[1]), .Z(n173)) /* synthesis lut_function=(!(A (C)+!A (B (C+!(D))+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_2_i173_3_lut_4_lut_4_lut_4_lut.init = 16'h0f1a;
    LUT4 mux_231_Mux_5_i954_3_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[1]), .Z(n954_adj_2969)) /* synthesis lut_function=(!(A (C)+!A (B+((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_5_i954_3_lut_4_lut_4_lut.init = 16'h0a1a;
    LUT4 mux_231_Mux_0_i46_3_lut_4_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[1]), .D(index_i[3]), .Z(n46_adj_2808)) /* synthesis lut_function=(A (D)+!A (B+(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_0_i46_3_lut_4_lut_4_lut_4_lut.init = 16'hfe55;
    LUT4 mux_231_Mux_8_i716_3_lut_4_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[1]), .D(index_i[3]), .Z(n716_adj_2988)) /* synthesis lut_function=(!(A (D)+!A !(B+(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_8_i716_3_lut_4_lut_4_lut_4_lut.init = 16'h55fe;
    LUT4 mux_231_Mux_9_i285_3_lut_3_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[1]), .Z(n285_adj_2885)) /* synthesis lut_function=(A (C)+!A !(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_9_i285_3_lut_3_lut_4_lut_4_lut.init = 16'ha0a1;
    LUT4 mux_231_Mux_2_i763_4_lut_4_lut (.A(index_i[0]), .B(n12034), .C(index_i[4]), 
         .D(n157_adj_2984), .Z(n763_adj_2869)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_2_i763_4_lut_4_lut.init = 16'hdfd0;
    LUT4 i11529_2_lut_rep_463_3_lut_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[1]), .Z(n27128)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11529_2_lut_rep_463_3_lut_4_lut.init = 16'hf0e0;
    LUT4 n172_bdd_2_lut_3_lut_3_lut_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[1]), .D(index_i[3]), .Z(n26080)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n172_bdd_2_lut_3_lut_3_lut_4_lut.init = 16'h00fe;
    LUT4 mux_231_Mux_2_i731_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n731_adj_2966)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_2_i731_3_lut_4_lut_4_lut.init = 16'h6cc6;
    LUT4 mux_231_Mux_7_i156_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n204)) /* synthesis lut_function=(!(A (B)+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_7_i156_3_lut_3_lut.init = 16'h6363;
    LUT4 mux_231_Mux_5_i356_3_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n325)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_5_i356_3_lut_4_lut_3_lut.init = 16'h6d6d;
    LUT4 mux_231_Mux_1_i882_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n882)) /* synthesis lut_function=(A ((C)+!B)+!A !((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_1_i882_3_lut_3_lut.init = 16'ha6a6;
    LUT4 mux_231_Mux_4_i14_3_lut_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n14)) /* synthesis lut_function=(!(A (B+(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_4_i14_3_lut_3_lut_3_lut.init = 16'h5656;
    LUT4 i22158_3_lut (.A(n109), .B(n124_adj_2849), .C(index_i[4]), .Z(n21829)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22158_3_lut.init = 16'hcaca;
    LUT4 i9668_3_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[4]), 
         .Z(n12157)) /* synthesis lut_function=(!(A (B)+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9668_3_lut_4_lut_3_lut.init = 16'h6262;
    LUT4 i9510_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n526)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+(D)))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9510_3_lut_4_lut_4_lut.init = 16'h666c;
    L6MUX21 i21073 (.D0(n23431), .D1(n23432), .SD(index_i[5]), .Z(n23447));
    L6MUX21 i21074 (.D0(n23433), .D1(n23434), .SD(index_i[5]), .Z(n23448));
    L6MUX21 i21075 (.D0(n23435), .D1(n23436), .SD(index_i[5]), .Z(n23449));
    L6MUX21 i21076 (.D0(n23437), .D1(n23438), .SD(index_i[5]), .Z(n23450));
    LUT4 i9524_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(n27318), .D(index_i[4]), .Z(n221_adj_2989)) /* synthesis lut_function=(!(A (B)+!A (B (C+(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9524_3_lut_4_lut_4_lut_4_lut.init = 16'h3336;
    L6MUX21 i21077 (.D0(n23439), .D1(n23440), .SD(index_i[5]), .Z(n23451));
    LUT4 n21650_bdd_3_lut_23969 (.A(n27368), .B(n27400), .C(index_i[3]), 
         .Z(n25681)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n21650_bdd_3_lut_23969.init = 16'hcaca;
    L6MUX21 i21078 (.D0(n23441), .D1(n23442), .SD(index_i[5]), .Z(n23452));
    L6MUX21 i21079 (.D0(n23443), .D1(n23444), .SD(index_i[5]), .Z(n23453));
    L6MUX21 i21080 (.D0(n23445), .D1(n23446), .SD(index_i[5]), .Z(n23454));
    PFUMX i19502 (.BLUT(n21855), .ALUT(n21856), .C0(index_i[5]), .Z(n21857));
    PFUMX i23604 (.BLUT(n25285), .ALUT(n25281), .C0(index_i[6]), .Z(n25286));
    PFUMX i19505 (.BLUT(n21858), .ALUT(n21859), .C0(index_i[5]), .Z(n21860));
    LUT4 mux_231_Mux_3_i507_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[4]), .D(n491), .Z(n507_adj_2976)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_3_i507_3_lut_4_lut.init = 16'h6f60;
    PFUMX i19508 (.BLUT(n21861), .ALUT(n21862), .C0(index_i[5]), .Z(n21863));
    LUT4 mux_231_Mux_6_i660_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n108)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_6_i660_3_lut_3_lut.init = 16'hc6c6;
    LUT4 n428_bdd_3_lut_24941_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n26192)) /* synthesis lut_function=(!(A (B)+!A !(B (C+(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n428_bdd_3_lut_24941_4_lut_4_lut_4_lut.init = 16'h6663;
    LUT4 i9627_3_lut_4_lut_4_lut (.A(index_i[0]), .B(n14), .C(index_i[4]), 
         .D(n27325), .Z(n12113)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B ((D)+!C)+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9627_3_lut_4_lut_4_lut.init = 16'h5c0c;
    LUT4 i9542_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[4]), .Z(n444_adj_2909)) /* synthesis lut_function=(!(A (B)+!A !(B (C (D))+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9542_3_lut_4_lut_4_lut_4_lut.init = 16'h6333;
    LUT4 mux_231_Mux_5_i828_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[4]), .D(n27336), .Z(n828_adj_2949)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_5_i828_4_lut_4_lut.init = 16'hc66c;
    LUT4 mux_231_Mux_0_i747_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n747_adj_2838)) /* synthesis lut_function=(!(A (B+!(C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_0_i747_3_lut_4_lut_4_lut_4_lut.init = 16'h6556;
    LUT4 i19518_3_lut_4_lut_4_lut (.A(index_i[0]), .B(n27379), .C(index_i[3]), 
         .D(n27372), .Z(n21873)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19518_3_lut_4_lut_4_lut.init = 16'hcfc5;
    LUT4 mux_231_Mux_5_i683_3_lut_4_lut_3_lut_rep_710 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27375)) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_5_i683_3_lut_4_lut_3_lut_rep_710.init = 16'h6b6b;
    LUT4 i20871_3_lut (.A(n23237), .B(n23238), .C(index_i[7]), .Z(n23245)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20871_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_5_i262_rep_711 (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .Z(n27376)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_5_i262_rep_711.init = 16'h6464;
    LUT4 mux_231_Mux_6_i141_3_lut_4_lut_3_lut_rep_712 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27377)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_6_i141_3_lut_4_lut_3_lut_rep_712.init = 16'hd6d6;
    LUT4 mux_231_Mux_5_i754_3_lut_4_lut_3_lut_rep_713 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27378)) /* synthesis lut_function=(!(A (B)+!A ((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_5_i754_3_lut_4_lut_3_lut_rep_713.init = 16'h2626;
    LUT4 mux_231_Mux_4_i70_3_lut_3_lut_rep_714 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27379)) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_4_i70_3_lut_3_lut_rep_714.init = 16'h6a6a;
    LUT4 mux_231_Mux_2_i491_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n491_adj_2990)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A !(B (C)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_2_i491_3_lut_4_lut_4_lut.init = 16'h6a5a;
    LUT4 i19617_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21972)) /* synthesis lut_function=(!(A (B)+!A (B (C+(D))+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19617_3_lut_3_lut_4_lut.init = 16'h3326;
    LUT4 i19519_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21874)) /* synthesis lut_function=(A (B (C)+!B !(C (D)+!C !(D)))+!A (B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19519_3_lut_4_lut_4_lut.init = 16'hd6a5;
    LUT4 n21650_bdd_3_lut_24026_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n25682)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C))+!A !(B (C+!(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n21650_bdd_3_lut_24026_4_lut_4_lut.init = 16'h5ad6;
    PFUMX mux_231_Mux_7_i190 (.BLUT(n22457), .ALUT(n173_adj_2986), .C0(index_i[5]), 
          .Z(n190)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 i19542_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21897)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19542_3_lut_4_lut.init = 16'h64cc;
    LUT4 mux_231_Mux_5_i460_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n460_adj_2932)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A !(B (C)+!B !(C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_5_i460_3_lut_4_lut_4_lut.init = 16'h6b5a;
    LUT4 mux_231_Mux_3_i94_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[4]), .D(n93_adj_2905), .Z(n94_adj_2973)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_3_i94_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_231_Mux_3_i62_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[4]), .D(n812_adj_2890), .Z(n62_adj_2981)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_3_i62_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_231_Mux_3_i796_3_lut_3_lut (.A(index_i[4]), .B(n412_adj_2844), 
         .C(index_i[2]), .Z(n796_adj_2979)) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam mux_231_Mux_3_i796_3_lut_3_lut.init = 16'he4e4;
    LUT4 mux_231_Mux_4_i142_3_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[3]), 
         .C(index_i[2]), .Z(n142_adj_2799)) /* synthesis lut_function=(A (B (C))+!A !(B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_4_i142_3_lut_4_lut_3_lut.init = 16'h9595;
    LUT4 i20660_4_lut_4_lut (.A(index_i[4]), .B(index_i[5]), .C(n27493), 
         .D(n908), .Z(n23034)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam i20660_4_lut_4_lut.init = 16'hd1c0;
    LUT4 i9496_4_lut_4_lut (.A(index_i[4]), .B(n22736), .C(n27515), .D(n27412), 
         .Z(n11982)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam i9496_4_lut_4_lut.init = 16'hf4b0;
    LUT4 n25744_bdd_3_lut (.A(n25744), .B(n25741), .C(index_i[4]), .Z(n21806)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n25744_bdd_3_lut.init = 16'hcaca;
    PFUMX mux_231_Mux_8_i764 (.BLUT(n716_adj_2988), .ALUT(n732_adj_2840), 
          .C0(n22640), .Z(n764)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    PFUMX i24532 (.BLUT(n26282), .ALUT(n26281), .C0(index_i[5]), .Z(n26283));
    PFUMX mux_231_Mux_8_i574 (.BLUT(n542), .ALUT(n11985), .C0(index_i[5]), 
          .Z(n574_adj_2831)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 i11598_4_lut (.A(n27204), .B(index_i[7]), .C(n892), .D(index_i[6]), 
         .Z(n1021)) /* synthesis lut_function=(A (B+(C (D)))+!A (B+(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11598_4_lut.init = 16'hfcdd;
    CCU2D unary_minus_10_add_3_13 (.A0(quarter_wave_sample_register_i[11]), 
          .B0(GND_net), .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[12]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17956), .COUT(n17957), 
          .S0(o_val_pipeline_i_0__15__N_2176[11]), .S1(o_val_pipeline_i_0__15__N_2176[12]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam unary_minus_10_add_3_13.INIT0 = 16'hf555;
    defparam unary_minus_10_add_3_13.INIT1 = 16'hf555;
    defparam unary_minus_10_add_3_13.INJECT1_0 = "NO";
    defparam unary_minus_10_add_3_13.INJECT1_1 = "NO";
    CCU2D unary_minus_10_add_3_11 (.A0(quarter_wave_sample_register_i[9]), 
          .B0(GND_net), .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[10]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17955), .COUT(n17956), 
          .S0(o_val_pipeline_i_0__15__N_2176[9]), .S1(o_val_pipeline_i_0__15__N_2176[10]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam unary_minus_10_add_3_11.INIT0 = 16'hf555;
    defparam unary_minus_10_add_3_11.INIT1 = 16'hf555;
    defparam unary_minus_10_add_3_11.INJECT1_0 = "NO";
    defparam unary_minus_10_add_3_11.INJECT1_1 = "NO";
    LUT4 i20971_3_lut_3_lut (.A(n27416), .B(index_i[3]), .C(n29957), .Z(n23345)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam i20971_3_lut_3_lut.init = 16'h7474;
    LUT4 i20864_3_lut (.A(n23223), .B(n26194), .C(index_i[6]), .Z(n23238)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20864_3_lut.init = 16'hcaca;
    LUT4 i19537_3_lut_3_lut (.A(n27416), .B(index_i[3]), .C(n38), .Z(n21892)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam i19537_3_lut_3_lut.init = 16'h7474;
    LUT4 i11544_4_lut (.A(n15304), .B(index_i[8]), .C(n765), .D(index_i[7]), 
         .Z(n1022)) /* synthesis lut_function=(A (B+(C (D)))+!A (B+(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11544_4_lut.init = 16'hfcdd;
    LUT4 mux_231_Mux_7_i379_3_lut_3_lut (.A(n27416), .B(index_i[3]), .C(n27408), 
         .Z(n379_adj_2846)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam mux_231_Mux_7_i379_3_lut_3_lut.init = 16'h7474;
    LUT4 mux_231_Mux_4_i668_3_lut_3_lut (.A(n27416), .B(index_i[3]), .C(n29957), 
         .Z(n668_adj_2918)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;
    defparam mux_231_Mux_4_i668_3_lut_3_lut.init = 16'hd1d1;
    PFUMX i20847 (.BLUT(n12114), .ALUT(n62_adj_2991), .C0(index_i[5]), 
          .Z(n23221));
    CCU2D unary_minus_10_add_3_9 (.A0(quarter_wave_sample_register_i[7]), 
          .B0(GND_net), .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[8]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17954), .COUT(n17955), 
          .S0(o_val_pipeline_i_0__15__N_2176[7]), .S1(o_val_pipeline_i_0__15__N_2176[8]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam unary_minus_10_add_3_9.INIT0 = 16'hf555;
    defparam unary_minus_10_add_3_9.INIT1 = 16'hf555;
    defparam unary_minus_10_add_3_9.INJECT1_0 = "NO";
    defparam unary_minus_10_add_3_9.INJECT1_1 = "NO";
    LUT4 mux_231_Mux_2_i507_3_lut_3_lut (.A(index_i[0]), .B(index_i[4]), 
         .C(n491_adj_2990), .Z(n507)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_2_i507_3_lut_3_lut.init = 16'h7474;
    LUT4 mux_231_Mux_6_i924_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[4]), .D(n762_adj_2957), .Z(n924)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_6_i924_3_lut_4_lut.init = 16'h6f60;
    LUT4 i20873_3_lut (.A(n23241), .B(n23242), .C(index_i[7]), .Z(n23247)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20873_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_2_i859_3_lut_4_lut_4_lut (.A(index_i[0]), .B(n27370), 
         .C(index_i[3]), .D(n27325), .Z(n859)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B ((D)+!C)+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_2_i859_3_lut_4_lut_4_lut.init = 16'h5c0c;
    LUT4 mux_231_Mux_7_i364_3_lut_3_lut (.A(n27416), .B(index_i[3]), .C(n27417), 
         .Z(n364_adj_2845)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;
    defparam mux_231_Mux_7_i364_3_lut_3_lut.init = 16'hd1d1;
    LUT4 i22236_3_lut (.A(n21915), .B(n21916), .C(index_i[4]), .Z(n21917)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22236_3_lut.init = 16'hcaca;
    LUT4 index_i_0__bdd_4_lut_25223 (.A(index_i[0]), .B(index_i[3]), .C(index_i[1]), 
         .D(index_i[2]), .Z(n27564)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C))+!A (B (C (D)+!C !(D))+!B !(C+!(D))))) */ ;
    defparam index_i_0__bdd_4_lut_25223.init = 16'h16d3;
    LUT4 mux_231_Mux_4_i221_3_lut_3_lut (.A(index_i[0]), .B(index_i[4]), 
         .C(n205_adj_2983), .Z(n221_adj_2953)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_4_i221_3_lut_3_lut.init = 16'h7474;
    LUT4 i20867_3_lut (.A(n26207), .B(n23230), .C(index_i[6]), .Z(n23241)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20867_3_lut.init = 16'hcaca;
    CCU2D unary_minus_10_add_3_7 (.A0(quarter_wave_sample_register_i[5]), 
          .B0(GND_net), .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[6]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17953), .COUT(n17954), 
          .S0(o_val_pipeline_i_0__15__N_2176[5]), .S1(o_val_pipeline_i_0__15__N_2176[6]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam unary_minus_10_add_3_7.INIT0 = 16'hf555;
    defparam unary_minus_10_add_3_7.INIT1 = 16'hf555;
    defparam unary_minus_10_add_3_7.INJECT1_0 = "NO";
    defparam unary_minus_10_add_3_7.INJECT1_1 = "NO";
    LUT4 i20668_3_lut (.A(n26047), .B(n23033), .C(index_i[6]), .Z(n23042)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20668_3_lut.init = 16'hcaca;
    LUT4 i19575_3_lut_4_lut_4_lut (.A(index_i[0]), .B(n27375), .C(index_i[3]), 
         .D(n27325), .Z(n21930)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19575_3_lut_4_lut_4_lut.init = 16'hc5c0;
    CCU2D unary_minus_10_add_3_5 (.A0(quarter_wave_sample_register_i[3]), 
          .B0(GND_net), .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[4]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17952), .COUT(n17953), 
          .S0(o_val_pipeline_i_0__15__N_2176[3]), .S1(o_val_pipeline_i_0__15__N_2176[4]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam unary_minus_10_add_3_5.INIT0 = 16'hf555;
    defparam unary_minus_10_add_3_5.INIT1 = 16'hf555;
    defparam unary_minus_10_add_3_5.INJECT1_0 = "NO";
    defparam unary_minus_10_add_3_5.INJECT1_1 = "NO";
    LUT4 mux_231_Mux_2_i349_3_lut_3_lut (.A(index_i[0]), .B(index_i[4]), 
         .C(n348_adj_2985), .Z(n349_adj_2861)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_2_i349_3_lut_3_lut.init = 16'hd1d1;
    LUT4 mux_231_Mux_1_i890_4_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[3]), 
         .C(n204), .D(index_i[4]), .Z(n890_adj_2980)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (D))+!A !((C+(D))+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_1_i890_4_lut_4_lut_4_lut_4_lut.init = 16'h55f3;
    L6MUX21 i24485 (.D0(n26206), .D1(n26203), .SD(index_i[5]), .Z(n26207));
    PFUMX i24483 (.BLUT(n26205), .ALUT(n26204), .C0(index_i[4]), .Z(n26206));
    LUT4 i21086_3_lut (.A(n23457), .B(n23458), .C(index_i[7]), .Z(n23460)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21086_3_lut.init = 16'hcaca;
    LUT4 i21085_3_lut (.A(n23455), .B(n23456), .C(index_i[7]), .Z(n23459)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21085_3_lut.init = 16'hcaca;
    LUT4 i12138_2_lut_3_lut_3_lut (.A(index_i[0]), .B(index_i[2]), .C(index_i[3]), 
         .Z(n14736)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12138_2_lut_3_lut_3_lut.init = 16'h4040;
    CCU2D unary_minus_10_add_3_3 (.A0(quarter_wave_sample_register_i[1]), 
          .B0(GND_net), .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[2]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17951), .COUT(n17952), 
          .S0(o_val_pipeline_i_0__15__N_2176[1]), .S1(o_val_pipeline_i_0__15__N_2176[2]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam unary_minus_10_add_3_3.INIT0 = 16'hf555;
    defparam unary_minus_10_add_3_3.INIT1 = 16'hf555;
    defparam unary_minus_10_add_3_3.INJECT1_0 = "NO";
    defparam unary_minus_10_add_3_3.INJECT1_1 = "NO";
    LUT4 i19491_3_lut_4_lut_4_lut (.A(n27221), .B(index_i[4]), .C(index_i[3]), 
         .D(n27225), .Z(n21846)) /* synthesis lut_function=(A (B (C)+!B !(C+!(D)))+!A (B (C)+!B (C+(D)))) */ ;
    defparam i19491_3_lut_4_lut_4_lut.init = 16'hd3d0;
    PFUMX i24480 (.BLUT(n26202), .ALUT(n27101), .C0(index_i[4]), .Z(n26203));
    L6MUX21 i24470 (.D0(n26193), .D1(n26191), .SD(index_i[4]), .Z(n26194));
    PFUMX i24468 (.BLUT(n27103), .ALUT(n26192), .C0(index_i[5]), .Z(n26193));
    LUT4 i22981_2_lut_rep_730 (.A(index_i[0]), .B(index_i[1]), .Z(n27395)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i22981_2_lut_rep_730.init = 16'h9999;
    LUT4 i9512_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n541_adj_2896)) /* synthesis lut_function=(A (B (C (D))+!B !(C (D)))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9512_3_lut_4_lut_4_lut_4_lut.init = 16'h9333;
    LUT4 mux_231_Mux_6_i573_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[4]), .D(n572_adj_2992), .Z(n573_adj_2978)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_6_i573_3_lut_4_lut.init = 16'hf909;
    LUT4 i12021_2_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n844)) /* synthesis lut_function=(A (B+!(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12021_2_lut_3_lut_4_lut.init = 16'h9ff9;
    PFUMX i24466 (.BLUT(n26190), .ALUT(n26189), .C0(index_i[5]), .Z(n26191));
    LUT4 i9540_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(n27318), .D(index_i[4]), .Z(n189_adj_2993)) /* synthesis lut_function=(A (B (C (D)))+!A !(B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9540_3_lut_4_lut_4_lut_4_lut.init = 16'h9555;
    LUT4 mux_231_Mux_5_i572_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n572_adj_2987)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A !(B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_5_i572_3_lut_4_lut_4_lut.init = 16'ha9a5;
    LUT4 i9528_3_lut_4_lut_4_lut (.A(index_i[0]), .B(n27379), .C(index_i[4]), 
         .D(index_i[3]), .Z(n605_adj_2946)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A !(B+(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9528_3_lut_4_lut_4_lut.init = 16'h555c;
    LUT4 i21055_3_lut (.A(n23426), .B(n23427), .C(index_i[7]), .Z(n23429)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21055_3_lut.init = 16'hcaca;
    LUT4 i19941_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n22296)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !(B (C+!(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19941_3_lut_4_lut_4_lut.init = 16'ha5a9;
    LUT4 mux_231_Mux_1_i93_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n93_adj_2921)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C+(D)))+!A !(B (C (D)+!C !(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_1_i93_3_lut_4_lut_4_lut_4_lut.init = 16'h955a;
    LUT4 i15935_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n18121)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i15935_3_lut_4_lut_4_lut_4_lut.init = 16'h3999;
    LUT4 mux_231_Mux_4_i187_3_lut_3_lut_rep_668_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27333)) /* synthesis lut_function=(A (B (C))+!A !(B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_4_i187_3_lut_3_lut_rep_668_3_lut.init = 16'h9595;
    LUT4 i12007_2_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n668)) /* synthesis lut_function=(!(A ((D)+!B)+!A (B ((D)+!C)+!B (C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12007_2_lut_4_lut_4_lut_4_lut.init = 16'h00c9;
    LUT4 i21054_3_lut (.A(n23424), .B(n23425), .C(index_i[7]), .Z(n23428)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21054_3_lut.init = 16'hcaca;
    LUT4 i15934_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n18120)) /* synthesis lut_function=(A (B)+!A !(B (C (D))+!B !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i15934_3_lut_4_lut_4_lut.init = 16'h9ccc;
    LUT4 mux_231_Mux_5_i109_3_lut_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .Z(n109_adj_2937)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_5_i109_3_lut_3_lut_3_lut.init = 16'h3939;
    LUT4 mux_231_Mux_6_i498_3_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n404)) /* synthesis lut_function=(A (B+!(C))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_6_i498_3_lut_4_lut_3_lut.init = 16'h9b9b;
    LUT4 mux_231_Mux_6_i356_3_lut_4_lut_3_lut_rep_731 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27396)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_6_i356_3_lut_4_lut_3_lut_rep_731.init = 16'h4949;
    LUT4 mux_231_Mux_4_i262_3_lut_3_lut_rep_732 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27397)) /* synthesis lut_function=(A (B+(C))+!A !(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_4_i262_3_lut_3_lut_rep_732.init = 16'ha9a9;
    LUT4 i19398_3_lut (.A(n25185), .B(n21776), .C(index_i[8]), .Z(n21753)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19398_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_3_i340_3_lut_3_lut_3_lut_rep_733 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27398)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_3_i340_3_lut_3_lut_3_lut_rep_733.init = 16'h9393;
    LUT4 n18302_bdd_4_lut_then_4_lut (.A(index_i[3]), .B(index_i[4]), .C(index_i[1]), 
         .D(index_i[2]), .Z(n27572)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B+(C (D)+!C !(D)))) */ ;
    defparam n18302_bdd_4_lut_then_4_lut.init = 16'hf44f;
    LUT4 n18302_bdd_4_lut_else_4_lut (.A(index_i[3]), .B(index_i[4]), .C(index_i[1]), 
         .D(index_i[2]), .Z(n27571)) /* synthesis lut_function=(!(A (B (D)+!B ((D)+!C))+!A !(B+!((D)+!C)))) */ ;
    defparam n18302_bdd_4_lut_else_4_lut.init = 16'h44fc;
    LUT4 mux_231_Mux_7_i77_3_lut_3_lut_rep_734 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27399)) /* synthesis lut_function=(A (B)+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_7_i77_3_lut_3_lut_rep_734.init = 16'h9c9c;
    LUT4 mux_231_Mux_6_i92_3_lut_4_lut_3_lut_rep_735 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27400)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_6_i92_3_lut_4_lut_3_lut_rep_735.init = 16'h6969;
    LUT4 mux_231_Mux_6_i250_3_lut_4_lut_3_lut_rep_736 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27401)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_6_i250_3_lut_4_lut_3_lut_rep_736.init = 16'h9696;
    LUT4 mux_231_Mux_3_i723_3_lut_4_lut_3_lut_rep_737 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27402)) /* synthesis lut_function=(A (B (C))+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_3_i723_3_lut_4_lut_3_lut_rep_737.init = 16'h9494;
    LUT4 mux_231_Mux_6_i564_3_lut_4_lut_3_lut_rep_738 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27403)) /* synthesis lut_function=(A (B)+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_6_i564_3_lut_4_lut_3_lut_rep_738.init = 16'hd9d9;
    LUT4 mux_231_Mux_6_i505_3_lut_rep_739 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27404)) /* synthesis lut_function=(A (B)+!A (B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_6_i505_3_lut_rep_739.init = 16'hc9c9;
    LUT4 mux_231_Mux_7_i116_3_lut_3_lut_rep_740 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27405)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_7_i116_3_lut_3_lut_rep_740.init = 16'h3939;
    LUT4 mux_231_Mux_1_i62_3_lut_4_lut (.A(index_i[0]), .B(index_i[3]), 
         .C(index_i[2]), .D(index_i[4]), .Z(n62_adj_2991)) /* synthesis lut_function=(A (B (D)+!B ((D)+!C))+!A !(B (D)+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_1_i62_3_lut_4_lut.init = 16'haa56;
    LUT4 mux_231_Mux_6_i389_3_lut_4_lut_3_lut_rep_741 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27406)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_6_i389_3_lut_4_lut_3_lut_rep_741.init = 16'h9292;
    LUT4 i19626_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21981)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C))+!A !(B ((D)+!C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19626_3_lut_4_lut_4_lut.init = 16'h925a;
    LUT4 mux_231_Mux_0_i812_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n812_adj_2847)) /* synthesis lut_function=(A (B (C+(D))+!B !(C))+!A (B (D)+!B !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_0_i812_3_lut_4_lut_4_lut_4_lut.init = 16'hcf92;
    LUT4 mux_231_Mux_2_i604_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n604_adj_2968)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)+!C !(D)))+!A (B (D)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_2_i604_3_lut_4_lut_4_lut_4_lut.init = 16'h39cf;
    LUT4 i20014_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n22369)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C+(D)))+!A (B (C)+!B !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20014_3_lut_4_lut_4_lut.init = 16'hc95a;
    PFUMX i20126 (.BLUT(n22479), .ALUT(n22480), .C0(index_i[4]), .Z(n22481));
    LUT4 mux_231_Mux_3_i444_3_lut_4_lut (.A(index_i[0]), .B(index_i[3]), 
         .C(n27372), .D(index_i[4]), .Z(n444_adj_2975)) /* synthesis lut_function=(!(A (B (D)+!B (C (D)))+!A !(B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_3_i444_3_lut_4_lut.init = 16'h46aa;
    LUT4 mux_231_Mux_6_i572_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n572_adj_2992)) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_6_i572_3_lut_4_lut.init = 16'hccd9;
    LUT4 n572_bdd_3_lut_24900_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n26202)) /* synthesis lut_function=(A (B (C+(D)))+!A (B ((D)+!C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n572_bdd_3_lut_24900_4_lut.init = 16'hcc94;
    LUT4 mux_231_Mux_4_i252_4_lut_4_lut (.A(index_i[0]), .B(index_i[3]), 
         .C(n27325), .D(index_i[4]), .Z(n252_adj_2954)) /* synthesis lut_function=(!(A (B (D)+!B !(D))+!A !(B ((D)+!C)+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_4_i252_4_lut_4_lut.init = 16'h669d;
    LUT4 mux_231_Mux_2_i653_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n653_adj_2967)) /* synthesis lut_function=(A (B (C+!(D))+!B !(D))+!A !(B (C+!(D))+!B !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_2_i653_3_lut_4_lut.init = 16'h94aa;
    LUT4 mux_231_Mux_3_i684_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[4]), .Z(n684_adj_2982)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A !(B ((D)+!C)+!B (C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_3_i684_3_lut_3_lut_4_lut.init = 16'h5594;
    LUT4 n715_bdd_3_lut_24482_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n26204)) /* synthesis lut_function=(A (B (C+(D))+!B ((D)+!C))+!A !(B (C+(D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n715_bdd_3_lut_24482_4_lut.init = 16'haa96;
    LUT4 mux_231_Mux_0_i142_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n142_adj_2820)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C))+!A !(B (C (D)+!C !(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_0_i142_3_lut_4_lut_4_lut.init = 16'ha569;
    LUT4 mux_231_Mux_3_i859_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n859_adj_2951)) /* synthesis lut_function=(!(A (B (D)+!B !(D))+!A (B (C+(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_3_i859_3_lut_3_lut_4_lut.init = 16'h339c;
    L6MUX21 i23529 (.D0(n25184), .D1(n27063), .SD(index_i[6]), .Z(n25185));
    LUT4 i20675_3_lut (.A(n23046), .B(n23047), .C(index_i[8]), .Z(n23049)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20675_3_lut.init = 16'hcaca;
    LUT4 i19986_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n22341)) /* synthesis lut_function=(A (B (C)+!B (C (D)+!C !(D)))+!A !(B (C+!(D))+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19986_3_lut_4_lut_4_lut.init = 16'ha593;
    LUT4 i19509_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21864)) /* synthesis lut_function=(A (B (C (D))+!B !(C (D)))+!A !(B (D)+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19509_3_lut_4_lut_4_lut.init = 16'h9366;
    PFUMX i23527 (.BLUT(n25183), .ALUT(n27083), .C0(index_i[7]), .Z(n25184));
    LUT4 i19569_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21924)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A !(B (D)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19569_3_lut_3_lut_4_lut.init = 16'ha955;
    LUT4 mux_231_Mux_3_i397_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n397_adj_2903)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !(B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_3_i397_3_lut_4_lut_4_lut.init = 16'ha95a;
    PFUMX i20132 (.BLUT(n22485), .ALUT(n22486), .C0(index_i[4]), .Z(n22487));
    LUT4 i19914_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n22269)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (D))+!A !(B (C (D))+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19914_3_lut_3_lut_4_lut.init = 16'h4933;
    LUT4 i11760_2_lut_rep_742 (.A(index_i[0]), .B(index_i[1]), .Z(n27407)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11760_2_lut_rep_742.init = 16'h8888;
    LUT4 i19554_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n21909)) /* synthesis lut_function=(!(A (B (D)+!B !(D))+!A (B ((D)+!C)+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19554_3_lut_4_lut_4_lut_4_lut.init = 16'h33c8;
    LUT4 i19624_3_lut_4_lut_4_lut (.A(index_i[2]), .B(n250), .C(index_i[3]), 
         .D(n27413), .Z(n21979)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19624_3_lut_4_lut_4_lut.init = 16'hc5c0;
    LUT4 i23048_2_lut_rep_481_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n27146)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i23048_2_lut_rep_481_3_lut_4_lut.init = 16'h0007;
    LUT4 i20963_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n23337)) /* synthesis lut_function=(A (B (D)+!B !(C (D)+!C !(D)))+!A !(B (C+!(D))+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20963_3_lut_4_lut_4_lut.init = 16'h8f30;
    LUT4 n300_bdd_3_lut_24313_4_lut_4_lut (.A(index_i[2]), .B(n77), .C(index_i[3]), 
         .D(n27413), .Z(n26044)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B ((D)+!C)+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n300_bdd_3_lut_24313_4_lut_4_lut.init = 16'h5c0c;
    LUT4 i19933_3_lut_4_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n22288)) /* synthesis lut_function=(!(A (B (D)+!B !((D)+!C))+!A (B (C+(D))+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19933_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'h338f;
    CCU2D unary_minus_10_add_3_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(quarter_wave_sample_register_i[0]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .COUT(n17951), .S1(o_val_pipeline_i_0__15__N_2176[0]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam unary_minus_10_add_3_1.INIT0 = 16'hF000;
    defparam unary_minus_10_add_3_1.INIT1 = 16'h0aaa;
    defparam unary_minus_10_add_3_1.INJECT1_0 = "NO";
    defparam unary_minus_10_add_3_1.INJECT1_1 = "NO";
    LUT4 i21404_3_lut (.A(n23773), .B(n23774), .C(index_i[7]), .Z(n23778)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21404_3_lut.init = 16'hcaca;
    LUT4 i20674_3_lut (.A(n23044), .B(n23045), .C(index_i[8]), .Z(n23048)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20674_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_4_i491_3_lut_4_lut_4_lut (.A(index_i[2]), .B(n27417), 
         .C(index_i[3]), .D(n27407), .Z(n491_adj_2950)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_4_i491_3_lut_4_lut_4_lut.init = 16'hfc5c;
    LUT4 i11610_2_lut_rep_438_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n27103)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11610_2_lut_rep_438_3_lut_4_lut.init = 16'hf080;
    L6MUX21 i23514 (.D0(n25169), .D1(n25167), .SD(index_i[6]), .Z(n25170));
    PFUMX i19571 (.BLUT(n21924), .ALUT(n21925), .C0(index_i[4]), .Z(n21926));
    PFUMX i23512 (.BLUT(n924_adj_2994), .ALUT(n25168), .C0(index_i[5]), 
          .Z(n25169));
    LUT4 index_i_0__bdd_4_lut_25332 (.A(index_i[0]), .B(index_i[3]), .C(index_i[1]), 
         .D(index_i[2]), .Z(n27577)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C (D)))+!A !(B (C+!(D))+!B !(C+(D))))) */ ;
    defparam index_i_0__bdd_4_lut_25332.init = 16'h4ae7;
    PFUMX i25165 (.BLUT(n27491), .ALUT(n27492), .C0(index_i[0]), .Z(n27493));
    LUT4 mux_231_Mux_7_i747_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n747_adj_2956)) /* synthesis lut_function=(A (B (C)+!B (C (D)+!C !(D)))+!A (B (C+!(D))+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_7_i747_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hf0c7;
    LUT4 i19558_3_lut (.A(n29957), .B(n27415), .C(index_i[3]), .Z(n21913)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19558_3_lut.init = 16'hcaca;
    LUT4 i20425_3_lut (.A(n22792), .B(n22793), .C(index_i[7]), .Z(n22799)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20425_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_7_i506_3_lut_4_lut_4_lut (.A(index_i[2]), .B(n27417), 
         .C(index_i[3]), .D(n27413), .Z(n506_adj_2959)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B ((D)+!C)+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_7_i506_3_lut_4_lut_4_lut.init = 16'h5c0c;
    LUT4 mux_231_Mux_3_i1002_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n20184)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (D))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_3_i1002_3_lut_3_lut_4_lut.init = 16'hf708;
    LUT4 mux_231_Mux_8_i635_3_lut_4_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n635_adj_2810)) /* synthesis lut_function=(!(A (B (C (D))+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_8_i635_3_lut_4_lut_3_lut_4_lut.init = 16'h0ff8;
    LUT4 n10642_bdd_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n26434)) /* synthesis lut_function=(A (B (C+!(D))+!B ((D)+!C))+!A (B (C (D)+!C !(D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n10642_bdd_3_lut_4_lut_4_lut_4_lut.init = 16'hf38f;
    LUT4 mux_231_Mux_7_i526_3_lut_4_lut_4_lut_3_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n526_adj_2970)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(D))+!A !(D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_7_i526_3_lut_4_lut_4_lut_3_lut_4_lut.init = 16'h887f;
    LUT4 i20424_3_lut (.A(n22790), .B(n22791), .C(index_i[7]), .Z(n22798)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20424_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_8_i526_3_lut_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n526_adj_2809)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_8_i526_3_lut_3_lut_3_lut_4_lut.init = 16'h0f70;
    LUT4 i20429_3_lut (.A(n22800), .B(n22801), .C(index_i[8]), .Z(n22803)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20429_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_1_i348_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n348_adj_2914)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A (B ((D)+!C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_1_i348_3_lut_4_lut_4_lut_4_lut.init = 16'h38f0;
    LUT4 mux_231_Mux_9_i316_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n316)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C+(D)))+!A (B (C (D)+!C !(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_9_i316_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h3ff8;
    LUT4 i19950_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n22305)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A (B (C)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19950_3_lut_4_lut_4_lut.init = 16'h3c8c;
    LUT4 index_i_6__bdd_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[6]), .D(n27336), .Z(n25742)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)+!C !(D)))+!A (B (C (D))+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam index_i_6__bdd_4_lut_4_lut_4_lut.init = 16'h0f7c;
    LUT4 i11678_2_lut_2_lut_3_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .Z(n14276)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11678_2_lut_2_lut_3_lut.init = 16'h0808;
    LUT4 mux_231_Mux_7_i491_3_lut_4_lut_4_lut_4_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[2]), .D(index_i[3]), .Z(n491_adj_2958)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A (B ((D)+!C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_7_i491_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'h3870;
    PFUMX i23510 (.BLUT(n25166), .ALUT(n27171), .C0(index_i[5]), .Z(n25167));
    LUT4 n10642_bdd_3_lut_24639_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n26431)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+!(D)))+!A (B (D)+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n10642_bdd_3_lut_24639_4_lut_4_lut_4_lut.init = 16'h30f7;
    LUT4 mux_231_Mux_9_i62_3_lut_4_lut_then_4_lut (.A(index_i[4]), .B(index_i[2]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n27579)) /* synthesis lut_function=(!(A (B (C+(D)))+!A (B+(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_9_i62_3_lut_4_lut_then_4_lut.init = 16'h222b;
    LUT4 mux_231_Mux_9_i62_3_lut_4_lut_else_4_lut (.A(index_i[4]), .B(index_i[2]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n27578)) /* synthesis lut_function=((B+(C (D)))+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_9_i62_3_lut_4_lut_else_4_lut.init = 16'hfddd;
    LUT4 i11652_3_lut_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n14250)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (D))+!A (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11652_3_lut_3_lut_3_lut_4_lut.init = 16'h00f7;
    LUT4 i11852_2_lut_rep_436_4_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n27101)) /* synthesis lut_function=(!(A (B (C+(D))+!B (C+!(D)))+!A (B+(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11852_2_lut_rep_436_4_lut_4_lut_4_lut_4_lut.init = 16'h0308;
    LUT4 n172_bdd_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n26081)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)+!C !(D)))+!A (B (C+!(D))+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n172_bdd_3_lut_4_lut_4_lut_4_lut.init = 16'h0f38;
    LUT4 mux_231_Mux_6_i812_3_lut_4_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n812_adj_2890)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(D))+!A !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_6_i812_3_lut_4_lut_3_lut_4_lut.init = 16'h7780;
    LUT4 mux_231_Mux_4_i1002_3_lut_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n1002_adj_2912)) /* synthesis lut_function=(A (B (C (D))+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_4_i1002_3_lut_3_lut_3_lut_4_lut.init = 16'hf007;
    LUT4 n308_bdd_3_lut_24937_3_lut_4_lut_4_lut_3_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n26190)) /* synthesis lut_function=(A (B (C)+!B !(D))+!A !(D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n308_bdd_3_lut_24937_3_lut_4_lut_4_lut_3_lut_4_lut.init = 16'h80f7;
    LUT4 i1_2_lut_rep_531_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n27196)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_2_lut_rep_531_3_lut_4_lut.init = 16'h8000;
    LUT4 mux_231_Mux_6_i781_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n781_adj_2876)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A (B (C (D)+!C !(D))+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_6_i781_3_lut_4_lut_4_lut_4_lut.init = 16'hc837;
    LUT4 i20987_3_lut (.A(n250), .B(n27337), .C(index_i[3]), .Z(n23361)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20987_3_lut.init = 16'hcaca;
    LUT4 i20986_3_lut (.A(n77), .B(n27417), .C(index_i[3]), .Z(n23360)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20986_3_lut.init = 16'hcaca;
    LUT4 i21396_3_lut (.A(n23757), .B(n25643), .C(index_i[6]), .Z(n23770)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21396_3_lut.init = 16'hcaca;
    LUT4 i21395_3_lut (.A(n25637), .B(n23756), .C(index_i[6]), .Z(n23769)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21395_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_7_i262_3_lut_rep_672_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27337)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_7_i262_3_lut_rep_672_3_lut.init = 16'h3838;
    LUT4 mux_231_Mux_7_i123_3_lut_3_lut_rep_743 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27408)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_7_i123_3_lut_3_lut_rep_743.init = 16'hc7c7;
    PFUMX i24350 (.BLUT(n26081), .ALUT(n26080), .C0(index_i[4]), .Z(n26082));
    LUT4 mux_231_Mux_8_i172_rep_747 (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .Z(n27412)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_8_i172_rep_747.init = 16'h7c7c;
    LUT4 n12154_bdd_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[4]), 
         .D(index_i[2]), .Z(n26579)) /* synthesis lut_function=(A (B)+!A !(B (D)+!B !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n12154_bdd_3_lut_4_lut.init = 16'h98cc;
    LUT4 mux_231_Mux_0_i762_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n762_adj_2839)) /* synthesis lut_function=(A (B+!((D)+!C))+!A !(B (D)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_0_i762_3_lut_4_lut_4_lut.init = 16'h98fc;
    LUT4 mux_231_Mux_5_i924_4_lut_3_lut (.A(index_i[2]), .B(n15075), .C(index_i[4]), 
         .Z(n924_adj_2994)) /* synthesis lut_function=(!(A (B+(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_5_i924_4_lut_3_lut.init = 16'h5656;
    LUT4 i21393_3_lut (.A(n25684), .B(n23752), .C(index_i[6]), .Z(n23767)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21393_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_8_i93_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n93_adj_2870)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C))+!A (B (C+!(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_8_i93_3_lut_3_lut_4_lut.init = 16'h0f83;
    LUT4 mux_231_Mux_7_i620_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n620_adj_2816)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B ((D)+!C)+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_7_i620_3_lut_4_lut_4_lut.init = 16'h83c3;
    LUT4 mux_231_Mux_5_i30_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n30_adj_2940)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A (B+!(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_5_i30_3_lut_4_lut.init = 16'hcc67;
    LUT4 i19632_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21987)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+(D)))+!A !(B (D)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19632_3_lut_4_lut_4_lut.init = 16'h99c7;
    LUT4 n123_bdd_3_lut_24853_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n26499)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C))+!A (B (C (D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n123_bdd_3_lut_24853_3_lut_4_lut.init = 16'h0fc7;
    LUT4 i11759_2_lut_rep_748 (.A(index_i[0]), .B(index_i[1]), .Z(n27413)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11759_2_lut_rep_748.init = 16'heeee;
    LUT4 i1_2_lut_rep_653 (.A(index_i[3]), .B(index_i[2]), .Z(n27318)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_2_lut_rep_653.init = 16'h8888;
    LUT4 mux_231_Mux_0_i333_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n333_adj_2826)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_0_i333_3_lut_3_lut_4_lut.init = 16'hf10e;
    PFUMX i23305 (.BLUT(n24895), .ALUT(n1022), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2145[12]));
    LUT4 i19557_3_lut (.A(n27416), .B(n77), .C(index_i[3]), .Z(n21912)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19557_3_lut.init = 16'hcaca;
    LUT4 i19623_3_lut_3_lut_4_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n21978)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19623_3_lut_3_lut_4_lut_3_lut_4_lut.init = 16'h11ef;
    LUT4 index_i_1__bdd_3_lut_4_lut (.A(index_i[3]), .B(index_i[2]), .C(index_i[4]), 
         .D(index_i[1]), .Z(n23284)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam index_i_1__bdd_3_lut_4_lut.init = 16'h878f;
    LUT4 mux_231_Mux_2_i716_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n716_adj_2965)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)+!C !(D)))+!A (B (D)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_2_i716_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h31cf;
    LUT4 i12562_2_lut_rep_479_3_lut (.A(index_i[3]), .B(index_i[2]), .C(index_i[1]), 
         .Z(n27144)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12562_2_lut_rep_479_3_lut.init = 16'h8080;
    LUT4 i19902_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n22257)) /* synthesis lut_function=(A (B (D)+!B ((D)+!C))+!A (B (D)+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19902_3_lut_4_lut_4_lut_4_lut.init = 16'hfe13;
    LUT4 i20985_3_lut (.A(n29917), .B(n27416), .C(index_i[3]), .Z(n23359)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20985_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_7_i924_3_lut_3_lut_4_lut (.A(index_i[3]), .B(index_i[2]), 
         .C(index_i[4]), .D(n27413), .Z(n924_adj_2974)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_7_i924_3_lut_3_lut_4_lut.init = 16'h878f;
    LUT4 i20984_3_lut (.A(n27337), .B(n27408), .C(index_i[3]), .Z(n23358)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20984_3_lut.init = 16'hcaca;
    LUT4 i12422_2_lut_rep_560_3_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .Z(n27225)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12422_2_lut_rep_560_3_lut.init = 16'he0e0;
    L6MUX21 i24329 (.D0(n26057), .D1(n26055), .SD(index_i[5]), .Z(n26058));
    PFUMX i24327 (.BLUT(n572_adj_2987), .ALUT(n26056), .C0(index_i[4]), 
          .Z(n26057));
    PFUMX i24324 (.BLUT(n26054), .ALUT(n26053), .C0(index_i[4]), .Z(n26055));
    LUT4 index_i_6__bdd_3_lut_4_lut (.A(index_i[3]), .B(index_i[2]), .C(n27407), 
         .D(index_i[6]), .Z(n25743)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(D))+!A !(D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam index_i_6__bdd_3_lut_4_lut.init = 16'h887f;
    LUT4 mux_231_Mux_7_i762_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n762_adj_2957)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A (B (C (D)+!C !(D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_7_i762_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h1cf0;
    LUT4 i11511_2_lut_rep_465_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n27130)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11511_2_lut_rep_465_3_lut_4_lut.init = 16'hfef0;
    LUT4 i11586_2_lut_rep_447_3_lut_4_lut (.A(index_i[3]), .B(index_i[2]), 
         .C(index_i[4]), .D(n27413), .Z(n27112)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11586_2_lut_rep_447_3_lut_4_lut.init = 16'hf8f0;
    LUT4 mux_231_Mux_4_i541_3_lut_4_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n541_adj_2864)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_4_i541_3_lut_4_lut_3_lut_4_lut.init = 16'h0ef0;
    LUT4 i20361_1_lut_2_lut (.A(index_i[3]), .B(index_i[2]), .Z(n22735)) /* synthesis lut_function=(!(A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20361_1_lut_2_lut.init = 16'h7777;
    LUT4 i19924_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n22279)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B ((D)+!C)+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19924_3_lut_4_lut_4_lut.init = 16'hfc1c;
    LUT4 mux_231_Mux_8_i397_3_lut_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n397_adj_2865)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_8_i397_3_lut_3_lut_3_lut_4_lut.init = 16'hf10f;
    LUT4 index_i_0__bdd_4_lut_25214 (.A(index_i[0]), .B(index_i[3]), .C(index_i[1]), 
         .D(index_i[2]), .Z(n27481)) /* synthesis lut_function=(A (B (C)+!B !(C+!(D)))+!A !(B ((D)+!C)+!B !(C (D)+!C !(D)))) */ ;
    defparam index_i_0__bdd_4_lut_25214.init = 16'h92c1;
    LUT4 i11553_2_lut_rep_454_3_lut_4_lut (.A(index_i[3]), .B(index_i[2]), 
         .C(index_i[4]), .D(n27407), .Z(n27119)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11553_2_lut_rep_454_3_lut_4_lut.init = 16'hf8f0;
    LUT4 n348_bdd_3_lut_25037_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n26042)) /* synthesis lut_function=(A (B (D)+!B (C+(D)))+!A (B (D)+!B !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n348_bdd_3_lut_25037_4_lut_4_lut.init = 16'hef30;
    L6MUX21 i24316 (.D0(n26046), .D1(n26043), .SD(index_i[5]), .Z(n26047));
    PFUMX i9508 (.BLUT(n12157), .ALUT(n12158), .C0(n22735), .Z(n11994));
    LUT4 i19951_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n22306)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)+!C !(D)))+!A (B (C+!(D))+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19951_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h0e30;
    PFUMX i24314 (.BLUT(n26045), .ALUT(n26044), .C0(index_i[4]), .Z(n26046));
    LUT4 mux_231_Mux_3_i157_3_lut_3_lut_rep_467_3_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n27132)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_3_i157_3_lut_3_lut_rep_467_3_lut_4_lut.init = 16'h1ff0;
    LUT4 mux_231_Mux_7_i250_3_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n250)) /* synthesis lut_function=(A ((C)+!B)+!A (B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_7_i250_3_lut_4_lut_3_lut.init = 16'he7e7;
    PFUMX i24311 (.BLUT(n27077), .ALUT(n26042), .C0(index_i[4]), .Z(n26043));
    PFUMX i23301 (.BLUT(n254_adj_2971), .ALUT(n24889), .C0(index_i[8]), 
          .Z(n24890));
    LUT4 i12088_2_lut_rep_495_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n27160)) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12088_2_lut_rep_495_3_lut_4_lut.init = 16'he000;
    LUT4 i11725_3_lut_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n14323)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11725_3_lut_3_lut_3_lut_4_lut.init = 16'h10ff;
    LUT4 i11856_2_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n635_adj_2794)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A (B (C+!(D))+!B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11856_2_lut_4_lut_4_lut.init = 16'hf1fc;
    LUT4 i19903_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n22258)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C+(D)))+!A (B (C (D)+!C !(D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19903_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h3ef0;
    LUT4 mux_231_Mux_7_i572_3_lut_rep_411_3_lut_3_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n27076)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_7_i572_3_lut_rep_411_3_lut_3_lut_4_lut.init = 16'hfe01;
    LUT4 mux_231_Mux_8_i101_3_lut_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n101)) /* synthesis lut_function=(!(A (B (C))+!A (B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_8_i101_3_lut_3_lut_3_lut.init = 16'h3e3e;
    LUT4 i12681_1_lut_rep_412_2_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n27077)) /* synthesis lut_function=(!(A (C+(D))+!A (B (C+(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12681_1_lut_rep_412_2_lut_3_lut_4_lut.init = 16'h010f;
    LUT4 mux_231_Mux_8_i46_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n46)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (D)+!B !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_8_i46_3_lut_4_lut_4_lut.init = 16'hcf10;
    LUT4 i21296_3_lut (.A(n23665), .B(n23666), .C(index_i[7]), .Z(n23670)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21296_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_3_i30_3_lut_3_lut_4_lut_3_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n30_adj_2877)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_3_i30_3_lut_3_lut_4_lut_3_lut_4_lut.init = 16'hfe11;
    PFUMX i25505 (.BLUT(n28004), .ALUT(n28003), .C0(index_i[3]), .Z(n28005));
    LUT4 i21197_3_lut (.A(n23564), .B(n23565), .C(index_i[7]), .Z(n23571)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21197_3_lut.init = 16'hcaca;
    LUT4 i21196_3_lut (.A(n23562), .B(n23563), .C(index_i[7]), .Z(n23570)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21196_3_lut.init = 16'hcaca;
    PFUMX i25503 (.BLUT(n28000), .ALUT(n27999), .C0(index_i[2]), .Z(n28001));
    LUT4 mux_231_Mux_5_i38_3_lut_4_lut_3_lut_rep_750 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27415)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_5_i38_3_lut_4_lut_3_lut_rep_750.init = 16'h1919;
    LUT4 mux_231_Mux_7_i29_3_lut_rep_751 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27416)) /* synthesis lut_function=(A (B+!(C))+!A !((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_7_i29_3_lut_rep_751.init = 16'h8e8e;
    LUT4 mux_231_Mux_7_i243_3_lut_rep_752 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27417)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_7_i243_3_lut_rep_752.init = 16'h1c1c;
    LUT4 mux_231_Mux_7_i60_3_lut_4_lut_3_lut_rep_753 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27418)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_7_i60_3_lut_4_lut_3_lut_rep_753.init = 16'h1818;
    LUT4 mux_231_Mux_6_i723_3_lut_rep_754 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27419)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_6_i723_3_lut_rep_754.init = 16'he3e3;
    LUT4 mux_231_Mux_6_i627_3_lut_4_lut_3_lut_rep_756 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27421)) /* synthesis lut_function=(A ((C)+!B)+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_6_i627_3_lut_4_lut_3_lut_rep_756.init = 16'he6e6;
    LUT4 mux_231_Mux_7_i691_3_lut_rep_757 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27422)) /* synthesis lut_function=(!(A (B (C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_7_i691_3_lut_rep_757.init = 16'h7e7e;
    LUT4 mux_231_Mux_8_i30_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n30)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A !(B ((D)+!C)+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_8_i30_3_lut_3_lut_4_lut.init = 16'h7e0f;
    LUT4 mux_231_Mux_6_i635_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n635)) /* synthesis lut_function=(A (B (C+(D))+!B !(D))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_6_i635_3_lut_4_lut.init = 16'hcce6;
    LUT4 n10642_bdd_3_lut_24640_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n26433)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C (D)+!C !(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n10642_bdd_3_lut_24640_3_lut_4_lut.init = 16'h0fc1;
    LUT4 mux_231_Mux_7_i541_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n541_adj_2856)) /* synthesis lut_function=(A (B (C)+!B ((D)+!C))+!A (B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_7_i541_3_lut_4_lut_4_lut.init = 16'he3c3;
    LUT4 mux_231_Mux_2_i557_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n557_adj_2887)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C+!(D))+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_2_i557_3_lut_3_lut_4_lut.init = 16'h0f18;
    LUT4 i19900_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n22255)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A (B (D)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19900_3_lut_4_lut.init = 16'h18cc;
    LUT4 i11562_2_lut_rep_659 (.A(index_i[3]), .B(index_i[4]), .Z(n27324)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11562_2_lut_rep_659.init = 16'h8888;
    LUT4 mux_231_Mux_0_i699_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n699_adj_2835)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (D))+!A (B (C+!(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_0_i699_3_lut_3_lut_4_lut.init = 16'h1c33;
    LUT4 i19995_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n22350)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C (D)))+!A (B (C+(D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19995_4_lut_4_lut_4_lut.init = 16'h301c;
    LUT4 i19564_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21919)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19564_3_lut_3_lut_4_lut.init = 16'h0f1c;
    LUT4 mux_231_Mux_0_i557_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n557)) /* synthesis lut_function=(A ((D)+!C)+!A !((D)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_0_i557_3_lut_4_lut.init = 16'haa4e;
    LUT4 i20433_3_lut_3_lut_4_lut (.A(index_i[3]), .B(index_i[4]), .C(n413), 
         .D(index_i[5]), .Z(n22807)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20433_3_lut_3_lut_4_lut.init = 16'h77f0;
    LUT4 i19563_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21918)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)))+!A !(B (C+!(D))+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19563_3_lut_3_lut_4_lut.init = 16'h71cc;
    PFUMX i23290 (.BLUT(n24870), .ALUT(n24868), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2145[10]));
    PFUMX i21241 (.BLUT(n221_adj_2989), .ALUT(n252_adj_2807), .C0(index_i[5]), 
          .Z(n23615));
    LUT4 i1_2_lut_rep_539_3_lut (.A(index_i[3]), .B(index_i[4]), .C(index_i[5]), 
         .Z(n27204)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_2_lut_rep_539_3_lut.init = 16'hf8f8;
    LUT4 i1_2_lut_3_lut (.A(index_i[3]), .B(index_i[4]), .C(index_i[5]), 
         .Z(n20892)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_2_lut_3_lut.init = 16'h8080;
    LUT4 i20142_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n22497)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(D))+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20142_3_lut_3_lut_4_lut.init = 16'h3319;
    LUT4 i20980_3_lut (.A(n27405), .B(n27408), .C(index_i[3]), .Z(n23354)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20980_3_lut.init = 16'hcaca;
    PFUMX i23288 (.BLUT(n21777), .ALUT(n24866), .C0(index_i[7]), .Z(n24867));
    LUT4 i12104_2_lut_3_lut_4_lut (.A(index_i[3]), .B(index_i[4]), .C(index_i[2]), 
         .D(n27407), .Z(n125_adj_2972)) /* synthesis lut_function=(A (B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12104_2_lut_3_lut_4_lut.init = 16'h8880;
    LUT4 i7499_2_lut_rep_660 (.A(index_i[1]), .B(index_i[2]), .Z(n27325)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i7499_2_lut_rep_660.init = 16'heeee;
    LUT4 mux_231_Mux_7_i716_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n716_adj_2960)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C+!(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_7_i716_3_lut_3_lut_4_lut.init = 16'h0f81;
    LUT4 i20979_3_lut (.A(n29917), .B(n108), .C(index_i[3]), .Z(n23353)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20979_3_lut.init = 16'hcaca;
    PFUMX i21271 (.BLUT(n158), .ALUT(n189_adj_2993), .C0(index_i[5]), 
          .Z(n23645));
    LUT4 n557_bdd_3_lut_23863_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[4]), .D(index_i[3]), .Z(n25574)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C+(D)))+!A (B (C (D)+!C !(D))+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n557_bdd_3_lut_23863_4_lut_4_lut_4_lut.init = 16'hc10f;
    FD1S3BX quarter_wave_sample_register_i_i14 (.D(quarter_wave_sample_register_i_15__N_2145[14]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_i[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_i_i14.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i13 (.D(quarter_wave_sample_register_i_15__N_2145[13]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_i[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_i_i13.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i12 (.D(quarter_wave_sample_register_i_15__N_2145[12]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_i[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_i_i12.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i11 (.D(quarter_wave_sample_register_i_15__N_2145[11]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_i[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_i_i11.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i10 (.D(quarter_wave_sample_register_i_15__N_2145[10]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_i[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_i_i10.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i9 (.D(quarter_wave_sample_register_i_15__N_2145[9]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_i[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_i_i9.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i8 (.D(quarter_wave_sample_register_i_15__N_2145[8]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_i[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_i_i8.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i7 (.D(quarter_wave_sample_register_i_15__N_2145[7]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_i[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_i_i7.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i6 (.D(quarter_wave_sample_register_i_15__N_2145[6]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_i[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_i_i6.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i5 (.D(quarter_wave_sample_register_i_15__N_2145[5]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_i[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_i_i5.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i4 (.D(quarter_wave_sample_register_i_15__N_2145[4]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_i[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_i_i4.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i3 (.D(quarter_wave_sample_register_i_15__N_2145[3]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_i[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_i_i3.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i2 (.D(quarter_wave_sample_register_i_15__N_2145[2]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_i[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_i_i2.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i1 (.D(quarter_wave_sample_register_i_15__N_2145[1]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_i[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_i_i1.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i32 (.D(n1087[15]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_i[0] [15])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i32.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i31 (.D(n1087[14]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_i[0] [14])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i31.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i30 (.D(n1087[13]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_i[0] [13])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i30.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i29 (.D(n1087[12]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_i[0] [12])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i29.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i28 (.D(n1087[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_i[0] [11])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i28.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i27 (.D(n1087[10]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_i[0] [10])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i27.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i26 (.D(n1087[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_i[0] [9])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i26.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i25 (.D(n1087[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_i[0] [8])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i25.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i24 (.D(n1087[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_i[0] [7])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i24.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i23 (.D(n1087[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_i[0] [6])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i23.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i22 (.D(n1087[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_i[0] [5])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i22.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i21 (.D(n1087[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_i[0] [4])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i21.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i20 (.D(n1087[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_i[0] [3])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i20.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i19 (.D(n1087[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_i[0] [2])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i19.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i18 (.D(n1087[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_i[0] [1])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i18.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i17 (.D(n1087[0]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_i[0] [0])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i17.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i16 (.D(\o_val_pipeline_i[0] [15]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(modulation_output[15])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i16.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i15 (.D(\o_val_pipeline_i[0] [14]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(modulation_output[14])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i15.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i14 (.D(\o_val_pipeline_i[0] [13]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(modulation_output[13])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i14.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i13 (.D(\o_val_pipeline_i[0] [12]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(modulation_output[12])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i13.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i12 (.D(\o_val_pipeline_i[0] [11]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(modulation_output[11])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i12.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i11 (.D(\o_val_pipeline_i[0] [10]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(modulation_output[10])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i11.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i10 (.D(\o_val_pipeline_i[0] [9]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(modulation_output[9])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i10.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i9 (.D(\o_val_pipeline_i[0] [8]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(modulation_output[8])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i9.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i8 (.D(\o_val_pipeline_i[0] [7]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(modulation_output[7])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i8.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i7 (.D(\o_val_pipeline_i[0] [6]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(modulation_output[6])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i7.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i6 (.D(\o_val_pipeline_i[0] [5]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(modulation_output[5])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i6.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i5 (.D(\o_val_pipeline_i[0] [4]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(modulation_output[4])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i5.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i4 (.D(\o_val_pipeline_i[0] [3]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(modulation_output[3])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i4.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i3 (.D(\o_val_pipeline_i[0] [2]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(modulation_output[2])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i3.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i2 (.D(\o_val_pipeline_i[0] [1]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(modulation_output[1])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i2.GSR = "DISABLED";
    FD1S3DX index_i_i9 (.D(index_i_9__N_2125[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(index_i[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam index_i_i9.GSR = "DISABLED";
    FD1S3DX index_i_i8 (.D(index_i_9__N_2125[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(index_i[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam index_i_i8.GSR = "DISABLED";
    FD1S3DX index_i_i7 (.D(index_i_9__N_2125[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(index_i[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam index_i_i7.GSR = "DISABLED";
    FD1S3DX index_i_i6 (.D(index_i_9__N_2125[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(index_i[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam index_i_i6.GSR = "DISABLED";
    FD1S3DX index_i_i5 (.D(index_i_9__N_2125[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(index_i[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam index_i_i5.GSR = "DISABLED";
    FD1S3DX index_i_i4 (.D(index_i_9__N_2125[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(index_i[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam index_i_i4.GSR = "DISABLED";
    FD1S3DX index_i_i3 (.D(index_i_9__N_2125[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(index_i[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam index_i_i3.GSR = "DISABLED";
    FD1S3DX index_i_i2 (.D(index_i_9__N_2125[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(index_i[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam index_i_i2.GSR = "DISABLED";
    FD1S3DX index_i_i1 (.D(index_i_9__N_2125[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(index_i[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam index_i_i1.GSR = "DISABLED";
    FD1S3DX phase_negation_i_i1 (.D(phase_negation_i[0]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(phase_negation_i[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam phase_negation_i_i1.GSR = "DISABLED";
    LUT4 i20978_3_lut (.A(n77), .B(n27416), .C(index_i[3]), .Z(n23352)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20978_3_lut.init = 16'hcaca;
    LUT4 mux_231_Mux_11_i766_3_lut (.A(n638), .B(n765), .C(index_i[7]), 
         .Z(n766)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_231_Mux_11_i766_3_lut.init = 16'h3a3a;
    
endmodule
//
// Verilog Description of module \nco(OW=12) 
//

module \nco(OW=12)  (dac_clk_p_c, i_sw0_c, increment, o_phase, GND_net) /* synthesis syn_module_defined=1 */ ;
    input dac_clk_p_c;
    input i_sw0_c;
    input [30:0]increment;
    output [11:0]o_phase;
    input GND_net;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[49:58])
    wire [31:0]n233;
    wire [31:0]n133;
    
    wire n17993, n17992, n17991, n17990, n17989, n17988, n17987, 
        n17986, n17985, n17984, n17983, n17982, n17981, n17980, 
        n17979;
    
    FD1S3DX phase_register_599__i0 (.D(n133[0]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[0])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_599__i0.GSR = "DISABLED";
    CCU2D phase_register_599_add_4_32 (.A0(increment[30]), .B0(o_phase[10]), 
          .C0(GND_net), .D0(GND_net), .A1(o_phase[11]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n17993), .S0(n133[30]), .S1(n133[31]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_599_add_4_32.INIT0 = 16'h5666;
    defparam phase_register_599_add_4_32.INIT1 = 16'hfaaa;
    defparam phase_register_599_add_4_32.INJECT1_0 = "NO";
    defparam phase_register_599_add_4_32.INJECT1_1 = "NO";
    CCU2D phase_register_599_add_4_30 (.A0(increment[28]), .B0(o_phase[8]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[29]), .B1(o_phase[9]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17992), .COUT(n17993), .S0(n133[28]), 
          .S1(n133[29]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_599_add_4_30.INIT0 = 16'h5666;
    defparam phase_register_599_add_4_30.INIT1 = 16'h5666;
    defparam phase_register_599_add_4_30.INJECT1_0 = "NO";
    defparam phase_register_599_add_4_30.INJECT1_1 = "NO";
    CCU2D phase_register_599_add_4_28 (.A0(increment[26]), .B0(o_phase[6]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[27]), .B1(o_phase[7]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17991), .COUT(n17992), .S0(n133[26]), 
          .S1(n133[27]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_599_add_4_28.INIT0 = 16'h5666;
    defparam phase_register_599_add_4_28.INIT1 = 16'h5666;
    defparam phase_register_599_add_4_28.INJECT1_0 = "NO";
    defparam phase_register_599_add_4_28.INJECT1_1 = "NO";
    CCU2D phase_register_599_add_4_26 (.A0(increment[24]), .B0(o_phase[4]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[25]), .B1(o_phase[5]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17990), .COUT(n17991), .S0(n133[24]), 
          .S1(n133[25]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_599_add_4_26.INIT0 = 16'h5666;
    defparam phase_register_599_add_4_26.INIT1 = 16'h5666;
    defparam phase_register_599_add_4_26.INJECT1_0 = "NO";
    defparam phase_register_599_add_4_26.INJECT1_1 = "NO";
    CCU2D phase_register_599_add_4_24 (.A0(increment[22]), .B0(o_phase[2]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[23]), .B1(o_phase[3]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17989), .COUT(n17990), .S0(n133[22]), 
          .S1(n133[23]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_599_add_4_24.INIT0 = 16'h5666;
    defparam phase_register_599_add_4_24.INIT1 = 16'h5666;
    defparam phase_register_599_add_4_24.INJECT1_0 = "NO";
    defparam phase_register_599_add_4_24.INJECT1_1 = "NO";
    LUT4 i15860_2_lut (.A(increment[0]), .B(n233[0]), .Z(n133[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i15860_2_lut.init = 16'h6666;
    CCU2D phase_register_599_add_4_22 (.A0(increment[20]), .B0(o_phase[0]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[21]), .B1(o_phase[1]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17988), .COUT(n17989), .S0(n133[20]), 
          .S1(n133[21]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_599_add_4_22.INIT0 = 16'h5666;
    defparam phase_register_599_add_4_22.INIT1 = 16'h5666;
    defparam phase_register_599_add_4_22.INJECT1_0 = "NO";
    defparam phase_register_599_add_4_22.INJECT1_1 = "NO";
    CCU2D phase_register_599_add_4_20 (.A0(increment[18]), .B0(n233[18]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[19]), .B1(n233[19]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17987), .COUT(n17988), .S0(n133[18]), 
          .S1(n133[19]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_599_add_4_20.INIT0 = 16'h5666;
    defparam phase_register_599_add_4_20.INIT1 = 16'h5666;
    defparam phase_register_599_add_4_20.INJECT1_0 = "NO";
    defparam phase_register_599_add_4_20.INJECT1_1 = "NO";
    CCU2D phase_register_599_add_4_18 (.A0(increment[16]), .B0(n233[16]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[17]), .B1(n233[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17986), .COUT(n17987), .S0(n133[16]), 
          .S1(n133[17]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_599_add_4_18.INIT0 = 16'h5666;
    defparam phase_register_599_add_4_18.INIT1 = 16'h5666;
    defparam phase_register_599_add_4_18.INJECT1_0 = "NO";
    defparam phase_register_599_add_4_18.INJECT1_1 = "NO";
    CCU2D phase_register_599_add_4_16 (.A0(increment[14]), .B0(n233[14]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[15]), .B1(n233[15]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17985), .COUT(n17986), .S0(n133[14]), 
          .S1(n133[15]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_599_add_4_16.INIT0 = 16'h5666;
    defparam phase_register_599_add_4_16.INIT1 = 16'h5666;
    defparam phase_register_599_add_4_16.INJECT1_0 = "NO";
    defparam phase_register_599_add_4_16.INJECT1_1 = "NO";
    CCU2D phase_register_599_add_4_14 (.A0(increment[12]), .B0(n233[12]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[13]), .B1(n233[13]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17984), .COUT(n17985), .S0(n133[12]), 
          .S1(n133[13]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_599_add_4_14.INIT0 = 16'h5666;
    defparam phase_register_599_add_4_14.INIT1 = 16'h5666;
    defparam phase_register_599_add_4_14.INJECT1_0 = "NO";
    defparam phase_register_599_add_4_14.INJECT1_1 = "NO";
    CCU2D phase_register_599_add_4_12 (.A0(increment[10]), .B0(n233[10]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[11]), .B1(n233[11]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17983), .COUT(n17984), .S0(n133[10]), 
          .S1(n133[11]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_599_add_4_12.INIT0 = 16'h5666;
    defparam phase_register_599_add_4_12.INIT1 = 16'h5666;
    defparam phase_register_599_add_4_12.INJECT1_0 = "NO";
    defparam phase_register_599_add_4_12.INJECT1_1 = "NO";
    CCU2D phase_register_599_add_4_10 (.A0(increment[8]), .B0(n233[8]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[9]), .B1(n233[9]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17982), .COUT(n17983), .S0(n133[8]), 
          .S1(n133[9]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_599_add_4_10.INIT0 = 16'h5666;
    defparam phase_register_599_add_4_10.INIT1 = 16'h5666;
    defparam phase_register_599_add_4_10.INJECT1_0 = "NO";
    defparam phase_register_599_add_4_10.INJECT1_1 = "NO";
    CCU2D phase_register_599_add_4_8 (.A0(increment[6]), .B0(n233[6]), .C0(GND_net), 
          .D0(GND_net), .A1(increment[7]), .B1(n233[7]), .C1(GND_net), 
          .D1(GND_net), .CIN(n17981), .COUT(n17982), .S0(n133[6]), .S1(n133[7]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_599_add_4_8.INIT0 = 16'h5666;
    defparam phase_register_599_add_4_8.INIT1 = 16'h5666;
    defparam phase_register_599_add_4_8.INJECT1_0 = "NO";
    defparam phase_register_599_add_4_8.INJECT1_1 = "NO";
    CCU2D phase_register_599_add_4_6 (.A0(increment[4]), .B0(n233[4]), .C0(GND_net), 
          .D0(GND_net), .A1(increment[5]), .B1(n233[5]), .C1(GND_net), 
          .D1(GND_net), .CIN(n17980), .COUT(n17981), .S0(n133[4]), .S1(n133[5]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_599_add_4_6.INIT0 = 16'h5666;
    defparam phase_register_599_add_4_6.INIT1 = 16'h5666;
    defparam phase_register_599_add_4_6.INJECT1_0 = "NO";
    defparam phase_register_599_add_4_6.INJECT1_1 = "NO";
    CCU2D phase_register_599_add_4_4 (.A0(increment[2]), .B0(n233[2]), .C0(GND_net), 
          .D0(GND_net), .A1(increment[3]), .B1(n233[3]), .C1(GND_net), 
          .D1(GND_net), .CIN(n17979), .COUT(n17980), .S0(n133[2]), .S1(n133[3]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_599_add_4_4.INIT0 = 16'h5666;
    defparam phase_register_599_add_4_4.INIT1 = 16'h5666;
    defparam phase_register_599_add_4_4.INJECT1_0 = "NO";
    defparam phase_register_599_add_4_4.INJECT1_1 = "NO";
    CCU2D phase_register_599_add_4_2 (.A0(increment[0]), .B0(n233[0]), .C0(GND_net), 
          .D0(GND_net), .A1(increment[1]), .B1(n233[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n17979), .S1(n133[1]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_599_add_4_2.INIT0 = 16'h7000;
    defparam phase_register_599_add_4_2.INIT1 = 16'h5666;
    defparam phase_register_599_add_4_2.INJECT1_0 = "NO";
    defparam phase_register_599_add_4_2.INJECT1_1 = "NO";
    FD1S3DX phase_register_599__i31 (.D(n133[31]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_phase[11])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_599__i31.GSR = "DISABLED";
    FD1S3DX phase_register_599__i30 (.D(n133[30]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_phase[10])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_599__i30.GSR = "DISABLED";
    FD1S3DX phase_register_599__i29 (.D(n133[29]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_phase[9])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_599__i29.GSR = "DISABLED";
    FD1S3DX phase_register_599__i28 (.D(n133[28]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_phase[8])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_599__i28.GSR = "DISABLED";
    FD1S3DX phase_register_599__i27 (.D(n133[27]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_phase[7])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_599__i27.GSR = "DISABLED";
    FD1S3DX phase_register_599__i26 (.D(n133[26]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_phase[6])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_599__i26.GSR = "DISABLED";
    FD1S3DX phase_register_599__i25 (.D(n133[25]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_phase[5])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_599__i25.GSR = "DISABLED";
    FD1S3DX phase_register_599__i24 (.D(n133[24]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_phase[4])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_599__i24.GSR = "DISABLED";
    FD1S3DX phase_register_599__i23 (.D(n133[23]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_phase[3])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_599__i23.GSR = "DISABLED";
    FD1S3DX phase_register_599__i22 (.D(n133[22]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_phase[2])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_599__i22.GSR = "DISABLED";
    FD1S3DX phase_register_599__i21 (.D(n133[21]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_phase[1])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_599__i21.GSR = "DISABLED";
    FD1S3DX phase_register_599__i20 (.D(n133[20]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_phase[0])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_599__i20.GSR = "DISABLED";
    FD1S3DX phase_register_599__i19 (.D(n133[19]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[19])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_599__i19.GSR = "DISABLED";
    FD1S3DX phase_register_599__i18 (.D(n133[18]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[18])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_599__i18.GSR = "DISABLED";
    FD1S3DX phase_register_599__i17 (.D(n133[17]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[17])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_599__i17.GSR = "DISABLED";
    FD1S3DX phase_register_599__i16 (.D(n133[16]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[16])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_599__i16.GSR = "DISABLED";
    FD1S3DX phase_register_599__i15 (.D(n133[15]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[15])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_599__i15.GSR = "DISABLED";
    FD1S3DX phase_register_599__i14 (.D(n133[14]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[14])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_599__i14.GSR = "DISABLED";
    FD1S3DX phase_register_599__i13 (.D(n133[13]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[13])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_599__i13.GSR = "DISABLED";
    FD1S3DX phase_register_599__i12 (.D(n133[12]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[12])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_599__i12.GSR = "DISABLED";
    FD1S3DX phase_register_599__i11 (.D(n133[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[11])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_599__i11.GSR = "DISABLED";
    FD1S3DX phase_register_599__i10 (.D(n133[10]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[10])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_599__i10.GSR = "DISABLED";
    FD1S3DX phase_register_599__i9 (.D(n133[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[9])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_599__i9.GSR = "DISABLED";
    FD1S3DX phase_register_599__i8 (.D(n133[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[8])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_599__i8.GSR = "DISABLED";
    FD1S3DX phase_register_599__i7 (.D(n133[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[7])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_599__i7.GSR = "DISABLED";
    FD1S3DX phase_register_599__i6 (.D(n133[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[6])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_599__i6.GSR = "DISABLED";
    FD1S3DX phase_register_599__i5 (.D(n133[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[5])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_599__i5.GSR = "DISABLED";
    FD1S3DX phase_register_599__i4 (.D(n133[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[4])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_599__i4.GSR = "DISABLED";
    FD1S3DX phase_register_599__i3 (.D(n133[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[3])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_599__i3.GSR = "DISABLED";
    FD1S3DX phase_register_599__i2 (.D(n133[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[2])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_599__i2.GSR = "DISABLED";
    FD1S3DX phase_register_599__i1 (.D(n133[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[1])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_599__i1.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module dds_U2
//

module dds_U2 (dac_clk_p_c, i_sw0_c, carrier_increment, dac_clk_p_c_enable_488, 
            o_dac_b_c_7, \o_sample_i[7] , \o_sample_i[15] , \o_sample_i[14] , 
            \o_sample_i[13] , \o_sample_i[12] , \o_sample_i[11] , \o_sample_i[10] , 
            \o_sample_i[9] , \o_sample_i[8] , GND_net, \quarter_wave_sample_register_q[15] , 
            n29968, o_dac_b_c_15, o_dac_b_c_14, o_dac_b_c_13, o_dac_b_c_12, 
            o_dac_b_c_11, o_dac_b_c_10, n3639, o_dac_b_c_8) /* synthesis syn_module_defined=1 */ ;
    input dac_clk_p_c;
    input i_sw0_c;
    input [30:0]carrier_increment;
    input dac_clk_p_c_enable_488;
    output o_dac_b_c_7;
    output \o_sample_i[7] ;
    output \o_sample_i[15] ;
    output \o_sample_i[14] ;
    output \o_sample_i[13] ;
    output \o_sample_i[12] ;
    output \o_sample_i[11] ;
    output \o_sample_i[10] ;
    output \o_sample_i[9] ;
    output \o_sample_i[8] ;
    input GND_net;
    output \quarter_wave_sample_register_q[15] ;
    input n29968;
    output o_dac_b_c_15;
    output o_dac_b_c_14;
    output o_dac_b_c_13;
    output o_dac_b_c_12;
    output o_dac_b_c_11;
    output o_dac_b_c_10;
    output n3639;
    output o_dac_b_c_8;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[49:58])
    wire o_dac_b_c_7 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire \o_sample_i[7]  /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[39:49])
    wire \o_sample_i[15]  /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[39:49])
    wire \o_sample_i[14]  /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[39:49])
    wire \o_sample_i[13]  /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[39:49])
    wire \o_sample_i[12]  /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[39:49])
    wire \o_sample_i[11]  /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[39:49])
    wire \o_sample_i[10]  /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[39:49])
    wire \o_sample_i[9]  /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[39:49])
    wire \o_sample_i[8]  /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[39:49])
    wire o_dac_b_c_15 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire o_dac_b_c_14 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire o_dac_b_c_13 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire o_dac_b_c_12 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire o_dac_b_c_11 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire o_dac_b_c_10 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire n3639 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire o_dac_b_c_8 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire [30:0]increment;   // d:/documents/git_local/fm_modulator/rtl/dds.v(14[31:40])
    wire [11:0]o_phase;   // d:/documents/git_local/fm_modulator/rtl/dds.v(18[26:33])
    
    FD1S3DX increment_i0 (.D(carrier_increment[0]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[0])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i0.GSR = "DISABLED";
    FD1S3DX increment_i30 (.D(carrier_increment[30]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(increment[30])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i30.GSR = "DISABLED";
    FD1S3DX increment_i29 (.D(carrier_increment[29]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(increment[29])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i29.GSR = "DISABLED";
    FD1S3DX increment_i28 (.D(carrier_increment[28]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(increment[28])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i28.GSR = "DISABLED";
    FD1S3DX increment_i27 (.D(carrier_increment[27]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(increment[27])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i27.GSR = "DISABLED";
    FD1S3DX increment_i26 (.D(carrier_increment[26]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(increment[26])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i26.GSR = "DISABLED";
    FD1S3DX increment_i25 (.D(carrier_increment[25]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(increment[25])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i25.GSR = "DISABLED";
    FD1S3DX increment_i24 (.D(carrier_increment[24]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(increment[24])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i24.GSR = "DISABLED";
    FD1S3DX increment_i23 (.D(carrier_increment[23]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(increment[23])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i23.GSR = "DISABLED";
    FD1S3DX increment_i22 (.D(carrier_increment[22]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(increment[22])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i22.GSR = "DISABLED";
    FD1S3DX increment_i21 (.D(carrier_increment[21]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(increment[21])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i21.GSR = "DISABLED";
    FD1S3DX increment_i20 (.D(carrier_increment[20]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(increment[20])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i20.GSR = "DISABLED";
    FD1S3DX increment_i19 (.D(carrier_increment[19]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(increment[19])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i19.GSR = "DISABLED";
    FD1S3DX increment_i18 (.D(carrier_increment[18]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(increment[18])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i18.GSR = "DISABLED";
    FD1S3DX increment_i17 (.D(carrier_increment[17]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(increment[17])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i17.GSR = "DISABLED";
    FD1S3DX increment_i16 (.D(carrier_increment[16]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(increment[16])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i16.GSR = "DISABLED";
    FD1S3DX increment_i15 (.D(carrier_increment[15]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(increment[15])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i15.GSR = "DISABLED";
    FD1S3DX increment_i14 (.D(carrier_increment[14]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(increment[14])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i14.GSR = "DISABLED";
    FD1S3DX increment_i13 (.D(carrier_increment[13]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(increment[13])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i13.GSR = "DISABLED";
    FD1S3DX increment_i12 (.D(carrier_increment[12]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(increment[12])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i12.GSR = "DISABLED";
    FD1S3DX increment_i11 (.D(carrier_increment[11]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(increment[11])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i11.GSR = "DISABLED";
    FD1S3DX increment_i10 (.D(carrier_increment[10]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(increment[10])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i10.GSR = "DISABLED";
    FD1S3DX increment_i9 (.D(carrier_increment[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[9])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i9.GSR = "DISABLED";
    FD1S3DX increment_i8 (.D(carrier_increment[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[8])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i8.GSR = "DISABLED";
    FD1S3DX increment_i7 (.D(carrier_increment[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[7])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i7.GSR = "DISABLED";
    FD1S3DX increment_i6 (.D(carrier_increment[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[6])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i6.GSR = "DISABLED";
    FD1S3DX increment_i5 (.D(carrier_increment[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[5])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i5.GSR = "DISABLED";
    FD1S3DX increment_i4 (.D(carrier_increment[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[4])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i4.GSR = "DISABLED";
    FD1S3DX increment_i3 (.D(carrier_increment[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[3])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i3.GSR = "DISABLED";
    FD1S3DX increment_i2 (.D(carrier_increment[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[2])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i2.GSR = "DISABLED";
    FD1S3DX increment_i1 (.D(carrier_increment[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[1])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i1.GSR = "DISABLED";
    quarter_wave_sine_lookup_U0 qtr_inst (.dac_clk_p_c(dac_clk_p_c), .dac_clk_p_c_enable_488(dac_clk_p_c_enable_488), 
            .o_phase({o_phase}), .o_dac_b_c_7(o_dac_b_c_7), .i_sw0_c(i_sw0_c), 
            .\o_sample_i[7] (\o_sample_i[7] ), .\o_sample_i[15] (\o_sample_i[15] ), 
            .\o_sample_i[14] (\o_sample_i[14] ), .\o_sample_i[13] (\o_sample_i[13] ), 
            .\o_sample_i[12] (\o_sample_i[12] ), .\o_sample_i[11] (\o_sample_i[11] ), 
            .\o_sample_i[10] (\o_sample_i[10] ), .\o_sample_i[9] (\o_sample_i[9] ), 
            .\o_sample_i[8] (\o_sample_i[8] ), .GND_net(GND_net), .\quarter_wave_sample_register_q[15] (\quarter_wave_sample_register_q[15] ), 
            .n29968(n29968), .o_dac_b_c_15(o_dac_b_c_15), .o_dac_b_c_14(o_dac_b_c_14), 
            .o_dac_b_c_13(o_dac_b_c_13), .o_dac_b_c_12(o_dac_b_c_12), .o_dac_b_c_11(o_dac_b_c_11), 
            .o_dac_b_c_10(o_dac_b_c_10), .n3639(n3639), .o_dac_b_c_8(o_dac_b_c_8)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(21[70:134])
    \nco(OW=12)_U1  nco_inst (.increment({increment}), .o_phase({o_phase}), 
            .GND_net(GND_net), .dac_clk_p_c(dac_clk_p_c), .i_sw0_c(i_sw0_c)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(20[49:100])
    
endmodule
//
// Verilog Description of module quarter_wave_sine_lookup_U0
//

module quarter_wave_sine_lookup_U0 (dac_clk_p_c, dac_clk_p_c_enable_488, 
            o_phase, o_dac_b_c_7, i_sw0_c, \o_sample_i[7] , \o_sample_i[15] , 
            \o_sample_i[14] , \o_sample_i[13] , \o_sample_i[12] , \o_sample_i[11] , 
            \o_sample_i[10] , \o_sample_i[9] , \o_sample_i[8] , GND_net, 
            \quarter_wave_sample_register_q[15] , n29968, o_dac_b_c_15, 
            o_dac_b_c_14, o_dac_b_c_13, o_dac_b_c_12, o_dac_b_c_11, 
            o_dac_b_c_10, n3639, o_dac_b_c_8) /* synthesis syn_module_defined=1 */ ;
    input dac_clk_p_c;
    input dac_clk_p_c_enable_488;
    input [11:0]o_phase;
    output o_dac_b_c_7;
    input i_sw0_c;
    output \o_sample_i[7] ;
    output \o_sample_i[15] ;
    output \o_sample_i[14] ;
    output \o_sample_i[13] ;
    output \o_sample_i[12] ;
    output \o_sample_i[11] ;
    output \o_sample_i[10] ;
    output \o_sample_i[9] ;
    output \o_sample_i[8] ;
    input GND_net;
    output \quarter_wave_sample_register_q[15] ;
    input n29968;
    output o_dac_b_c_15;
    output o_dac_b_c_14;
    output o_dac_b_c_13;
    output o_dac_b_c_12;
    output o_dac_b_c_11;
    output o_dac_b_c_10;
    output n3639;
    output o_dac_b_c_8;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[49:58])
    wire o_dac_b_c_7 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire [15:0]\o_val_pipeline_q[0]  /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(16[24:40])
    wire \o_sample_i[7]  /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[39:49])
    wire [15:0]\o_val_pipeline_i[0]  /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(15[24:40])
    wire \o_sample_i[15]  /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[39:49])
    wire \o_sample_i[14]  /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[39:49])
    wire \o_sample_i[13]  /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[39:49])
    wire \o_sample_i[12]  /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[39:49])
    wire \o_sample_i[11]  /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[39:49])
    wire \o_sample_i[10]  /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[39:49])
    wire \o_sample_i[9]  /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[39:49])
    wire \o_sample_i[8]  /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[39:49])
    wire o_dac_b_c_15 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire o_dac_b_c_14 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire o_dac_b_c_13 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire o_dac_b_c_12 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire o_dac_b_c_11 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire o_dac_b_c_10 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire n3639 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire o_dac_b_c_8 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire [9:0]index_q;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(31[26:33])
    
    wire n27424, n27297, n29934, n364, n29958, n23380, n668, n23218, 
        n23219;
    wire [14:0]quarter_wave_sample_register_q_15__N_2160;
    
    wire n939, n954;
    wire [9:0]index_i;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(31[17:24])
    
    wire n23537, n22008, n22009, n22010, n26658, n157, n27429, 
        n27162, n25796, n25795, n25797, n22011, n22012, n22013, 
        n716, n14102, n142, n25779, n25776, n21815, n908, n412, 
        n22348, n22017, n22018, n22019, n22363, n27381, n20714, 
        n25785, n25783, n21818, n22020, n22021, n22022, n22893, 
        n22894;
    wire [14:0]quarter_wave_sample_register_i_15__N_2145;
    
    wire n25784, n62, n25010, n25007, n27219, n27174, n189, n971, 
        n986, n23538, n25782, n25781;
    wire [11:0]phase_q;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(12[17:24])
    
    wire n22032, n22033, n22034, n25009, n25008, n29935, n379, 
        n205, n26220, n25778, n25777, n27538, n22035, n22036, 
        n22037, n28892, n22984, n22985, n22987, n22955, n22956, 
        n29955, n27279, n22248, n27339, n22982, n22983, n22986, 
        n22249, n22250, n158, n23676, n22038, n22039, n22040, 
        n27274, n27277, n1002, n1017, n23539;
    wire [1:0]phase_negation_i;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(23[12:28])
    wire [11:0]phase_i;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(11[17:24])
    wire [1:0]phase_negation_q;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(23[30:46])
    wire [9:0]index_i_9__N_2125;
    wire [9:0]index_q_9__N_2135;
    wire [15:0]quarter_wave_sample_register_q;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(22[56:86])
    wire [15:0]quarter_wave_sample_register_i;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(22[24:54])
    
    wire n29913, n204, n397, n348, n349, n25761, n25759, n21809, 
        n25760, n62_adj_2269, n38, n14, n22245, n27348, n29944, 
        n506, n27200, n27123, n637, n18112, n22041, n22042, n22043, 
        n25758, n25757, n574, n637_adj_2270, n21786, n27255, n21756, 
        n21757, n29914, n27388, n15, n23187, n23188, n22246, n22247, 
        n22047, n22048, n22049, n404, o_val_pipeline_i_0__15__N_2175, 
        o_val_pipeline_i_0__15__N_2177, n23698, n23699, n23702, o_val_pipeline_i_0__15__N_2179, 
        o_val_pipeline_i_0__15__N_2181, o_val_pipeline_i_0__15__N_2183, 
        o_val_pipeline_i_0__15__N_2185, o_val_pipeline_i_0__15__N_2187, 
        n23748, n23749, o_val_pipeline_i_0__15__N_2189, o_val_pipeline_i_0__15__N_2191, 
        n557, n511, n20675, n17892;
    wire [15:0]o_val_pipeline_q_0__15__N_2208;
    
    wire n716_adj_2271, n27477, n27478, n27479, n22137, n22138, 
        n931, n23523, n23554, n23492, n23819, n851, n859, n25006, 
        n22923, n22843, n22844, n22847, n22862, n22863, n333, 
        n511_adj_2272, n20536, n27385, n27435, n875, n22671, n286, 
        n317, n22776, n27278, n29919, n22237, n27159, n21018, 
        n27125, n27299, n22030, n251, n26451, n29922, n27352, 
        n61, n29912, n270;
    wire [14:0]n1790;
    
    wire n23011, n23012, n23016, n23552, n23553;
    wire [11:0]phase_q_11__N_2251;
    
    wire n635, n21693, n21694, n21695, n21696, n21697, n21698, 
        n23059, n23060, n23063, n17891, n23061, n23062, n23064, 
        n22065, n22066, n476, n23150, n23151, n23155, n23212, 
        n23213, n23217, n17890, n588, n15_adj_2273, n27350, n27346, 
        n348_adj_2274, n652, n660, n684, n23267, n23268, n23271, 
        n23269, n23270, n23272, n23690, n23691, n27474, n27475, 
        n27476, n23692, n23693, n17889, n27296, n22504, n27673, 
        n27672, n27674, n620, n635_adj_2275, n636, n21708, n21709, 
        n21710, n26661, n25718, n25715, n22787, n27669, n27668, 
        n27670, n844, n12112, n23799, n27574, n27575, n27576, 
        n27256, n22308, n27386, n22835, n22836, n25717, n25716, 
        n18092, n653, n349_adj_2276, n29925, n985, n22837, n22838, 
        n27275, n985_adj_2277, n986_adj_2278, n22095, n22096, n22097, 
        n27340, n21711, n21712, n21713, n27568, n27569, n27570, 
        n29928, n971_adj_2279, n27257, n22029, n22031, n27214, n22347, 
        n27471, n27472, n27473, n23817, n23818, n27224, n25714, 
        n25713, n491, n21744, n25711, n25708, n25712, n332, n21714, 
        n21715, n21716, n26195, n15_adj_2280, n25710, n25709, n22949, 
        n22950, n22954, n27565, n27566, n27567, n23490, n23491, 
        n23521, n23522, n23001, n23002, n23007, n23008, n23014, 
        n18105, n18106, n18107, n46, n29923, n27439, n27238, n22027, 
        n27425, n684_adj_2281, n875_adj_2282, n890, n891, n23055, 
        n23056, n23057, n23058, n27436, n27537, n844_adj_2283, n859_adj_2284, 
        n860, n27561, n27562, n27563, n21717, n21718, n21719, 
        n14095, n25707, n25706, n23082, n23083, n23090, n954_adj_2285, 
        n27071, n23084, n23085, n23091, n23581, n23582, n23583, 
        n285, n142_adj_2286, n27438, n173, n27126, n27166, n23372, 
        n23373, n23376, n27558, n27559, n27560, n27440, n23140, 
        n23141, n23144, n23145, n23152, n23146, n23147, n23153, 
        n23177, n23178, n23184, n21723, n21724, n21725, n23154, 
        n23157, n23179, n23180, n23185, n23181, n23182, n23186, 
        n27467, n27468, n11955, n17888, n29951, n27345, n25816, 
        n29926, n22174, n27442, n24994, n24991, n22225, n27218, 
        n316, n23296, n26359, n9630, n765, n747, n29952, n27347, 
        n25824, n890_adj_2287, n891_adj_2288, n23156, n557_adj_2289, 
        n14_adj_2290, n22000, n23094, n27387, n25827, n93, n21967, 
        n17887, n23200, n23201, n23211, n498, n27342, n25830, 
        n23202, n23203, n22210, n25831, n23208, n23209, n23215, 
        n443, n26167, n308, n21999, n27389, n348_adj_2291, n29916, 
        n173_adj_2292, n541, n251_adj_2293, n27220, n412_adj_2294, 
        n23302, n574_adj_2295, n21795, n747_adj_2296, n762, n763, 
        n27358, n25834, n27147, n23304, n413, n908_adj_2297, n157_adj_2298, 
        n828, n25838, n157_adj_2299, n25839, n444, n27317, n221, 
        n18125, n1017_adj_2300, n381, n27172, n252, n22345, n142_adj_2301, 
        n716_adj_2302, n762_adj_2303, n781, n506_adj_2304, n23374, 
        n23375, n23377, n26387, n22281, n716_adj_2305, n604, n635_adj_2306, 
        n26165, n526, n428, n444_adj_2307, n21783, n21784, n21785, 
        n25794, n21824, n22026, n22028, n17886, n541_adj_2308, n29936, 
        n653_adj_2309, n23015, n23018, n557_adj_2310, n24993, n24992, 
        n397_adj_2311, n443_adj_2312, n23013, n23017, n844_adj_2313, 
        n11927, n23534, n11924, n875_adj_2314, n526_adj_2315, n316_adj_2316, 
        n653_adj_2317, n23263, n23264, n635_adj_2318, n26778, n251_adj_2319, 
        n844_adj_2320, n27316, n221_adj_2321, n18118, n781_adj_2322, 
        n23265, n23266, n716_adj_2323, n428_adj_2324, n844_adj_2325, 
        n22192, n762_adj_2326, n24843, n26094, n26091, n475, n684_adj_2327, 
        n23694, n23695, n23700, n21738, n21739, n476_adj_2328, n27349, 
        n21705, n475_adj_2329, n747_adj_2330, n21726, n23740, n23741, 
        n23746, n18091, n23742, n23743, n23747, n954_adj_2331, n22282, 
        n24844, n24849, n812, n27464, n27465, n27466, n27074, 
        n955, n27068, n701, n24851, n27253, n939_adj_2332, n22357, 
        n22788, n24854, n21792, n21793, n21794, n22782, n24855, 
        n252_adj_2333, n699, n890_adj_2334, n22116, n22780, n22781, 
        n27096, n251_adj_2335, n23558, n23379, n23383, n699_adj_2336, 
        n109, n460, n23556, n22401, n27156, n413_adj_2337, n27229, 
        n252_adj_2338, n828_adj_2339, n26358, n25917, n25918, n22185, 
        n22186, n22187, n22024, n22267, n22398, n381_adj_2340, n15_adj_2341, 
        n23557, n27488, n27097, n22191, n22193, n22839, n22840, 
        n22845, n22854, n22855, n22860, n22856, n22857, n22861, 
        n251_adj_2342, n684_adj_2343, n27383, n23608, n443_adj_2344, 
        n379_adj_2345, n443_adj_2346, n23607, n22889, n22890, n23606, 
        n379_adj_2347, n27432, n23605, n22881, n22882, n412_adj_2348, 
        n22242, n25921, n27392, n23601, n22883, n22884, n27549, 
        n27550, n27551, n15350, n252_adj_2349, n24876, n890_adj_2350, 
        n890_adj_2351, n699_adj_2352, n22939, n22940, n23600, n109_adj_2353, 
        n460_adj_2354, n22943, n22944, n22951, n890_adj_2355, n604_adj_2356, 
        n22444, n445, n716_adj_2357, n27271, n22945, n22946, n22952, 
        n22976, n22977, n26484, n27248, n445_adj_2358, n252_adj_2359, 
        n27461, n27462, n27463, n716_adj_2360, n23599, n27213, n891_adj_2361, 
        n22978, n22979, n22980, n22981, n25978, n25979, n173_adj_2362, 
        n27623, n23381, n23382, n23384, n29931, n923, n24877, 
        n24882, n25980, n25983, n23598, n27252, n27291, n25516, 
        n348_adj_2363, n356, n890_adj_2364, n29945, n22999, n23000, 
        n23010, n23003, n23004, n22290, n23594, n1001, n23593, 
        n23591, n23386, n23387, n23390, n18089, n18088, n27322, 
        n635_adj_2365, n22150, n526_adj_2366, n542, n27301, n700, 
        n23388, n23389, n23391, n27334, n526_adj_2367, n542_adj_2368, 
        n21964, n557_adj_2369, n124, n21949, n526_adj_2370, n541_adj_2371, 
        n23789, n22052, n22112, n23054, n22505, n22118, n93_adj_2372, 
        n23464, n22121, n22124, n22447, n22127, n892, n29953, 
        n142_adj_2373, n157_adj_2374, n158_adj_2375, n605, n526_adj_2376, 
        n541_adj_2377, n23524, n27263, n475_adj_2378, n491_adj_2379, 
        n29229, n189_adj_2380, n27458, n27459, n27460, n22947, n22948, 
        n22953, n22937, n22938, n27434, n22402, n859_adj_2381, n285_adj_2382, 
        n27624, n27625, n27540, n27541, n27542, n27394, n908_adj_2383, 
        n526_adj_2384, n23393, n23394, n23397, n716_adj_2385, n557_adj_2386, 
        n572, n23790, n900, n22525, n29929, n23066, n23067, n23068, 
        n23069, n23070, n23071, n23072, n23073, n23074, n23075, 
        n23086, n23078, n23079, n23088, n23577, n23578, n173_adj_2387, 
        n25150, n23097, n23098, n23113, n25649, n27052, n638, 
        n23099, n23100, n23114, n23395, n23396, n23398, n23101, 
        n23102, n23115, n25648, n25647, n589, n23791, n46_adj_2388, 
        n23105, n23106, n23117, n23107, n23108, n23118, n23579, 
        n23580, n22848, n22846, n23076, n23077, n23087, n25417, 
        n23176, n23183, n27305, n700_adj_2389, n620_adj_2390, n635_adj_2391, 
        n23792, n23109, n23110, n23119, n23111, n23112, n23120, 
        n27293, n27307, n15348, n25630, n25627, n509, n25629, 
        n25628, n541_adj_2392, n26093, n25626, n25625, n27539, n26119, 
        n27494, n124_adj_2393, n25411, n699_adj_2394, n23463, n526_adj_2395, 
        n25413, n22090, n26128, n22239, n10667, n797, n26130, 
        n1021, n26983, n26984, n653_adj_2396, n668_adj_2397, n23793, 
        n23128, n23129, n23130, n23131, n23132, n23133, n23134, 
        n23135, n23136, n23137, n23148, n23142, n23143, n28896, 
        n12079, n731, n732, n356_adj_2398, n21751, n23161, n23162, 
        n23163, n23164, n23165, n23166, n23167, n23168, n23169, 
        n23170, n21750, n21752, n684_adj_2399, n23794, n27267, n475_adj_2400, 
        n27426, n491_adj_2401, n732_adj_2402, n763_adj_2403, n124_adj_2404, 
        n22244, n891_adj_2405, n23190, n23191, n23206, n23194, n23195, 
        n23196, n23197, n23316, n573, n23204, n23205, n716_adj_2406, 
        n731_adj_2407, n23795, n29959, n109_adj_2408, n573_adj_2409, 
        n27195, n27179, n25198, n397_adj_2410, n573_adj_2411, n22203, 
        n22204, n22205, n125;
    wire [15:0]o_val_pipeline_i_0__15__N_2176;
    
    wire n27269, n29941, n668_adj_2412, n23597, n23604, n23259, 
        n762_adj_2413, n22172, n22181, n23262, n747_adj_2414, n763_adj_2415, 
        n29918, n22190, n22199, n22208, n22217, n29938, n22220, 
        n892_adj_2416, n220, n23468, n747_adj_2417, n23796, n26164, 
        n27302, n15218, n189_adj_2418, n508, n27086, n27120, n638_adj_2419, 
        n27064, n27382, n924, n27498, n23682, n23683, n22875, 
        n22876, n22886, n22389, n22390, n22391, n27288, n26173, 
        n23684, n23685, n23686, n23687, n23696, n23688, n23689, 
        n23697, n20112, n29964, n22381, n22382, n27185, n27165, 
        n25220, n796, n23797, n23703, n23701, n25984, n22975, 
        n22209, n22211, n541_adj_2420, n348_adj_2421, n349_adj_2422, 
        n22353, n22354, n22355, n812_adj_2423, n12109, n23798, n364_adj_2424, 
        n23299, n23300, n23301, n22212, n22213, n22214, n254, 
        n27066, n875_adj_2425, n23800, n23306, n23307, n23308, n22195, 
        n22224, n22226, n93_adj_2426, n94, n23801, n27087, n27116, 
        n638_adj_2427, n12043, n21953, n23737, n954_adj_2428, n23802, 
        n254_adj_2429, n21959, n21962, n23739, n23320, n23321, n382, 
        n574_adj_2430, n21965, n21968, n764, n27320, n20603, n22868, 
        n23803, n27455, n27456, n1002_adj_2431, n23804, n221_adj_2432, 
        n619, n939_adj_2433, n27430, n25264, n22230, n22231, n22232, 
        n747_adj_2434, n22777, n22236, n22238, n27321, n444_adj_2435, 
        n22778, n22779, n22240, n22241, n29940, n27499, n236, 
        n23500, n27353, n25813, n668_adj_2436, n22243, n397_adj_2437, 
        n21947, n21950, n23736, n763_adj_2438, n892_adj_2439, n23493, 
        n22785, n22786, n29911, n27500, n22309, n190, n26535, 
        n23052, n14724, n27502, n23399, n21971, n23053, n731_adj_2440, 
        n22399, n251_adj_2441, n11265, n26219, n731_adj_2442, n732_adj_2443, 
        n25833, n669, n142_adj_2444, n604_adj_2445, n605_adj_2446, 
        n684_adj_2447, n700_adj_2448, n22327, n22328, n22320, n22321, 
        n22322, n397_adj_2449, n413_adj_2450, n316_adj_2451, n317_adj_2452, 
        n25601, n27053, n23315, n270_adj_2453, n653_adj_2454, n286_adj_2455, 
        n25644, n30, n31, n20166, n1018, n190_adj_2456, n253, 
        n23260, n29924, n62_adj_2457, n27098, n31_adj_2458, n23611, 
        n22160, n23261, n653_adj_2459, n30_adj_2460, n31_adj_2461, 
        n22045, n25600, n25599, n11977, n11978, n189_adj_2462, n684_adj_2463, 
        n26096, n23378, n23738, n15_adj_2464, n30_adj_2465, n31_adj_2466, 
        n27208, n61_adj_2467, n62_adj_2468, n15_adj_2469, n27158, 
        n31_adj_2470, n25596, n30_adj_2471, n31_adj_2472, n796_adj_2473, 
        n12103, n12104, n29231, n158_adj_2474, n29946, n22101, n62_adj_2475, 
        n28686, n27501, n27450, n28684, n22827, n22828, n28687, 
        n892_adj_2476, n22829, n22830, n29947, n22831, n22832, n22841, 
        n22833, n22834, n22842, n684_adj_2477, n27193, n23469, n22266, 
        n22268, n12124, n22136, n22851, n27622, n23116, n24930, 
        n22145, n22148, n22853, n574_adj_2478, n22151, n860_adj_2479, 
        n22154, n764_adj_2480, n29960, n23462, n46_adj_2481, n21946, 
        n684_adj_2482, n28766, n22299, n22301, n28767, n924_adj_2483, 
        n22865, n22866, n890_adj_2484, n891_adj_2485, n22867, n22869, 
        n22870, n29948, n669_adj_2486, n11965, n22871, n22872, n22873, 
        n22874, n22885, n22877, n22878, n22887, n23805, n23806, 
        n23813, n23807, n23808, n23814, n23809, n23810, n23815, 
        n23811, n23812, n23816, n22283, n22896, n22897, n22912, 
        n22898, n22899, n22913, n22900, n22901, n22914, n316_adj_2487, 
        n23317, n460_adj_2488, n285_adj_2489, n476_adj_2490, n22904, 
        n22905, n22916, n22906, n22907, n22917, n413_adj_2491, n22234, 
        n22908, n22909, n22918, n26390, n23561, n22852, n22910, 
        n22911, n22919, n93_adj_2492, n286_adj_2493, n24928, n158_adj_2494, 
        n797_adj_2495, n29949, n109_adj_2496, n125_adj_2497, n22200, 
        n22927, n22928, n124_adj_2498, n22929, n22930, n28893, n28895, 
        n1002_adj_2499, n908_adj_2500, n860_adj_2501, n892_adj_2502, 
        n15_adj_2503, n860_adj_2504, n22931, n22932, n29233, n23481, 
        n23487, n21747, n21748, n21749, n28898, n23483, n23488, 
        n22933, n22934, n21745, n21746, n22935, n22936, n22941, 
        n22942, n23511, n23512, n23518, n26729, n23514, n23519, 
        n475_adj_2505, n124_adj_2506, n318, n700_adj_2507, n668_adj_2508, 
        n669_adj_2509, n318_adj_2510, n24931, n542_adj_2511, n27152, 
        n27505, n189_adj_2512, n508_adj_2513, n29950, n27323, n27276, 
        n444_adj_2514, n286_adj_2515, n157_adj_2516, n27280, n27504, 
        n27449, n859_adj_2517, n23478, n23479, n23486, n27355, n94_adj_2518, 
        n23385, n23392, n23051, n491_adj_2519, n491_adj_2520, n23484, 
        n23485, n23489, n158_adj_2521, n29921, n24990, n23785, n732_adj_2522, 
        n22001, n22960, n22961, n22962, n22963, n22964, n22965, 
        n890_adj_2523, n891_adj_2524, n22966, n22967, n860_adj_2525, 
        n23509, n23510, n23517, n27124, n22968, n22969, n23515, 
        n23516, n23520, n27528, n27529, n27530, n26986, n21720, 
        n21721, n21722, n22356, n29915, n22130, n22133, n22850, 
        n700_adj_2526, n22291, n22292, n157_adj_2527, n27212, n636_adj_2528, 
        n18093, n26982, n507, n460_adj_2529, n475_adj_2530, n476_adj_2531, 
        n20198, n1018_adj_2532, n413_adj_2533, n732_adj_2534, n763_adj_2535, 
        n27371, n23295, n22403, n891_adj_2536, n22989, n22990, n23005, 
        n22113, n573_adj_2537, n573_adj_2538, n27525, n27526, n27527, 
        n397_adj_2539, n573_adj_2540, n18117, n18119, n109_adj_2541, 
        n124_adj_2542, n125_adj_2543, n653_adj_2544, n94_adj_2545, n29166, 
        n29167, n23297, n27522, n27523, n27524, n12047, n30_adj_2546, 
        n22993, n22994, n27626, n23540, n23541, n23548, n22995, 
        n22996, n22056, n23542, n23543, n23549, n23544, n23545, 
        n23550, n23546, n23547, n23551, n173_adj_2547, n747_adj_2548, 
        n908_adj_2549, n22216, n15204, n22215, n93_adj_2550, n22207, 
        n620_adj_2551, n653_adj_2552, n22206, n29228, n78, n891_adj_2553, 
        n812_adj_2554, n14070, n828_adj_2555, n844_adj_2556, n25353, 
        n25354, n797_adj_2557, n668_adj_2558, n669_adj_2559, n526_adj_2560, 
        n542_adj_2561, n26452, n526_adj_2562, n22188, n22189, n475_adj_2563, 
        n26454, n26455, n21703, n23494, n15103, n25357, n22197, 
        n286_adj_2564, n397_adj_2565, n22179, n348_adj_2566, n443_adj_2567, 
        n22171, n781_adj_2568, n22170, n25266, n22892, n21702, n23207, 
        n23214, n22284, n860_adj_2569, n491_adj_2570, n23192, n26169, 
        n364_adj_2571, n22159, n23210, n23216, n333_adj_2572, n22158, 
        n23559, n23560, n26175, n23199, n22503, n27508, n348_adj_2573, 
        n491_adj_2574, n22147, n220_adj_2575, n23499, n956, n20671, 
        n475_adj_2576, n22146, n27131, n23586, n22003, n221_adj_2577, 
        n22144, n22143, n93_adj_2578, n23495, n27507, n30_adj_2579, 
        n94_adj_2580, n125_adj_2581, n23318, n18126, n12128, n22131, 
        n22128, n413_adj_2582, n668_adj_2583, n24945, n22123, n15090, 
        n22122, n476_adj_2584, n507_adj_2585, n18113, n573_adj_2586, 
        n22344, n22346, n890_adj_2587, n605_adj_2588, n636_adj_2589, 
        n22349, n93_adj_2590, n22120, n22119, n22046, n700_adj_2591, 
        n25412, n797_adj_2592, n828_adj_2593, n397_adj_2594, n22110, 
        n26531, n860_adj_2595, n891_adj_2596, n27155, n860_adj_2597, 
        n892_adj_2598, n22891, n25416, n12145, n22397, n22388, n173_adj_2599, 
        n94_adj_2600, n22055, n21945, n348_adj_2601, n443_adj_2602, 
        n22051, n21948, n731_adj_2603, n22050, n24947, n22057, n221_adj_2604, 
        n252_adj_2605, n22362, n22364, n286_adj_2606, n22058, n22061, 
        n22365, n22366, n22367, n29966, n923_adj_2607, n21957, n21958, 
        n22858, n22859, n29965, n22371, n22372, n22373, n27111, 
        n27117, n669_adj_2608, n700_adj_2609, n22098, n22526, n22152, 
        n22044, n27127, n27183, n22073, n828_adj_2610, n22374, n22375, 
        n22376, n29956, n27113, n27118, n860_adj_2611, n22076, n22285, 
        n716_adj_2612, n27627, n22317, n21960, n21961, n27072, n27335, 
        n653_adj_2613, n26779, n26777, n26780, n21963, n27108, n25262, 
        n26776, n26775, n27629, n24948, n620_adj_2614, n572_adj_2615, 
        n573_adj_2616, n589_adj_2617, n364_adj_2618, n21014, n12127, 
        n796_adj_2619, n21966, n572_adj_2620, n732_adj_2621, n22714, 
        n22449, n15004, n22450, n22451, n22446, n22448, n94_adj_2622, 
        n125_adj_2623, n22149, n158_adj_2624, n23592, n78_adj_2625, 
        n891_adj_2626, n286_adj_2627, n22085, n812_adj_2628, n14376, 
        n828_adj_2629, n27075, n797_adj_2630, n349_adj_2631, n22088, 
        n333_adj_2632, n23472, n653_adj_2633, n668_adj_2634, n669_adj_2635, 
        n413_adj_2636, n444_adj_2637, n12053, n476_adj_2638, n507_adj_2639, 
        n22383, n22384, n22385, n26662, n542_adj_2640, n397_adj_2641, 
        n25148, n22730, n15358, n23473, n22155, n188, n27328, 
        n22091, n26659, n27104, n15412, n12091, n22094, n669_adj_2642, 
        n700_adj_2643, n23138, n364_adj_2644, n12046, n26196, n124_adj_2645, 
        n23496, n397_adj_2646, n23474, n27393, n731_adj_2647, n23139, 
        n26703, n860_adj_2648, n891_adj_2649, n27351, n22339, n26728, 
        n26725, n924_adj_2650, n22100, n26727, n26726, n25515, n22103, 
        n23475, n21969, n21970, n747_adj_2651, n23595, n23596, n158_adj_2652, 
        n22392, n22393, n22394, n25525, n25522, n25526, n25524, 
        n475_adj_2653, n221_adj_2654, n22109, n924_adj_2655, n22395, 
        n22396, n27628, n286_adj_2656, n317_adj_2657, n22233, n22235, 
        n25518, n349_adj_2658, n22115, n348_adj_2659, n349_adj_2660, 
        n22724, n22194, n22196, n14081, n413_adj_2661, n22157, n636_adj_2662, 
        n26724, n22163, n507_adj_2663, n22169, n93_adj_2664, n94_adj_2665, 
        n25521, n23476, n605_adj_2666, n22175, n26705, n669_adj_2667, 
        n732_adj_2668, n763_adj_2669, n27084, n731_adj_2670, n653_adj_2671, 
        n23172, n22400, n142_adj_2672, n604_adj_2673, n23602, n23603, 
        n22168, n22161, n22162, n397_adj_2674, n23609, n23610, n316_adj_2675, 
        n491_adj_2676, n11325, n23477, n270_adj_2677, n653_adj_2678, 
        n491_adj_2679, n26706, n26704, n26707, n27289, n572_adj_2680, 
        n14388, n333_adj_2681, n27470, n908_adj_2682, n22387, n22386, 
        n22184, n22089, n460_adj_2683, n285_adj_2684, n397_adj_2685, 
        n506_adj_2686, n27310, n93_adj_2687, n15111, n859_adj_2688, 
        n25519, n25517, n25520, n875_adj_2689, n27311, n317_adj_2690, 
        n26702, n22202, n1002_adj_2691, n270_adj_2692, n491_adj_2693, 
        n29967, n27181, n987, n890_adj_2694, n891_adj_2695, n108, 
        n684_adj_2696, n22071, n22072, n22524, n542_adj_2697, n859_adj_2698, 
        n860_adj_2699, n29963, n27503, n15_adj_2700, n763_adj_2701, 
        n27309, n348_adj_2702, n27085, n22358, n124_adj_2703, n23465, 
        n22431, n22432, n22433, n301, n908_adj_2704, n317_adj_2705, 
        n27427, n27211, n732_adj_2706, n900_adj_2707, n18111, n573_adj_2708, 
        n460_adj_2709, n26663, n26660, n26664, n22340, n18124, n635_adj_2710, 
        n142_adj_2711, n157_adj_2712, n23497, n986_adj_2713, n22329, 
        n22330, n22331, n24949, n24946, n605_adj_2714, n27182, n766, 
        n23498, n924_adj_2715, n22318, n22319, n924_adj_2716, n956_adj_2717, 
        n684_adj_2718, n701_adj_2719, n22312, n22311, n22313, n348_adj_2720, 
        n23503, n22310, n364_adj_2721, n23504, n15194, n27060, n23675, 
        n27178, n1021_adj_2722, n27069, n27451, n23505, n23679, 
        n12055, n23680, n573_adj_2723, n636_adj_2724, n23506, n22294, 
        n22293, n22295, n28689, n22972, n15104, n27062, n700_adj_2725, 
        n23507, n732_adj_2726, n20896, n254_adj_2727, n22286, n20888, 
        n254_adj_2728, n11368, n23508, n173_adj_2729, n22276, n22275, 
        n22277, n22273, n22272, n22274, n924_adj_2730, n22443, n22445, 
        n924_adj_2731, n955_adj_2732, n22201, n205_adj_2733, n25840, 
        n732_adj_2734, n684_adj_2735, n700_adj_2736, n20711, n20187, 
        n986_adj_2737, n23525, n26221, n23526, n26486, n22219, n635_adj_2738, 
        n23527, n23298, n22740, n22092, n20213, n23255, n491_adj_2739, 
        n23528, n14725, n23303, n23529, n23305, n23530, n23173, 
        n26132, n762_adj_2740, n23531, n828_adj_2741, n25203, n797_adj_2742, 
        n23532, n23319, n812_adj_2743, n23533, n796_adj_2744, n27506, 
        n27509, n94_adj_2745, n875_adj_2746, n23535, n23006, n22991, 
        n23009, n22997, n22998, n23536, n62_adj_2747, n700_adj_2748, 
        n27070, n27264, n26534, n26532, n26533, n882, n890_adj_2749, 
        n27268, n22915, n620_adj_2750, n22111, n22117, n908_adj_2751, 
        n22129, n22132, n23149, n22053, n22054, n317_adj_2752, n348_adj_2753, 
        n349_adj_2754, n26170, n507_adj_2755, n12165, n22153, n205_adj_2756, 
        n221_adj_2757, n26485, n11969, n763_adj_2758, n17900, n14744, 
        n301_adj_2759, n26385, n22180, n491_adj_2760, n26360, n22126, 
        n25814, n444_adj_2761, n26172, n23744, n23745, n252_adj_2762, 
        n26453, n26388, n62_adj_2763, n27480, n22820, n18090, n22824, 
        n11931, n22825, n605_adj_2764, n636_adj_2765, n24932, n24929, 
        n27285, n21704, n29232, n29230, n860_adj_2766, n22198, n22183, 
        n22971, n22074, n572_adj_2767, n22093, n812_adj_2768, n491_adj_2769, 
        n14743, n26389, n26386, n620_adj_2770, n14788, n12095, n27384, 
        n25825, n700_adj_2771, n12129, n765_adj_2772, n1022, n828_adj_2773, 
        n1022_adj_2774, n22156, n27247, n507_adj_2775, n21728, n21731, 
        n15146, n21734, n491_adj_2776, n506_adj_2777, n22173, n27081, 
        n12048, n27675, n25837, n28897, n28894, n189_adj_2778, n252_adj_2779, 
        n882_adj_2780, n349_adj_2781, n22107, n26116, n21733, n21732, 
        n25265, n25263, n12166, n27107, n21727, n21730, n21729, 
        n924_adj_2782, n28688, n28685, n25201, n25152, n23093, n26121, 
        n62_adj_2783, n23092, n23095, n62_adj_2784, n26127, n12172, 
        n25225, n221_adj_2785, n573_adj_2786, n17899, n987_adj_2787, 
        n14372, n22114, n21707, n17898, n23124, n506_adj_2788, n12152, 
        n22108, n12151, n12173, n25224, n572_adj_2789, n17897, n22099, 
        n23555, n26174, n26171, n26118, n25836, n25829, n26168, 
        n26166, n25202, n25819, n27671, n26131, n26129, n924_adj_2790, 
        n17896, n22087, n29961, n22086, n26120, n26117, n29962, 
        n22743, n26095, n26092, n25151, n25149, n22084, n22083, 
        n24852, n24853, n22729, n21706, n22075, n20713, n766_adj_2791, 
        n93_adj_2792, n22060, n22059, n17895, n17894, n25835, n25832, 
        n25828, n25826, n25818, n25815;
    
    LUT4 i12491_2_lut_rep_759 (.A(index_q[2]), .B(index_q[0]), .Z(n27424)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i12491_2_lut_rep_759.init = 16'heeee;
    LUT4 mux_230_Mux_7_i364_3_lut_3_lut (.A(n27297), .B(index_q[3]), .C(n29934), 
         .Z(n364)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;
    defparam mux_230_Mux_7_i364_3_lut_3_lut.init = 16'hd1d1;
    LUT4 i21006_3_lut_3_lut (.A(n27297), .B(index_q[3]), .C(n29958), .Z(n23380)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam i21006_3_lut_3_lut.init = 16'h7474;
    LUT4 mux_230_Mux_4_i668_3_lut_3_lut (.A(n27297), .B(index_q[3]), .C(n29958), 
         .Z(n668)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;
    defparam mux_230_Mux_4_i668_3_lut_3_lut.init = 16'hd1d1;
    PFUMX i20846 (.BLUT(n23218), .ALUT(n23219), .C0(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_2160[1]));
    PFUMX i21163 (.BLUT(n939), .ALUT(n954), .C0(index_i[4]), .Z(n23537));
    PFUMX i19655 (.BLUT(n22008), .ALUT(n22009), .C0(index_q[4]), .Z(n22010));
    LUT4 index_i_5__bdd_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n26658)) /* synthesis lut_function=(A (B (C)+!B (C+(D)))+!A (B (C)+!B !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam index_i_5__bdd_3_lut_4_lut_4_lut_4_lut.init = 16'he3f0;
    LUT4 mux_229_Mux_3_i157_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n157)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_3_i157_3_lut_3_lut_4_lut.init = 16'h1ff0;
    LUT4 i1_3_lut_rep_497_4_lut (.A(index_i[3]), .B(index_i[4]), .C(index_i[2]), 
         .D(n27429), .Z(n27162)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_3_lut_rep_497_4_lut.init = 16'hfffe;
    PFUMX i24086 (.BLUT(n25796), .ALUT(n25795), .C0(index_i[5]), .Z(n25797));
    PFUMX i19658 (.BLUT(n22011), .ALUT(n22012), .C0(index_q[4]), .Z(n22013));
    LUT4 mux_229_Mux_2_i716_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n716)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)+!C !(D)))+!A (B (D)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_2_i716_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h31cf;
    LUT4 i11505_3_lut_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n14102)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11505_3_lut_3_lut_3_lut_4_lut.init = 16'h10ff;
    LUT4 mux_229_Mux_4_i142_3_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[3]), 
         .C(index_i[2]), .Z(n142)) /* synthesis lut_function=(A (B (C))+!A !(B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_4_i142_3_lut_4_lut_3_lut.init = 16'h9595;
    LUT4 n25779_bdd_3_lut (.A(n25779), .B(n25776), .C(index_q[4]), .Z(n21815)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n25779_bdd_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_0_i908_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n908)) /* synthesis lut_function=(!(A (B (C (D))+!B !(D))+!A (B+((D)+!C)))) */ ;
    defparam mux_230_Mux_0_i908_3_lut_4_lut_4_lut.init = 16'h2a98;
    LUT4 mux_229_Mux_0_i412_3_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[1]), .D(index_i[3]), .Z(n412)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C (D)))+!A (B (C+!(D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_0_i412_3_lut_4_lut_4_lut.init = 16'hf14c;
    LUT4 i19993_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n22348)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C+(D)))+!A (B (C (D)+!C !(D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19993_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h3ef0;
    PFUMX i19664 (.BLUT(n22017), .ALUT(n22018), .C0(index_q[4]), .Z(n22019));
    LUT4 i20008_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n22363)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B ((D)+!C)+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20008_3_lut_4_lut_4_lut.init = 16'hfc1c;
    LUT4 i1_3_lut_4_lut (.A(index_i[3]), .B(index_i[4]), .C(index_i[5]), 
         .D(n27381), .Z(n20714)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_3_lut_4_lut.init = 16'hfffe;
    L6MUX21 i24075 (.D0(n25785), .D1(n25783), .SD(index_i[6]), .Z(n21818));
    PFUMX i19667 (.BLUT(n22020), .ALUT(n22021), .C0(index_q[4]), .Z(n22022));
    PFUMX i20521 (.BLUT(n22893), .ALUT(n22894), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2145[5]));
    PFUMX i24073 (.BLUT(n25784), .ALUT(n62), .C0(index_i[5]), .Z(n25785));
    L6MUX21 i23408 (.D0(n25010), .D1(n25007), .SD(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2145[4]));
    LUT4 mux_230_Mux_3_i189_3_lut_3_lut_4_lut (.A(n27219), .B(index_q[3]), 
         .C(index_q[4]), .D(n27174), .Z(n189)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_3_i189_3_lut_3_lut_4_lut.init = 16'h08f8;
    PFUMX i21164 (.BLUT(n971), .ALUT(n986), .C0(index_i[4]), .Z(n23538));
    PFUMX i24071 (.BLUT(n25782), .ALUT(n25781), .C0(index_i[5]), .Z(n25783));
    FD1P3AX phase_q__i1 (.D(o_phase[0]), .SP(dac_clk_p_c_enable_488), .CK(dac_clk_p_c), 
            .Q(phase_q[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam phase_q__i1.GSR = "DISABLED";
    PFUMX i19679 (.BLUT(n22032), .ALUT(n22033), .C0(index_q[4]), .Z(n22034));
    PFUMX i23406 (.BLUT(n25009), .ALUT(n25008), .C0(index_i[8]), .Z(n25010));
    LUT4 mux_230_Mux_7_i379_3_lut_3_lut (.A(n27297), .B(index_q[3]), .C(n29935), 
         .Z(n379)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam mux_230_Mux_7_i379_3_lut_3_lut.init = 16'h7474;
    LUT4 n251_bdd_3_lut_4_lut (.A(index_q[0]), .B(index_q[2]), .C(index_q[4]), 
         .D(n205), .Z(n26220)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam n251_bdd_3_lut_4_lut.init = 16'h6f60;
    PFUMX i24068 (.BLUT(n25778), .ALUT(n25777), .C0(index_q[5]), .Z(n25779));
    LUT4 i23669_then_4_lut (.A(index_q[0]), .B(index_q[4]), .C(index_q[1]), 
         .D(index_q[3]), .Z(n27538)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam i23669_then_4_lut.init = 16'h3c69;
    PFUMX i19682 (.BLUT(n22035), .ALUT(n22036), .C0(index_q[4]), .Z(n22037));
    LUT4 n581_bdd_3_lut_26341_4_lut (.A(index_q[2]), .B(index_q[1]), .C(index_q[0]), 
         .D(index_q[5]), .Z(n28892)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(D))+!A (B (D)+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam n581_bdd_3_lut_26341_4_lut.init = 16'h33c4;
    LUT4 i20613_3_lut (.A(n22984), .B(n22985), .C(index_i[8]), .Z(n22987)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20613_3_lut.init = 16'hcaca;
    PFUMX i20583 (.BLUT(n22955), .ALUT(n22956), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2145[3]));
    LUT4 i19893_3_lut (.A(n29955), .B(n27279), .C(index_q[3]), .Z(n22248)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19893_3_lut.init = 16'hcaca;
    LUT4 i2765_2_lut_rep_674 (.A(index_i[0]), .B(index_i[2]), .Z(n27339)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i2765_2_lut_rep_674.init = 16'h6666;
    LUT4 i20612_3_lut (.A(n22982), .B(n22983), .C(index_i[8]), .Z(n22986)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20612_3_lut.init = 16'hcaca;
    LUT4 i22304_3_lut (.A(n22248), .B(n22249), .C(index_q[4]), .Z(n22250)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22304_3_lut.init = 16'hcaca;
    LUT4 i21302_3_lut_4_lut (.A(index_q[0]), .B(index_q[2]), .C(index_q[5]), 
         .D(n158), .Z(n23676)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i21302_3_lut_4_lut.init = 16'h6f60;
    PFUMX i19685 (.BLUT(n22038), .ALUT(n22039), .C0(index_q[4]), .Z(n22040));
    LUT4 i19677_3_lut (.A(n27274), .B(n27277), .C(index_q[3]), .Z(n22032)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19677_3_lut.init = 16'hcaca;
    PFUMX i21165 (.BLUT(n1002), .ALUT(n1017), .C0(index_i[4]), .Z(n23539));
    FD1S3DX o_val_pipeline_q_1__i1 (.D(\o_val_pipeline_q[0] [7]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(o_dac_b_c_7)) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_q_1__i1.GSR = "DISABLED";
    FD1S3DX phase_negation_i_i0 (.D(phase_i[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(phase_negation_i[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam phase_negation_i_i0.GSR = "DISABLED";
    FD1S3DX phase_negation_q_i0 (.D(phase_q[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(phase_negation_q[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam phase_negation_q_i0.GSR = "DISABLED";
    FD1S3DX index_i_i0 (.D(index_i_9__N_2125[0]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(index_i[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam index_i_i0.GSR = "DISABLED";
    FD1S3DX index_q_i0 (.D(index_q_9__N_2135[0]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(index_q[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam index_q_i0.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i0 (.D(quarter_wave_sample_register_q_15__N_2160[0]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_q[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_q_i0.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i1 (.D(\o_val_pipeline_i[0] [7]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(\o_sample_i[7] )) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i1.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i0 (.D(quarter_wave_sample_register_i_15__N_2145[0]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_i[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_i_i0.GSR = "DISABLED";
    LUT4 mux_229_Mux_5_i397_3_lut (.A(n29913), .B(n204), .C(index_i[3]), 
         .Z(n397)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_5_i397_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_4_i349_3_lut_4_lut (.A(index_q[0]), .B(index_q[2]), 
         .C(index_q[4]), .D(n348), .Z(n349)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_4_i349_3_lut_4_lut.init = 16'hf606;
    L6MUX21 i24049 (.D0(n25761), .D1(n25759), .SD(index_q[6]), .Z(n21809));
    PFUMX i24047 (.BLUT(n25760), .ALUT(n62_adj_2269), .C0(index_q[5]), 
          .Z(n25761));
    LUT4 i19890_3_lut (.A(n38), .B(n14), .C(index_q[3]), .Z(n22245)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19890_3_lut.init = 16'hcaca;
    FD1S3BX quarter_wave_sample_register_i_i14 (.D(quarter_wave_sample_register_i_15__N_2145[14]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_i[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_i_i14.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i13 (.D(quarter_wave_sample_register_i_15__N_2145[13]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_i[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_i_i13.GSR = "DISABLED";
    LUT4 mux_229_Mux_5_i506_3_lut (.A(n27348), .B(n29944), .C(index_i[3]), 
         .Z(n506)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_5_i506_3_lut.init = 16'hcaca;
    FD1S3BX quarter_wave_sample_register_i_i12 (.D(quarter_wave_sample_register_i_15__N_2145[12]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_i[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_i_i12.GSR = "DISABLED";
    LUT4 mux_229_Mux_10_i637_3_lut_4_lut_4_lut (.A(n27200), .B(index_i[4]), 
         .C(index_i[5]), .D(n27123), .Z(n637)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_10_i637_3_lut_4_lut_4_lut.init = 16'h1f1c;
    FD1S3BX quarter_wave_sample_register_i_i11 (.D(quarter_wave_sample_register_i_15__N_2145[11]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_i[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_i_i11.GSR = "DISABLED";
    LUT4 i15926_3_lut_3_lut (.A(index_q[0]), .B(index_q[2]), .C(index_q[3]), 
         .Z(n18112)) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i15926_3_lut_3_lut.init = 16'h6a6a;
    FD1S3BX quarter_wave_sample_register_i_i10 (.D(quarter_wave_sample_register_i_15__N_2145[10]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_i[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_i_i10.GSR = "DISABLED";
    PFUMX i19688 (.BLUT(n22041), .ALUT(n22042), .C0(index_q[4]), .Z(n22043));
    PFUMX i24045 (.BLUT(n25758), .ALUT(n25757), .C0(index_q[5]), .Z(n25759));
    FD1S3BX quarter_wave_sample_register_i_i9 (.D(quarter_wave_sample_register_i_15__N_2145[9]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_i[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_i_i9.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i8 (.D(quarter_wave_sample_register_i_15__N_2145[8]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_i[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_i_i8.GSR = "DISABLED";
    LUT4 i22927_3_lut (.A(n574), .B(n637_adj_2270), .C(index_q[6]), .Z(n21786)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22927_3_lut.init = 16'hcaca;
    FD1S3BX quarter_wave_sample_register_i_i7 (.D(quarter_wave_sample_register_i_15__N_2145[7]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_i[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_i_i7.GSR = "DISABLED";
    LUT4 i11358_2_lut_rep_590 (.A(index_i[0]), .B(index_i[1]), .Z(n27255)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11358_2_lut_rep_590.init = 16'h4444;
    PFUMX i19403 (.BLUT(n21756), .ALUT(n21757), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2145[11]));
    FD1S3BX quarter_wave_sample_register_i_i6 (.D(quarter_wave_sample_register_i_15__N_2145[6]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_i[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_i_i6.GSR = "DISABLED";
    LUT4 mux_229_Mux_5_i15_3_lut (.A(n29914), .B(n27388), .C(index_i[3]), 
         .Z(n15)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_5_i15_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_554_3_lut (.A(index_q[2]), .B(index_q[0]), .C(index_q[1]), 
         .Z(n27219)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_554_3_lut.init = 16'hfefe;
    FD1S3BX quarter_wave_sample_register_i_i5 (.D(quarter_wave_sample_register_i_15__N_2145[5]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_i[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_i_i5.GSR = "DISABLED";
    PFUMX i20815 (.BLUT(n23187), .ALUT(n23188), .C0(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_2160[2]));
    FD1S3BX quarter_wave_sample_register_i_i4 (.D(quarter_wave_sample_register_i_15__N_2145[4]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_i[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_i_i4.GSR = "DISABLED";
    LUT4 i22306_3_lut (.A(n22245), .B(n22246), .C(index_q[4]), .Z(n22247)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22306_3_lut.init = 16'hcaca;
    FD1S3BX quarter_wave_sample_register_i_i3 (.D(quarter_wave_sample_register_i_15__N_2145[3]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_i[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_i_i3.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i2 (.D(quarter_wave_sample_register_i_15__N_2145[2]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_i[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_i_i2.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i1 (.D(quarter_wave_sample_register_i_15__N_2145[1]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_i[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_i_i1.GSR = "DISABLED";
    PFUMX i19694 (.BLUT(n22047), .ALUT(n22048), .C0(index_q[4]), .Z(n22049));
    LUT4 mux_230_Mux_6_i498_3_lut_4_lut_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n404)) /* synthesis lut_function=(A (B+!(C))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_6_i498_3_lut_4_lut_3_lut.init = 16'h9b9b;
    FD1S3DX o_val_pipeline_i_1__i18 (.D(o_val_pipeline_i_0__15__N_2175), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(\o_val_pipeline_i[0] [15])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i18.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i17 (.D(o_val_pipeline_i_0__15__N_2177), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(\o_val_pipeline_i[0] [14])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i17.GSR = "DISABLED";
    L6MUX21 i21328 (.D0(n23698), .D1(n23699), .SD(index_q[8]), .Z(n23702));
    FD1S3DX o_val_pipeline_i_1__i16 (.D(o_val_pipeline_i_0__15__N_2179), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(\o_val_pipeline_i[0] [13])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i16.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i15 (.D(o_val_pipeline_i_0__15__N_2181), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(\o_val_pipeline_i[0] [12])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i15.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i14 (.D(o_val_pipeline_i_0__15__N_2183), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(\o_val_pipeline_i[0] [11])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i14.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i13 (.D(o_val_pipeline_i_0__15__N_2185), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(\o_val_pipeline_i[0] [10])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i13.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i12 (.D(o_val_pipeline_i_0__15__N_2187), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(\o_val_pipeline_i[0] [9])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i12.GSR = "DISABLED";
    PFUMX i21376 (.BLUT(n23748), .ALUT(n23749), .C0(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_2160[8]));
    FD1S3DX o_val_pipeline_i_1__i11 (.D(o_val_pipeline_i_0__15__N_2189), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(\o_val_pipeline_i[0] [8])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i11.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i10 (.D(o_val_pipeline_i_0__15__N_2191), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(\o_val_pipeline_i[0] [7])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i10.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i9 (.D(\o_val_pipeline_i[0] [15]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(\o_sample_i[15] )) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i9.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i8 (.D(\o_val_pipeline_i[0] [14]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(\o_sample_i[14] )) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i8.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i7 (.D(\o_val_pipeline_i[0] [13]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(\o_sample_i[13] )) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i7.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i6 (.D(\o_val_pipeline_i[0] [12]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(\o_sample_i[12] )) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i6.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i5 (.D(\o_val_pipeline_i[0] [11]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(\o_sample_i[11] )) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i5.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i4 (.D(\o_val_pipeline_i[0] [10]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(\o_sample_i[10] )) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i4.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i3 (.D(\o_val_pipeline_i[0] [9]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(\o_sample_i[9] )) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i3.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i2 (.D(\o_val_pipeline_i[0] [8]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(\o_sample_i[8] )) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i2.GSR = "DISABLED";
    LUT4 mux_229_Mux_1_i557_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n557)) /* synthesis lut_function=(A (B (C+(D)))+!A (B ((D)+!C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_1_i557_3_lut_4_lut.init = 16'hcc94;
    PFUMX mux_229_Mux_14_i1023 (.BLUT(n511), .ALUT(n20675), .C0(index_i[9]), 
          .Z(quarter_wave_sample_register_i_15__N_2145[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 mux_229_Mux_0_i954_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n954)) /* synthesis lut_function=(A (D)+!A !(B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_0_i954_3_lut_4_lut_4_lut.init = 16'haf40;
    CCU2D add_418_15 (.A0(quarter_wave_sample_register_q[14]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(\quarter_wave_sample_register_q[15] ), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17892), .S0(o_val_pipeline_q_0__15__N_2208[14]), 
          .S1(o_val_pipeline_q_0__15__N_2208[15]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(81[29:60])
    defparam add_418_15.INIT0 = 16'hf555;
    defparam add_418_15.INIT1 = 16'hf555;
    defparam add_418_15.INJECT1_0 = "NO";
    defparam add_418_15.INJECT1_1 = "NO";
    LUT4 mux_230_Mux_8_i716_3_lut_4_lut_4_lut_4_lut (.A(index_q[2]), .B(index_q[0]), 
         .C(index_q[1]), .D(index_q[3]), .Z(n716_adj_2271)) /* synthesis lut_function=(!(A (D)+!A !(B+(C+(D))))) */ ;
    defparam mux_230_Mux_8_i716_3_lut_4_lut_4_lut_4_lut.init = 16'h55fe;
    PFUMX i25158 (.BLUT(n27477), .ALUT(n27478), .C0(index_i[0]), .Z(n27479));
    PFUMX i19784 (.BLUT(n22137), .ALUT(n22138), .C0(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_2160[11]));
    LUT4 mux_229_Mux_2_i931_3_lut_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n931)) /* synthesis lut_function=(!(A (B (C))+!A (B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_2_i931_3_lut_3_lut_3_lut.init = 16'h3e3e;
    L6MUX21 i13250362_i1 (.D0(n23523), .D1(n23554), .SD(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2145[0]));
    L6MUX21 i13244359_i1 (.D0(n23492), .D1(n23819), .SD(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_2160[0]));
    LUT4 mux_229_Mux_5_i859_3_lut (.A(n851), .B(n29914), .C(index_i[3]), 
         .Z(n859)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_5_i859_3_lut.init = 16'hcaca;
    PFUMX i23403 (.BLUT(n25006), .ALUT(n22923), .C0(index_i[8]), .Z(n25007));
    FD1S3BX quarter_wave_sample_register_q_i15 (.D(n29968), .CK(dac_clk_p_c), 
            .PD(i_sw0_c), .Q(\quarter_wave_sample_register_q[15] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_q_i15.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i14 (.D(quarter_wave_sample_register_q_15__N_2160[14]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_q[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_q_i14.GSR = "DISABLED";
    L6MUX21 i20473 (.D0(n22843), .D1(n22844), .SD(index_i[8]), .Z(n22847));
    PFUMX i20490 (.BLUT(n22862), .ALUT(n22863), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2145[8]));
    LUT4 mux_229_Mux_0_i333_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n333)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_0_i333_3_lut_3_lut_4_lut.init = 16'hf10e;
    PFUMX mux_230_Mux_14_i1023 (.BLUT(n511_adj_2272), .ALUT(n20536), .C0(index_q[9]), 
          .Z(quarter_wave_sample_register_q_15__N_2160[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 mux_229_Mux_5_i875_3_lut (.A(n27385), .B(n27435), .C(index_i[3]), 
         .Z(n875)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_5_i875_3_lut.init = 16'hcaca;
    LUT4 i23114_2_lut (.A(index_q[5]), .B(index_q[4]), .Z(n22671)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i23114_2_lut.init = 16'heeee;
    LUT4 i22592_3_lut (.A(n286), .B(n317), .C(index_q[5]), .Z(n22776)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22592_3_lut.init = 16'hcaca;
    LUT4 i19882_3_lut (.A(n27278), .B(n29919), .C(index_q[3]), .Z(n22237)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19882_3_lut.init = 16'hcaca;
    LUT4 i11960_2_lut_rep_494_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n27159)) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11960_2_lut_rep_494_3_lut_4_lut.init = 16'he000;
    LUT4 i1_3_lut (.A(index_q[0]), .B(index_q[4]), .C(index_q[2]), .Z(n21018)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i1_3_lut.init = 16'hfefe;
    LUT4 i11574_2_lut_rep_460_3_lut_4_lut (.A(index_q[2]), .B(index_q[0]), 
         .C(index_q[3]), .D(index_q[1]), .Z(n27125)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;
    defparam i11574_2_lut_rep_460_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i19675_3_lut (.A(n27299), .B(n29958), .C(index_q[3]), .Z(n22030)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19675_3_lut.init = 16'hcaca;
    LUT4 index_i_5__bdd_3_lut_24845_4_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(n251), .D(index_i[5]), .Z(n26451)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam index_i_5__bdd_3_lut_24845_4_lut.init = 16'hf066;
    LUT4 mux_229_Mux_4_i61_3_lut (.A(n29922), .B(n27352), .C(index_i[3]), 
         .Z(n61)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_4_i61_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_4_i270_3_lut (.A(n29912), .B(n27348), .C(index_i[3]), 
         .Z(n270)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_4_i270_3_lut.init = 16'hcaca;
    FD1S3BX quarter_wave_sample_register_q_i13 (.D(quarter_wave_sample_register_q_15__N_2160[13]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_q[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_q_i13.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i12 (.D(quarter_wave_sample_register_q_15__N_2160[12]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_q[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_q_i12.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i11 (.D(quarter_wave_sample_register_q_15__N_2160[11]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_q[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_q_i11.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i10 (.D(quarter_wave_sample_register_q_15__N_2160[10]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_q[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_q_i10.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i9 (.D(quarter_wave_sample_register_q_15__N_2160[9]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_q[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_q_i9.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i8 (.D(quarter_wave_sample_register_q_15__N_2160[8]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_q[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_q_i8.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i7 (.D(quarter_wave_sample_register_q_15__N_2160[7]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_q[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_q_i7.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i6 (.D(quarter_wave_sample_register_q_15__N_2160[6]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_q[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_q_i6.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i5 (.D(quarter_wave_sample_register_q_15__N_2160[5]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_q[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_q_i5.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i4 (.D(quarter_wave_sample_register_q_15__N_2160[4]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_q[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_q_i4.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i3 (.D(quarter_wave_sample_register_q_15__N_2160[3]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_q[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_q_i3.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i2 (.D(quarter_wave_sample_register_q_15__N_2160[2]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_q[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_q_i2.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i1 (.D(quarter_wave_sample_register_q_15__N_2160[1]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_q[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_q_i1.GSR = "DISABLED";
    FD1S3DX index_q_i9 (.D(index_q_9__N_2135[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(index_q[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam index_q_i9.GSR = "DISABLED";
    FD1S3DX index_q_i8 (.D(index_q_9__N_2135[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(index_q[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam index_q_i8.GSR = "DISABLED";
    PFUMX i20614 (.BLUT(n22986), .ALUT(n22987), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2145[2]));
    FD1S3DX index_q_i7 (.D(index_q_9__N_2135[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(index_q[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam index_q_i7.GSR = "DISABLED";
    FD1S3DX index_q_i6 (.D(index_q_9__N_2135[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(index_q[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam index_q_i6.GSR = "DISABLED";
    FD1S3DX index_q_i5 (.D(index_q_9__N_2135[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(index_q[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam index_q_i5.GSR = "DISABLED";
    FD1S3DX index_q_i4 (.D(index_q_9__N_2135[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(index_q[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam index_q_i4.GSR = "DISABLED";
    FD1S3DX index_q_i3 (.D(index_q_9__N_2135[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(index_q[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam index_q_i3.GSR = "DISABLED";
    FD1S3DX index_q_i2 (.D(index_q_9__N_2135[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(index_q[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam index_q_i2.GSR = "DISABLED";
    FD1S3DX index_q_i1 (.D(index_q_9__N_2135[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(index_q[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam index_q_i1.GSR = "DISABLED";
    FD1S3DX index_i_i9 (.D(index_i_9__N_2125[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(index_i[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam index_i_i9.GSR = "DISABLED";
    FD1S3DX index_i_i8 (.D(index_i_9__N_2125[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(index_i[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam index_i_i8.GSR = "DISABLED";
    FD1S3DX index_i_i7 (.D(index_i_9__N_2125[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(index_i[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam index_i_i7.GSR = "DISABLED";
    FD1S3DX index_i_i6 (.D(index_i_9__N_2125[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(index_i[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam index_i_i6.GSR = "DISABLED";
    FD1S3DX index_i_i5 (.D(index_i_9__N_2125[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(index_i[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam index_i_i5.GSR = "DISABLED";
    FD1S3DX index_i_i4 (.D(index_i_9__N_2125[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(index_i[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam index_i_i4.GSR = "DISABLED";
    FD1S3DX index_i_i3 (.D(index_i_9__N_2125[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(index_i[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam index_i_i3.GSR = "DISABLED";
    FD1S3DX index_i_i2 (.D(index_i_9__N_2125[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(index_i[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam index_i_i2.GSR = "DISABLED";
    FD1S3DX index_i_i1 (.D(index_i_9__N_2125[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(index_i[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam index_i_i1.GSR = "DISABLED";
    FD1S3DX phase_negation_q_i1 (.D(phase_negation_q[0]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(phase_negation_q[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam phase_negation_q_i1.GSR = "DISABLED";
    FD1S3DX phase_negation_i_i1 (.D(phase_negation_i[0]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(phase_negation_i[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam phase_negation_i_i1.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i18 (.D(n1790[14]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_q[0] [15])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_q_1__i18.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i17 (.D(n1790[13]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_q[0] [14])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_q_1__i17.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i16 (.D(n1790[12]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_q[0] [13])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_q_1__i16.GSR = "DISABLED";
    L6MUX21 i20642 (.D0(n23011), .D1(n23012), .SD(index_i[7]), .Z(n23016));
    FD1S3DX o_val_pipeline_q_1__i15 (.D(n1790[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_q[0] [12])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_q_1__i15.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i14 (.D(n1790[10]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_q[0] [11])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_q_1__i14.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i13 (.D(n1790[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_q[0] [10])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_q_1__i13.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i12 (.D(n1790[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_q[0] [9])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_q_1__i12.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i11 (.D(n1790[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_q[0] [8])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_q_1__i11.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i10 (.D(n1790[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_q[0] [7])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_q_1__i10.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i9 (.D(\o_val_pipeline_q[0] [15]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(o_dac_b_c_15)) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_q_1__i9.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i8 (.D(\o_val_pipeline_q[0] [14]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(o_dac_b_c_14)) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_q_1__i8.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i7 (.D(\o_val_pipeline_q[0] [13]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(o_dac_b_c_13)) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_q_1__i7.GSR = "DISABLED";
    PFUMX i21180 (.BLUT(n23552), .ALUT(n23553), .C0(index_i[8]), .Z(n23554));
    FD1S3DX o_val_pipeline_q_1__i6 (.D(\o_val_pipeline_q[0] [12]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(o_dac_b_c_12)) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_q_1__i6.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i5 (.D(\o_val_pipeline_q[0] [11]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(o_dac_b_c_11)) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_q_1__i5.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i4 (.D(\o_val_pipeline_q[0] [10]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(o_dac_b_c_10)) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_q_1__i4.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i3 (.D(\o_val_pipeline_q[0] [9]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(n3639)) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_q_1__i3.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i2 (.D(\o_val_pipeline_q[0] [8]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(o_dac_b_c_8)) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_q_1__i2.GSR = "DISABLED";
    FD1P3AX phase_q__i11 (.D(phase_q_11__N_2251[11]), .SP(dac_clk_p_c_enable_488), 
            .CK(dac_clk_p_c), .Q(phase_q[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam phase_q__i11.GSR = "DISABLED";
    LUT4 i11546_2_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n635)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A (B (C+!(D))+!B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11546_2_lut_4_lut_4_lut.init = 16'hf1fc;
    PFUMX i19340 (.BLUT(n21693), .ALUT(n21694), .C0(index_i[4]), .Z(n21695));
    PFUMX i19343 (.BLUT(n21696), .ALUT(n21697), .C0(index_i[4]), .Z(n21698));
    PFUMX i20689 (.BLUT(n23059), .ALUT(n23060), .C0(index_q[8]), .Z(n23063));
    CCU2D add_418_13 (.A0(quarter_wave_sample_register_q[12]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_q[13]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17891), .COUT(n17892), 
          .S0(o_val_pipeline_q_0__15__N_2208[12]), .S1(o_val_pipeline_q_0__15__N_2208[13]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(81[29:60])
    defparam add_418_13.INIT0 = 16'hf555;
    defparam add_418_13.INIT1 = 16'hf555;
    defparam add_418_13.INJECT1_0 = "NO";
    defparam add_418_13.INJECT1_1 = "NO";
    L6MUX21 i20690 (.D0(n23061), .D1(n23062), .SD(index_q[8]), .Z(n23064));
    PFUMX i19712 (.BLUT(n22065), .ALUT(n22066), .C0(index_q[4]), .Z(n476));
    L6MUX21 i20781 (.D0(n23150), .D1(n23151), .SD(index_q[7]), .Z(n23155));
    L6MUX21 i20843 (.D0(n23212), .D1(n23213), .SD(index_q[7]), .Z(n23217));
    CCU2D add_418_11 (.A0(quarter_wave_sample_register_q[10]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_q[11]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17890), .COUT(n17891), 
          .S0(o_val_pipeline_q_0__15__N_2208[10]), .S1(o_val_pipeline_q_0__15__N_2208[11]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(81[29:60])
    defparam add_418_11.INIT0 = 16'hf555;
    defparam add_418_11.INIT1 = 16'hf555;
    defparam add_418_11.INJECT1_0 = "NO";
    defparam add_418_11.INJECT1_1 = "NO";
    LUT4 mux_229_Mux_4_i15_3_lut (.A(n29944), .B(n588), .C(index_i[3]), 
         .Z(n15_adj_2273)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_4_i15_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_4_i348_3_lut (.A(n27350), .B(n27346), .C(index_i[3]), 
         .Z(n348_adj_2274)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_4_i348_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_4_i684_3_lut (.A(n652), .B(n660), .C(index_i[3]), 
         .Z(n684)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_4_i684_3_lut.init = 16'hcaca;
    PFUMX i20897 (.BLUT(n23267), .ALUT(n23268), .C0(index_i[8]), .Z(n23271));
    L6MUX21 i20898 (.D0(n23269), .D1(n23270), .SD(index_i[8]), .Z(n23272));
    PFUMX i21324 (.BLUT(n23690), .ALUT(n23691), .C0(index_q[7]), .Z(n23698));
    PFUMX i25156 (.BLUT(n27474), .ALUT(n27475), .C0(index_i[1]), .Z(n27476));
    FD1P3AX phase_q__i10 (.D(o_phase[9]), .SP(dac_clk_p_c_enable_488), .CK(dac_clk_p_c), 
            .Q(phase_q[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam phase_q__i10.GSR = "DISABLED";
    FD1P3AX phase_q__i9 (.D(o_phase[8]), .SP(dac_clk_p_c_enable_488), .CK(dac_clk_p_c), 
            .Q(phase_q[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam phase_q__i9.GSR = "DISABLED";
    FD1P3AX phase_q__i8 (.D(o_phase[7]), .SP(dac_clk_p_c_enable_488), .CK(dac_clk_p_c), 
            .Q(phase_q[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam phase_q__i8.GSR = "DISABLED";
    FD1P3AX phase_q__i7 (.D(o_phase[6]), .SP(dac_clk_p_c_enable_488), .CK(dac_clk_p_c), 
            .Q(phase_q[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam phase_q__i7.GSR = "DISABLED";
    FD1P3AX phase_q__i6 (.D(o_phase[5]), .SP(dac_clk_p_c_enable_488), .CK(dac_clk_p_c), 
            .Q(phase_q[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam phase_q__i6.GSR = "DISABLED";
    FD1P3AX phase_q__i5 (.D(o_phase[4]), .SP(dac_clk_p_c_enable_488), .CK(dac_clk_p_c), 
            .Q(phase_q[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam phase_q__i5.GSR = "DISABLED";
    PFUMX i21325 (.BLUT(n23692), .ALUT(n23693), .C0(index_q[7]), .Z(n23699));
    FD1P3AX phase_q__i4 (.D(o_phase[3]), .SP(dac_clk_p_c_enable_488), .CK(dac_clk_p_c), 
            .Q(phase_q[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam phase_q__i4.GSR = "DISABLED";
    FD1P3AX phase_q__i3 (.D(o_phase[2]), .SP(dac_clk_p_c_enable_488), .CK(dac_clk_p_c), 
            .Q(phase_q[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam phase_q__i3.GSR = "DISABLED";
    FD1P3AX phase_q__i2 (.D(o_phase[1]), .SP(dac_clk_p_c_enable_488), .CK(dac_clk_p_c), 
            .Q(phase_q[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam phase_q__i2.GSR = "DISABLED";
    CCU2D add_418_9 (.A0(quarter_wave_sample_register_q[8]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_q[9]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17889), .COUT(n17890), 
          .S0(o_val_pipeline_q_0__15__N_2208[8]), .S1(o_val_pipeline_q_0__15__N_2208[9]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(81[29:60])
    defparam add_418_9.INIT0 = 16'hf555;
    defparam add_418_9.INIT1 = 16'hf555;
    defparam add_418_9.INJECT1_0 = "NO";
    defparam add_418_9.INJECT1_1 = "NO";
    LUT4 i20149_3_lut_4_lut_4_lut_4_lut (.A(n27296), .B(index_q[2]), .C(index_q[3]), 
         .D(index_q[4]), .Z(n22504)) /* synthesis lut_function=(A (B)+!A (B (C (D))+!B !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i20149_3_lut_4_lut_4_lut_4_lut.init = 16'hc999;
    PFUMX i25279 (.BLUT(n27673), .ALUT(n27672), .C0(index_q[3]), .Z(n27674));
    PFUMX mux_230_Mux_1_i636 (.BLUT(n620), .ALUT(n635_adj_2275), .C0(index_q[4]), 
          .Z(n636)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    PFUMX i19355 (.BLUT(n21708), .ALUT(n21709), .C0(index_i[4]), .Z(n21710));
    LUT4 n627_bdd_1_lut_2_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n26661)) /* synthesis lut_function=(!(A (C+(D))+!A (B (C+(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n627_bdd_1_lut_2_lut_3_lut_4_lut.init = 16'h010f;
    L6MUX21 i24007 (.D0(n25718), .D1(n25715), .SD(index_q[6]), .Z(n22787));
    PFUMX i25277 (.BLUT(n27669), .ALUT(n27668), .C0(index_q[2]), .Z(n27670));
    PFUMX i21425 (.BLUT(n844), .ALUT(n12112), .C0(index_q[4]), .Z(n23799));
    PFUMX i25221 (.BLUT(n27574), .ALUT(n27575), .C0(index_i[8]), .Z(n27576));
    LUT4 mux_229_Mux_5_i739_rep_591 (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .Z(n27256)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_5_i739_rep_591.init = 16'h6464;
    LUT4 i19953_3_lut_3_lut_4_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n22308)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19953_3_lut_3_lut_4_lut_3_lut_4_lut.init = 16'h11ef;
    LUT4 mux_229_Mux_0_i14_3_lut_rep_721_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27386)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_0_i14_3_lut_rep_721_3_lut.init = 16'he3e3;
    PFUMX i20469 (.BLUT(n22835), .ALUT(n22836), .C0(index_i[7]), .Z(n22843));
    PFUMX i24005 (.BLUT(n25717), .ALUT(n25716), .C0(index_q[5]), .Z(n25718));
    LUT4 i15906_3_lut_3_lut (.A(index_i[0]), .B(index_i[2]), .C(index_i[3]), 
         .Z(n18092)) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i15906_3_lut_3_lut.init = 16'h6a6a;
    LUT4 mux_229_Mux_2_i653_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n653)) /* synthesis lut_function=(A (B (C+!(D))+!B !(D))+!A !(B (C+!(D))+!B !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_2_i653_3_lut_4_lut.init = 16'h94aa;
    LUT4 mux_229_Mux_4_i349_3_lut_4_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[4]), .D(n348_adj_2274), .Z(n349_adj_2276)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_4_i349_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_229_Mux_0_i986_3_lut (.A(n29925), .B(n985), .C(index_i[3]), 
         .Z(n986)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_0_i986_3_lut.init = 16'hcaca;
    PFUMX i20470 (.BLUT(n22837), .ALUT(n22838), .C0(index_i[7]), .Z(n22844));
    LUT4 mux_230_Mux_0_i986_3_lut (.A(n27275), .B(n985_adj_2277), .C(index_q[3]), 
         .Z(n986_adj_2278)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_0_i986_3_lut.init = 16'hcaca;
    PFUMX i19742 (.BLUT(n22095), .ALUT(n22096), .C0(index_q[4]), .Z(n22097));
    LUT4 i12392_2_lut_rep_675 (.A(index_i[2]), .B(index_i[0]), .Z(n27340)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12392_2_lut_rep_675.init = 16'heeee;
    PFUMX i19358 (.BLUT(n21711), .ALUT(n21712), .C0(index_i[4]), .Z(n21713));
    PFUMX i25217 (.BLUT(n27568), .ALUT(n27569), .C0(index_q[1]), .Z(n27570));
    LUT4 mux_230_Mux_0_i971_3_lut (.A(n27277), .B(n29928), .C(index_q[3]), 
         .Z(n971_adj_2279)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_0_i971_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_6_i347_3_lut_4_lut_3_lut_rep_592 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27257)) /* synthesis lut_function=(!(A (B+!(C))+!A ((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_6_i347_3_lut_4_lut_3_lut_rep_592.init = 16'h2424;
    LUT4 mux_229_Mux_5_i851_3_lut_3_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n851)) /* synthesis lut_function=(A ((C)+!B)+!A (B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_5_i851_3_lut_3_lut_4_lut_3_lut.init = 16'he7e7;
    LUT4 i22007_3_lut (.A(n22029), .B(n22030), .C(index_q[4]), .Z(n22031)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22007_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_549_3_lut (.A(index_i[2]), .B(index_i[0]), .C(index_i[1]), 
         .Z(n27214)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_2_lut_rep_549_3_lut.init = 16'hfefe;
    LUT4 i19992_3_lut_4_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n22347)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))+!A (B (C)+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19992_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'hf1e3;
    PFUMX i25154 (.BLUT(n27471), .ALUT(n27472), .C0(index_q[0]), .Z(n27473));
    PFUMX i21445 (.BLUT(n23817), .ALUT(n23818), .C0(index_q[8]), .Z(n23819));
    LUT4 i12403_2_lut_rep_559_3_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .Z(n27224)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12403_2_lut_rep_559_3_lut.init = 16'he0e0;
    LUT4 i11495_2_lut_rep_458_3_lut_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[1]), .Z(n27123)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11495_2_lut_rep_458_3_lut_4_lut.init = 16'hf0e0;
    PFUMX i24003 (.BLUT(n25714), .ALUT(n25713), .C0(index_q[5]), .Z(n25715));
    LUT4 mux_229_Mux_0_i491_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n491)) /* synthesis lut_function=(!(A (B (D)+!B !(C+!(D)))+!A ((C+!(D))+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_0_i491_3_lut_4_lut.init = 16'h24aa;
    LUT4 i19389_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21744)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19389_3_lut_4_lut.init = 16'h64cc;
    L6MUX21 i24001 (.D0(n25711), .D1(n25708), .SD(index_q[5]), .Z(n25712));
    LUT4 mux_230_Mux_6_i332_3_lut_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n332)) /* synthesis lut_function=(!(A (C)+!A !((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_6_i332_3_lut_3_lut.init = 16'h5b5b;
    PFUMX i19361 (.BLUT(n21714), .ALUT(n21715), .C0(index_i[4]), .Z(n21716));
    LUT4 n903_bdd_3_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .Z(n26195)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n903_bdd_3_lut_4_lut_3_lut.init = 16'h6161;
    LUT4 mux_229_Mux_0_i15_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n15_adj_2280)) /* synthesis lut_function=(A (B (D)+!B (C+!(D)))+!A (B (D)+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_0_i15_3_lut_4_lut_4_lut_4_lut.init = 16'hec33;
    PFUMX i23999 (.BLUT(n25710), .ALUT(n25709), .C0(index_q[4]), .Z(n25711));
    LUT4 mux_229_Mux_3_i533_3_lut_rep_770 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27435)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_3_i533_3_lut_rep_770.init = 16'h1c1c;
    L6MUX21 i20580 (.D0(n22949), .D1(n22950), .SD(index_i[7]), .Z(n22954));
    PFUMX i25215 (.BLUT(n27565), .ALUT(n27566), .C0(index_i[2]), .Z(n27567));
    PFUMX i21118 (.BLUT(n23490), .ALUT(n23491), .C0(index_q[8]), .Z(n23492));
    PFUMX i21149 (.BLUT(n23521), .ALUT(n23522), .C0(index_i[8]), .Z(n23523));
    L6MUX21 i20637 (.D0(n23001), .D1(n23002), .SD(index_i[6]), .Z(n23011));
    L6MUX21 i20640 (.D0(n23007), .D1(n23008), .SD(index_i[7]), .Z(n23014));
    PFUMX i15921 (.BLUT(n18105), .ALUT(n18106), .C0(index_q[4]), .Z(n18107));
    LUT4 mux_230_Mux_0_i46_3_lut_4_lut_4_lut_4_lut (.A(index_q[2]), .B(index_q[0]), 
         .C(index_q[1]), .D(index_q[3]), .Z(n46)) /* synthesis lut_function=(A (D)+!A (B+(C+!(D)))) */ ;
    defparam mux_230_Mux_0_i46_3_lut_4_lut_4_lut_4_lut.init = 16'hfe55;
    LUT4 mux_229_Mux_0_i971_3_lut (.A(n29923), .B(n27439), .C(index_i[3]), 
         .Z(n971)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_0_i971_3_lut.init = 16'hcaca;
    LUT4 i19672_3_lut_4_lut (.A(n27296), .B(index_q[2]), .C(index_q[3]), 
         .D(n27238), .Z(n22027)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i19672_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_230_Mux_2_i684_3_lut_4_lut (.A(n27296), .B(index_q[2]), .C(index_q[3]), 
         .D(n27425), .Z(n684_adj_2281)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_2_i684_3_lut_4_lut.init = 16'h6f60;
    PFUMX mux_230_Mux_2_i891 (.BLUT(n875_adj_2282), .ALUT(n890), .C0(index_q[4]), 
          .Z(n891)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    L6MUX21 i20687 (.D0(n23055), .D1(n23056), .SD(index_q[7]), .Z(n23061));
    L6MUX21 i20688 (.D0(n23057), .D1(n23058), .SD(index_q[7]), .Z(n23062));
    LUT4 mux_229_Mux_5_i70_3_lut_4_lut_3_lut_rep_771 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27436)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_5_i70_3_lut_4_lut_3_lut_rep_771.init = 16'h1919;
    LUT4 i23669_else_4_lut (.A(index_q[0]), .B(index_q[4]), .C(index_q[1]), 
         .D(index_q[3]), .Z(n27537)) /* synthesis lut_function=(!(A (B (C)+!B !(C (D)+!C !(D)))+!A (B ((D)+!C)+!B !((D)+!C)))) */ ;
    defparam i23669_else_4_lut.init = 16'h394b;
    PFUMX mux_230_Mux_2_i860 (.BLUT(n844_adj_2283), .ALUT(n859_adj_2284), 
          .C0(index_q[4]), .Z(n860)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    PFUMX i25212 (.BLUT(n27561), .ALUT(n27562), .C0(index_q[8]), .Z(n27563));
    PFUMX i19364 (.BLUT(n21717), .ALUT(n21718), .C0(index_i[4]), .Z(n21719));
    LUT4 i11498_3_lut (.A(index_i[3]), .B(index_i[1]), .C(index_i[0]), 
         .Z(n14095)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11498_3_lut.init = 16'hc8c8;
    PFUMX i23996 (.BLUT(n25707), .ALUT(n25706), .C0(index_q[4]), .Z(n25708));
    L6MUX21 i20716 (.D0(n23082), .D1(n23083), .SD(index_q[7]), .Z(n23090));
    LUT4 mux_230_Mux_5_i954_3_lut_4_lut_4_lut (.A(index_q[2]), .B(index_q[0]), 
         .C(index_q[3]), .D(index_q[1]), .Z(n954_adj_2285)) /* synthesis lut_function=(!(A (C)+!A (B+((D)+!C)))) */ ;
    defparam mux_230_Mux_5_i954_3_lut_4_lut_4_lut.init = 16'h0a1a;
    LUT4 mux_229_Mux_6_i796_3_lut_rep_406_3_lut_3_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n27071)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_6_i796_3_lut_rep_406_3_lut_3_lut_4_lut.init = 16'hfe01;
    L6MUX21 i20717 (.D0(n23084), .D1(n23085), .SD(index_q[7]), .Z(n23091));
    L6MUX21 i21209 (.D0(n23581), .D1(n23582), .SD(index_i[7]), .Z(n23583));
    LUT4 mux_230_Mux_9_i285_3_lut_3_lut_4_lut_4_lut (.A(index_q[2]), .B(index_q[0]), 
         .C(index_q[3]), .D(index_q[1]), .Z(n285)) /* synthesis lut_function=(A (C)+!A !(B+(C+(D)))) */ ;
    defparam mux_230_Mux_9_i285_3_lut_3_lut_4_lut_4_lut.init = 16'ha0a1;
    LUT4 mux_229_Mux_2_i142_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n142_adj_2286)) /* synthesis lut_function=(!(A (B (D)+!B (C (D)+!C !(D)))+!A (B (D)+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_2_i142_3_lut_4_lut_4_lut_4_lut.init = 16'h03ec;
    LUT4 mux_229_Mux_6_i627_3_lut_4_lut_3_lut_rep_773 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27438)) /* synthesis lut_function=(A ((C)+!B)+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_6_i627_3_lut_4_lut_3_lut_rep_773.init = 16'he6e6;
    LUT4 mux_230_Mux_2_i173_3_lut_4_lut_4_lut_4_lut (.A(index_q[2]), .B(index_q[0]), 
         .C(index_q[3]), .D(index_q[1]), .Z(n173)) /* synthesis lut_function=(!(A (C)+!A (B (C+!(D))+!B (C (D)+!C !(D))))) */ ;
    defparam mux_230_Mux_2_i173_3_lut_4_lut_4_lut_4_lut.init = 16'h0f1a;
    LUT4 n699_bdd_4_lut (.A(n27126), .B(index_q[6]), .C(n27166), .D(index_q[5]), 
         .Z(n25776)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C+!(D))+!B (D))) */ ;
    defparam n699_bdd_4_lut.init = 16'hd1cc;
    PFUMX i21002 (.BLUT(n23372), .ALUT(n23373), .C0(index_q[4]), .Z(n23376));
    LUT4 mux_229_Mux_0_i970_3_lut_rep_774 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27439)) /* synthesis lut_function=(!(A (B (C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_0_i970_3_lut_rep_774.init = 16'h7e7e;
    PFUMX i25210 (.BLUT(n27558), .ALUT(n27559), .C0(index_i[1]), .Z(n27560));
    LUT4 mux_229_Mux_6_i691_3_lut_rep_775 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27440)) /* synthesis lut_function=(A (B+!(C))+!A !((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_6_i691_3_lut_rep_775.init = 16'h8e8e;
    L6MUX21 i20776 (.D0(n23140), .D1(n23141), .SD(index_q[6]), .Z(n23150));
    L6MUX21 i20778 (.D0(n23144), .D1(n23145), .SD(index_q[7]), .Z(n23152));
    L6MUX21 i20779 (.D0(n23146), .D1(n23147), .SD(index_q[7]), .Z(n23153));
    L6MUX21 i20810 (.D0(n23177), .D1(n23178), .SD(index_q[7]), .Z(n23184));
    PFUMX i19370 (.BLUT(n21723), .ALUT(n21724), .C0(index_i[4]), .Z(n21725));
    LUT4 i20783_3_lut (.A(n23154), .B(n23155), .C(index_q[8]), .Z(n23157)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20783_3_lut.init = 16'hcaca;
    L6MUX21 i20811 (.D0(n23179), .D1(n23180), .SD(index_q[7]), .Z(n23185));
    PFUMX i20812 (.BLUT(n23181), .ALUT(n23182), .C0(index_q[7]), .Z(n23186));
    PFUMX i25152 (.BLUT(n27467), .ALUT(n27468), .C0(index_i[3]), .Z(n62));
    LUT4 i9469_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n11955)) /* synthesis lut_function=(!(A (B (C)+!B ((D)+!C))+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9469_3_lut_4_lut_4_lut.init = 16'h4969;
    CCU2D add_418_7 (.A0(quarter_wave_sample_register_q[6]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_q[7]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17888), .COUT(n17889), 
          .S1(o_val_pipeline_q_0__15__N_2208[7]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(81[29:60])
    defparam add_418_7.INIT0 = 16'hf555;
    defparam add_418_7.INIT1 = 16'hf555;
    defparam add_418_7.INJECT1_0 = "NO";
    defparam add_418_7.INJECT1_1 = "NO";
    LUT4 n21655_bdd_3_lut_24104 (.A(n29951), .B(n27345), .C(index_i[3]), 
         .Z(n25816)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n21655_bdd_3_lut_24104.init = 16'hcaca;
    LUT4 mux_230_Mux_7_i134_3_lut_3_lut_4_lut_3_lut_rep_799 (.A(index_q[0]), 
         .B(index_q[1]), .C(index_q[2]), .Z(n29926)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B+!(C)))) */ ;
    defparam mux_230_Mux_7_i134_3_lut_3_lut_4_lut_3_lut_rep_799.init = 16'h1818;
    LUT4 i19819_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n22174)) /* synthesis lut_function=(A (C+(D))+!A !(B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i19819_3_lut_4_lut_4_lut.init = 16'haba5;
    LUT4 mux_229_Mux_0_i180_3_lut_4_lut_3_lut_rep_777 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27442)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_0_i180_3_lut_4_lut_3_lut_rep_777.init = 16'h1818;
    L6MUX21 i23393 (.D0(n24994), .D1(n24991), .SD(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_2160[9]));
    LUT4 i19870_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .D(index_q[0]), .Z(n22225)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B (C+!(D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i19870_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h1c18;
    LUT4 i20922_3_lut_3_lut_4_lut (.A(n27218), .B(index_q[3]), .C(n316), 
         .D(index_q[4]), .Z(n23296)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i20922_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 n172_bdd_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .D(index_q[0]), .Z(n26359)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam n172_bdd_3_lut_4_lut_4_lut_4_lut.init = 16'h1e1c;
    LUT4 i11624_3_lut_4_lut (.A(n27218), .B(index_q[3]), .C(n9630), .D(index_q[6]), 
         .Z(n765)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i11624_3_lut_4_lut.init = 16'hffe0;
    LUT4 mux_230_Mux_10_i317_3_lut_3_lut_4_lut (.A(n27218), .B(index_q[3]), 
         .C(n27174), .D(index_q[4]), .Z(n317)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_10_i317_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 mux_230_Mux_7_i747_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), 
         .B(index_q[2]), .C(index_q[3]), .D(index_q[0]), .Z(n747)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))+!A (B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_7_i747_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'he1e3;
    LUT4 n347_bdd_3_lut_24112 (.A(n29952), .B(index_i[3]), .C(n27347), 
         .Z(n25824)) /* synthesis lut_function=(A (B+(C))+!A !(B+!(C))) */ ;
    defparam n347_bdd_3_lut_24112.init = 16'hb8b8;
    LUT4 mux_230_Mux_7_i891_3_lut_4_lut (.A(n27218), .B(index_q[3]), .C(index_q[4]), 
         .D(n890_adj_2287), .Z(n891_adj_2288)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_7_i891_3_lut_4_lut.init = 16'hfe0e;
    LUT4 i20782_3_lut (.A(n23152), .B(n23153), .C(index_q[8]), .Z(n23156)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20782_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_2_i557_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n557_adj_2289)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C+!(D))+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_2_i557_3_lut_3_lut_4_lut.init = 16'h0f18;
    LUT4 i19645_3_lut (.A(n29934), .B(n14_adj_2290), .C(index_q[3]), .Z(n22000)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19645_3_lut.init = 16'hcaca;
    LUT4 i20720_3_lut (.A(n23090), .B(n23091), .C(index_q[8]), .Z(n23094)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20720_3_lut.init = 16'hcaca;
    LUT4 n285_bdd_3_lut (.A(n27387), .B(n29952), .C(index_i[3]), .Z(n25827)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n285_bdd_3_lut.init = 16'hcaca;
    LUT4 n124_bdd_3_lut_4_lut (.A(n27218), .B(index_q[3]), .C(index_q[4]), 
         .D(n93), .Z(n25758)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam n124_bdd_3_lut_4_lut.init = 16'hfe0e;
    LUT4 i19612_3_lut_3_lut_4_lut (.A(n27218), .B(index_q[3]), .C(n93), 
         .D(index_q[4]), .Z(n21967)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i19612_3_lut_3_lut_4_lut.init = 16'h11f0;
    CCU2D add_418_5 (.A0(quarter_wave_sample_register_q[4]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_q[5]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17887), .COUT(n17888));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(81[29:60])
    defparam add_418_5.INIT0 = 16'hf555;
    defparam add_418_5.INIT1 = 16'hf555;
    defparam add_418_5.INJECT1_0 = "NO";
    defparam add_418_5.INJECT1_1 = "NO";
    L6MUX21 i20837 (.D0(n23200), .D1(n23201), .SD(index_q[6]), .Z(n23211));
    LUT4 n498_bdd_3_lut_24119 (.A(n498), .B(n27342), .C(index_i[3]), .Z(n25830)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n498_bdd_3_lut_24119.init = 16'hcaca;
    L6MUX21 i20838 (.D0(n23202), .D1(n23203), .SD(index_q[6]), .Z(n23212));
    LUT4 i19855_3_lut_4_lut_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[0]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n22210)) /* synthesis lut_function=(!(A (B (C)+!B (C+(D)))+!A !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i19855_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'h585f;
    LUT4 n498_bdd_3_lut_24664 (.A(index_i[3]), .B(n29925), .C(n29923), 
         .Z(n25831)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam n498_bdd_3_lut_24664.init = 16'he4e4;
    L6MUX21 i20841 (.D0(n23208), .D1(n23209), .SD(index_q[7]), .Z(n23215));
    LUT4 mux_230_Mux_0_i443_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[0]), .D(index_q[3]), .Z(n443)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C (D))+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_0_i443_3_lut_4_lut_4_lut_4_lut.init = 16'h0ed5;
    LUT4 n526_bdd_3_lut_24981_4_lut_3_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .D(index_q[0]), .Z(n26167)) /* synthesis lut_function=(!(A (B (D)+!B ((D)+!C))+!A !(B (D)+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam n526_bdd_3_lut_24981_4_lut_3_lut_4_lut.init = 16'h55a9;
    LUT4 i19644_3_lut (.A(n29926), .B(n308), .C(index_q[3]), .Z(n21999)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19644_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_3_i348_3_lut (.A(n27389), .B(n27342), .C(index_i[3]), 
         .Z(n348_adj_2291)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_3_i348_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_7_i173_3_lut (.A(n29916), .B(n14_adj_2290), .C(index_q[3]), 
         .Z(n173_adj_2292)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_7_i173_3_lut.init = 16'hcaca;
    LUT4 i20998_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[3]), 
         .C(index_q[2]), .D(index_q[0]), .Z(n23372)) /* synthesis lut_function=(A (B (C (D))+!B (C))+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i20998_3_lut_4_lut_4_lut_4_lut.init = 16'hb434;
    LUT4 i9573_3_lut_4_lut_3_lut_4_lut (.A(index_q[1]), .B(index_q[3]), 
         .C(index_q[2]), .D(index_q[0]), .Z(n541)) /* synthesis lut_function=(A (B (C (D)))+!A !(B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i9573_3_lut_4_lut_3_lut_4_lut.init = 16'h9555;
    LUT4 mux_230_Mux_0_i251_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[0]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n251_adj_2293)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A !(B ((D)+!C)+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_0_i251_3_lut_4_lut_4_lut_4_lut.init = 16'h543c;
    LUT4 i20928_3_lut_3_lut_4_lut (.A(n27220), .B(index_q[3]), .C(n412_adj_2294), 
         .D(index_q[4]), .Z(n23302)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i20928_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 i22938_3_lut (.A(n574_adj_2295), .B(n637), .C(index_i[6]), .Z(n21795)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22938_3_lut.init = 16'hcaca;
    PFUMX mux_230_Mux_3_i763 (.BLUT(n747_adj_2296), .ALUT(n762), .C0(index_q[4]), 
          .Z(n763)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 n803_bdd_3_lut (.A(n27358), .B(n27389), .C(index_i[3]), .Z(n25834)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n803_bdd_3_lut.init = 16'hacac;
    LUT4 i20930_3_lut_4_lut (.A(n27220), .B(index_q[3]), .C(index_q[4]), 
         .D(n27147), .Z(n23304)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i20930_3_lut_4_lut.init = 16'hfe0e;
    LUT4 mux_230_Mux_10_i413_3_lut_3_lut_4_lut (.A(n27220), .B(index_q[3]), 
         .C(n27174), .D(index_q[4]), .Z(n413)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_10_i413_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 mux_230_Mux_1_i908_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[3]), 
         .C(index_q[2]), .D(index_q[0]), .Z(n908_adj_2297)) /* synthesis lut_function=(!(A (B+(C))+!A !(B+(C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_1_i908_3_lut_4_lut_4_lut_4_lut.init = 16'h5647;
    LUT4 mux_230_Mux_3_i828_3_lut_3_lut_4_lut (.A(n27220), .B(index_q[3]), 
         .C(n157_adj_2298), .D(index_q[4]), .Z(n828)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_3_i828_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 n25838_bdd_3_lut (.A(n25838), .B(n157_adj_2299), .C(index_i[4]), 
         .Z(n25839)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n25838_bdd_3_lut.init = 16'hcaca;
    LUT4 i9603_3_lut_4_lut_3_lut_4_lut (.A(index_q[1]), .B(index_q[3]), 
         .C(index_q[4]), .D(index_q[0]), .Z(n444)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A !(((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i9603_3_lut_4_lut_3_lut_4_lut.init = 16'h5595;
    LUT4 i9585_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[0]), 
         .C(index_q[4]), .D(n27317), .Z(n221)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A !(B+(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i9585_3_lut_4_lut_4_lut_4_lut.init = 16'h5556;
    LUT4 i15939_3_lut_4_lut_3_lut_4_lut (.A(index_q[1]), .B(index_q[3]), 
         .C(index_q[2]), .D(index_q[0]), .Z(n18125)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(D))+!A !(B (C+!(D))+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i15939_3_lut_4_lut_3_lut_4_lut.init = 16'h6a55;
    LUT4 mux_230_Mux_0_i1017_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .D(index_q[0]), .Z(n1017_adj_2300)) /* synthesis lut_function=(A (B (C)+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_0_i1017_4_lut_4_lut_4_lut.init = 16'hd7d0;
    LUT4 i12745_1_lut_2_lut_3_lut_4_lut (.A(n27220), .B(index_q[3]), .C(index_q[5]), 
         .D(index_q[4]), .Z(n381)) /* synthesis lut_function=(!(A (C+(D))+!A (B (C+(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i12745_1_lut_2_lut_3_lut_4_lut.init = 16'h010f;
    LUT4 mux_230_Mux_10_i252_3_lut_4_lut_4_lut (.A(n27220), .B(index_q[3]), 
         .C(index_q[4]), .D(n27172), .Z(n252)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B (C (D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_10_i252_3_lut_4_lut_4_lut.init = 16'h3efe;
    LUT4 i19990_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n22345)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A (B (D)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19990_3_lut_4_lut.init = 16'h18cc;
    LUT4 i19388_else_4_lut (.A(index_i[2]), .B(index_i[1]), .C(index_i[4]), 
         .D(index_i[3]), .Z(n27477)) /* synthesis lut_function=(!(A (B (C)+!B (C+(D)))+!A !(B (C (D)+!C !(D))+!B (C+!(D))))) */ ;
    defparam i19388_else_4_lut.init = 16'h581f;
    LUT4 mux_230_Mux_2_i142_3_lut_4_lut_4_lut_4_lut_4_lut (.A(index_q[1]), 
         .B(index_q[2]), .C(index_q[0]), .D(index_q[3]), .Z(n142_adj_2301)) /* synthesis lut_function=(!(A (B)+!A (B (D)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_2_i142_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'h3266;
    LUT4 mux_230_Mux_2_i716_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), 
         .B(index_q[2]), .C(index_q[3]), .D(index_q[0]), .Z(n716_adj_2302)) /* synthesis lut_function=(!(A (B)+!A !(B (C+!(D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_2_i716_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h6367;
    LUT4 i9481_3_lut_3_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[0]), .D(index_i[1]), .Z(n762_adj_2303)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C (D)+!C !(D)))+!A !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9481_3_lut_3_lut_4_lut_4_lut.init = 16'h700f;
    LUT4 mux_230_Mux_0_i781_4_lut_4_lut_4_lut (.A(index_q[2]), .B(index_q[3]), 
         .C(index_q[1]), .D(index_q[0]), .Z(n781)) /* synthesis lut_function=(!(A (B+!((D)+!C))+!A !(B (C)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_0_i781_4_lut_4_lut_4_lut.init = 16'h6252;
    LUT4 mux_230_Mux_8_i506_3_lut_4_lut_3_lut_4_lut (.A(index_q[2]), .B(index_q[3]), 
         .C(index_q[0]), .D(index_q[1]), .Z(n506_adj_2304)) /* synthesis lut_function=(!(A (B+!(C+(D)))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_8_i506_3_lut_4_lut_3_lut_4_lut.init = 16'h6664;
    PFUMX i21003 (.BLUT(n23374), .ALUT(n23375), .C0(index_q[4]), .Z(n23377));
    LUT4 n15000_bdd_3_lut_24608_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n26387)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C (D)+!C !(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n15000_bdd_3_lut_24608_3_lut_4_lut.init = 16'h0fc1;
    LUT4 i19926_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n22281)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)))+!A !(B (C+!(D))+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19926_3_lut_3_lut_4_lut.init = 16'h71cc;
    LUT4 mux_230_Mux_7_i716_3_lut_3_lut_4_lut (.A(index_q[2]), .B(index_q[3]), 
         .C(index_q[0]), .D(index_q[1]), .Z(n716_adj_2305)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A !(B+!(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_7_i716_3_lut_3_lut_4_lut.init = 16'h6445;
    LUT4 mux_230_Mux_0_i604_3_lut_4_lut_4_lut_4_lut (.A(index_q[2]), .B(index_q[0]), 
         .C(index_q[1]), .D(index_q[3]), .Z(n604)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A !(B (D)+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_0_i604_3_lut_4_lut_4_lut_4_lut.init = 16'h5439;
    LUT4 mux_230_Mux_8_i635_3_lut_4_lut_3_lut_4_lut (.A(index_q[2]), .B(index_q[3]), 
         .C(index_q[0]), .D(index_q[1]), .Z(n635_adj_2306)) /* synthesis lut_function=(!(A (B)+!A !(B+(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_8_i635_3_lut_4_lut_3_lut_4_lut.init = 16'h7666;
    LUT4 n250_bdd_3_lut_24977_3_lut_4_lut_4_lut_3_lut_4_lut (.A(index_q[2]), 
         .B(index_q[3]), .C(index_q[0]), .D(index_q[1]), .Z(n26165)) /* synthesis lut_function=(A (B (C (D)))+!A (B+!(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam n250_bdd_3_lut_24977_3_lut_4_lut_4_lut_3_lut_4_lut.init = 16'hc555;
    LUT4 mux_230_Mux_7_i526_3_lut_3_lut_4_lut_4_lut_3_lut_4_lut (.A(index_q[2]), 
         .B(index_q[3]), .C(index_q[0]), .D(index_q[1]), .Z(n526)) /* synthesis lut_function=(A (C (D))+!A !(B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_7_i526_3_lut_3_lut_4_lut_4_lut_3_lut_4_lut.init = 16'hb555;
    LUT4 mux_230_Mux_0_i428_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_q[2]), 
         .B(index_q[0]), .C(index_q[1]), .D(index_q[3]), .Z(n428)) /* synthesis lut_function=(A (B (C+!(D))+!B !((D)+!C))+!A (B (D)+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_0_i428_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hd5a9;
    LUT4 i9477_3_lut_4_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[3]), 
         .C(index_i[4]), .D(index_i[0]), .Z(n444_adj_2307)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A !(((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9477_3_lut_4_lut_3_lut_4_lut.init = 16'h5595;
    L6MUX21 i19430 (.D0(n21783), .D1(n21784), .SD(index_q[7]), .Z(n21785));
    LUT4 n25797_bdd_3_lut (.A(n25797), .B(n25794), .C(index_i[4]), .Z(n21824)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n25797_bdd_3_lut.init = 16'hcaca;
    LUT4 i22253_3_lut (.A(n22026), .B(n22027), .C(index_q[4]), .Z(n22028)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22253_3_lut.init = 16'hcaca;
    CCU2D add_418_3 (.A0(quarter_wave_sample_register_q[2]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_q[3]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17886), .COUT(n17887));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(81[29:60])
    defparam add_418_3.INIT0 = 16'hf555;
    defparam add_418_3.INIT1 = 16'hf555;
    defparam add_418_3.INJECT1_0 = "NO";
    defparam add_418_3.INJECT1_1 = "NO";
    LUT4 i9449_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n541_adj_2308)) /* synthesis lut_function=(A (B (C (D)))+!A !(B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9449_3_lut_4_lut_4_lut_4_lut.init = 16'h9555;
    LUT4 mux_230_Mux_7_i653_3_lut_4_lut (.A(n27296), .B(index_q[2]), .C(index_q[3]), 
         .D(n29936), .Z(n653_adj_2309)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_7_i653_3_lut_4_lut.init = 16'hf606;
    LUT4 i20644_3_lut (.A(n23015), .B(n23016), .C(index_i[8]), .Z(n23018)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20644_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_0_i557_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n557_adj_2310)) /* synthesis lut_function=(A ((D)+!C)+!A !((D)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_0_i557_3_lut_4_lut.init = 16'haa4e;
    CCU2D add_418_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(quarter_wave_sample_register_q[0]), .B1(quarter_wave_sample_register_q[1]), 
          .C1(GND_net), .D1(GND_net), .COUT(n17886));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(81[29:60])
    defparam add_418_1.INIT0 = 16'hF000;
    defparam add_418_1.INIT1 = 16'ha666;
    defparam add_418_1.INJECT1_0 = "NO";
    defparam add_418_1.INJECT1_1 = "NO";
    PFUMX i23391 (.BLUT(n24993), .ALUT(n24992), .C0(index_q[8]), .Z(n24994));
    LUT4 mux_229_Mux_3_i397_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n397_adj_2311)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !(B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_3_i397_3_lut_4_lut_4_lut.init = 16'ha95a;
    LUT4 mux_229_Mux_0_i443_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n443_adj_2312)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(D))+!A (B (D)+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_0_i443_3_lut_4_lut_4_lut_4_lut.init = 16'h32d5;
    LUT4 i20643_3_lut (.A(n23013), .B(n23014), .C(index_i[8]), .Z(n23017)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20643_3_lut.init = 16'hcaca;
    PFUMX i21160 (.BLUT(n844_adj_2313), .ALUT(n11927), .C0(index_i[4]), 
          .Z(n23534));
    LUT4 i9438_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n11924)) /* synthesis lut_function=(A (B (D)+!B !((D)+!C))+!A (((D)+!C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9438_3_lut_4_lut_4_lut_4_lut.init = 16'hdd35;
    LUT4 i9488_3_lut_4_lut_3_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n875_adj_2314)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(D))+!A (B (C+!(D))+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9488_3_lut_4_lut_3_lut_3_lut_4_lut.init = 16'hc07f;
    LUT4 mux_229_Mux_4_i526_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n526_adj_2315)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A !(B ((D)+!C)+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_4_i526_3_lut_3_lut_4_lut.init = 16'h7e0f;
    LUT4 mux_229_Mux_0_i316_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[3]), 
         .C(index_i[2]), .D(index_i[0]), .Z(n316_adj_2316)) /* synthesis lut_function=(!(A (B+(C))+!A !(B+(C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_0_i316_3_lut_4_lut_4_lut_4_lut.init = 16'h5647;
    LUT4 mux_230_Mux_4_i653_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), 
         .B(index_q[2]), .C(index_q[3]), .D(index_q[0]), .Z(n653_adj_2317)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+(D)))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_4_i653_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h9993;
    L6MUX21 i20895 (.D0(n23263), .D1(n23264), .SD(index_i[7]), .Z(n23269));
    LUT4 mux_229_Mux_6_i635_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n635_adj_2318)) /* synthesis lut_function=(A (B (C+(D))+!B !(D))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_6_i635_3_lut_4_lut.init = 16'hcce6;
    LUT4 n205_bdd_3_lut_25101_4_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n26778)) /* synthesis lut_function=(!(A (B (D)+!B ((D)+!C))+!A !(B (D)+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n205_bdd_3_lut_25101_4_lut_3_lut_4_lut.init = 16'h55a9;
    LUT4 mux_229_Mux_0_i251_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n251_adj_2319)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A !(B ((D)+!C)+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_0_i251_3_lut_4_lut_4_lut_4_lut.init = 16'h543c;
    LUT4 i9486_3_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[3]), .C(index_i[0]), 
         .D(index_i[1]), .Z(n844_adj_2320)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9486_3_lut_4_lut_4_lut.init = 16'hf00e;
    LUT4 i9461_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[4]), .D(n27316), .Z(n221_adj_2321)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A !(B+(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9461_3_lut_4_lut_4_lut_4_lut.init = 16'h5556;
    LUT4 i15932_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n18118)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A !((C (D))+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i15932_3_lut_4_lut_4_lut_4_lut.init = 16'h5999;
    LUT4 mux_229_Mux_0_i781_4_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n781_adj_2322)) /* synthesis lut_function=(!(A (B+!((D)+!C))+!A !(B (C)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_0_i781_4_lut_4_lut_4_lut.init = 16'h6252;
    L6MUX21 i20896 (.D0(n23265), .D1(n23266), .SD(index_i[7]), .Z(n23270));
    LUT4 mux_229_Mux_7_i716_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n716_adj_2323)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C+!(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_7_i716_3_lut_3_lut_4_lut.init = 16'h0f81;
    LUT4 mux_229_Mux_0_i428_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[2]), 
         .B(index_i[0]), .C(index_i[1]), .D(index_i[3]), .Z(n428_adj_2324)) /* synthesis lut_function=(A (B (C+!(D))+!B !((D)+!C))+!A (B (D)+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_0_i428_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hd5a9;
    LUT4 mux_230_Mux_6_i844_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n844_adj_2325)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (B (C)+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_6_i844_3_lut_4_lut_4_lut.init = 16'hc1e0;
    LUT4 i19837_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .D(index_q[0]), .Z(n22192)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B (C+(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i19837_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h7c78;
    LUT4 mux_230_Mux_7_i762_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), 
         .B(index_q[2]), .C(index_q[3]), .D(index_q[0]), .Z(n762_adj_2326)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B ((D)+!C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_7_i762_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h3878;
    LUT4 n254_bdd_4_lut_25077 (.A(index_i[5]), .B(index_i[3]), .C(index_i[6]), 
         .D(index_i[4]), .Z(n24843)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;
    defparam n254_bdd_4_lut_25077.init = 16'hf8f0;
    LUT4 n45_bdd_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .D(index_q[0]), .Z(n26094)) /* synthesis lut_function=(A (B (C)+!B ((D)+!C))+!A (B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam n45_bdd_3_lut_4_lut_4_lut_4_lut.init = 16'he7c7;
    LUT4 n78_bdd_3_lut_24820_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .D(index_q[0]), .Z(n26091)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A !((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam n78_bdd_3_lut_24820_4_lut_4_lut_4_lut.init = 16'h7173;
    LUT4 mux_230_Mux_9_i316_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), 
         .B(index_q[2]), .C(index_q[3]), .D(index_q[0]), .Z(n316)) /* synthesis lut_function=(!(A (B (C)+!B !(C+(D)))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_9_i316_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h7e7c;
    LUT4 i19656_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[2]), 
         .C(index_q[3]), .D(index_q[1]), .Z(n22011)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+!(D)))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i19656_3_lut_4_lut_4_lut_4_lut.init = 16'h9399;
    LUT4 mux_230_Mux_5_i475_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[2]), 
         .C(index_q[3]), .D(index_q[1]), .Z(n475)) /* synthesis lut_function=(A (B ((D)+!C))+!A (B (C)+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_5_i475_3_lut_4_lut_4_lut.init = 16'hd949;
    LUT4 mux_230_Mux_1_i684_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n684_adj_2327)) /* synthesis lut_function=(A (B ((D)+!C)+!B !((D)+!C))+!A !(B (C+(D))+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_1_i684_3_lut_4_lut_4_lut.init = 16'h992d;
    L6MUX21 i21326 (.D0(n23694), .D1(n23695), .SD(index_q[7]), .Z(n23700));
    LUT4 i9626_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n12112)) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B ((D)+!C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i9626_3_lut_4_lut_4_lut.init = 16'hcdad;
    PFUMX i19385 (.BLUT(n21738), .ALUT(n21739), .C0(index_i[4]), .Z(n476_adj_2328));
    LUT4 mux_229_Mux_4_i236_3_lut_4_lut_4_lut_3_lut_rep_684_4_lut (.A(index_i[0]), 
         .B(index_i[3]), .C(index_i[1]), .D(index_i[2]), .Z(n27349)) /* synthesis lut_function=(A (B)+!A !(B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_4_i236_3_lut_4_lut_4_lut_3_lut_rep_684_4_lut.init = 16'h999d;
    LUT4 i19350_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21705)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(D))+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19350_3_lut_3_lut_4_lut.init = 16'h3319;
    LUT4 mux_230_Mux_7_i475_3_lut_3_lut_4_lut (.A(n27296), .B(index_q[2]), 
         .C(n29935), .D(index_q[3]), .Z(n475_adj_2329)) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))+!A !(B ((D)+!C)+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_7_i475_3_lut_3_lut_4_lut.init = 16'h99f0;
    LUT4 mux_229_Mux_0_i747_3_lut_4_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[1]), .Z(n747_adj_2330)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C+(D)))+!A !(B ((D)+!C)+!B (C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_0_i747_3_lut_4_lut_3_lut_4_lut.init = 16'h5596;
    LUT4 i19371_3_lut_4_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[3]), 
         .C(index_i[1]), .D(index_i[2]), .Z(n21726)) /* synthesis lut_function=(!(A (B)+!A !(B (C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19371_3_lut_4_lut_3_lut_4_lut.init = 16'h6662;
    L6MUX21 i21372 (.D0(n23740), .D1(n23741), .SD(index_q[7]), .Z(n23746));
    LUT4 i15905_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[1]), .Z(n18091)) /* synthesis lut_function=(A (B (C (D))+!B !(C))+!A (B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i15905_3_lut_4_lut_4_lut_4_lut.init = 16'hd656;
    LUT4 i9441_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n11927)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D))+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9441_3_lut_4_lut_4_lut_4_lut.init = 16'hcadd;
    PFUMX i21373 (.BLUT(n23742), .ALUT(n23743), .C0(index_q[7]), .Z(n23747));
    LUT4 mux_229_Mux_5_i954_3_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[1]), .Z(n954_adj_2331)) /* synthesis lut_function=(!(A (C)+!A (B+((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_5_i954_3_lut_4_lut_4_lut.init = 16'h0a1a;
    LUT4 i19927_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n22282)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19927_3_lut_3_lut_4_lut.init = 16'h0f1c;
    LUT4 n24848_bdd_3_lut (.A(n27576), .B(n24844), .C(index_i[7]), .Z(n24849)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n24848_bdd_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_4_i812_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[4]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n812)) /* synthesis lut_function=(A (B (C+(D)))+!A !(B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_4_i812_3_lut_3_lut_4_lut.init = 16'h9995;
    PFUMX i25150 (.BLUT(n27464), .ALUT(n27465), .C0(index_q[1]), .Z(n27466));
    LUT4 mux_230_Mux_6_i955_3_lut_4_lut (.A(n27219), .B(index_q[3]), .C(index_q[4]), 
         .D(n27074), .Z(n955)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_6_i955_3_lut_4_lut.init = 16'h8f80;
    LUT4 n21786_bdd_3_lut_25074 (.A(n27068), .B(n701), .C(index_q[6]), 
         .Z(n24851)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n21786_bdd_3_lut_25074.init = 16'hacac;
    LUT4 mux_230_Mux_0_i939_4_lut (.A(n14), .B(n27253), .C(index_q[3]), 
         .D(index_q[2]), .Z(n939_adj_2332)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_0_i939_4_lut.init = 16'hfaca;
    LUT4 i20002_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n22357)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(D))+!A (B (D)+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20002_3_lut_4_lut_4_lut_4_lut.init = 16'hd52b;
    LUT4 n22782_bdd_3_lut (.A(n22787), .B(n22788), .C(index_q[7]), .Z(n24854)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n22782_bdd_3_lut.init = 16'hcaca;
    L6MUX21 i19439 (.D0(n21792), .D1(n21793), .SD(index_i[7]), .Z(n21794));
    LUT4 n24854_bdd_3_lut (.A(n24854), .B(n22782), .C(index_q[8]), .Z(n24855)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n24854_bdd_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_5_i252_3_lut_4_lut (.A(index_i[1]), .B(index_i[3]), 
         .C(index_i[0]), .D(index_i[4]), .Z(n252_adj_2333)) /* synthesis lut_function=(A (B (C+(D))+!B (C (D)))+!A !(B (C+(D))+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_5_i252_3_lut_4_lut.init = 16'ha995;
    LUT4 mux_229_Mux_7_i699_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n699)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C+!(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_7_i699_3_lut_4_lut_4_lut.init = 16'hf07e;
    LUT4 mux_229_Mux_6_i890_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[2]), .D(index_i[3]), .Z(n890_adj_2334)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !((D)+!C))+!A !(B ((D)+!C)+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_6_i890_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h7e07;
    LUT4 i19761_4_lut_4_lut_4_lut (.A(n27296), .B(index_q[2]), .C(index_q[4]), 
         .D(index_q[3]), .Z(n22116)) /* synthesis lut_function=(A (B)+!A !(B (C+(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i19761_4_lut_4_lut_4_lut.init = 16'h999c;
    L6MUX21 i20408 (.D0(n22780), .D1(n22781), .SD(index_q[7]), .Z(n22782));
    LUT4 mux_229_Mux_6_i859_3_lut_rep_431_4_lut_4_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[2]), .D(index_i[3]), .Z(n27096)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A (B (C)+!B !((D)+!C))) */ ;
    defparam mux_229_Mux_6_i859_3_lut_rep_431_4_lut_4_lut_4_lut.init = 16'he0f8;
    LUT4 mux_229_Mux_8_i251_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[2]), .D(index_i[3]), .Z(n251_adj_2335)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B (C+!(D))))) */ ;
    defparam mux_229_Mux_8_i251_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h07e0;
    LUT4 i21184_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n23558)) /* synthesis lut_function=(A (B (C+!(D))+!B !((D)+!C))+!A !(B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;
    defparam i21184_3_lut_4_lut_4_lut.init = 16'h81f8;
    PFUMX i21009 (.BLUT(n23379), .ALUT(n23380), .C0(index_q[4]), .Z(n23383));
    LUT4 mux_229_Mux_0_i699_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n699_adj_2336)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (D))+!A (B (C+!(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_0_i699_3_lut_3_lut_4_lut.init = 16'h1c33;
    LUT4 mux_229_Mux_8_i109_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n109)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C+!(D)))+!A (B (C (D)+!C !(D))+!B (C))) */ ;
    defparam mux_229_Mux_8_i109_3_lut_4_lut_4_lut.init = 16'hf83e;
    LUT4 mux_229_Mux_0_i460_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n460)) /* synthesis lut_function=(A (B+(C (D)+!C !(D)))+!A (B (C)+!B (C (D)+!C !(D)))) */ ;
    defparam mux_229_Mux_0_i460_3_lut_4_lut_4_lut.init = 16'hf8cb;
    LUT4 i21182_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n23556)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B (C+!(D)))) */ ;
    defparam i21182_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hf81f;
    LUT4 i20046_3_lut_4_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n22401)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B+(C+(D))))) */ ;
    defparam i20046_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'h2aab;
    LUT4 mux_229_Mux_10_i413_3_lut_4_lut (.A(n27224), .B(index_i[3]), .C(index_i[4]), 
         .D(n27156), .Z(n413_adj_2337)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_10_i413_3_lut_4_lut.init = 16'hf101;
    LUT4 mux_229_Mux_10_i252_3_lut_4_lut_4_lut (.A(n27224), .B(index_i[3]), 
         .C(index_i[4]), .D(n27229), .Z(n252_adj_2338)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B (C (D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_10_i252_3_lut_4_lut_4_lut.init = 16'h3efe;
    LUT4 mux_229_Mux_3_i828_3_lut_3_lut_4_lut (.A(n27224), .B(index_i[3]), 
         .C(n157), .D(index_i[4]), .Z(n828_adj_2339)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_3_i828_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 n172_bdd_2_lut_3_lut_3_lut_4_lut (.A(index_q[2]), .B(index_q[0]), 
         .C(index_q[1]), .D(index_q[3]), .Z(n26358)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B ((D)+!C)))) */ ;
    defparam n172_bdd_2_lut_3_lut_3_lut_4_lut.init = 16'h00fe;
    LUT4 n476_bdd_3_lut_24256 (.A(n476_adj_2328), .B(n25917), .C(index_i[5]), 
         .Z(n25918)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n476_bdd_3_lut_24256.init = 16'hcaca;
    PFUMX i19832 (.BLUT(n22185), .ALUT(n22186), .C0(index_q[4]), .Z(n22187));
    LUT4 i19669_3_lut (.A(n404), .B(n29919), .C(index_q[3]), .Z(n22024)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19669_3_lut.init = 16'hcaca;
    LUT4 i19912_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n22267)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C))+!A (B (C)+!B !((D)+!C))) */ ;
    defparam i19912_3_lut_4_lut_4_lut_4_lut.init = 16'he078;
    LUT4 i20043_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n22398)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C (D)))+!A (B (C+(D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20043_4_lut_4_lut_4_lut.init = 16'h301c;
    LUT4 i12524_1_lut_2_lut_3_lut_4_lut (.A(n27224), .B(index_i[3]), .C(index_i[5]), 
         .D(index_i[4]), .Z(n381_adj_2340)) /* synthesis lut_function=(!(A (C+(D))+!A (B (C+(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12524_1_lut_2_lut_3_lut_4_lut.init = 16'h010f;
    LUT4 mux_229_Mux_8_i15_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n15_adj_2341)) /* synthesis lut_function=(A (B (C)+!B !(C (D)+!C !(D)))+!A !(B ((D)+!C)+!B (C+!(D)))) */ ;
    defparam mux_229_Mux_8_i15_3_lut_4_lut_4_lut.init = 16'h83e0;
    LUT4 i21183_3_lut_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n23557)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C+!(D))+!B !((D)+!C)))) */ ;
    defparam i21183_3_lut_3_lut_4_lut_4_lut.init = 16'h1f81;
    LUT4 index_i_1__bdd_4_lut_25169 (.A(index_i[1]), .B(index_i[0]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n27488)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A !(B ((D)+!C)+!B (D))) */ ;
    defparam index_i_1__bdd_4_lut_25169.init = 16'h8a51;
    LUT4 mux_230_Mux_8_i61_3_lut_rep_432_4_lut_4_lut_4_lut (.A(index_q[0]), 
         .B(index_q[1]), .C(index_q[2]), .D(index_q[3]), .Z(n27097)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A (B (C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_8_i61_3_lut_rep_432_4_lut_4_lut_4_lut.init = 16'he0f8;
    PFUMX i19838 (.BLUT(n22191), .ALUT(n22192), .C0(index_q[4]), .Z(n22193));
    L6MUX21 i20471 (.D0(n22839), .D1(n22840), .SD(index_i[7]), .Z(n22845));
    LUT4 i21000_3_lut_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n23374)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C+!(D))+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i21000_3_lut_3_lut_4_lut_4_lut.init = 16'h1f81;
    L6MUX21 i20486 (.D0(n22854), .D1(n22855), .SD(index_i[7]), .Z(n22860));
    PFUMX i20487 (.BLUT(n22856), .ALUT(n22857), .C0(index_i[7]), .Z(n22861));
    LUT4 i20999_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n23373)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i20999_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hf81f;
    LUT4 mux_230_Mux_8_i251_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), 
         .B(index_q[1]), .C(index_q[2]), .D(index_q[3]), .Z(n251_adj_2342)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_8_i251_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h07e0;
    LUT4 mux_229_Mux_1_i684_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n684_adj_2343)) /* synthesis lut_function=(A (B ((D)+!C)+!B !((D)+!C))+!A !(B (C+(D))+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_1_i684_3_lut_4_lut_4_lut.init = 16'h992d;
    LUT4 i21234_3_lut (.A(n851), .B(n27383), .C(index_i[3]), .Z(n23608)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21234_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_8_i443_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n443_adj_2344)) /* synthesis lut_function=(A (B (C+!(D))+!B !((D)+!C))+!A !(B (D)+!B ((D)+!C))) */ ;
    defparam mux_230_Mux_8_i443_3_lut_4_lut_4_lut.init = 16'h80fc;
    LUT4 mux_230_Mux_0_i379_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n379_adj_2345)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !((D)+!C))+!A !(B ((D)+!C)+!B (D))) */ ;
    defparam mux_230_Mux_0_i379_3_lut_4_lut_4_lut.init = 16'h8079;
    LUT4 mux_229_Mux_8_i443_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n443_adj_2346)) /* synthesis lut_function=(A (B (C+!(D))+!B !((D)+!C))+!A !(B (D)+!B ((D)+!C))) */ ;
    defparam mux_229_Mux_8_i443_3_lut_4_lut_4_lut.init = 16'h80fc;
    LUT4 i21233_3_lut (.A(n652), .B(n27435), .C(index_i[3]), .Z(n23607)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21233_3_lut.init = 16'hcaca;
    LUT4 i20519_3_lut (.A(n22889), .B(n22890), .C(index_i[8]), .Z(n22893)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20519_3_lut.init = 16'hcaca;
    LUT4 i21232_3_lut (.A(n27388), .B(n27440), .C(index_i[3]), .Z(n23606)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21232_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_0_i379_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n379_adj_2347)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !((D)+!C))+!A !(B ((D)+!C)+!B (D))) */ ;
    defparam mux_229_Mux_0_i379_3_lut_4_lut_4_lut.init = 16'h8079;
    LUT4 i21231_3_lut (.A(n27383), .B(n27432), .C(index_i[3]), .Z(n23605)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21231_3_lut.init = 16'hcaca;
    L6MUX21 i20515 (.D0(n22881), .D1(n22882), .SD(index_i[7]), .Z(n22889));
    LUT4 mux_230_Mux_0_i412_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n412_adj_2348)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(D))+!A (B (D)+!B !(C+!(D)))) */ ;
    defparam mux_230_Mux_0_i412_3_lut_4_lut_4_lut.init = 16'hcd2a;
    LUT4 i19887_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n22242)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B+(C+(D))))) */ ;
    defparam i19887_3_lut_4_lut_4_lut_4_lut.init = 16'h2aab;
    LUT4 n25920_bdd_3_lut (.A(n27567), .B(n444_adj_2307), .C(index_i[5]), 
         .Z(n25921)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n25920_bdd_3_lut.init = 16'hcaca;
    LUT4 i21227_3_lut (.A(n27392), .B(n27432), .C(index_i[3]), .Z(n23601)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21227_3_lut.init = 16'hcaca;
    L6MUX21 i20516 (.D0(n22883), .D1(n22884), .SD(index_i[7]), .Z(n22890));
    PFUMX i25204 (.BLUT(n27549), .ALUT(n27550), .C0(index_q[0]), .Z(n27551));
    LUT4 mux_230_Mux_3_i252_3_lut_4_lut (.A(n27219), .B(index_q[3]), .C(index_q[4]), 
         .D(n15350), .Z(n252_adj_2349)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_3_i252_3_lut_4_lut.init = 16'h08f8;
    LUT4 n254_bdd_4_lut_25054 (.A(index_q[5]), .B(index_q[3]), .C(index_q[6]), 
         .D(index_q[4]), .Z(n24876)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;
    defparam n254_bdd_4_lut_25054.init = 16'hf8f0;
    LUT4 mux_230_Mux_0_i890_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n890_adj_2350)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)+!C !(D)))+!A !(B (C)+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_0_i890_3_lut_4_lut_4_lut.init = 16'h70ca;
    LUT4 mux_230_Mux_6_i890_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), 
         .B(index_q[1]), .C(index_q[2]), .D(index_q[3]), .Z(n890_adj_2351)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !((D)+!C))+!A !(B ((D)+!C)+!B (C (D)+!C !(D))))) */ ;
    defparam mux_230_Mux_6_i890_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h7e07;
    LUT4 mux_230_Mux_7_i699_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n699_adj_2352)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (D))) */ ;
    defparam mux_230_Mux_7_i699_3_lut_4_lut_4_lut_4_lut.init = 16'hf70e;
    L6MUX21 i20575 (.D0(n22939), .D1(n22940), .SD(index_i[6]), .Z(n22949));
    LUT4 i21001_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n23375)) /* synthesis lut_function=(A (B (C+!(D))+!B !((D)+!C))+!A !(B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;
    defparam i21001_3_lut_4_lut_4_lut_4_lut.init = 16'h81f8;
    LUT4 i21226_3_lut (.A(n27388), .B(n660), .C(index_i[3]), .Z(n23600)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21226_3_lut.init = 16'hcaca;
    LUT4 i19894_3_lut_4_lut_3_lut (.A(index_q[1]), .B(index_q[3]), .C(index_q[2]), 
         .Z(n22249)) /* synthesis lut_function=(A (B)+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i19894_3_lut_4_lut_3_lut.init = 16'hd9d9;
    LUT4 mux_230_Mux_8_i109_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n109_adj_2353)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C+!(D)))+!A (B (C (D)+!C !(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_8_i109_3_lut_4_lut_4_lut.init = 16'hf83e;
    LUT4 mux_230_Mux_0_i460_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n460_adj_2354)) /* synthesis lut_function=(A (B+(C (D)+!C !(D)))+!A (B (C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_0_i460_3_lut_4_lut_4_lut.init = 16'hf8cb;
    L6MUX21 i20577 (.D0(n22943), .D1(n22944), .SD(index_i[7]), .Z(n22951));
    LUT4 mux_229_Mux_0_i890_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n890_adj_2355)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)+!C !(D)))+!A !(B (C)+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_0_i890_3_lut_4_lut_4_lut.init = 16'h70ca;
    LUT4 mux_229_Mux_0_i604_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n604_adj_2356)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)+!C !(D)))+!A (B (C (D))+!B (C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_0_i604_3_lut_4_lut_4_lut.init = 16'h0e65;
    LUT4 i20089_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n22444)) /* synthesis lut_function=(A (C)+!A !(B (C)+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20089_3_lut_4_lut_4_lut.init = 16'hb4b5;
    LUT4 mux_229_Mux_11_i445_3_lut_4_lut_4_lut_4_lut (.A(index_i[3]), .B(index_i[4]), 
         .C(index_i[5]), .D(n27224), .Z(n445)) /* synthesis lut_function=(!(A (B (C))+!A !(B+(C+(D))))) */ ;
    defparam mux_229_Mux_11_i445_3_lut_4_lut_4_lut_4_lut.init = 16'h7f7e;
    LUT4 i19657_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n22012)) /* synthesis lut_function=(A (C)+!A !(B (C)+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i19657_3_lut_4_lut_4_lut.init = 16'hb4b5;
    LUT4 mux_230_Mux_1_i716_3_lut_4_lut_4_lut (.A(index_q[2]), .B(index_q[0]), 
         .C(index_q[1]), .D(index_q[3]), .Z(n716_adj_2357)) /* synthesis lut_function=(!(A (B (D)+!B !(C))+!A !(B (C (D))+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_1_i716_3_lut_4_lut_4_lut.init = 16'h70a9;
    LUT4 i19666_3_lut (.A(n404), .B(n27271), .C(index_q[3]), .Z(n22021)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19666_3_lut.init = 16'hcaca;
    L6MUX21 i20578 (.D0(n22945), .D1(n22946), .SD(index_i[7]), .Z(n22952));
    L6MUX21 i20609 (.D0(n22976), .D1(n22977), .SD(index_i[7]), .Z(n22983));
    LUT4 n172_bdd_2_lut_3_lut_3_lut_4_lut_adj_77 (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[1]), .D(index_i[3]), .Z(n26484)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n172_bdd_2_lut_3_lut_3_lut_4_lut_adj_77.init = 16'h00fe;
    LUT4 mux_229_Mux_0_i939_4_lut (.A(n588), .B(n27248), .C(index_i[3]), 
         .D(index_i[2]), .Z(n939)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_0_i939_4_lut.init = 16'hfaca;
    LUT4 mux_230_Mux_11_i445_3_lut_4_lut_4_lut_4_lut (.A(index_q[3]), .B(index_q[4]), 
         .C(index_q[5]), .D(n27220), .Z(n445_adj_2358)) /* synthesis lut_function=(!(A (B (C))+!A !(B+(C+(D))))) */ ;
    defparam mux_230_Mux_11_i445_3_lut_4_lut_4_lut_4_lut.init = 16'h7f7e;
    LUT4 mux_230_Mux_5_i252_3_lut_4_lut (.A(index_q[1]), .B(index_q[3]), 
         .C(index_q[0]), .D(index_q[4]), .Z(n252_adj_2359)) /* synthesis lut_function=(A (B (C+(D))+!B (C (D)))+!A !(B (C+(D))+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_5_i252_3_lut_4_lut.init = 16'ha995;
    PFUMX i25148 (.BLUT(n27461), .ALUT(n27462), .C0(index_q[0]), .Z(n27463));
    LUT4 mux_229_Mux_1_i716_3_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[1]), .D(index_i[3]), .Z(n716_adj_2360)) /* synthesis lut_function=(!(A (B (D)+!B !(C))+!A !(B (C (D))+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_1_i716_3_lut_4_lut_4_lut.init = 16'h70a9;
    LUT4 i21225_3_lut (.A(n652), .B(n27440), .C(index_i[3]), .Z(n23599)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21225_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_7_i891_3_lut_4_lut_4_lut (.A(n27229), .B(index_i[3]), 
         .C(n27213), .D(index_i[4]), .Z(n891_adj_2361)) /* synthesis lut_function=(A (B (C+!(D))+!B !((D)+!C))+!A (B (C+!(D))+!B (C+(D)))) */ ;
    defparam mux_229_Mux_7_i891_3_lut_4_lut_4_lut.init = 16'hd1fc;
    L6MUX21 i20610 (.D0(n22978), .D1(n22979), .SD(index_i[7]), .Z(n22984));
    PFUMX i20611 (.BLUT(n22980), .ALUT(n22981), .C0(index_i[7]), .Z(n22985));
    LUT4 n25978_bdd_3_lut (.A(n25978), .B(n476_adj_2328), .C(index_i[5]), 
         .Z(n25979)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n25978_bdd_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_2_i173_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[2]), 
         .B(index_i[0]), .C(index_i[3]), .D(index_i[1]), .Z(n173_adj_2362)) /* synthesis lut_function=(!(A (C)+!A (B (C+!(D))+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_2_i173_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h0f1a;
    LUT4 index_i_6__bdd_4_lut_25255 (.A(index_i[6]), .B(index_i[5]), .C(index_i[1]), 
         .D(index_i[0]), .Z(n27623)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C))+!A (B (C)+!B !(C)))) */ ;
    defparam index_i_6__bdd_4_lut_25255.init = 16'h3cbc;
    PFUMX i21010 (.BLUT(n23381), .ALUT(n23382), .C0(index_q[4]), .Z(n23384));
    LUT4 mux_230_Mux_0_i923_3_lut (.A(n29931), .B(n29935), .C(index_q[3]), 
         .Z(n923)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_0_i923_3_lut.init = 16'hcaca;
    LUT4 n24881_bdd_3_lut (.A(n27563), .B(n24877), .C(index_q[7]), .Z(n24882)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n24881_bdd_3_lut.init = 16'hcaca;
    LUT4 n25982_bdd_3_lut (.A(n27560), .B(n25980), .C(index_i[5]), .Z(n25983)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n25982_bdd_3_lut.init = 16'hcaca;
    LUT4 i21224_3_lut (.A(n27385), .B(n29914), .C(index_i[3]), .Z(n23598)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21224_3_lut.init = 16'hcaca;
    LUT4 n269_bdd_3_lut_24395_4_lut (.A(n27252), .B(index_q[2]), .C(index_q[3]), 
         .D(n27291), .Z(n25516)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam n269_bdd_3_lut_24395_4_lut.init = 16'hf606;
    LUT4 mux_230_Mux_0_i348_3_lut_4_lut (.A(n27252), .B(index_q[2]), .C(index_q[3]), 
         .D(n27425), .Z(n348_adj_2363)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_0_i348_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_230_Mux_6_i205_3_lut_4_lut (.A(n27252), .B(index_q[2]), .C(index_q[3]), 
         .D(n332), .Z(n205)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_6_i205_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_230_Mux_3_i890_3_lut_4_lut (.A(n27252), .B(index_q[2]), .C(index_q[3]), 
         .D(n356), .Z(n890_adj_2364)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_3_i890_3_lut_4_lut.init = 16'h6f60;
    LUT4 i19654_3_lut_4_lut (.A(n27252), .B(index_q[2]), .C(index_q[3]), 
         .D(n29945), .Z(n22009)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i19654_3_lut_4_lut.init = 16'hf606;
    L6MUX21 i20636 (.D0(n22999), .D1(n23000), .SD(index_i[6]), .Z(n23010));
    L6MUX21 i20638 (.D0(n23003), .D1(n23004), .SD(index_i[6]), .Z(n23012));
    LUT4 i19935_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n22290)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A !(B (D)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19935_3_lut_3_lut_4_lut.init = 16'ha955;
    LUT4 mux_229_Mux_2_i262_3_lut_3_lut_rep_787 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29914)) /* synthesis lut_function=(A (B)+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_2_i262_3_lut_3_lut_rep_787.init = 16'h9c9c;
    LUT4 i21220_3_lut (.A(n27432), .B(n27442), .C(index_i[3]), .Z(n23594)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21220_3_lut.init = 16'hcaca;
    LUT4 i21219_3_lut (.A(n1001), .B(n27392), .C(index_i[3]), .Z(n23593)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21219_3_lut.init = 16'hcaca;
    LUT4 i21217_3_lut (.A(n27442), .B(n27385), .C(index_i[3]), .Z(n23591)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21217_3_lut.init = 16'hcaca;
    PFUMX i21016 (.BLUT(n23386), .ALUT(n23387), .C0(index_q[4]), .Z(n23390));
    LUT4 i15903_3_lut (.A(n27257), .B(n29913), .C(index_i[3]), .Z(n18089)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15903_3_lut.init = 16'hcaca;
    LUT4 i15902_3_lut (.A(n29913), .B(n27346), .C(index_i[3]), .Z(n18088)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15902_3_lut.init = 16'hcaca;
    LUT4 i19795_3_lut_4_lut (.A(n27322), .B(index_i[3]), .C(index_i[4]), 
         .D(n635_adj_2365), .Z(n22150)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19795_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_229_Mux_8_i542_3_lut_4_lut (.A(n27322), .B(index_i[3]), .C(index_i[4]), 
         .D(n526_adj_2366), .Z(n542)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_8_i542_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_229_Mux_1_i700_3_lut_4_lut (.A(n27301), .B(index_i[3]), .C(index_i[4]), 
         .D(n684_adj_2343), .Z(n700)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_1_i700_3_lut_4_lut.init = 16'hefe0;
    PFUMX i21017 (.BLUT(n23388), .ALUT(n23389), .C0(index_q[4]), .Z(n23391));
    LUT4 mux_230_Mux_8_i542_3_lut_4_lut (.A(n27334), .B(index_q[3]), .C(index_q[4]), 
         .D(n526_adj_2367), .Z(n542_adj_2368)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_8_i542_3_lut_4_lut.init = 16'h6f60;
    LUT4 i19609_3_lut_4_lut (.A(n27334), .B(index_q[3]), .C(index_q[4]), 
         .D(n635_adj_2306), .Z(n21964)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i19609_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_230_Mux_2_i557_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n557_adj_2369)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C+!(D))+!B (C (D)+!C !(D))))) */ ;
    defparam mux_230_Mux_2_i557_3_lut_3_lut_4_lut.init = 16'h0f18;
    LUT4 i22414_3_lut (.A(n109_adj_2353), .B(n124), .C(index_q[4]), .Z(n21949)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22414_3_lut.init = 16'hcaca;
    PFUMX i21415 (.BLUT(n526_adj_2370), .ALUT(n541_adj_2371), .C0(index_q[4]), 
          .Z(n23789));
    L6MUX21 i20680 (.D0(n22052), .D1(n22112), .SD(index_q[6]), .Z(n23054));
    L6MUX21 i20681 (.D0(n22505), .D1(n22118), .SD(index_q[6]), .Z(n23055));
    LUT4 i21090_3_lut_3_lut_4_lut (.A(n27172), .B(index_q[3]), .C(n93_adj_2372), 
         .D(index_q[4]), .Z(n23464)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i21090_3_lut_3_lut_4_lut.init = 16'hf077;
    L6MUX21 i20682 (.D0(n22121), .D1(n22124), .SD(index_q[6]), .Z(n23056));
    LUT4 i20092_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n22447)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C+(D)))+!A (B (C)+!B !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20092_3_lut_4_lut_4_lut.init = 16'hc95a;
    PFUMX i20683 (.BLUT(n22127), .ALUT(n892), .C0(index_q[6]), .Z(n23057));
    LUT4 i19665_3_lut (.A(n29953), .B(n356), .C(index_q[3]), .Z(n22020)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19665_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_4_i158_3_lut (.A(n142_adj_2373), .B(n157_adj_2374), 
         .C(index_q[4]), .Z(n158_adj_2375)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_4_i158_3_lut.init = 16'hcaca;
    LUT4 i9465_3_lut_4_lut_4_lut (.A(index_i[0]), .B(n29922), .C(index_i[4]), 
         .D(index_i[3]), .Z(n605)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A !(B+(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9465_3_lut_4_lut_4_lut.init = 16'h555c;
    PFUMX i21150 (.BLUT(n526_adj_2376), .ALUT(n541_adj_2377), .C0(index_i[4]), 
          .Z(n23524));
    LUT4 mux_229_Mux_0_i475_3_lut_4_lut (.A(n27263), .B(index_i[1]), .C(index_i[3]), 
         .D(n27229), .Z(n475_adj_2378)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_0_i475_3_lut_4_lut.init = 16'h4f40;
    LUT4 mux_229_Mux_3_i491_3_lut_4_lut (.A(n27263), .B(index_i[1]), .C(index_i[3]), 
         .D(n27389), .Z(n491_adj_2379)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_3_i491_3_lut_4_lut.init = 16'h4f40;
    LUT4 n27298_bdd_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[5]), .Z(n29229)) /* synthesis lut_function=(!(A (B (C (D))+!B (D))+!A (B+!(C (D))))) */ ;
    defparam n27298_bdd_3_lut_4_lut.init = 16'h18aa;
    LUT4 i9475_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[4]), .D(n27316), .Z(n189_adj_2380)) /* synthesis lut_function=(A (B (C (D)))+!A !(B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9475_3_lut_4_lut_4_lut_4_lut.init = 16'h9555;
    LUT4 mux_230_Mux_7_i77_3_lut_3_lut_rep_789 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29916)) /* synthesis lut_function=(A (B)+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_7_i77_3_lut_3_lut_rep_789.init = 16'h9c9c;
    LUT4 i19693_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n22048)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A (B (C (D)+!C !(D))+!B (D))) */ ;
    defparam i19693_3_lut_4_lut.init = 16'hd926;
    PFUMX i25146 (.BLUT(n27458), .ALUT(n27459), .C0(index_q[1]), .Z(n27460));
    LUT4 i20579_3_lut (.A(n22947), .B(n22948), .C(index_i[7]), .Z(n22953)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20579_3_lut.init = 16'hcaca;
    LUT4 i19663_3_lut (.A(n29953), .B(n27271), .C(index_q[3]), .Z(n22018)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19663_3_lut.init = 16'hcaca;
    LUT4 i20574_3_lut (.A(n22937), .B(n22938), .C(index_i[6]), .Z(n22948)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20574_3_lut.init = 16'hcaca;
    LUT4 i20047_3_lut_4_lut (.A(n27434), .B(index_i[2]), .C(index_i[3]), 
         .D(n27342), .Z(n22402)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20047_3_lut_4_lut.init = 16'hdfd0;
    LUT4 mux_230_Mux_3_i859_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n859_adj_2381)) /* synthesis lut_function=(!(A (B (D)+!B !(D))+!A (B (C+(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_3_i859_3_lut_3_lut_4_lut.init = 16'h339c;
    LUT4 mux_229_Mux_9_i285_3_lut_3_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[1]), .Z(n285_adj_2382)) /* synthesis lut_function=(A (C)+!A !(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_9_i285_3_lut_3_lut_4_lut_4_lut.init = 16'ha0a1;
    LUT4 index_i_5__bdd_3_lut_26114 (.A(index_i[5]), .B(n27624), .C(index_i[3]), 
         .Z(n27625)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam index_i_5__bdd_3_lut_26114.init = 16'hcaca;
    LUT4 i19369_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21724)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A (B (C (D)+!C !(D))+!B (D))) */ ;
    defparam i19369_3_lut_4_lut.init = 16'hd926;
    PFUMX i25198 (.BLUT(n27540), .ALUT(n27541), .C0(index_i[0]), .Z(n27542));
    LUT4 mux_230_Mux_4_i525_3_lut_rep_801 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29928)) /* synthesis lut_function=(!(A (B (C))+!A !(B+(C)))) */ ;
    defparam mux_230_Mux_4_i525_3_lut_rep_801.init = 16'h7e7e;
    LUT4 mux_229_Mux_3_i908_3_lut (.A(n27394), .B(n27352), .C(index_i[3]), 
         .Z(n908_adj_2383)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_3_i908_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_4_i526_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n526_adj_2384)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A !(B ((D)+!C)+!B (C (D)+!C !(D))))) */ ;
    defparam mux_230_Mux_4_i526_3_lut_3_lut_4_lut.init = 16'h7e0f;
    LUT4 i19662_3_lut (.A(n356), .B(n332), .C(index_q[3]), .Z(n22017)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19662_3_lut.init = 16'hcaca;
    PFUMX i21023 (.BLUT(n23393), .ALUT(n23394), .C0(index_q[4]), .Z(n23397));
    LUT4 mux_229_Mux_8_i716_3_lut_4_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[1]), .D(index_i[3]), .Z(n716_adj_2385)) /* synthesis lut_function=(!(A (D)+!A !(B+(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_8_i716_3_lut_4_lut_4_lut_4_lut.init = 16'h55fe;
    PFUMX i21416 (.BLUT(n557_adj_2386), .ALUT(n572), .C0(index_q[4]), 
          .Z(n23790));
    LUT4 i20170_3_lut (.A(n900), .B(n356), .C(index_q[3]), .Z(n22525)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20170_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_6_i645_3_lut_4_lut_3_lut_rep_802 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29929)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B))) */ ;
    defparam mux_230_Mux_6_i645_3_lut_4_lut_3_lut_rep_802.init = 16'h1919;
    LUT4 i19674_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n22029)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(D))+!A (B))) */ ;
    defparam i19674_3_lut_3_lut_4_lut.init = 16'h3319;
    L6MUX21 i20708 (.D0(n23066), .D1(n23067), .SD(index_q[6]), .Z(n23082));
    L6MUX21 i20709 (.D0(n23068), .D1(n23069), .SD(index_q[6]), .Z(n23083));
    L6MUX21 i20710 (.D0(n23070), .D1(n23071), .SD(index_q[6]), .Z(n23084));
    L6MUX21 i20711 (.D0(n23072), .D1(n23073), .SD(index_q[6]), .Z(n23085));
    L6MUX21 i20712 (.D0(n23074), .D1(n23075), .SD(index_q[6]), .Z(n23086));
    L6MUX21 i20714 (.D0(n23078), .D1(n23079), .SD(index_q[6]), .Z(n23088));
    PFUMX i21207 (.BLUT(n23577), .ALUT(n23578), .C0(index_i[6]), .Z(n23581));
    LUT4 n70_bdd_4_lut (.A(n29936), .B(n173_adj_2387), .C(index_q[4]), 
         .D(index_q[3]), .Z(n25150)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D)))) */ ;
    defparam n70_bdd_4_lut.init = 16'hcacc;
    LUT4 i12397_3_lut (.A(index_i[2]), .B(index_i[1]), .C(index_i[0]), 
         .Z(n1001)) /* synthesis lut_function=(A (B)+!A (B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12397_3_lut.init = 16'hdcdc;
    LUT4 i6479_2_lut (.A(phase_q[0]), .B(phase_i[10]), .Z(index_i_9__N_2125[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(60[14] 63[8])
    defparam i6479_2_lut.init = 16'h6666;
    L6MUX21 i20739 (.D0(n23097), .D1(n23098), .SD(index_q[6]), .Z(n23113));
    L6MUX21 i23940 (.D0(n25649), .D1(n27052), .SD(index_i[6]), .Z(n638));
    L6MUX21 i20740 (.D0(n23099), .D1(n23100), .SD(index_q[6]), .Z(n23114));
    PFUMX i21024 (.BLUT(n23395), .ALUT(n23396), .C0(index_q[4]), .Z(n23398));
    L6MUX21 i20741 (.D0(n23101), .D1(n23102), .SD(index_q[6]), .Z(n23115));
    LUT4 i22941_2_lut (.A(phase_q[0]), .B(phase_i[10]), .Z(index_q_9__N_2135[0])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(60[14] 63[8])
    defparam i22941_2_lut.init = 16'h9999;
    PFUMX i23938 (.BLUT(n25648), .ALUT(n25647), .C0(index_i[5]), .Z(n25649));
    PFUMX i21417 (.BLUT(n589), .ALUT(n604), .C0(index_q[4]), .Z(n23791));
    LUT4 mux_229_Mux_0_i46_3_lut_4_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[1]), .D(index_i[3]), .Z(n46_adj_2388)) /* synthesis lut_function=(A (D)+!A (B+(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_0_i46_3_lut_4_lut_4_lut_4_lut.init = 16'hfe55;
    PFUMX i20743 (.BLUT(n23105), .ALUT(n23106), .C0(index_q[6]), .Z(n23117));
    LUT4 i20899_3_lut (.A(n23271), .B(n23272), .C(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2145[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20899_3_lut.init = 16'hcaca;
    L6MUX21 i20744 (.D0(n23107), .D1(n23108), .SD(index_q[6]), .Z(n23118));
    PFUMX i21208 (.BLUT(n23579), .ALUT(n23580), .C0(index_i[6]), .Z(n23582));
    LUT4 i20475_3_lut (.A(n22847), .B(n22848), .C(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2145[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20475_3_lut.init = 16'hcaca;
    LUT4 i20474_3_lut (.A(n22845), .B(n22846), .C(index_i[8]), .Z(n22848)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20474_3_lut.init = 16'hcaca;
    LUT4 i20713_3_lut (.A(n23076), .B(n23077), .C(index_q[6]), .Z(n23087)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20713_3_lut.init = 16'hcaca;
    LUT4 i20809_3_lut (.A(n25417), .B(n23176), .C(index_q[7]), .Z(n23183)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20809_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_1_i700_3_lut_4_lut (.A(n27305), .B(index_q[3]), .C(index_q[4]), 
         .D(n684_adj_2327), .Z(n700_adj_2389)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_1_i700_3_lut_4_lut.init = 16'hefe0;
    PFUMX i21418 (.BLUT(n620_adj_2390), .ALUT(n635_adj_2391), .C0(index_q[4]), 
          .Z(n23792));
    L6MUX21 i20745 (.D0(n23109), .D1(n23110), .SD(index_q[6]), .Z(n23119));
    LUT4 i7209_2_lut (.A(index_q[4]), .B(index_q[5]), .Z(n9630)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i7209_2_lut.init = 16'h8888;
    PFUMX i20746 (.BLUT(n23111), .ALUT(n23112), .C0(index_q[6]), .Z(n23120));
    LUT4 mux_230_Mux_8_i763_3_lut_4_lut (.A(n27293), .B(n27307), .C(index_q[4]), 
         .D(n27166), .Z(n15348)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam mux_230_Mux_8_i763_3_lut_4_lut.init = 16'hfe0e;
    L6MUX21 i23918 (.D0(n25630), .D1(n25627), .SD(index_i[4]), .Z(n509));
    PFUMX i23916 (.BLUT(n25629), .ALUT(n25628), .C0(index_i[5]), .Z(n25630));
    LUT4 mux_230_Mux_7_i404_3_lut_rep_804 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29931)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C)+!B !(C))) */ ;
    defparam mux_230_Mux_7_i404_3_lut_rep_804.init = 16'he3e3;
    LUT4 mux_230_Mux_7_i541_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n541_adj_2392)) /* synthesis lut_function=(A (B (C)+!B ((D)+!C))+!A (B (C)+!B !(C))) */ ;
    defparam mux_230_Mux_7_i541_3_lut_4_lut_4_lut.init = 16'he3c3;
    LUT4 n45_bdd_3_lut_24361_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n26093)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C (D)+!C !(D))+!B (C)))) */ ;
    defparam n45_bdd_3_lut_24361_3_lut_4_lut.init = 16'h0fc1;
    PFUMX i23914 (.BLUT(n25626), .ALUT(n25625), .C0(index_i[6]), .Z(n25627));
    PFUMX i25196 (.BLUT(n27537), .ALUT(n27538), .C0(index_q[2]), .Z(n27539));
    LUT4 n300_bdd_3_lut_24403 (.A(n27291), .B(n27277), .C(index_q[3]), 
         .Z(n26119)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n300_bdd_3_lut_24403.init = 16'hcaca;
    LUT4 index_i_0__bdd_4_lut_26060 (.A(index_i[0]), .B(index_i[3]), .C(index_i[1]), 
         .D(index_i[2]), .Z(n27494)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C))+!A (B (C (D)+!C !(D))+!B !(C+!(D))))) */ ;
    defparam index_i_0__bdd_4_lut_26060.init = 16'h16d3;
    LUT4 n476_bdd_3_lut_24573_3_lut (.A(index_q[1]), .B(index_q[4]), .C(n124_adj_2393), 
         .Z(n25411)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam n476_bdd_3_lut_24573_3_lut.init = 16'hd1d1;
    LUT4 mux_230_Mux_7_i243_3_lut_rep_807 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29934)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B (C)+!B !(C)))) */ ;
    defparam mux_230_Mux_7_i243_3_lut_rep_807.init = 16'h1c1c;
    LUT4 mux_230_Mux_0_i699_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n699_adj_2394)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (D))+!A (B (C+!(D))+!B !(C+!(D))))) */ ;
    defparam mux_230_Mux_0_i699_3_lut_3_lut_4_lut.init = 16'h1c33;
    LUT4 i21089_3_lut_4_lut (.A(n27172), .B(index_q[3]), .C(index_q[4]), 
         .D(n46), .Z(n23463)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i21089_3_lut_4_lut.init = 16'h8f80;
    LUT4 n22105_bdd_3_lut_3_lut (.A(index_q[1]), .B(n526_adj_2395), .C(index_q[4]), 
         .Z(n25413)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam n22105_bdd_3_lut_3_lut.init = 16'h5c5c;
    LUT4 i19735_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n22090)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B (C (D)+!C !(D))))) */ ;
    defparam i19735_3_lut_3_lut_4_lut.init = 16'h0f1c;
    LUT4 n442_bdd_3_lut_24409 (.A(n27274), .B(n29958), .C(index_q[3]), 
         .Z(n26128)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n442_bdd_3_lut_24409.init = 16'hcaca;
    LUT4 i19884_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n22239)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C (D)))+!A (B (C+(D))+!B !(C)))) */ ;
    defparam i19884_4_lut_4_lut_4_lut.init = 16'h301c;
    LUT4 i8246_2_lut (.A(index_i[4]), .B(index_i[5]), .Z(n10667)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i8246_2_lut.init = 16'h8888;
    LUT4 mux_230_Mux_7_i123_3_lut_3_lut_3_lut_rep_808 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29935)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (B+!(C))) */ ;
    defparam mux_230_Mux_7_i123_3_lut_3_lut_3_lut_rep_808.init = 16'hc7c7;
    PFUMX i20766 (.BLUT(n797), .ALUT(n828), .C0(index_q[5]), .Z(n23140));
    LUT4 n300_bdd_3_lut_24999 (.A(n27291), .B(n14), .C(index_q[3]), .Z(n26130)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n300_bdd_3_lut_24999.init = 16'hacac;
    LUT4 n26983_bdd_3_lut_3_lut (.A(n1021), .B(index_i[8]), .C(n26983), 
         .Z(n26984)) /* synthesis lut_function=(A (B+(C))+!A !(B+!(C))) */ ;
    defparam n26983_bdd_3_lut_3_lut.init = 16'hb8b8;
    PFUMX i21419 (.BLUT(n653_adj_2396), .ALUT(n668_adj_2397), .C0(index_q[4]), 
          .Z(n23793));
    L6MUX21 i20770 (.D0(n23128), .D1(n23129), .SD(index_q[6]), .Z(n23144));
    L6MUX21 i20771 (.D0(n23130), .D1(n23131), .SD(index_q[6]), .Z(n23145));
    L6MUX21 i20772 (.D0(n23132), .D1(n23133), .SD(index_q[6]), .Z(n23146));
    L6MUX21 i20773 (.D0(n23134), .D1(n23135), .SD(index_q[6]), .Z(n23147));
    L6MUX21 i20774 (.D0(n23136), .D1(n23137), .SD(index_q[6]), .Z(n23148));
    L6MUX21 i20777 (.D0(n23142), .D1(n23143), .SD(index_q[6]), .Z(n23151));
    LUT4 n27294_bdd_3_lut_26323_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n28896)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C))+!A (B (C (D))+!B (C)))) */ ;
    defparam n27294_bdd_3_lut_26323_4_lut.init = 16'h0fc7;
    PFUMX mux_230_Mux_5_i732 (.BLUT(n12079), .ALUT(n731), .C0(index_q[4]), 
          .Z(n732)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 i19396_3_lut (.A(n27387), .B(n356_adj_2398), .C(index_i[3]), 
         .Z(n21751)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19396_3_lut.init = 16'hcaca;
    L6MUX21 i20802 (.D0(n23161), .D1(n23162), .SD(index_q[6]), .Z(n23176));
    L6MUX21 i20803 (.D0(n23163), .D1(n23164), .SD(index_q[6]), .Z(n23177));
    L6MUX21 i20804 (.D0(n23165), .D1(n23166), .SD(index_q[6]), .Z(n23178));
    L6MUX21 i20805 (.D0(n23167), .D1(n23168), .SD(index_q[6]), .Z(n23179));
    L6MUX21 i20806 (.D0(n23169), .D1(n23170), .SD(index_q[6]), .Z(n23180));
    LUT4 i22065_3_lut (.A(n21750), .B(n21751), .C(index_i[4]), .Z(n21752)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22065_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_8_i172_rep_809 (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .Z(n29936)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B+(C)))) */ ;
    defparam mux_230_Mux_8_i172_rep_809.init = 16'h7c7c;
    PFUMX i21420 (.BLUT(n684_adj_2399), .ALUT(n699_adj_2394), .C0(index_q[4]), 
          .Z(n23794));
    LUT4 mux_230_Mux_0_i475_3_lut_4_lut (.A(n27267), .B(index_q[1]), .C(index_q[3]), 
         .D(n27172), .Z(n475_adj_2400)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_0_i475_3_lut_4_lut.init = 16'h4f40;
    LUT4 mux_230_Mux_3_i491_3_lut_4_lut (.A(n27267), .B(index_q[1]), .C(index_q[3]), 
         .D(n27426), .Z(n491_adj_2401)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_3_i491_3_lut_4_lut.init = 16'h4f40;
    PFUMX i20827 (.BLUT(n732_adj_2402), .ALUT(n763_adj_2403), .C0(index_q[5]), 
          .Z(n23201));
    LUT4 n124_bdd_3_lut_24070_4_lut (.A(n27381), .B(index_i[3]), .C(index_i[4]), 
         .D(n124_adj_2404), .Z(n25781)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n124_bdd_3_lut_24070_4_lut.init = 16'hf101;
    L6MUX21 i20829 (.D0(n22244), .D1(n891_adj_2405), .SD(index_q[5]), 
            .Z(n23203));
    LUT4 mux_230_Mux_8_i124_3_lut_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n124)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C+!(D)))+!A (B (C (D)+!C !(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_8_i124_3_lut_3_lut_4_lut_4_lut.init = 16'h07c1;
    L6MUX21 i20832 (.D0(n23190), .D1(n23191), .SD(index_q[6]), .Z(n23206));
    L6MUX21 i20834 (.D0(n23194), .D1(n23195), .SD(index_q[6]), .Z(n23208));
    L6MUX21 i20835 (.D0(n23196), .D1(n23197), .SD(index_q[6]), .Z(n23209));
    LUT4 i20942_3_lut_4_lut (.A(n27381), .B(index_i[3]), .C(index_i[4]), 
         .D(n285_adj_2382), .Z(n23316)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20942_3_lut_4_lut.init = 16'hfe0e;
    LUT4 mux_229_Mux_2_i573_3_lut_3_lut_4_lut (.A(n27381), .B(index_i[3]), 
         .C(n557_adj_2289), .D(index_i[4]), .Z(n573)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_2_i573_3_lut_3_lut_4_lut.init = 16'h11f0;
    L6MUX21 i20839 (.D0(n23204), .D1(n23205), .SD(index_q[6]), .Z(n23213));
    PFUMX i21421 (.BLUT(n716_adj_2406), .ALUT(n731_adj_2407), .C0(index_q[4]), 
          .Z(n23795));
    LUT4 index_q_0__bdd_4_lut (.A(index_q[0]), .B(index_q[3]), .C(index_q[1]), 
         .D(index_q[2]), .Z(n29959)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C (D)))+!A !(B (C+!(D))+!B !(C+(D))))) */ ;
    defparam index_q_0__bdd_4_lut.init = 16'h4ae7;
    LUT4 mux_230_Mux_5_i109_3_lut_4_lut_3_lut (.A(index_q[1]), .B(index_q[3]), 
         .C(index_q[0]), .Z(n109_adj_2408)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_5_i109_3_lut_4_lut_3_lut.init = 16'h6565;
    LUT4 mux_229_Mux_4_i573_3_lut_3_lut_4_lut_4_lut (.A(n27381), .B(index_i[3]), 
         .C(index_i[4]), .D(n27224), .Z(n573_adj_2409)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_4_i573_3_lut_3_lut_4_lut_4_lut.init = 16'h1f1c;
    LUT4 index_q_4__bdd_4_lut_24239 (.A(index_q[4]), .B(n27195), .C(index_q[7]), 
         .D(n27179), .Z(n25198)) /* synthesis lut_function=(A (C+!(D))+!A (B+!(C))) */ ;
    defparam index_q_4__bdd_4_lut_24239.init = 16'he5ef;
    LUT4 mux_229_Mux_3_i573_3_lut_3_lut_4_lut (.A(n27381), .B(index_i[3]), 
         .C(n397_adj_2410), .D(index_i[4]), .Z(n573_adj_2411)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_3_i573_3_lut_3_lut_4_lut.init = 16'h11f0;
    PFUMX i19850 (.BLUT(n22203), .ALUT(n22204), .C0(index_q[4]), .Z(n22205));
    LUT4 mux_229_Mux_10_i125_3_lut_4_lut_4_lut (.A(n27381), .B(index_i[3]), 
         .C(index_i[4]), .D(n27229), .Z(n125)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B (C (D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_10_i125_3_lut_4_lut_4_lut.init = 16'h3efe;
    LUT4 quarter_wave_sample_register_i_15__I_0_3_lut (.A(\quarter_wave_sample_register_q[15] ), 
         .B(o_val_pipeline_i_0__15__N_2176[15]), .C(phase_negation_i[1]), 
         .Z(o_val_pipeline_i_0__15__N_2175)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(76[14] 78[8])
    defparam quarter_wave_sample_register_i_15__I_0_3_lut.init = 16'hcaca;
    LUT4 quarter_wave_sample_register_i_14__I_0_3_lut (.A(quarter_wave_sample_register_i[14]), 
         .B(o_val_pipeline_i_0__15__N_2176[14]), .C(phase_negation_i[1]), 
         .Z(o_val_pipeline_i_0__15__N_2177)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(76[14] 78[8])
    defparam quarter_wave_sample_register_i_14__I_0_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_7_i14_3_lut_4_lut_3_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[0]), .Z(n14_adj_2290)) /* synthesis lut_function=(!(A ((C)+!B)+!A !((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_7_i14_3_lut_4_lut_3_lut.init = 16'h5959;
    LUT4 quarter_wave_sample_register_i_13__I_0_3_lut (.A(quarter_wave_sample_register_i[13]), 
         .B(o_val_pipeline_i_0__15__N_2176[13]), .C(phase_negation_i[1]), 
         .Z(o_val_pipeline_i_0__15__N_2179)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(76[14] 78[8])
    defparam quarter_wave_sample_register_i_13__I_0_3_lut.init = 16'hcaca;
    LUT4 quarter_wave_sample_register_i_12__I_0_3_lut (.A(quarter_wave_sample_register_i[12]), 
         .B(o_val_pipeline_i_0__15__N_2176[12]), .C(phase_negation_i[1]), 
         .Z(o_val_pipeline_i_0__15__N_2181)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(76[14] 78[8])
    defparam quarter_wave_sample_register_i_12__I_0_3_lut.init = 16'hcaca;
    LUT4 quarter_wave_sample_register_i_11__I_0_3_lut (.A(quarter_wave_sample_register_i[11]), 
         .B(o_val_pipeline_i_0__15__N_2176[11]), .C(phase_negation_i[1]), 
         .Z(o_val_pipeline_i_0__15__N_2183)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(76[14] 78[8])
    defparam quarter_wave_sample_register_i_11__I_0_3_lut.init = 16'hcaca;
    LUT4 n53_bdd_3_lut_23995_4_lut (.A(n27269), .B(index_q[2]), .C(n29941), 
         .D(index_q[3]), .Z(n25706)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam n53_bdd_3_lut_23995_4_lut.init = 16'hf066;
    LUT4 mux_230_Mux_3_i668_3_lut_4_lut (.A(n27269), .B(index_q[2]), .C(index_q[3]), 
         .D(n29953), .Z(n668_adj_2412)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_3_i668_3_lut_4_lut.init = 16'h6f60;
    LUT4 quarter_wave_sample_register_i_10__I_0_3_lut (.A(quarter_wave_sample_register_i[10]), 
         .B(o_val_pipeline_i_0__15__N_2176[10]), .C(phase_negation_i[1]), 
         .Z(o_val_pipeline_i_0__15__N_2185)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(76[14] 78[8])
    defparam quarter_wave_sample_register_i_10__I_0_3_lut.init = 16'hcaca;
    L6MUX21 i20885 (.D0(n23597), .D1(n23604), .SD(index_i[6]), .Z(n23259));
    LUT4 mux_230_Mux_0_i762_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n762_adj_2413)) /* synthesis lut_function=(A (B+!((D)+!C))+!A !(B (D)+!B !(C))) */ ;
    defparam mux_230_Mux_0_i762_3_lut_4_lut_4_lut.init = 16'h98fc;
    L6MUX21 i20888 (.D0(n22172), .D1(n22181), .SD(index_i[6]), .Z(n23262));
    LUT4 quarter_wave_sample_register_i_9__I_0_3_lut (.A(quarter_wave_sample_register_i[9]), 
         .B(o_val_pipeline_i_0__15__N_2176[9]), .C(phase_negation_i[1]), 
         .Z(o_val_pipeline_i_0__15__N_2187)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(76[14] 78[8])
    defparam quarter_wave_sample_register_i_9__I_0_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_4_i763_3_lut_4_lut (.A(n27269), .B(index_q[2]), .C(index_q[4]), 
         .D(n747_adj_2414), .Z(n763_adj_2415)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_4_i763_3_lut_4_lut.init = 16'h6f60;
    LUT4 quarter_wave_sample_register_i_8__I_0_3_lut (.A(quarter_wave_sample_register_i[8]), 
         .B(o_val_pipeline_i_0__15__N_2176[8]), .C(phase_negation_i[1]), 
         .Z(o_val_pipeline_i_0__15__N_2189)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(76[14] 78[8])
    defparam quarter_wave_sample_register_i_8__I_0_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_3_i396_3_lut_3_lut_rep_791 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29918)) /* synthesis lut_function=(A (B+(C))+!A !(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_3_i396_3_lut_3_lut_rep_791.init = 16'ha9a9;
    L6MUX21 i20889 (.D0(n22190), .D1(n22199), .SD(index_i[6]), .Z(n23263));
    LUT4 quarter_wave_sample_register_i_7__I_0_3_lut (.A(quarter_wave_sample_register_i[7]), 
         .B(o_val_pipeline_i_0__15__N_2176[7]), .C(phase_negation_i[1]), 
         .Z(o_val_pipeline_i_0__15__N_2191)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(76[14] 78[8])
    defparam quarter_wave_sample_register_i_7__I_0_3_lut.init = 16'hcaca;
    L6MUX21 i20890 (.D0(n22208), .D1(n22217), .SD(index_i[6]), .Z(n23264));
    LUT4 mux_230_Mux_6_i420_3_lut_4_lut_3_lut_rep_811 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29938)) /* synthesis lut_function=(A (B+!(C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_6_i420_3_lut_4_lut_3_lut_rep_811.init = 16'hdbdb;
    PFUMX i20891 (.BLUT(n22220), .ALUT(n892_adj_2416), .C0(index_i[6]), 
          .Z(n23265));
    LUT4 i21094_3_lut_4_lut (.A(n27172), .B(index_q[3]), .C(index_q[4]), 
         .D(n220), .Z(n23468)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i21094_3_lut_4_lut.init = 16'hf808;
    PFUMX i21422 (.BLUT(n747_adj_2417), .ALUT(n762_adj_2413), .C0(index_q[4]), 
          .Z(n23796));
    LUT4 n250_bdd_3_lut_24438 (.A(n29945), .B(n27277), .C(index_q[3]), 
         .Z(n26164)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n250_bdd_3_lut_24438.init = 16'hacac;
    LUT4 n890_bdd_3_lut_23913_4_lut (.A(n27429), .B(n27302), .C(index_i[5]), 
         .D(n27316), .Z(n25625)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;
    defparam n890_bdd_3_lut_23913_4_lut.init = 16'hf101;
    LUT4 mux_229_Mux_8_i763_3_lut_4_lut (.A(n27429), .B(n27302), .C(index_i[4]), 
         .D(n27159), .Z(n15218)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam mux_229_Mux_8_i763_3_lut_4_lut.init = 16'hfe0e;
    LUT4 mux_229_Mux_2_i189_3_lut_3_lut_4_lut (.A(index_i[1]), .B(n27316), 
         .C(n173_adj_2362), .D(index_i[4]), .Z(n189_adj_2418)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(C+(D)))) */ ;
    defparam mux_229_Mux_2_i189_3_lut_3_lut_4_lut.init = 16'h77f0;
    LUT4 i11895_2_lut_3_lut_4_lut (.A(index_i[1]), .B(n27316), .C(index_i[5]), 
         .D(index_i[4]), .Z(n508)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;
    defparam i11895_2_lut_3_lut_4_lut.init = 16'hf080;
    LUT4 mux_229_Mux_11_i638_4_lut_4_lut (.A(n27086), .B(index_i[5]), .C(index_i[6]), 
         .D(n27120), .Z(n638_adj_2419)) /* synthesis lut_function=(A (B (C (D))+!B !(C))+!A (B ((D)+!C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_11_i638_4_lut_4_lut.init = 16'hc707;
    LUT4 i11605_3_lut_4_lut (.A(n27064), .B(index_q[7]), .C(index_q[8]), 
         .D(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_2160[14])) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i11605_3_lut_4_lut.init = 16'hffe0;
    LUT4 mux_229_Mux_1_i924_3_lut (.A(n316_adj_2316), .B(n27382), .C(index_i[4]), 
         .Z(n924)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_1_i924_3_lut.init = 16'hcaca;
    LUT4 index_i_1__bdd_4_lut_25170 (.A(index_i[1]), .B(index_i[3]), .C(index_i[2]), 
         .D(index_i[0]), .Z(n27498)) /* synthesis lut_function=(!(A (B (C (D))+!B (C+!(D)))+!A !(B (C (D)+!C !(D))+!B ((D)+!C)))) */ ;
    defparam index_i_1__bdd_4_lut_25170.init = 16'h5b8d;
    L6MUX21 i21320 (.D0(n23682), .D1(n23683), .SD(index_q[6]), .Z(n23694));
    LUT4 i20512_3_lut (.A(n22875), .B(n22876), .C(index_i[6]), .Z(n22886)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20512_3_lut.init = 16'hcaca;
    LUT4 i21945_3_lut (.A(n22389), .B(n22390), .C(index_i[4]), .Z(n22391)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21945_3_lut.init = 16'hcaca;
    LUT4 n284_bdd_3_lut_24881 (.A(n27297), .B(n27288), .C(index_q[3]), 
         .Z(n26173)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n284_bdd_3_lut_24881.init = 16'hcaca;
    L6MUX21 i21321 (.D0(n23684), .D1(n23685), .SD(index_q[6]), .Z(n23695));
    L6MUX21 i21322 (.D0(n23686), .D1(n23687), .SD(index_q[6]), .Z(n23696));
    PFUMX i21323 (.BLUT(n23688), .ALUT(n23689), .C0(index_q[6]), .Z(n23697));
    LUT4 i1_2_lut (.A(index_q[6]), .B(index_q[7]), .Z(n20112)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i21949_3_lut (.A(n29964), .B(n22381), .C(index_i[4]), .Z(n22382)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21949_3_lut.init = 16'hcaca;
    LUT4 index_i_4__bdd_4_lut_24281 (.A(index_i[4]), .B(n27185), .C(index_i[7]), 
         .D(n27165), .Z(n25220)) /* synthesis lut_function=(A (C+!(D))+!A (B+!(C))) */ ;
    defparam index_i_4__bdd_4_lut_24281.init = 16'he5ef;
    PFUMX i21423 (.BLUT(n781), .ALUT(n796), .C0(index_q[4]), .Z(n23797));
    LUT4 i20691_3_lut (.A(n23063), .B(n23064), .C(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_2160[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20691_3_lut.init = 16'hcaca;
    LUT4 i21330_3_lut (.A(n23702), .B(n23703), .C(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_2160[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21330_3_lut.init = 16'hcaca;
    LUT4 i21329_3_lut (.A(n23700), .B(n23701), .C(index_q[8]), .Z(n23703)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21329_3_lut.init = 16'hcaca;
    LUT4 i22943_2_lut (.A(phase_q[9]), .B(phase_i[10]), .Z(index_q_9__N_2135[9])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(60[14] 63[8])
    defparam i22943_2_lut.init = 16'h9999;
    LUT4 i22945_2_lut (.A(phase_q[8]), .B(phase_i[10]), .Z(index_q_9__N_2135[8])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(60[14] 63[8])
    defparam i22945_2_lut.init = 16'h9999;
    LUT4 i20608_3_lut (.A(n25984), .B(n22975), .C(index_i[7]), .Z(n22982)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20608_3_lut.init = 16'hcaca;
    LUT4 i22947_2_lut (.A(phase_q[7]), .B(phase_i[10]), .Z(index_q_9__N_2135[7])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(60[14] 63[8])
    defparam i22947_2_lut.init = 16'h9999;
    PFUMX i19856 (.BLUT(n22209), .ALUT(n22210), .C0(index_q[4]), .Z(n22211));
    LUT4 mux_229_Mux_1_i349_3_lut (.A(n541_adj_2420), .B(n348_adj_2421), 
         .C(index_i[4]), .Z(n349_adj_2422)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_1_i349_3_lut.init = 16'hcaca;
    LUT4 i22949_2_lut (.A(phase_q[6]), .B(phase_i[10]), .Z(index_q_9__N_2135[6])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(60[14] 63[8])
    defparam i22949_2_lut.init = 16'h9999;
    LUT4 i21955_3_lut (.A(n22353), .B(n22354), .C(index_i[4]), .Z(n22355)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21955_3_lut.init = 16'hcaca;
    LUT4 i22951_2_lut (.A(phase_q[5]), .B(phase_i[10]), .Z(index_q_9__N_2135[5])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(60[14] 63[8])
    defparam i22951_2_lut.init = 16'h9999;
    PFUMX i21424 (.BLUT(n812_adj_2423), .ALUT(n12109), .C0(index_q[4]), 
          .Z(n23798));
    LUT4 mux_230_Mux_0_i364_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n364_adj_2424)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A ((C+!(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_0_i364_3_lut_3_lut_4_lut.init = 16'hdb55;
    L6MUX21 i20927 (.D0(n23299), .D1(n23300), .SD(index_q[6]), .Z(n23301));
    PFUMX i19859 (.BLUT(n22212), .ALUT(n22213), .C0(index_q[4]), .Z(n22214));
    LUT4 i22953_2_lut (.A(phase_q[4]), .B(phase_i[10]), .Z(index_q_9__N_2135[4])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(60[14] 63[8])
    defparam i22953_2_lut.init = 16'h9999;
    LUT4 i22955_2_lut (.A(phase_q[3]), .B(phase_i[10]), .Z(index_q_9__N_2135[3])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(60[14] 63[8])
    defparam i22955_2_lut.init = 16'h9999;
    LUT4 mux_230_Mux_14_i511_4_lut_4_lut (.A(n27064), .B(index_q[7]), .C(index_q[8]), 
         .D(n254), .Z(n511_adj_2272)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (B (C+!(D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_14_i511_4_lut_4_lut.init = 16'h1c10;
    LUT4 i22957_2_lut (.A(phase_q[2]), .B(phase_i[10]), .Z(index_q_9__N_2135[2])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(60[14] 63[8])
    defparam i22957_2_lut.init = 16'h9999;
    LUT4 i11874_3_lut_4_lut (.A(n27066), .B(index_i[7]), .C(index_i[8]), 
         .D(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2145[14])) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11874_3_lut_4_lut.init = 16'hffe0;
    PFUMX i21426 (.BLUT(n875_adj_2425), .ALUT(n890_adj_2350), .C0(index_q[4]), 
          .Z(n23800));
    LUT4 i22959_2_lut (.A(phase_q[1]), .B(phase_i[10]), .Z(index_q_9__N_2135[1])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(60[14] 63[8])
    defparam i22959_2_lut.init = 16'h9999;
    LUT4 i6501_2_lut (.A(phase_q[9]), .B(phase_i[10]), .Z(index_i_9__N_2125[9])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(60[14] 63[8])
    defparam i6501_2_lut.init = 16'h6666;
    LUT4 i6502_2_lut (.A(phase_q[8]), .B(phase_i[10]), .Z(index_i_9__N_2125[8])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(60[14] 63[8])
    defparam i6502_2_lut.init = 16'h6666;
    L6MUX21 i20934 (.D0(n23306), .D1(n23307), .SD(index_q[6]), .Z(n23308));
    LUT4 i19840_3_lut_4_lut (.A(index_q[0]), .B(n27334), .C(index_q[3]), 
         .D(n29941), .Z(n22195)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i19840_3_lut_4_lut.init = 16'hfb0b;
    PFUMX i19871 (.BLUT(n22224), .ALUT(n22225), .C0(index_q[4]), .Z(n22226));
    LUT4 i6503_2_lut (.A(phase_q[7]), .B(phase_i[10]), .Z(index_i_9__N_2125[7])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(60[14] 63[8])
    defparam i6503_2_lut.init = 16'h6666;
    LUT4 i6504_2_lut (.A(phase_q[6]), .B(phase_i[10]), .Z(index_i_9__N_2125[6])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(60[14] 63[8])
    defparam i6504_2_lut.init = 16'h6666;
    LUT4 i6505_2_lut (.A(phase_q[5]), .B(phase_i[10]), .Z(index_i_9__N_2125[5])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(60[14] 63[8])
    defparam i6505_2_lut.init = 16'h6666;
    LUT4 i6506_2_lut (.A(phase_q[4]), .B(phase_i[10]), .Z(index_i_9__N_2125[4])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(60[14] 63[8])
    defparam i6506_2_lut.init = 16'h6666;
    LUT4 i6507_2_lut (.A(phase_q[3]), .B(phase_i[10]), .Z(index_i_9__N_2125[3])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(60[14] 63[8])
    defparam i6507_2_lut.init = 16'h6666;
    LUT4 i6508_2_lut (.A(phase_q[2]), .B(phase_i[10]), .Z(index_i_9__N_2125[2])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(60[14] 63[8])
    defparam i6508_2_lut.init = 16'h6666;
    LUT4 i6509_2_lut (.A(phase_q[1]), .B(phase_i[10]), .Z(index_i_9__N_2125[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(60[14] 63[8])
    defparam i6509_2_lut.init = 16'h6666;
    LUT4 mux_458_i9_3_lut (.A(\quarter_wave_sample_register_q[15] ), .B(o_val_pipeline_q_0__15__N_2208[15]), 
         .C(phase_negation_q[1]), .Z(n1790[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(81[29:60])
    defparam mux_458_i9_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_1_i94_3_lut (.A(index_i[0]), .B(n93_adj_2426), .C(index_i[4]), 
         .Z(n94)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_1_i94_3_lut.init = 16'hcaca;
    LUT4 mux_458_i8_3_lut (.A(quarter_wave_sample_register_q[14]), .B(o_val_pipeline_q_0__15__N_2208[14]), 
         .C(phase_negation_q[1]), .Z(n1790[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(81[29:60])
    defparam mux_458_i8_3_lut.init = 16'hcaca;
    LUT4 mux_458_i7_3_lut (.A(quarter_wave_sample_register_q[13]), .B(o_val_pipeline_q_0__15__N_2208[13]), 
         .C(phase_negation_q[1]), .Z(n1790[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(81[29:60])
    defparam mux_458_i7_3_lut.init = 16'hcaca;
    LUT4 mux_458_i6_3_lut (.A(quarter_wave_sample_register_q[12]), .B(o_val_pipeline_q_0__15__N_2208[12]), 
         .C(phase_negation_q[1]), .Z(n1790[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(81[29:60])
    defparam mux_458_i6_3_lut.init = 16'hcaca;
    LUT4 mux_458_i5_3_lut (.A(quarter_wave_sample_register_q[11]), .B(o_val_pipeline_q_0__15__N_2208[11]), 
         .C(phase_negation_q[1]), .Z(n1790[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(81[29:60])
    defparam mux_458_i5_3_lut.init = 16'hcaca;
    LUT4 mux_458_i4_3_lut (.A(quarter_wave_sample_register_q[10]), .B(o_val_pipeline_q_0__15__N_2208[10]), 
         .C(phase_negation_q[1]), .Z(n1790[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(81[29:60])
    defparam mux_458_i4_3_lut.init = 16'hcaca;
    LUT4 mux_458_i3_3_lut (.A(quarter_wave_sample_register_q[9]), .B(o_val_pipeline_q_0__15__N_2208[9]), 
         .C(phase_negation_q[1]), .Z(n1790[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(81[29:60])
    defparam mux_458_i3_3_lut.init = 16'hcaca;
    PFUMX i21427 (.BLUT(n908), .ALUT(n923), .C0(index_q[4]), .Z(n23801));
    LUT4 mux_458_i2_3_lut (.A(quarter_wave_sample_register_q[8]), .B(o_val_pipeline_q_0__15__N_2208[8]), 
         .C(phase_negation_q[1]), .Z(n1790[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(81[29:60])
    defparam mux_458_i2_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_11_i638_4_lut_4_lut (.A(n27087), .B(index_q[5]), .C(index_q[6]), 
         .D(n27116), .Z(n638_adj_2427)) /* synthesis lut_function=(A (B (C (D))+!B !(C))+!A (B ((D)+!C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_11_i638_4_lut_4_lut.init = 16'hc707;
    PFUMX i21363 (.BLUT(n12043), .ALUT(n21953), .C0(index_q[6]), .Z(n23737));
    LUT4 mux_458_i1_3_lut (.A(quarter_wave_sample_register_q[7]), .B(o_val_pipeline_q_0__15__N_2208[7]), 
         .C(phase_negation_q[1]), .Z(n1790[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(81[29:60])
    defparam mux_458_i1_3_lut.init = 16'hcaca;
    PFUMX i21428 (.BLUT(n939_adj_2332), .ALUT(n954_adj_2428), .C0(index_q[4]), 
          .Z(n23802));
    LUT4 mux_229_Mux_14_i511_4_lut_4_lut (.A(n27066), .B(index_i[7]), .C(index_i[8]), 
         .D(n254_adj_2429), .Z(n511)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (B (C+!(D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_14_i511_4_lut_4_lut.init = 16'h1c10;
    L6MUX21 i21365 (.D0(n21959), .D1(n21962), .SD(index_q[6]), .Z(n23739));
    L6MUX21 i20948 (.D0(n23320), .D1(n23321), .SD(index_i[6]), .Z(n382));
    L6MUX21 i21366 (.D0(n574_adj_2430), .D1(n21965), .SD(index_q[6]), 
            .Z(n23740));
    L6MUX21 i21367 (.D0(n21968), .D1(n764), .SD(index_q[6]), .Z(n23741));
    LUT4 i1_3_lut_4_lut_adj_78 (.A(n27087), .B(index_q[5]), .C(index_q[8]), 
         .D(n20112), .Z(n20536)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i1_3_lut_4_lut_adj_78.init = 16'hfff8;
    LUT4 i1_3_lut_4_lut_adj_79 (.A(n27434), .B(n27316), .C(index_i[4]), 
         .D(n27320), .Z(n20603)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;
    defparam i1_3_lut_4_lut_adj_79.init = 16'hfff8;
    PFUMX i20494 (.BLUT(n221_adj_2321), .ALUT(n252_adj_2333), .C0(index_i[5]), 
          .Z(n22868));
    PFUMX i21429 (.BLUT(n971_adj_2279), .ALUT(n986_adj_2278), .C0(index_q[4]), 
          .Z(n23803));
    PFUMX i25144 (.BLUT(n27455), .ALUT(n27456), .C0(index_q[3]), .Z(n62_adj_2269));
    PFUMX i21430 (.BLUT(n1002_adj_2431), .ALUT(n1017_adj_2300), .C0(index_q[4]), 
          .Z(n23804));
    LUT4 mux_230_Mux_3_i221_3_lut_4_lut (.A(n27172), .B(index_q[3]), .C(index_q[4]), 
         .D(n27195), .Z(n221_adj_2432)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_3_i221_3_lut_4_lut.init = 16'h08f8;
    LUT4 i11770_3_lut_3_lut (.A(index_q[1]), .B(index_q[0]), .C(index_q[2]), 
         .Z(n619)) /* synthesis lut_function=(!(A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i11770_3_lut_3_lut.init = 16'h7575;
    LUT4 n939_bdd_4_lut (.A(n939_adj_2433), .B(n27430), .C(index_i[4]), 
         .D(index_i[3]), .Z(n25264)) /* synthesis lut_function=(A (B+(C+!(D)))+!A !((C+!(D))+!B)) */ ;
    defparam n939_bdd_4_lut.init = 16'hacaa;
    PFUMX i19877 (.BLUT(n22230), .ALUT(n22231), .C0(index_q[4]), .Z(n22232));
    LUT4 i1_2_lut_adj_80 (.A(o_phase[11]), .B(o_phase[10]), .Z(phase_q_11__N_2251[11])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i1_2_lut_adj_80.init = 16'h9999;
    LUT4 mux_229_Mux_4_i747_3_lut_4_lut (.A(n27248), .B(index_i[2]), .C(index_i[3]), 
         .D(n27387), .Z(n747_adj_2434)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_4_i747_3_lut_4_lut.init = 16'hf606;
    PFUMX i20406 (.BLUT(n22776), .ALUT(n22777), .C0(index_q[6]), .Z(n22780));
    LUT4 i19740_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n22095)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A !(B (D)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i19740_3_lut_3_lut_4_lut.init = 16'ha955;
    PFUMX i19883 (.BLUT(n22236), .ALUT(n22237), .C0(index_q[4]), .Z(n22238));
    LUT4 mux_229_Mux_6_i157_3_lut_4_lut (.A(n27248), .B(index_i[2]), .C(index_i[3]), 
         .D(n27348), .Z(n157_adj_2299)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_6_i157_3_lut_4_lut.init = 16'hf606;
    LUT4 i9463_3_lut_4_lut (.A(n27248), .B(index_i[2]), .C(n27321), .D(n27347), 
         .Z(n444_adj_2435)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9463_3_lut_4_lut.init = 16'h6f60;
    PFUMX i20407 (.BLUT(n22778), .ALUT(n22779), .C0(index_q[6]), .Z(n22781));
    LUT4 mux_229_Mux_6_i251_3_lut_4_lut (.A(n27248), .B(index_i[2]), .C(index_i[3]), 
         .D(n27347), .Z(n251)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_6_i251_3_lut_4_lut.init = 16'hf606;
    PFUMX i19886 (.BLUT(n22239), .ALUT(n22240), .C0(index_q[4]), .Z(n22241));
    LUT4 mux_230_Mux_6_i38_3_lut_3_lut_rep_813 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29940)) /* synthesis lut_function=(A (B+(C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_6_i38_3_lut_3_lut_rep_813.init = 16'hadad;
    LUT4 index_i_1__bdd_4_lut_26242 (.A(index_i[1]), .B(index_i[0]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n27499)) /* synthesis lut_function=(!(A (B (D)+!B (C+!(D)))+!A !(B (C (D)+!C !(D))+!B !((D)+!C)))) */ ;
    defparam index_i_1__bdd_4_lut_26242.init = 16'h429c;
    LUT4 i21126_3_lut (.A(n236), .B(n251_adj_2319), .C(index_i[4]), .Z(n23500)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21126_3_lut.init = 16'hcaca;
    LUT4 n123_bdd_3_lut_24101_4_lut (.A(n27255), .B(index_i[2]), .C(n27353), 
         .D(index_i[3]), .Z(n25813)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n123_bdd_3_lut_24101_4_lut.init = 16'hf066;
    LUT4 i11843_2_lut_rep_587 (.A(index_q[0]), .B(index_q[1]), .Z(n27252)) /* synthesis lut_function=(A+!(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i11843_2_lut_rep_587.init = 16'hbbbb;
    LUT4 mux_229_Mux_3_i668_3_lut_4_lut (.A(n27255), .B(index_i[2]), .C(index_i[3]), 
         .D(n27346), .Z(n668_adj_2436)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_3_i668_3_lut_4_lut.init = 16'h6f60;
    PFUMX i19889 (.BLUT(n22242), .ALUT(n22243), .C0(index_q[4]), .Z(n22244));
    LUT4 mux_230_Mux_3_i397_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n397_adj_2437)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !(B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_3_i397_3_lut_4_lut_4_lut.init = 16'ha95a;
    L6MUX21 i21362 (.D0(n21947), .D1(n21950), .SD(index_q[6]), .Z(n23736));
    LUT4 mux_229_Mux_4_i763_3_lut_4_lut (.A(n27255), .B(index_i[2]), .C(index_i[4]), 
         .D(n747_adj_2434), .Z(n763_adj_2438)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_4_i763_3_lut_4_lut.init = 16'h6f60;
    LUT4 i11916_3_lut_4_lut (.A(index_i[4]), .B(n27316), .C(index_i[5]), 
         .D(n27434), .Z(n892_adj_2439)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11916_3_lut_4_lut.init = 16'hf8f0;
    LUT4 mux_230_Mux_0_i796_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n796)) /* synthesis lut_function=(A (B (C+(D))+!B (C (D)))+!A !(B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_0_i796_3_lut_4_lut_4_lut.init = 16'hadc0;
    LUT4 i21119_3_lut (.A(n15_adj_2280), .B(n27488), .C(index_i[4]), .Z(n23493)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21119_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_6_i505_3_lut_rep_792 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29919)) /* synthesis lut_function=(A (B)+!A (B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_6_i505_3_lut_rep_792.init = 16'hc9c9;
    PFUMX i20414 (.BLUT(n22785), .ALUT(n22786), .C0(index_q[6]), .Z(n22788));
    LUT4 i19891_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n22246)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C+(D)))+!A (B (C)+!B !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i19891_3_lut_4_lut_4_lut.init = 16'hc95a;
    LUT4 mux_229_Mux_2_i308_3_lut_4_lut_3_lut_rep_784 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29911)) /* synthesis lut_function=(A (B (C))+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_2_i308_3_lut_4_lut_3_lut_rep_784.init = 16'h9494;
    LUT4 n53_bdd_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n25707)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam n53_bdd_3_lut_4_lut_4_lut.init = 16'ha5ad;
    LUT4 mux_230_Mux_6_i7_3_lut_4_lut_3_lut_rep_814 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29941)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_6_i7_3_lut_4_lut_3_lut_rep_814.init = 16'hd6d6;
    LUT4 index_q_0__bdd_4_lut_25636 (.A(index_q[0]), .B(index_q[3]), .C(index_q[1]), 
         .D(index_q[2]), .Z(n27500)) /* synthesis lut_function=(A (B (C)+!B !(C+!(D)))+!A !(B ((D)+!C)+!B !(C (D)+!C !(D)))) */ ;
    defparam index_q_0__bdd_4_lut_25636.init = 16'h92c1;
    LUT4 i19954_3_lut_4_lut (.A(n27434), .B(index_i[2]), .C(index_i[3]), 
         .D(n851), .Z(n22309)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19954_3_lut_4_lut.init = 16'hf202;
    LUT4 i20678_3_lut (.A(n190), .B(n26535), .C(index_q[6]), .Z(n23052)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20678_3_lut.init = 16'hcaca;
    LUT4 i12126_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[4]), 
         .C(n27317), .D(index_q[0]), .Z(n14724)) /* synthesis lut_function=(!(A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i12126_3_lut_4_lut_4_lut_4_lut.init = 16'h55d5;
    LUT4 i19597_3_lut_then_4_lut (.A(index_q[4]), .B(index_q[2]), .C(index_q[3]), 
         .D(index_q[0]), .Z(n27502)) /* synthesis lut_function=(!(A (B (C)+!B ((D)+!C))+!A !((C)+!B))) */ ;
    defparam i19597_3_lut_then_4_lut.init = 16'h5979;
    LUT4 i20679_3_lut (.A(n23399), .B(n21971), .C(index_q[6]), .Z(n23053)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20679_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_0_i731_3_lut_4_lut (.A(n27429), .B(index_i[2]), .C(index_i[3]), 
         .D(n27435), .Z(n731_adj_2440)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_0_i731_3_lut_4_lut.init = 16'h4f40;
    LUT4 i20044_3_lut_4_lut (.A(n27429), .B(index_i[2]), .C(index_i[3]), 
         .D(n29925), .Z(n22399)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20044_3_lut_4_lut.init = 16'hf404;
    LUT4 n251_bdd_4_lut_26461 (.A(n251_adj_2441), .B(n11265), .C(index_q[2]), 
         .D(index_q[4]), .Z(n26219)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C+(D)))+!A !(B (C+(D))+!B ((D)+!C))) */ ;
    defparam n251_bdd_4_lut_26461.init = 16'haa3c;
    LUT4 i12500_3_lut (.A(index_q[2]), .B(index_q[1]), .C(index_q[0]), 
         .Z(n38)) /* synthesis lut_function=(A (B)+!A (B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i12500_3_lut.init = 16'hdcdc;
    LUT4 i21982_3_lut (.A(n716), .B(n731_adj_2442), .C(index_i[4]), .Z(n732_adj_2443)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21982_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_2_i669_3_lut (.A(n653), .B(n25833), .C(index_i[4]), 
         .Z(n669)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_2_i669_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_2_i605_3_lut (.A(n142_adj_2444), .B(n604_adj_2445), 
         .C(index_i[4]), .Z(n605_adj_2446)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_2_i605_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_2_i700_3_lut_4_lut (.A(index_i[1]), .B(n27302), .C(index_i[4]), 
         .D(n684_adj_2447), .Z(n700_adj_2448)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam mux_229_Mux_2_i700_3_lut_4_lut.init = 16'hefe0;
    LUT4 i21987_3_lut (.A(n27498), .B(n22327), .C(index_i[4]), .Z(n22328)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21987_3_lut.init = 16'hcaca;
    LUT4 i21989_3_lut (.A(n22320), .B(n22321), .C(index_i[4]), .Z(n22322)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21989_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_2_i413_3_lut (.A(n397_adj_2449), .B(n954_adj_2331), 
         .C(index_i[4]), .Z(n413_adj_2450)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_2_i413_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_2_i317_3_lut (.A(n668_adj_2436), .B(n316_adj_2451), 
         .C(index_i[4]), .Z(n317_adj_2452)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_2_i317_3_lut.init = 16'hcaca;
    L6MUX21 i23890 (.D0(n25601), .D1(n27053), .SD(index_q[6]), .Z(n23315));
    LUT4 mux_229_Mux_2_i286_3_lut (.A(n270_adj_2453), .B(n653_adj_2454), 
         .C(index_i[4]), .Z(n286_adj_2455)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_2_i286_3_lut.init = 16'hcaca;
    LUT4 n954_bdd_4_lut (.A(n27123), .B(index_i[4]), .C(n25644), .D(index_i[5]), 
         .Z(n27052)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (B (C (D))+!B (C+!(D)))) */ ;
    defparam n954_bdd_4_lut.init = 16'hf099;
    LUT4 mux_229_Mux_5_i31_3_lut (.A(n15), .B(n30), .C(index_i[4]), .Z(n31)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_5_i31_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_3_i1018_3_lut_4_lut (.A(index_i[1]), .B(n27302), .C(index_i[4]), 
         .D(n20166), .Z(n1018)) /* synthesis lut_function=(A (C+!(D))+!A (B (C+!(D))+!B !(C+(D)))) */ ;
    defparam mux_229_Mux_3_i1018_3_lut_4_lut.init = 16'he0ef;
    LUT4 i20886_3_lut (.A(n190_adj_2456), .B(n253), .C(index_i[6]), .Z(n23260)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20886_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_4_i62_4_lut (.A(n29924), .B(n61), .C(index_i[4]), 
         .D(index_i[3]), .Z(n62_adj_2457)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_4_i62_4_lut.init = 16'hc5ca;
    LUT4 mux_229_Mux_4_i31_4_lut (.A(n15_adj_2273), .B(n27098), .C(index_i[4]), 
         .D(index_i[3]), .Z(n31_adj_2458)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_4_i31_4_lut.init = 16'h3aca;
    LUT4 i20887_3_lut (.A(n23611), .B(n22160), .C(index_i[6]), .Z(n23261)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20887_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_3_i31_3_lut (.A(n653_adj_2459), .B(n30_adj_2460), .C(index_i[4]), 
         .Z(n31_adj_2461)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_3_i31_3_lut.init = 16'hcaca;
    LUT4 i19690_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n22045)) /* synthesis lut_function=(A (B (C)+!B !(C (D)+!C !(D)))+!A (B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i19690_3_lut_4_lut_4_lut.init = 16'hd6a5;
    PFUMX i23888 (.BLUT(n25600), .ALUT(n25599), .C0(index_q[5]), .Z(n25601));
    LUT4 i9492_3_lut (.A(n11977), .B(n29912), .C(index_i[3]), .Z(n11978)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9492_3_lut.init = 16'hcaca;
    LUT4 i9601_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[4]), .D(n27317), .Z(n189_adj_2462)) /* synthesis lut_function=(A (B (C (D)))+!A !(B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i9601_3_lut_4_lut_4_lut_4_lut.init = 16'h9555;
    LUT4 mux_229_Mux_0_i684_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n684_adj_2463)) /* synthesis lut_function=(!(A ((D)+!B)+!A !(B (D)+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_0_i684_3_lut_4_lut_4_lut_4_lut.init = 16'h5498;
    LUT4 i21364_3_lut (.A(n26096), .B(n23378), .C(index_q[6]), .Z(n23738)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21364_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_5_i31_3_lut (.A(n15_adj_2464), .B(n30_adj_2465), .C(index_q[4]), 
         .Z(n31_adj_2466)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_5_i31_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_4_i62_4_lut (.A(n27208), .B(n61_adj_2467), .C(index_q[4]), 
         .D(index_q[3]), .Z(n62_adj_2468)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_4_i62_4_lut.init = 16'hc5ca;
    LUT4 mux_230_Mux_4_i31_4_lut (.A(n15_adj_2469), .B(n27158), .C(index_q[4]), 
         .D(index_q[3]), .Z(n31_adj_2470)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_4_i31_4_lut.init = 16'h3aca;
    LUT4 n557_bdd_4_lut (.A(n27125), .B(index_q[4]), .C(n25596), .D(index_q[5]), 
         .Z(n27053)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (B (C (D))+!B (C+!(D)))) */ ;
    defparam n557_bdd_4_lut.init = 16'hf099;
    LUT4 mux_230_Mux_3_i31_3_lut (.A(n653_adj_2317), .B(n30_adj_2471), .C(index_q[4]), 
         .Z(n31_adj_2472)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_3_i31_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_0_i851_3_lut_4_lut_3_lut_rep_817 (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[1]), .Z(n29944)) /* synthesis lut_function=(A (B+(C))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_0_i851_3_lut_4_lut_3_lut_rep_817.init = 16'hb9b9;
    LUT4 mux_229_Mux_0_i796_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[1]), .D(index_i[3]), .Z(n796_adj_2473)) /* synthesis lut_function=(A (B (C+(D))+!B (C (D)))+!A !(B ((D)+!C)+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_0_i796_3_lut_4_lut_4_lut.init = 16'hb9c0;
    LUT4 mux_230_Mux_6_i29_3_lut_4_lut_3_lut_rep_818 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29945)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_6_i29_3_lut_4_lut_3_lut_rep_818.init = 16'h6969;
    LUT4 i9618_3_lut (.A(n12103), .B(n29918), .C(index_q[3]), .Z(n12104)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i9618_3_lut.init = 16'hcaca;
    LUT4 n173_bdd_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n29231)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C))+!A !(B (C (D)+!C !(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam n173_bdd_4_lut_4_lut.init = 16'ha569;
    LUT4 i22016_3_lut (.A(n142_adj_2286), .B(n14102), .C(index_i[4]), 
         .Z(n158_adj_2474)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22016_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_3_i963_3_lut_4_lut_3_lut_rep_819 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29946)) /* synthesis lut_function=(!(A (B)+!A ((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_3_i963_3_lut_4_lut_3_lut_rep_819.init = 16'h2626;
    LUT4 i19746_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n22101)) /* synthesis lut_function=(!(A (B)+!A (B (C+(D))+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i19746_3_lut_3_lut_4_lut.init = 16'h3326;
    LUT4 n62_bdd_3_lut_26407 (.A(n62_adj_2475), .B(n125), .C(index_i[6]), 
         .Z(n28686)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n62_bdd_3_lut_26407.init = 16'hcaca;
    LUT4 i19597_3_lut_else_4_lut (.A(index_q[4]), .B(index_q[2]), .C(index_q[3]), 
         .D(index_q[0]), .Z(n27501)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A !(B (C+!(D))+!B !(C)))) */ ;
    defparam i19597_3_lut_else_4_lut.init = 16'h6965;
    LUT4 i24099_then_4_lut (.A(index_i[0]), .B(index_i[4]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n27450)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)+!C !(D))+!B (C (D)))) */ ;
    defparam i24099_then_4_lut.init = 16'hda0e;
    LUT4 n23586_bdd_4_lut_26404 (.A(n252_adj_2338), .B(n27185), .C(index_i[4]), 
         .D(index_i[5]), .Z(n28684)) /* synthesis lut_function=(A (B (D)+!B ((D)+!C))+!A !(B+(C+(D)))) */ ;
    defparam n23586_bdd_4_lut_26404.init = 16'haa03;
    L6MUX21 i20465 (.D0(n22827), .D1(n22828), .SD(index_i[6]), .Z(n22839));
    LUT4 n62_bdd_4_lut_26408 (.A(n27302), .B(n27165), .C(index_i[6]), 
         .D(index_i[4]), .Z(n28687)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C+(D)))+!A (B ((D)+!C)+!B !(C)))) */ ;
    defparam n62_bdd_4_lut_26408.init = 16'h3af0;
    LUT4 i11673_3_lut_4_lut (.A(index_q[4]), .B(n27317), .C(index_q[5]), 
         .D(n27296), .Z(n892_adj_2476)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i11673_3_lut_4_lut.init = 16'hf8f0;
    L6MUX21 i20466 (.D0(n22829), .D1(n22830), .SD(index_i[6]), .Z(n22840));
    LUT4 mux_230_Mux_3_i676_3_lut_4_lut_3_lut_rep_820 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29947)) /* synthesis lut_function=(A (B (C))+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_3_i676_3_lut_4_lut_3_lut_rep_820.init = 16'h9494;
    L6MUX21 i20467 (.D0(n22831), .D1(n22832), .SD(index_i[6]), .Z(n22841));
    PFUMX i20468 (.BLUT(n22833), .ALUT(n22834), .C0(index_i[6]), .Z(n22842));
    LUT4 mux_230_Mux_3_i684_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[4]), .Z(n684_adj_2477)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A !(B ((D)+!C)+!B (C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_3_i684_3_lut_3_lut_4_lut.init = 16'h5594;
    LUT4 i21095_3_lut (.A(n27193), .B(n251_adj_2293), .C(index_q[4]), 
         .Z(n23469)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21095_3_lut.init = 16'hcaca;
    PFUMX i19913 (.BLUT(n22266), .ALUT(n22267), .C0(index_i[4]), .Z(n22268));
    PFUMX i20477 (.BLUT(n12124), .ALUT(n22136), .C0(index_i[6]), .Z(n22851));
    LUT4 index_i_6__bdd_1_lut (.A(index_i[5]), .Z(n27622)) /* synthesis lut_function=(!(A)) */ ;
    defparam index_i_6__bdd_1_lut.init = 16'h5555;
    LUT4 n23116_bdd_3_lut_23332 (.A(n23116), .B(n23115), .C(index_q[7]), 
         .Z(n24930)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n23116_bdd_3_lut_23332.init = 16'hacac;
    L6MUX21 i20479 (.D0(n22145), .D1(n22148), .SD(index_i[6]), .Z(n22853));
    L6MUX21 i20480 (.D0(n574_adj_2478), .D1(n22151), .SD(index_i[6]), 
            .Z(n22854));
    LUT4 mux_230_Mux_6_i860_3_lut_3_lut (.A(n27097), .B(index_q[4]), .C(n844_adj_2325), 
         .Z(n860_adj_2479)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam mux_230_Mux_6_i860_3_lut_3_lut.init = 16'h7474;
    L6MUX21 i20481 (.D0(n22154), .D1(n764_adj_2480), .SD(index_i[6]), 
            .Z(n22855));
    LUT4 i21088_3_lut (.A(n541_adj_2392), .B(n29960), .C(index_q[4]), 
         .Z(n23462)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21088_3_lut.init = 16'hcaca;
    LUT4 i19591_3_lut_3_lut (.A(n27097), .B(index_q[4]), .C(n46_adj_2481), 
         .Z(n21946)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam i19591_3_lut_3_lut.init = 16'h7474;
    LUT4 i20405_3_lut_4_lut_4_lut (.A(n27147), .B(index_q[4]), .C(index_q[5]), 
         .D(n27174), .Z(n22779)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C)+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i20405_3_lut_4_lut_4_lut.init = 16'h0434;
    LUT4 mux_229_Mux_3_i684_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[4]), .Z(n684_adj_2482)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A !(B ((D)+!C)+!B (C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_3_i684_3_lut_3_lut_4_lut.init = 16'h5594;
    LUT4 index_q_1__bdd_4_lut_26138 (.A(index_q[1]), .B(index_q[3]), .C(index_q[0]), 
         .D(index_q[2]), .Z(n28766)) /* synthesis lut_function=(A (B (C+(D))+!B (C (D)))+!A !(B (C)+!B !(C+(D)))) */ ;
    defparam index_q_1__bdd_4_lut_26138.init = 16'hbd94;
    LUT4 i22031_3_lut (.A(n22299), .B(n27494), .C(index_i[4]), .Z(n22301)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22031_3_lut.init = 16'hcaca;
    LUT4 n28766_bdd_3_lut (.A(n28766), .B(index_q[1]), .C(index_q[4]), 
         .Z(n28767)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n28766_bdd_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_3_i924_3_lut (.A(n908_adj_2383), .B(index_i[0]), .C(index_i[4]), 
         .Z(n924_adj_2483)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_3_i924_3_lut.init = 16'hcaca;
    L6MUX21 i20507 (.D0(n22865), .D1(n22866), .SD(index_i[6]), .Z(n22881));
    LUT4 mux_229_Mux_3_i891_3_lut (.A(n541_adj_2308), .B(n890_adj_2484), 
         .C(index_i[4]), .Z(n891_adj_2485)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_3_i891_3_lut.init = 16'hcaca;
    L6MUX21 i20508 (.D0(n22867), .D1(n22868), .SD(index_i[6]), .Z(n22882));
    L6MUX21 i20509 (.D0(n22869), .D1(n22870), .SD(index_i[6]), .Z(n22883));
    LUT4 mux_230_Mux_6_i269_rep_821 (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .Z(n29948)) /* synthesis lut_function=(A (C)+!A !((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_6_i269_rep_821.init = 16'ha4a4;
    LUT4 mux_229_Mux_3_i669_3_lut (.A(n653_adj_2454), .B(n668_adj_2436), 
         .C(index_i[4]), .Z(n669_adj_2486)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_3_i669_3_lut.init = 16'hcaca;
    LUT4 i9479_4_lut (.A(n27381), .B(n27229), .C(index_i[3]), .D(index_i[4]), 
         .Z(n11965)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B ((D)+!C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9479_4_lut.init = 16'h3afa;
    L6MUX21 i20510 (.D0(n22871), .D1(n22872), .SD(index_i[6]), .Z(n22884));
    L6MUX21 i20511 (.D0(n22873), .D1(n22874), .SD(index_i[6]), .Z(n22885));
    L6MUX21 i20513 (.D0(n22877), .D1(n22878), .SD(index_i[6]), .Z(n22887));
    L6MUX21 i21439 (.D0(n23805), .D1(n23806), .SD(index_q[6]), .Z(n23813));
    L6MUX21 i21440 (.D0(n23807), .D1(n23808), .SD(index_q[6]), .Z(n23814));
    L6MUX21 i21441 (.D0(n23809), .D1(n23810), .SD(index_q[6]), .Z(n23815));
    L6MUX21 i21442 (.D0(n23811), .D1(n23812), .SD(index_q[6]), .Z(n23816));
    LUT4 mux_230_Mux_0_i220_3_lut (.A(n27238), .B(n27426), .C(index_q[3]), 
         .Z(n220)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_0_i220_3_lut.init = 16'hcaca;
    LUT4 i22042_3_lut (.A(n22281), .B(n22282), .C(index_i[4]), .Z(n22283)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22042_3_lut.init = 16'hcaca;
    L6MUX21 i20538 (.D0(n22896), .D1(n22897), .SD(index_i[6]), .Z(n22912));
    L6MUX21 i20539 (.D0(n22898), .D1(n22899), .SD(index_i[6]), .Z(n22913));
    L6MUX21 i20540 (.D0(n22900), .D1(n22901), .SD(index_i[6]), .Z(n22914));
    LUT4 i20943_3_lut_3_lut_4_lut (.A(n27213), .B(index_i[3]), .C(n316_adj_2487), 
         .D(index_i[4]), .Z(n23317)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20943_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 mux_229_Mux_3_i476_3_lut (.A(n460_adj_2488), .B(n285_adj_2489), 
         .C(index_i[4]), .Z(n476_adj_2490)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_3_i476_3_lut.init = 16'hcaca;
    PFUMX i20542 (.BLUT(n22904), .ALUT(n22905), .C0(index_i[6]), .Z(n22916));
    L6MUX21 i20543 (.D0(n22906), .D1(n22907), .SD(index_i[6]), .Z(n22917));
    LUT4 mux_229_Mux_3_i413_3_lut (.A(n397_adj_2311), .B(n27349), .C(index_i[4]), 
         .Z(n413_adj_2491)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_3_i413_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_7_i890_3_lut_4_lut (.A(n27293), .B(index_q[2]), .C(index_q[3]), 
         .D(n27218), .Z(n890_adj_2287)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_7_i890_3_lut_4_lut.init = 16'hf101;
    LUT4 i19879_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n22234)) /* synthesis lut_function=(!(A ((D)+!C)+!A !(B ((D)+!C)+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i19879_3_lut_3_lut_4_lut.init = 16'h55a4;
    L6MUX21 i20544 (.D0(n22908), .D1(n22909), .SD(index_i[6]), .Z(n22918));
    LUT4 i20478_3_lut (.A(n26390), .B(n23561), .C(index_i[6]), .Z(n22852)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20478_3_lut.init = 16'hcaca;
    PFUMX i20545 (.BLUT(n22910), .ALUT(n22911), .C0(index_i[6]), .Z(n22919));
    LUT4 mux_229_Mux_3_i286_4_lut (.A(n93_adj_2492), .B(index_i[2]), .C(index_i[4]), 
         .D(n14095), .Z(n286_adj_2493)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_3_i286_4_lut.init = 16'h3aca;
    LUT4 n23124_bdd_3_lut (.A(n23117), .B(n23118), .C(index_q[7]), .Z(n24928)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n23124_bdd_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_3_i158_3_lut (.A(n142_adj_2444), .B(n157), .C(index_i[4]), 
         .Z(n158_adj_2494)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_3_i158_3_lut.init = 16'hcaca;
    PFUMX i20565 (.BLUT(n797_adj_2495), .ALUT(n828_adj_2339), .C0(index_i[5]), 
          .Z(n22939));
    LUT4 mux_230_Mux_6_i356_3_lut_4_lut_3_lut_rep_822 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29949)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_6_i356_3_lut_4_lut_3_lut_rep_822.init = 16'h4949;
    LUT4 mux_229_Mux_3_i125_3_lut (.A(n109_adj_2496), .B(n526_adj_2315), 
         .C(index_i[4]), .Z(n125_adj_2497)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_3_i125_3_lut.init = 16'hcaca;
    LUT4 i19845_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n22200)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (D))+!A !(B (C (D))+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i19845_3_lut_3_lut_4_lut.init = 16'h4933;
    L6MUX21 i20569 (.D0(n22927), .D1(n22928), .SD(index_i[6]), .Z(n22943));
    LUT4 mux_229_Mux_8_i124_3_lut_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n124_adj_2498)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C+!(D)))+!A (B (C (D)+!C !(D))+!B (C)))) */ ;
    defparam mux_229_Mux_8_i124_3_lut_3_lut_4_lut_4_lut.init = 16'h07c1;
    L6MUX21 i20570 (.D0(n22929), .D1(n22930), .SD(index_i[6]), .Z(n22944));
    LUT4 n581_bdd_4_lut_26342 (.A(index_q[2]), .B(index_q[1]), .C(index_q[0]), 
         .D(index_q[5]), .Z(n28893)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A !(B+!(C (D)+!C !(D))))) */ ;
    defparam n581_bdd_4_lut_26342.init = 16'h657e;
    LUT4 n27294_bdd_4_lut_26322 (.A(index_q[2]), .B(index_q[1]), .C(index_q[0]), 
         .D(index_q[3]), .Z(n28895)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)+!C !(D)))+!A (B (C (D))+!B (C+!(D))))) */ ;
    defparam n27294_bdd_4_lut_26322.init = 16'h0f64;
    LUT4 i20537_4_lut (.A(n22268), .B(n1002_adj_2499), .C(index_i[5]), 
         .D(index_i[4]), .Z(n22911)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;
    defparam i20537_4_lut.init = 16'hfaca;
    LUT4 mux_229_Mux_0_i908_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n908_adj_2500)) /* synthesis lut_function=(!(A (B (C (D))+!B !(D))+!A (B+((D)+!C)))) */ ;
    defparam mux_229_Mux_0_i908_3_lut_4_lut_4_lut.init = 16'h2a98;
    LUT4 mux_230_Mux_8_i892_3_lut_4_lut (.A(n27147), .B(index_q[4]), .C(index_q[5]), 
         .D(n860_adj_2501), .Z(n892_adj_2502)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_8_i892_3_lut_4_lut.init = 16'h4f40;
    LUT4 mux_229_Mux_4_i860_3_lut (.A(n506), .B(n15_adj_2503), .C(index_i[4]), 
         .Z(n860_adj_2504)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_4_i860_3_lut.init = 16'hcaca;
    L6MUX21 i20571 (.D0(n22931), .D1(n22932), .SD(index_i[6]), .Z(n22945));
    LUT4 i21113_3_lut (.A(n29233), .B(n23481), .C(index_q[6]), .Z(n23487)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21113_3_lut.init = 16'hcaca;
    LUT4 i22068_3_lut (.A(n21747), .B(n21748), .C(index_i[4]), .Z(n21749)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22068_3_lut.init = 16'hcaca;
    LUT4 i21114_3_lut (.A(n28898), .B(n23483), .C(index_q[6]), .Z(n23488)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21114_3_lut.init = 16'hcaca;
    L6MUX21 i20572 (.D0(n22933), .D1(n22934), .SD(index_i[6]), .Z(n22946));
    LUT4 i22070_3_lut (.A(n21744), .B(n21745), .C(index_i[4]), .Z(n21746)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22070_3_lut.init = 16'hcaca;
    L6MUX21 i20573 (.D0(n22935), .D1(n22936), .SD(index_i[6]), .Z(n22947));
    L6MUX21 i20576 (.D0(n22941), .D1(n22942), .SD(index_i[6]), .Z(n22950));
    LUT4 i21144_3_lut (.A(n23511), .B(n23512), .C(index_i[6]), .Z(n23518)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21144_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_0_i1002_3_lut_3_lut_4_lut (.A(n27293), .B(index_q[2]), 
         .C(n38), .D(index_q[3]), .Z(n1002_adj_2431)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_0_i1002_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 i21145_3_lut (.A(n26729), .B(n23514), .C(index_i[6]), .Z(n23519)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21145_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_8_i475_3_lut_3_lut_4_lut (.A(n27293), .B(index_q[2]), 
         .C(n27219), .D(index_q[3]), .Z(n475_adj_2505)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_8_i475_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 mux_230_Mux_9_i124_3_lut_3_lut_4_lut (.A(n27293), .B(index_q[2]), 
         .C(n27219), .D(index_q[3]), .Z(n124_adj_2506)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_9_i124_3_lut_3_lut_4_lut.init = 16'h11f0;
    PFUMX i19437 (.BLUT(n318), .ALUT(n381_adj_2340), .C0(index_i[6]), 
          .Z(n21792));
    LUT4 mux_229_Mux_4_i700_3_lut (.A(n684), .B(index_i[1]), .C(index_i[4]), 
         .Z(n700_adj_2507)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_4_i700_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_4_i669_3_lut (.A(n653_adj_2459), .B(n668_adj_2508), 
         .C(index_i[4]), .Z(n669_adj_2509)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_4_i669_3_lut.init = 16'hcaca;
    PFUMX i19428 (.BLUT(n318_adj_2510), .ALUT(n381), .C0(index_q[6]), 
          .Z(n21783));
    LUT4 n23116_bdd_3_lut_24682 (.A(n23113), .B(n23114), .C(index_q[7]), 
         .Z(n24931)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n23116_bdd_3_lut_24682.init = 16'hcaca;
    LUT4 mux_229_Mux_4_i542_3_lut (.A(n526_adj_2315), .B(n541_adj_2420), 
         .C(index_i[4]), .Z(n542_adj_2511)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_4_i542_3_lut.init = 16'hcaca;
    LUT4 i20531_4_lut (.A(n27152), .B(n27479), .C(index_i[5]), .D(index_i[4]), 
         .Z(n22905)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam i20531_4_lut.init = 16'hc5ca;
    LUT4 i9681_3_lut_then_4_lut (.A(index_i[4]), .B(index_i[0]), .C(index_i[1]), 
         .D(index_i[2]), .Z(n27505)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C+(D)))+!A (B (C+(D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9681_3_lut_then_4_lut.init = 16'hd54a;
    LUT4 mux_230_Mux_2_i189_3_lut_3_lut_4_lut (.A(index_q[1]), .B(n27317), 
         .C(n173), .D(index_q[4]), .Z(n189_adj_2512)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(C+(D)))) */ ;
    defparam mux_230_Mux_2_i189_3_lut_3_lut_4_lut.init = 16'h77f0;
    LUT4 i11637_2_lut_3_lut_4_lut (.A(index_q[1]), .B(n27317), .C(index_q[5]), 
         .D(index_q[4]), .Z(n508_adj_2513)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;
    defparam i11637_2_lut_3_lut_4_lut.init = 16'hf080;
    LUT4 mux_230_Mux_6_i22_rep_823 (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .Z(n29950)) /* synthesis lut_function=(!(A (C)+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_6_i22_rep_823.init = 16'h4a4a;
    LUT4 i9587_3_lut_4_lut (.A(n27253), .B(index_q[2]), .C(n27323), .D(n27276), 
         .Z(n444_adj_2514)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i9587_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_230_Mux_6_i251_3_lut_4_lut (.A(n27253), .B(index_q[2]), .C(index_q[3]), 
         .D(n27276), .Z(n251_adj_2441)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_6_i251_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_229_Mux_4_i286_3_lut (.A(n270), .B(n15_adj_2273), .C(index_i[4]), 
         .Z(n286_adj_2515)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_4_i286_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_6_i157_3_lut_4_lut (.A(n27253), .B(index_q[2]), .C(index_q[3]), 
         .D(n29955), .Z(n157_adj_2516)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_6_i157_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_230_Mux_4_i747_3_lut_4_lut (.A(n27253), .B(index_q[2]), .C(index_q[3]), 
         .D(n27280), .Z(n747_adj_2414)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_4_i747_3_lut_4_lut.init = 16'hf606;
    LUT4 i11405_2_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n844_adj_2313)) /* synthesis lut_function=(A (B+!(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11405_2_lut_3_lut_4_lut.init = 16'h9ff9;
    LUT4 i9681_3_lut_else_4_lut (.A(index_i[4]), .B(index_i[0]), .C(index_i[1]), 
         .D(index_i[2]), .Z(n27504)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A !(B (D)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9681_3_lut_else_4_lut.init = 16'ha955;
    LUT4 i24099_else_4_lut (.A(index_i[0]), .B(index_i[4]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n27449)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C))+!A (B (C)+!B (C+(D)))) */ ;
    defparam i24099_else_4_lut.init = 16'hf178;
    LUT4 mux_229_Mux_6_i378_3_lut_4_lut_3_lut_rep_786 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29913)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_6_i378_3_lut_4_lut_3_lut_rep_786.init = 16'h4949;
    LUT4 mux_229_Mux_3_i859_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n859_adj_2517)) /* synthesis lut_function=(!(A (B (D)+!B !(D))+!A (B (C+(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_3_i859_3_lut_3_lut_4_lut.init = 16'h339c;
    L6MUX21 i21112 (.D0(n23478), .D1(n23479), .SD(index_q[6]), .Z(n23486));
    LUT4 mux_229_Mux_4_i94_3_lut (.A(n61), .B(n27355), .C(index_i[4]), 
         .Z(n94_adj_2518)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_4_i94_3_lut.init = 16'hcaca;
    L6MUX21 i20677 (.D0(n23385), .D1(n23392), .SD(index_q[6]), .Z(n23051));
    LUT4 mux_230_Mux_5_i491_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n491_adj_2519)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A !(B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_5_i491_3_lut_4_lut_4_lut.init = 16'ha54a;
    LUT4 mux_229_Mux_5_i483_rep_824 (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .Z(n29951)) /* synthesis lut_function=(!(A (C)+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_5_i483_rep_824.init = 16'h4a4a;
    LUT4 mux_229_Mux_4_i262_3_lut_3_lut_rep_785 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29912)) /* synthesis lut_function=(A (B+(C))+!A !(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_4_i262_3_lut_3_lut_rep_785.init = 16'ha9a9;
    LUT4 mux_229_Mux_5_i491_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n491_adj_2520)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A !(B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_5_i491_3_lut_4_lut_4_lut.init = 16'ha54a;
    L6MUX21 i21115 (.D0(n23484), .D1(n23485), .SD(index_q[6]), .Z(n23489));
    LUT4 i19999_3_lut_4_lut_4_lut (.A(n27322), .B(n27353), .C(index_i[3]), 
         .D(index_i[0]), .Z(n22354)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C))) */ ;
    defparam i19999_3_lut_4_lut_4_lut.init = 16'hcfc5;
    PFUMX i20524 (.BLUT(n158_adj_2521), .ALUT(n189_adj_2380), .C0(index_i[5]), 
          .Z(n22898));
    LUT4 mux_229_Mux_0_i708_3_lut_4_lut_3_lut_rep_794 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29921)) /* synthesis lut_function=(!(A (B)+!A ((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_0_i708_3_lut_4_lut_3_lut_rep_794.init = 16'h2626;
    PFUMX i23388 (.BLUT(n24990), .ALUT(n23785), .C0(index_q[8]), .Z(n24991));
    LUT4 mux_229_Mux_6_i315_rep_825 (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .Z(n29952)) /* synthesis lut_function=(A (C)+!A !((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_6_i315_rep_825.init = 16'ha4a4;
    LUT4 mux_230_Mux_8_i732_3_lut (.A(index_q[3]), .B(n15348), .C(index_q[5]), 
         .Z(n732_adj_2522)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_8_i732_3_lut.init = 16'h3a3a;
    LUT4 i19885_3_lut_4_lut (.A(n27293), .B(index_q[2]), .C(index_q[3]), 
         .D(n27275), .Z(n22240)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i19885_3_lut_4_lut.init = 16'hf404;
    LUT4 i22095_3_lut (.A(n21999), .B(n22000), .C(index_q[4]), .Z(n22001)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i22095_3_lut.init = 16'hcaca;
    LUT4 i20035_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n22390)) /* synthesis lut_function=(!(A ((D)+!C)+!A !(B ((D)+!C)+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20035_3_lut_3_lut_4_lut.init = 16'h55a4;
    LUT4 mux_230_Mux_6_i340_3_lut_4_lut_3_lut_rep_826 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29953)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_6_i340_3_lut_4_lut_3_lut_rep_826.init = 16'h9292;
    L6MUX21 i20601 (.D0(n22960), .D1(n22961), .SD(index_i[6]), .Z(n22975));
    L6MUX21 i20602 (.D0(n22962), .D1(n22963), .SD(index_i[6]), .Z(n22976));
    LUT4 mux_230_Mux_0_i731_3_lut_4_lut (.A(n27293), .B(index_q[2]), .C(index_q[3]), 
         .D(n29934), .Z(n731_adj_2407)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_0_i731_3_lut_4_lut.init = 16'h4f40;
    L6MUX21 i20603 (.D0(n22964), .D1(n22965), .SD(index_i[6]), .Z(n22977));
    LUT4 mux_229_Mux_5_i891_3_lut (.A(n875), .B(n890_adj_2523), .C(index_i[4]), 
         .Z(n891_adj_2524)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_5_i891_3_lut.init = 16'hcaca;
    L6MUX21 i20604 (.D0(n22966), .D1(n22967), .SD(index_i[6]), .Z(n22978));
    LUT4 mux_229_Mux_5_i860_3_lut (.A(n15), .B(n859), .C(index_i[4]), 
         .Z(n860_adj_2525)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_5_i860_3_lut.init = 16'hcaca;
    L6MUX21 i21143 (.D0(n23509), .D1(n23510), .SD(index_i[6]), .Z(n23517));
    LUT4 i20460_3_lut_4_lut (.A(n27152), .B(n27124), .C(index_i[4]), .D(index_i[5]), 
         .Z(n22834)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (B+((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20460_3_lut_4_lut.init = 16'hffc5;
    L6MUX21 i20605 (.D0(n22968), .D1(n22969), .SD(index_i[6]), .Z(n22979));
    L6MUX21 i21146 (.D0(n23515), .D1(n23516), .SD(index_i[6]), .Z(n23520));
    PFUMX i25190 (.BLUT(n27528), .ALUT(n27529), .C0(index_i[0]), .Z(n27530));
    PFUMX i25090 (.BLUT(n26986), .ALUT(n26984), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2145[10]));
    LUT4 i22101_3_lut (.A(n21720), .B(n21721), .C(index_i[4]), .Z(n21722)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22101_3_lut.init = 16'hcaca;
    LUT4 i20001_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n22356)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (D))+!A !(B (C (D))+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20001_3_lut_3_lut_4_lut.init = 16'h4933;
    LUT4 i22963_2_lut_rep_788 (.A(index_i[0]), .B(index_i[1]), .Z(n29915)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i22963_2_lut_rep_788.init = 16'h9999;
    L6MUX21 i20476 (.D0(n22130), .D1(n22133), .SD(index_i[6]), .Z(n22850));
    LUT4 mux_230_Mux_2_i700_3_lut_4_lut (.A(index_q[1]), .B(n27307), .C(index_q[4]), 
         .D(n684_adj_2281), .Z(n700_adj_2526)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_2_i700_3_lut_4_lut.init = 16'hefe0;
    PFUMX i19937 (.BLUT(n22290), .ALUT(n22291), .C0(index_i[4]), .Z(n22292));
    LUT4 mux_229_Mux_5_i636_4_lut (.A(n157_adj_2527), .B(n27212), .C(index_i[4]), 
         .D(index_i[3]), .Z(n636_adj_2528)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_5_i636_4_lut.init = 16'h3aca;
    LUT4 i22105_3_lut (.A(n18091), .B(n18092), .C(index_i[4]), .Z(n18093)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22105_3_lut.init = 16'hcaca;
    PFUMX i25088 (.BLUT(n21795), .ALUT(n26982), .C0(index_i[7]), .Z(n26983));
    LUT4 mux_229_Mux_5_i507_3_lut (.A(n491_adj_2520), .B(n506), .C(index_i[4]), 
         .Z(n507)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_5_i507_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_5_i476_3_lut (.A(n460_adj_2529), .B(n475_adj_2530), 
         .C(index_i[4]), .Z(n476_adj_2531)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_5_i476_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_3_i1018_3_lut_4_lut (.A(index_q[1]), .B(n27307), .C(index_q[4]), 
         .D(n20198), .Z(n1018_adj_2532)) /* synthesis lut_function=(A (C+!(D))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_3_i1018_3_lut_4_lut.init = 16'he0ef;
    LUT4 mux_229_Mux_5_i413_3_lut (.A(n397), .B(n251), .C(index_i[4]), 
         .Z(n413_adj_2533)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_5_i413_3_lut.init = 16'hcaca;
    LUT4 n986_bdd_4_lut (.A(n27124), .B(index_i[6]), .C(n27159), .D(index_i[5]), 
         .Z(n25794)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C+!(D))+!B (D))) */ ;
    defparam n986_bdd_4_lut.init = 16'hd1cc;
    PFUMX i20626 (.BLUT(n732_adj_2534), .ALUT(n763_adj_2535), .C0(index_i[5]), 
          .Z(n23000));
    LUT4 n124_bdd_3_lut_24044_4_lut (.A(n27371), .B(index_q[3]), .C(index_q[4]), 
         .D(n124_adj_2506), .Z(n25757)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam n124_bdd_3_lut_24044_4_lut.init = 16'hf101;
    LUT4 i20921_3_lut_4_lut (.A(n27371), .B(index_q[3]), .C(index_q[4]), 
         .D(n285), .Z(n23295)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i20921_3_lut_4_lut.init = 16'hfe0e;
    L6MUX21 i20628 (.D0(n22403), .D1(n891_adj_2536), .SD(index_i[5]), 
            .Z(n23002));
    L6MUX21 i20631 (.D0(n22989), .D1(n22990), .SD(index_i[6]), .Z(n23005));
    LUT4 n526_bdd_3_lut_24010_4_lut_4_lut (.A(n27371), .B(index_q[3]), .C(index_q[4]), 
         .D(n27172), .Z(n25713)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B (C (D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam n526_bdd_3_lut_24010_4_lut_4_lut.init = 16'h3efe;
    LUT4 mux_230_Mux_0_i812_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n812_adj_2423)) /* synthesis lut_function=(A (B (C+(D))+!B !(C))+!A (B (D)+!B !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_0_i812_3_lut_4_lut_4_lut_4_lut.init = 16'hcf92;
    LUT4 i19758_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n22113)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C))+!A !(B ((D)+!C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i19758_3_lut_4_lut_4_lut.init = 16'h925a;
    LUT4 mux_230_Mux_4_i573_3_lut_3_lut_4_lut_4_lut (.A(n27371), .B(index_q[3]), 
         .C(index_q[4]), .D(n27220), .Z(n573_adj_2537)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_4_i573_3_lut_3_lut_4_lut_4_lut.init = 16'h1f1c;
    LUT4 mux_230_Mux_2_i573_3_lut_3_lut_4_lut (.A(n27371), .B(index_q[3]), 
         .C(n557_adj_2369), .D(index_q[4]), .Z(n573_adj_2538)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_2_i573_3_lut_3_lut_4_lut.init = 16'h11f0;
    PFUMX i25188 (.BLUT(n27525), .ALUT(n27526), .C0(index_i[0]), .Z(n27527));
    LUT4 mux_230_Mux_3_i573_3_lut_3_lut_4_lut (.A(n27371), .B(index_q[3]), 
         .C(n397_adj_2539), .D(index_q[4]), .Z(n573_adj_2540)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_3_i573_3_lut_3_lut_4_lut.init = 16'h11f0;
    LUT4 i15933_3_lut (.A(n18117), .B(n18118), .C(index_i[4]), .Z(n18119)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15933_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_5_i125_3_lut (.A(n109_adj_2541), .B(n124_adj_2542), 
         .C(index_i[4]), .Z(n125_adj_2543)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_5_i125_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_5_i94_3_lut (.A(n653_adj_2544), .B(n635_adj_2318), 
         .C(index_i[4]), .Z(n94_adj_2545)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_5_i94_3_lut.init = 16'hcaca;
    LUT4 n29166_bdd_3_lut (.A(n29166), .B(index_i[1]), .C(index_i[4]), 
         .Z(n29167)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n29166_bdd_3_lut.init = 16'hcaca;
    LUT4 index_i_1__bdd_4_lut_26727 (.A(index_i[1]), .B(index_i[3]), .C(index_i[2]), 
         .D(index_i[0]), .Z(n29166)) /* synthesis lut_function=(A (B (C+(D))+!B (C (D)))+!A !(B (D)+!B !(C+(D)))) */ ;
    defparam index_i_1__bdd_4_lut_26727.init = 16'hb9d4;
    LUT4 i20923_3_lut_3_lut_4_lut_4_lut (.A(n27334), .B(index_q[3]), .C(index_q[4]), 
         .D(n27220), .Z(n23297)) /* synthesis lut_function=(!(A (B (C)+!B ((D)+!C))+!A (B+((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i20923_3_lut_3_lut_4_lut_4_lut.init = 16'h0838;
    LUT4 i19944_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n22299)) /* synthesis lut_function=(!(A (B)+!A (B (C+(D))+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19944_3_lut_3_lut_4_lut.init = 16'h3326;
    PFUMX i25186 (.BLUT(n27522), .ALUT(n27523), .C0(index_q[1]), .Z(n27524));
    LUT4 i9561_3_lut_4_lut_4_lut (.A(n27334), .B(index_q[3]), .C(index_q[5]), 
         .D(n27218), .Z(n12047)) /* synthesis lut_function=(A (B+(C (D)))+!A (B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i9561_3_lut_4_lut_4_lut.init = 16'hf8c8;
    LUT4 n62_bdd_3_lut_4_lut (.A(n27334), .B(index_q[3]), .C(index_q[4]), 
         .D(n30_adj_2546), .Z(n25760)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam n62_bdd_3_lut_4_lut.init = 16'hf808;
    LUT4 n557_bdd_3_lut_23912_4_lut_4_lut (.A(n27334), .B(index_q[3]), .C(index_q[4]), 
         .D(n27172), .Z(n25600)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C))+!A !(B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam n557_bdd_3_lut_23912_4_lut_4_lut.init = 16'h838f;
    L6MUX21 i20633 (.D0(n22993), .D1(n22994), .SD(index_i[6]), .Z(n23007));
    LUT4 n27434_bdd_3_lut_26388 (.A(n27213), .B(index_i[6]), .C(index_i[5]), 
         .Z(n27626)) /* synthesis lut_function=(!(A (B)+!A (C))) */ ;
    defparam n27434_bdd_3_lut_26388.init = 16'h2727;
    L6MUX21 i21174 (.D0(n23540), .D1(n23541), .SD(index_i[6]), .Z(n23548));
    L6MUX21 i20634 (.D0(n22995), .D1(n22996), .SD(index_i[6]), .Z(n23008));
    LUT4 i19701_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n22056)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A !(B (C+!(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i19701_3_lut_4_lut_4_lut.init = 16'ha52b;
    L6MUX21 i21175 (.D0(n23542), .D1(n23543), .SD(index_i[6]), .Z(n23549));
    L6MUX21 i21176 (.D0(n23544), .D1(n23545), .SD(index_i[6]), .Z(n23550));
    L6MUX21 i21177 (.D0(n23546), .D1(n23547), .SD(index_i[6]), .Z(n23551));
    LUT4 index_i_2__bdd_4_lut (.A(index_i[2]), .B(index_i[0]), .C(index_i[3]), 
         .D(index_i[1]), .Z(n29964)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B ((D)+!C)+!B !(C (D)+!C !(D)))) */ ;
    defparam index_i_2__bdd_4_lut.init = 16'hed34;
    LUT4 mux_230_Mux_6_i156_3_lut_rep_828 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29955)) /* synthesis lut_function=(!(A (B+(C))+!A !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_6_i156_3_lut_rep_828.init = 16'h5252;
    LUT4 mux_229_Mux_7_i892_3_lut (.A(n62), .B(n891_adj_2361), .C(index_i[5]), 
         .Z(n892_adj_2416)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_7_i892_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_0_i173_3_lut_4_lut (.A(n27340), .B(index_i[1]), .C(index_i[3]), 
         .D(n27346), .Z(n173_adj_2547)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_0_i173_3_lut_4_lut.init = 16'hdfd0;
    LUT4 i19861_3_lut (.A(n747_adj_2548), .B(n908_adj_2549), .C(index_i[4]), 
         .Z(n22216)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19861_3_lut.init = 16'hcaca;
    LUT4 i19860_3_lut (.A(n716_adj_2323), .B(n15204), .C(index_i[4]), 
         .Z(n22215)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19860_3_lut.init = 16'hcaca;
    LUT4 i19653_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n22008)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C))+!A !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i19653_3_lut_4_lut_4_lut.init = 16'h5a52;
    LUT4 i19852_3_lut (.A(n93_adj_2550), .B(n699), .C(index_i[4]), .Z(n22207)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19852_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_1_i620_3_lut_4_lut (.A(n27340), .B(index_i[1]), .C(index_i[3]), 
         .D(n29912), .Z(n620_adj_2551)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_1_i620_3_lut_4_lut.init = 16'hdfd0;
    LUT4 i19851_3_lut (.A(n653_adj_2552), .B(n27096), .C(index_i[4]), 
         .Z(n22206)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19851_3_lut.init = 16'hcaca;
    LUT4 i19354_3_lut_4_lut (.A(n27340), .B(index_i[1]), .C(index_i[3]), 
         .D(n498), .Z(n21709)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19354_3_lut_4_lut.init = 16'hdfd0;
    LUT4 n27298_bdd_4_lut (.A(index_q[5]), .B(index_q[0]), .C(index_q[1]), 
         .D(index_q[2]), .Z(n29228)) /* synthesis lut_function=(!(A (B (C (D))+!B (C (D)+!C !(D)))+!A !(B (C (D))+!B (C+(D))))) */ ;
    defparam n27298_bdd_4_lut.init = 16'h5bb8;
    LUT4 mux_229_Mux_6_i891_3_lut (.A(n78), .B(n890_adj_2334), .C(index_i[4]), 
         .Z(n891_adj_2553)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_6_i891_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_6_i828_4_lut (.A(n812_adj_2554), .B(n14070), .C(index_i[4]), 
         .D(index_i[2]), .Z(n828_adj_2555)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_6_i828_4_lut.init = 16'hfaca;
    LUT4 mux_229_Mux_6_i844_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n844_adj_2556)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (B (C)+!B !(C+!(D)))) */ ;
    defparam mux_229_Mux_6_i844_3_lut_4_lut_4_lut.init = 16'hc1e0;
    LUT4 n476_bdd_3_lut_23707 (.A(n476), .B(n25353), .C(index_q[5]), .Z(n25354)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n476_bdd_3_lut_23707.init = 16'hcaca;
    LUT4 mux_229_Mux_6_i797_3_lut (.A(n653_adj_2459), .B(n27071), .C(index_i[4]), 
         .Z(n797_adj_2557)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_6_i797_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_6_i669_3_lut (.A(n653_adj_2544), .B(n668_adj_2558), 
         .C(index_i[4]), .Z(n669_adj_2559)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_6_i669_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_6_i542_3_lut (.A(n526_adj_2560), .B(n541_adj_2308), 
         .C(index_i[4]), .Z(n542_adj_2561)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_6_i542_3_lut.init = 16'hcaca;
    LUT4 index_i_5__bdd_4_lut_24653 (.A(index_i[2]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[0]), .Z(n26452)) /* synthesis lut_function=(A (B (C+!(D))+!B !(D))+!A !(B (C+!(D))+!B !(D))) */ ;
    defparam index_i_5__bdd_4_lut_24653.init = 16'h95aa;
    LUT4 i19888_3_lut_4_lut (.A(n27296), .B(index_q[2]), .C(index_q[3]), 
         .D(n29919), .Z(n22243)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i19888_3_lut_4_lut.init = 16'hdfd0;
    LUT4 i19833_3_lut (.A(n526_adj_2562), .B(n15_adj_2280), .C(index_i[4]), 
         .Z(n22188)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19833_3_lut.init = 16'hcaca;
    LUT4 i19834_3_lut_4_lut_4_lut_4_lut (.A(n27434), .B(index_i[2]), .C(index_i[3]), 
         .D(index_i[4]), .Z(n22189)) /* synthesis lut_function=(A (B)+!A (B (C (D))+!B !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19834_3_lut_4_lut_4_lut_4_lut.init = 16'hc999;
    LUT4 mux_229_Mux_7_i475_3_lut_3_lut_4_lut (.A(n27434), .B(index_i[2]), 
         .C(n27432), .D(index_i[3]), .Z(n475_adj_2563)) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))+!A !(B ((D)+!C)+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_7_i475_3_lut_3_lut_4_lut.init = 16'h99f0;
    LUT4 n26454_bdd_3_lut (.A(n26454), .B(n26451), .C(index_i[4]), .Z(n26455)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n26454_bdd_3_lut.init = 16'hcaca;
    LUT4 i19348_3_lut_4_lut (.A(n27434), .B(index_i[2]), .C(index_i[3]), 
         .D(n27383), .Z(n21703)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19348_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_229_Mux_7_i653_3_lut_4_lut (.A(n27434), .B(index_i[2]), .C(index_i[3]), 
         .D(n27430), .Z(n653_adj_2552)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_7_i653_3_lut_4_lut.init = 16'hf606;
    LUT4 i21120_3_lut_4_lut (.A(n27229), .B(index_i[3]), .C(index_i[4]), 
         .D(n46_adj_2388), .Z(n23494)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21120_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_229_Mux_2_i684_3_lut_4_lut (.A(n27434), .B(index_i[2]), .C(index_i[3]), 
         .D(n27388), .Z(n684_adj_2447)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_2_i684_3_lut_4_lut.init = 16'h6f60;
    LUT4 i19858_3_lut (.A(n29940), .B(n27276), .C(index_q[3]), .Z(n22213)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19858_3_lut.init = 16'hcaca;
    LUT4 i12496_3_lut (.A(index_q[3]), .B(index_q[1]), .C(index_q[0]), 
         .Z(n15103)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i12496_3_lut.init = 16'hecec;
    LUT4 n25356_bdd_3_lut (.A(n27539), .B(n444), .C(index_q[5]), .Z(n25357)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n25356_bdd_3_lut.init = 16'hcaca;
    LUT4 i19842_4_lut_4_lut_4_lut (.A(n27434), .B(index_i[2]), .C(index_i[4]), 
         .D(index_i[3]), .Z(n22197)) /* synthesis lut_function=(A (B)+!A !(B (C+(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19842_4_lut_4_lut_4_lut.init = 16'h999c;
    LUT4 i15950_4_lut (.A(index_i[0]), .B(index_i[4]), .C(index_i[1]), 
         .D(n27302), .Z(n286_adj_2564)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i15950_4_lut.init = 16'hccc8;
    LUT4 i19824_3_lut (.A(n397_adj_2565), .B(n475_adj_2563), .C(index_i[4]), 
         .Z(n22179)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19824_3_lut.init = 16'hcaca;
    LUT4 i19816_3_lut (.A(n348_adj_2566), .B(n443_adj_2567), .C(index_i[4]), 
         .Z(n22171)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19816_3_lut.init = 16'hcaca;
    LUT4 i19815_3_lut (.A(n397_adj_2565), .B(n781_adj_2568), .C(index_i[4]), 
         .Z(n22170)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19815_3_lut.init = 16'hcaca;
    LUT4 i20518_3_lut (.A(n22887), .B(n25266), .C(index_i[7]), .Z(n22892)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20518_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_7_i443_3_lut_4_lut (.A(n27429), .B(index_i[2]), .C(index_i[3]), 
         .D(n27386), .Z(n443_adj_2567)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_7_i443_3_lut_4_lut.init = 16'h6f60;
    LUT4 i19347_3_lut_3_lut_4_lut (.A(n27429), .B(index_i[2]), .C(n27386), 
         .D(index_i[3]), .Z(n21702)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19347_3_lut_3_lut_4_lut.init = 16'hf099;
    LUT4 i20840_3_lut (.A(n23206), .B(n23207), .C(index_q[7]), .Z(n23214)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20840_3_lut.init = 16'hcaca;
    LUT4 i19929_3_lut_3_lut_4_lut (.A(n27429), .B(index_i[2]), .C(n27385), 
         .D(index_i[3]), .Z(n22284)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19929_3_lut_3_lut_4_lut.init = 16'hf099;
    LUT4 mux_229_Mux_3_i860_3_lut_4_lut (.A(n27429), .B(index_i[2]), .C(index_i[4]), 
         .D(n859_adj_2517), .Z(n860_adj_2569)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_3_i860_3_lut_4_lut.init = 16'hf606;
    LUT4 n476_bdd_3_lut_24205_3_lut_4_lut (.A(n27429), .B(index_i[2]), .C(n491_adj_2570), 
         .D(index_i[4]), .Z(n25917)) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))+!A !(B ((D)+!C)+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n476_bdd_3_lut_24205_3_lut_4_lut.init = 16'h99f0;
    LUT4 i20833_3_lut (.A(n23192), .B(n26169), .C(index_q[6]), .Z(n23207)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20833_3_lut.init = 16'hcaca;
    LUT4 i19804_3_lut (.A(n364_adj_2571), .B(n890_adj_2523), .C(index_i[4]), 
         .Z(n22159)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19804_3_lut.init = 16'hcaca;
    LUT4 i20842_3_lut (.A(n23210), .B(n23211), .C(index_q[7]), .Z(n23216)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20842_3_lut.init = 16'hcaca;
    LUT4 i19803_3_lut (.A(n333_adj_2572), .B(n348_adj_2566), .C(index_i[4]), 
         .Z(n22158)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19803_3_lut.init = 16'hcaca;
    L6MUX21 i21187 (.D0(n23559), .D1(n23560), .SD(index_i[5]), .Z(n23561));
    LUT4 i20836_3_lut (.A(n26175), .B(n23199), .C(index_q[6]), .Z(n23210)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20836_3_lut.init = 16'hcaca;
    PFUMX i20150 (.BLUT(n22503), .ALUT(n22504), .C0(index_q[5]), .Z(n22505));
    LUT4 mux_229_Mux_2_i955_then_4_lut (.A(index_i[4]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n27508)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B (C+!(D))+!B !(C (D)))) */ ;
    defparam mux_229_Mux_2_i955_then_4_lut.init = 16'he95d;
    LUT4 mux_230_Mux_2_i348_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n348_adj_2573)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_2_i348_3_lut_4_lut_4_lut.init = 16'h52a5;
    LUT4 i19792_3_lut (.A(n491_adj_2574), .B(n541_adj_2420), .C(index_i[4]), 
         .Z(n22147)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19792_3_lut.init = 16'hcaca;
    LUT4 i21125_3_lut_4_lut (.A(n27229), .B(index_i[3]), .C(index_i[4]), 
         .D(n220_adj_2575), .Z(n23499)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21125_3_lut_4_lut.init = 16'hf808;
    PFUMX i20684 (.BLUT(n956), .ALUT(n20671), .C0(index_q[6]), .Z(n23058));
    LUT4 i19791_3_lut (.A(n397_adj_2410), .B(n475_adj_2576), .C(index_i[4]), 
         .Z(n22146)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19791_3_lut.init = 16'hcaca;
    LUT4 i21212_4_lut_4_lut (.A(n27131), .B(n27200), .C(index_i[5]), .D(index_i[4]), 
         .Z(n23586)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C+(D))+!B !(C (D)+!C !(D)))) */ ;
    defparam i21212_4_lut_4_lut.init = 16'hcf50;
    LUT4 i19648_3_lut (.A(n29934), .B(n308), .C(index_q[3]), .Z(n22003)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19648_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_3_i221_3_lut_4_lut (.A(n27229), .B(index_i[3]), .C(index_i[4]), 
         .D(n27185), .Z(n221_adj_2577)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_3_i221_3_lut_4_lut.init = 16'h08f8;
    LUT4 i19789_3_lut (.A(n251_adj_2335), .B(n443_adj_2346), .C(index_i[4]), 
         .Z(n22144)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19789_3_lut.init = 16'hcaca;
    LUT4 i19788_3_lut (.A(n397_adj_2410), .B(n15204), .C(index_i[4]), 
         .Z(n22143)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;
    defparam i19788_3_lut.init = 16'h3a3a;
    LUT4 i21121_3_lut_3_lut_4_lut (.A(n27229), .B(index_i[3]), .C(n93_adj_2578), 
         .D(index_i[4]), .Z(n23495)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21121_3_lut_3_lut_4_lut.init = 16'hf077;
    LUT4 mux_229_Mux_2_i955_else_4_lut (.A(index_i[4]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n27507)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+(D)))+!A !(B (C+!(D))+!B !(C+!(D))))) */ ;
    defparam mux_229_Mux_2_i955_else_4_lut.init = 16'h49c6;
    LUT4 n557_bdd_3_lut_24212_3_lut_4_lut (.A(n27229), .B(index_i[3]), .C(index_i[6]), 
         .D(n27156), .Z(n25628)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n557_bdd_3_lut_24212_3_lut_4_lut.init = 16'h08f8;
    LUT4 i22543_3_lut (.A(n27527), .B(n27530), .C(index_i[5]), .Z(n22136)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22543_3_lut.init = 16'hcaca;
    LUT4 n62_bdd_3_lut_4_lut_adj_81 (.A(n27322), .B(index_i[3]), .C(index_i[4]), 
         .D(n30_adj_2579), .Z(n25784)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n62_bdd_3_lut_4_lut_adj_81.init = 16'hf808;
    PFUMX i20693 (.BLUT(n94_adj_2580), .ALUT(n125_adj_2581), .C0(index_q[5]), 
          .Z(n23067));
    LUT4 i20944_3_lut_3_lut_4_lut_4_lut (.A(n27322), .B(index_i[3]), .C(index_i[4]), 
         .D(n27224), .Z(n23318)) /* synthesis lut_function=(!(A (B (C)+!B ((D)+!C))+!A (B+((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20944_3_lut_3_lut_4_lut_4_lut.init = 16'h0838;
    PFUMX i20694 (.BLUT(n18126), .ALUT(n14724), .C0(index_q[5]), .Z(n23068));
    LUT4 i9642_3_lut_4_lut_4_lut (.A(n27322), .B(index_i[3]), .C(index_i[5]), 
         .D(n27213), .Z(n12128)) /* synthesis lut_function=(A (B+(C (D)))+!A (B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9642_3_lut_4_lut_4_lut.init = 16'hf8c8;
    LUT4 i19776_3_lut (.A(n78), .B(n93_adj_2550), .C(index_i[4]), .Z(n22131)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19776_3_lut.init = 16'hcaca;
    LUT4 i19773_3_lut (.A(n15_adj_2341), .B(n526_adj_2315), .C(index_i[4]), 
         .Z(n22128)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19773_3_lut.init = 16'hcaca;
    L6MUX21 i20696 (.D0(n22034), .D1(n22037), .SD(index_q[5]), .Z(n23070));
    L6MUX21 i20697 (.D0(n22040), .D1(n22043), .SD(index_q[5]), .Z(n23071));
    PFUMX i20698 (.BLUT(n413_adj_2582), .ALUT(n444_adj_2514), .C0(index_q[5]), 
          .Z(n23072));
    LUT4 n954_bdd_3_lut_24160_4_lut_4_lut (.A(n27322), .B(index_i[3]), .C(index_i[4]), 
         .D(n27229), .Z(n25648)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C))+!A !(B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n954_bdd_3_lut_24160_4_lut_4_lut.init = 16'h838f;
    LUT4 i11401_2_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n668_adj_2583)) /* synthesis lut_function=(!(A ((D)+!B)+!A (B ((D)+!C)+!B (C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11401_2_lut_4_lut_4_lut_4_lut.init = 16'h00c9;
    LUT4 n638_bdd_3_lut_24474 (.A(n638), .B(n21824), .C(index_i[7]), .Z(n24945)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n638_bdd_3_lut_24474.init = 16'hcaca;
    LUT4 mux_230_Mux_7_i892_3_lut (.A(n62_adj_2269), .B(n891_adj_2288), 
         .C(index_q[5]), .Z(n892)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_7_i892_3_lut.init = 16'hcaca;
    LUT4 i19768_3_lut (.A(n747), .B(n762_adj_2326), .C(index_q[4]), .Z(n22123)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19768_3_lut.init = 16'hcaca;
    LUT4 i19767_3_lut (.A(n716_adj_2305), .B(n15090), .C(index_q[4]), 
         .Z(n22122)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19767_3_lut.init = 16'hcaca;
    PFUMX i20699 (.BLUT(n476_adj_2584), .ALUT(n507_adj_2585), .C0(index_q[5]), 
          .Z(n23073));
    PFUMX i20700 (.BLUT(n18113), .ALUT(n573_adj_2586), .C0(index_q[5]), 
          .Z(n23074));
    PFUMX i19991 (.BLUT(n22344), .ALUT(n22345), .C0(index_i[4]), .Z(n22346));
    LUT4 mux_229_Mux_1_i890_4_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[4]), 
         .C(n27385), .D(index_i[3]), .Z(n890_adj_2587)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A !(B+(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_1_i890_4_lut_4_lut_4_lut_4_lut.init = 16'h7477;
    PFUMX i20701 (.BLUT(n605_adj_2588), .ALUT(n636_adj_2589), .C0(index_q[5]), 
          .Z(n23075));
    PFUMX i19994 (.BLUT(n22347), .ALUT(n22348), .C0(index_i[4]), .Z(n22349));
    LUT4 i19765_3_lut (.A(n93_adj_2590), .B(n699_adj_2352), .C(index_q[4]), 
         .Z(n22120)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19765_3_lut.init = 16'hcaca;
    LUT4 i19764_3_lut (.A(n653_adj_2309), .B(n27097), .C(index_q[4]), 
         .Z(n22119)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19764_3_lut.init = 16'hcaca;
    PFUMX i20702 (.BLUT(n22046), .ALUT(n700_adj_2591), .C0(index_q[5]), 
          .Z(n23076));
    L6MUX21 i20703 (.D0(n732), .D1(n22049), .SD(index_q[5]), .Z(n23077));
    LUT4 n25411_bdd_3_lut (.A(n25411), .B(n476), .C(index_q[5]), .Z(n25412)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n25411_bdd_3_lut.init = 16'hcaca;
    PFUMX i20704 (.BLUT(n797_adj_2592), .ALUT(n828_adj_2593), .C0(index_q[5]), 
          .Z(n23078));
    LUT4 i19755_3_lut (.A(n397_adj_2594), .B(n475_adj_2329), .C(index_q[4]), 
         .Z(n22110)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19755_3_lut.init = 16'hcaca;
    LUT4 i15952_4_lut (.A(index_q[0]), .B(index_q[4]), .C(index_q[1]), 
         .D(n27307), .Z(n286)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i15952_4_lut.init = 16'hccc8;
    LUT4 n22003_bdd_3_lut (.A(n29916), .B(n29931), .C(index_q[3]), .Z(n26531)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n22003_bdd_3_lut.init = 16'hcaca;
    PFUMX i20705 (.BLUT(n860_adj_2595), .ALUT(n891_adj_2596), .C0(index_q[5]), 
          .Z(n23079));
    LUT4 mux_229_Mux_8_i892_3_lut_4_lut (.A(n27155), .B(index_i[4]), .C(index_i[5]), 
         .D(n860_adj_2597), .Z(n892_adj_2598)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_8_i892_3_lut_4_lut.init = 16'h4f40;
    LUT4 i21206_3_lut_4_lut_4_lut (.A(n27155), .B(index_i[4]), .C(index_i[5]), 
         .D(n27156), .Z(n23580)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C)+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21206_3_lut_4_lut_4_lut.init = 16'h0434;
    LUT4 i20517_3_lut (.A(n22885), .B(n22886), .C(index_i[7]), .Z(n22891)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20517_3_lut.init = 16'hcaca;
    LUT4 n25415_bdd_3_lut_25007 (.A(n27524), .B(n25413), .C(index_q[5]), 
         .Z(n25416)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n25415_bdd_3_lut_25007.init = 16'hcaca;
    L6MUX21 mux_229_Mux_7_i253 (.D0(n12145), .D1(n22397), .SD(index_i[5]), 
            .Z(n253)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    PFUMX mux_229_Mux_7_i190 (.BLUT(n22388), .ALUT(n173_adj_2599), .C0(index_i[5]), 
          .Z(n190_adj_2456)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 i22925_3_lut (.A(n22891), .B(n22892), .C(index_i[8]), .Z(n22894)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22925_3_lut.init = 16'hcaca;
    PFUMX i20724 (.BLUT(n94_adj_2600), .ALUT(n22055), .C0(index_q[5]), 
          .Z(n23098));
    PFUMX i19592 (.BLUT(n21945), .ALUT(n21946), .C0(index_q[5]), .Z(n21947));
    LUT4 i19696_3_lut (.A(n348_adj_2601), .B(n443_adj_2602), .C(index_q[4]), 
         .Z(n22051)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19696_3_lut.init = 16'hcaca;
    PFUMX i19595 (.BLUT(n21948), .ALUT(n21949), .C0(index_q[5]), .Z(n21950));
    LUT4 i19695_3_lut (.A(n397_adj_2594), .B(n731_adj_2603), .C(index_q[4]), 
         .Z(n22050)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19695_3_lut.init = 16'hcaca;
    LUT4 n21818_bdd_3_lut_23349 (.A(n382), .B(n509), .C(index_i[7]), .Z(n24947)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n21818_bdd_3_lut_23349.init = 16'hcaca;
    LUT4 i11848_2_lut_rep_588 (.A(index_q[0]), .B(index_q[1]), .Z(n27253)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i11848_2_lut_rep_588.init = 16'h2222;
    LUT4 i19702_3_lut (.A(n29941), .B(n29955), .C(index_q[3]), .Z(n22057)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19702_3_lut.init = 16'hcaca;
    PFUMX i20726 (.BLUT(n221_adj_2604), .ALUT(n252_adj_2605), .C0(index_q[5]), 
          .Z(n23100));
    LUT4 i21204_3_lut_4_lut_4_lut (.A(n27159), .B(index_i[4]), .C(index_i[5]), 
         .D(n27131), .Z(n23578)) /* synthesis lut_function=(A ((C+!(D))+!B)+!A (B (C+!(D))+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21204_3_lut_4_lut_4_lut.init = 16'he3ef;
    PFUMX i20009 (.BLUT(n22362), .ALUT(n22363), .C0(index_i[4]), .Z(n22364));
    PFUMX i20727 (.BLUT(n286_adj_2606), .ALUT(n22058), .C0(index_q[5]), 
          .Z(n23101));
    PFUMX i20728 (.BLUT(n349), .ALUT(n22061), .C0(index_q[5]), .Z(n23102));
    PFUMX i20012 (.BLUT(n22365), .ALUT(n22366), .C0(index_i[4]), .Z(n22367));
    LUT4 mux_229_Mux_2_i270_3_lut (.A(n29914), .B(n27392), .C(index_i[3]), 
         .Z(n270_adj_2453)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_2_i270_3_lut.init = 16'hcaca;
    LUT4 i9671_3_lut_then_4_lut (.A(index_q[4]), .B(index_q[0]), .C(index_q[1]), 
         .D(index_q[2]), .Z(n29966)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C+(D)))+!A (B (C+(D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i9671_3_lut_then_4_lut.init = 16'hd54a;
    LUT4 mux_229_Mux_0_i923_3_lut (.A(n27386), .B(n27432), .C(index_i[3]), 
         .Z(n923_adj_2607)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_0_i923_3_lut.init = 16'hcaca;
    LUT4 i9617_3_lut_4_lut (.A(index_q[0]), .B(n27334), .C(index_q[4]), 
         .D(n14), .Z(n12103)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i9617_3_lut_4_lut.init = 16'h4f40;
    PFUMX i19604 (.BLUT(n21957), .ALUT(n21958), .C0(index_q[5]), .Z(n21959));
    LUT4 i22884_3_lut (.A(n22858), .B(n22859), .C(index_i[8]), .Z(n22862)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22884_3_lut.init = 16'hcaca;
    LUT4 i9671_3_lut_else_4_lut (.A(index_q[4]), .B(index_q[0]), .C(index_q[1]), 
         .D(index_q[2]), .Z(n29965)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A !(B (D)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i9671_3_lut_else_4_lut.init = 16'ha955;
    PFUMX i20018 (.BLUT(n22371), .ALUT(n22372), .C0(index_i[4]), .Z(n22373));
    LUT4 i20483_3_lut_4_lut (.A(n27111), .B(n27117), .C(index_i[5]), .D(index_i[6]), 
         .Z(n22857)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (B+((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20483_3_lut_4_lut.init = 16'hffc5;
    PFUMX i20733 (.BLUT(n669_adj_2608), .ALUT(n700_adj_2609), .C0(index_q[5]), 
          .Z(n23107));
    LUT4 mux_230_Mux_2_i859_3_lut_4_lut (.A(index_q[0]), .B(n27334), .C(index_q[3]), 
         .D(n29948), .Z(n859_adj_2284)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_2_i859_3_lut_4_lut.init = 16'h4f40;
    LUT4 i19743_3_lut_4_lut (.A(index_q[0]), .B(n27334), .C(index_q[3]), 
         .D(n27279), .Z(n22098)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i19743_3_lut_4_lut.init = 16'hf404;
    PFUMX i20734 (.BLUT(n22526), .ALUT(n763_adj_2415), .C0(index_q[5]), 
          .Z(n23108));
    LUT4 i19797_3_lut_4_lut_4_lut (.A(n27213), .B(index_i[4]), .C(index_i[3]), 
         .D(n27224), .Z(n22152)) /* synthesis lut_function=(A (B (C)+!B !(C+!(D)))+!A (B (C)+!B (C+(D)))) */ ;
    defparam i19797_3_lut_4_lut_4_lut.init = 16'hd3d0;
    LUT4 i19689_3_lut_4_lut (.A(index_q[0]), .B(n27371), .C(index_q[3]), 
         .D(n27278), .Z(n22044)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A ((D)+!C)) */ ;
    defparam i19689_3_lut_4_lut.init = 16'hfd0d;
    LUT4 i20411_4_lut_4_lut (.A(n27127), .B(n27183), .C(index_q[5]), .D(index_q[4]), 
         .Z(n22785)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C+(D))+!B !(C (D)+!C !(D)))) */ ;
    defparam i20411_4_lut_4_lut.init = 16'hcf50;
    PFUMX i20735 (.BLUT(n22073), .ALUT(n828_adj_2610), .C0(index_q[5]), 
          .Z(n23109));
    PFUMX i20021 (.BLUT(n22374), .ALUT(n22375), .C0(index_i[4]), .Z(n22376));
    LUT4 i12391_3_lut_rep_829 (.A(index_i[2]), .B(index_i[1]), .C(index_i[0]), 
         .Z(n29956)) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12391_3_lut_rep_829.init = 16'hc4c4;
    LUT4 i21369_3_lut_4_lut (.A(n27113), .B(n27118), .C(index_q[5]), .D(index_q[6]), 
         .Z(n23743)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (B+((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i21369_3_lut_4_lut.init = 16'hffc5;
    PFUMX i20736 (.BLUT(n860_adj_2611), .ALUT(n22076), .C0(index_q[5]), 
          .Z(n23110));
    LUT4 i19930_3_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[1]), .C(index_i[0]), 
         .D(index_i[3]), .Z(n22285)) /* synthesis lut_function=(A (B (C)+!B !(C+!(D)))+!A (B (C+!(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19930_3_lut_4_lut_4_lut.init = 16'hc3c4;
    LUT4 mux_229_Mux_0_i716_3_lut (.A(n29921), .B(n27352), .C(index_i[3]), 
         .Z(n716_adj_2612)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_0_i716_3_lut.init = 16'hcaca;
    LUT4 n27434_bdd_4_lut_25557 (.A(n27434), .B(index_i[6]), .C(index_i[2]), 
         .D(index_i[5]), .Z(n27627)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A !(B (C+(D))+!B (D)))) */ ;
    defparam n27434_bdd_4_lut_25557.init = 16'h5fe0;
    LUT4 i20403_3_lut_4_lut_4_lut (.A(n27166), .B(index_q[4]), .C(index_q[5]), 
         .D(n27127), .Z(n22777)) /* synthesis lut_function=(A ((C+!(D))+!B)+!A (B (C+!(D))+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i20403_3_lut_4_lut_4_lut.init = 16'he3ef;
    LUT4 i19962_3_lut_3_lut_4_lut (.A(index_i[0]), .B(n27381), .C(n27214), 
         .D(index_i[3]), .Z(n22317)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(C+(D)))) */ ;
    defparam i19962_3_lut_3_lut_4_lut.init = 16'h77f0;
    PFUMX i19607 (.BLUT(n21960), .ALUT(n21961), .C0(index_q[5]), .Z(n21962));
    LUT4 mux_229_Mux_6_i939_3_lut_rep_407_3_lut_4_lut (.A(index_i[0]), .B(n27381), 
         .C(n27224), .D(index_i[3]), .Z(n27072)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(C+(D)))) */ ;
    defparam mux_229_Mux_6_i939_3_lut_rep_407_3_lut_4_lut.init = 16'h77f0;
    LUT4 i11892_3_lut_4_lut (.A(index_i[0]), .B(n27381), .C(n27335), .D(index_i[5]), 
         .Z(n318)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (C (D))) */ ;
    defparam i11892_3_lut_4_lut.init = 16'hf800;
    LUT4 mux_229_Mux_0_i653_3_lut (.A(n27385), .B(n27348), .C(index_i[3]), 
         .Z(n653_adj_2613)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_0_i653_3_lut.init = 16'hcaca;
    L6MUX21 i24954 (.D0(n26779), .D1(n26777), .SD(index_i[4]), .Z(n26780));
    PFUMX i19610 (.BLUT(n21963), .ALUT(n21964), .C0(index_q[5]), .Z(n21965));
    PFUMX i24952 (.BLUT(n27108), .ALUT(n26778), .C0(index_i[5]), .Z(n26779));
    LUT4 i20010_3_lut_3_lut_4_lut (.A(index_i[0]), .B(n27381), .C(index_i[3]), 
         .D(n27214), .Z(n22365)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A !(C+(D))) */ ;
    defparam i20010_3_lut_3_lut_4_lut.init = 16'h808f;
    LUT4 n986_bdd_4_lut_24083_4_lut_4_lut (.A(index_i[0]), .B(n27381), .C(index_i[4]), 
         .D(index_i[3]), .Z(n25262)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (D))+!A (B (C (D)+!C !(D))+!B (D)))) */ ;
    defparam n986_bdd_4_lut_24083_4_lut_4_lut.init = 16'h0c73;
    PFUMX i24950 (.BLUT(n26776), .ALUT(n26775), .C0(index_i[5]), .Z(n26777));
    LUT4 n21818_bdd_3_lut (.A(n21818), .B(n27629), .C(index_i[7]), .Z(n24948)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n21818_bdd_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_0_i620_3_lut (.A(n27435), .B(n29912), .C(index_i[3]), 
         .Z(n620_adj_2614)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_0_i620_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_6_i573_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[4]), .D(n572_adj_2615), .Z(n573_adj_2616)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_6_i573_3_lut_4_lut.init = 16'hf909;
    LUT4 mux_229_Mux_0_i589_3_lut (.A(n27432), .B(n588), .C(index_i[3]), 
         .Z(n589_adj_2617)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_0_i589_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_9_i124_3_lut_3_lut_4_lut (.A(n27340), .B(index_i[1]), 
         .C(index_i[3]), .D(n27229), .Z(n124_adj_2404)) /* synthesis lut_function=(!(A (C (D))+!A (B (C (D))+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_9_i124_3_lut_3_lut_4_lut.init = 16'h0efe;
    LUT4 mux_229_Mux_9_i364_3_lut_3_lut_4_lut (.A(n27340), .B(index_i[1]), 
         .C(index_i[3]), .D(n27224), .Z(n364_adj_2618)) /* synthesis lut_function=(!(A (C (D))+!A (B (C (D))+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_9_i364_3_lut_3_lut_4_lut.init = 16'h0efe;
    LUT4 i9641_4_lut_4_lut (.A(n27340), .B(index_i[1]), .C(index_i[3]), 
         .D(n21014), .Z(n12127)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A (B (C)+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9641_4_lut_4_lut.init = 16'h0e3e;
    LUT4 mux_230_Mux_3_i796_3_lut (.A(index_q[2]), .B(n731_adj_2603), .C(index_q[4]), 
         .Z(n796_adj_2619)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_3_i796_3_lut.init = 16'hacac;
    LUT4 mux_230_Mux_6_i731_3_lut (.A(n29931), .B(n27238), .C(index_q[3]), 
         .Z(n731_adj_2603)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_6_i731_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_5_i124_3_lut (.A(n14_adj_2290), .B(n27299), .C(index_q[3]), 
         .Z(n124_adj_2393)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_5_i124_3_lut.init = 16'hcaca;
    PFUMX i19613 (.BLUT(n21966), .ALUT(n21967), .C0(index_q[5]), .Z(n21968));
    LUT4 mux_229_Mux_0_i572_3_lut_4_lut (.A(n27340), .B(index_i[1]), .C(index_i[3]), 
         .D(n29923), .Z(n572_adj_2620)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_0_i572_3_lut_4_lut.init = 16'hefe0;
    LUT4 i19392_3_lut (.A(n588), .B(n29922), .C(index_i[3]), .Z(n21747)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19392_3_lut.init = 16'hcaca;
    PFUMX mux_229_Mux_8_i764 (.BLUT(n716_adj_2385), .ALUT(n732_adj_2621), 
          .C0(n22714), .Z(n764_adj_2480)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 i11889_2_lut_rep_421_3_lut_4_lut (.A(n27340), .B(index_i[1]), .C(index_i[4]), 
         .D(index_i[3]), .Z(n27086)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11889_2_lut_rep_421_3_lut_4_lut.init = 16'hfef0;
    LUT4 i20094_3_lut (.A(n27348), .B(n27394), .C(index_i[3]), .Z(n22449)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20094_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_3_i251_3_lut_4_lut (.A(n27340), .B(index_i[1]), .C(index_i[3]), 
         .D(n27224), .Z(n15004)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_3_i251_3_lut_4_lut.init = 16'hfe0e;
    LUT4 i21936_3_lut (.A(n22449), .B(n22450), .C(index_i[4]), .Z(n22451)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21936_3_lut.init = 16'hcaca;
    LUT4 n954_bdd_3_lut_23937_3_lut_4_lut (.A(n27340), .B(index_i[1]), .C(index_i[4]), 
         .D(index_i[3]), .Z(n25647)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n954_bdd_3_lut_23937_3_lut_4_lut.init = 16'hf10f;
    LUT4 i20091_3_lut (.A(n1001), .B(n588), .C(index_i[3]), .Z(n22446)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20091_3_lut.init = 16'hcaca;
    LUT4 i21938_3_lut (.A(n22446), .B(n22447), .C(index_i[4]), .Z(n22448)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21938_3_lut.init = 16'hcaca;
    PFUMX i20755 (.BLUT(n94_adj_2622), .ALUT(n125_adj_2623), .C0(index_q[5]), 
          .Z(n23129));
    LUT4 i19794_4_lut_4_lut_3_lut_4_lut (.A(n27340), .B(index_i[1]), .C(index_i[4]), 
         .D(index_i[3]), .Z(n22149)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19794_4_lut_4_lut_3_lut_4_lut.init = 16'h11ef;
    LUT4 mux_229_Mux_8_i475_3_lut_3_lut_4_lut (.A(n27340), .B(index_i[1]), 
         .C(index_i[3]), .D(n27229), .Z(n475_adj_2576)) /* synthesis lut_function=(A (C+!(D))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_8_i475_3_lut_3_lut_4_lut.init = 16'he0ef;
    PFUMX i20756 (.BLUT(n158_adj_2624), .ALUT(n189), .C0(index_q[5]), 
          .Z(n23130));
    LUT4 i21218_3_lut_3_lut (.A(n27440), .B(index_i[3]), .C(n29956), .Z(n23592)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam i21218_3_lut_3_lut.init = 16'h7474;
    LUT4 i19384_3_lut_3_lut (.A(n27440), .B(index_i[3]), .C(n1001), .Z(n21739)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam i19384_3_lut_3_lut.init = 16'h7474;
    LUT4 mux_229_Mux_7_i364_3_lut_3_lut (.A(n27440), .B(index_i[3]), .C(n27435), 
         .Z(n364_adj_2571)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;
    defparam mux_229_Mux_7_i364_3_lut_3_lut.init = 16'hd1d1;
    PFUMX i20757 (.BLUT(n221_adj_2432), .ALUT(n252_adj_2349), .C0(index_q[5]), 
          .Z(n23131));
    LUT4 mux_230_Mux_6_i891_3_lut (.A(n78_adj_2625), .B(n890_adj_2351), 
         .C(index_q[4]), .Z(n891_adj_2626)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_6_i891_3_lut.init = 16'hcaca;
    PFUMX i20758 (.BLUT(n286_adj_2627), .ALUT(n22085), .C0(index_q[5]), 
          .Z(n23132));
    LUT4 i15931_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n18117)) /* synthesis lut_function=(A (B)+!A !(B (C (D))+!B !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i15931_3_lut_4_lut_4_lut.init = 16'h9ccc;
    LUT4 mux_230_Mux_6_i828_4_lut (.A(n812_adj_2628), .B(n14376), .C(index_q[4]), 
         .D(index_q[2]), .Z(n828_adj_2629)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_6_i828_4_lut.init = 16'hfaca;
    LUT4 mux_230_Mux_6_i797_3_lut (.A(n653_adj_2317), .B(n27075), .C(index_q[4]), 
         .Z(n797_adj_2630)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_6_i797_3_lut.init = 16'hcaca;
    PFUMX i20759 (.BLUT(n349_adj_2631), .ALUT(n22088), .C0(index_q[5]), 
          .Z(n23133));
    PFUMX i21098 (.BLUT(n333_adj_2632), .ALUT(n348_adj_2363), .C0(index_q[4]), 
          .Z(n23472));
    LUT4 mux_229_Mux_5_i890_3_lut_3_lut (.A(n27440), .B(index_i[3]), .C(n27432), 
         .Z(n890_adj_2523)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam mux_229_Mux_5_i890_3_lut_3_lut.init = 16'h7474;
    LUT4 mux_230_Mux_6_i669_3_lut (.A(n653_adj_2633), .B(n668_adj_2634), 
         .C(index_q[4]), .Z(n669_adj_2635)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_6_i669_3_lut.init = 16'hcaca;
    PFUMX i20760 (.BLUT(n413_adj_2636), .ALUT(n444_adj_2637), .C0(index_q[5]), 
          .Z(n23134));
    LUT4 mux_229_Mux_4_i668_3_lut_3_lut (.A(n27440), .B(index_i[3]), .C(n29956), 
         .Z(n668_adj_2508)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;
    defparam mux_229_Mux_4_i668_3_lut_3_lut.init = 16'hd1d1;
    LUT4 mux_230_Mux_6_i158_3_lut (.A(n12053), .B(n157_adj_2516), .C(index_q[4]), 
         .Z(n158)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_6_i158_3_lut.init = 16'hcaca;
    PFUMX i20761 (.BLUT(n476_adj_2638), .ALUT(n507_adj_2639), .C0(index_q[5]), 
          .Z(n23135));
    PFUMX i20030 (.BLUT(n22383), .ALUT(n22384), .C0(index_i[4]), .Z(n22385));
    LUT4 n627_bdd_3_lut_24893 (.A(n27350), .B(n29923), .C(index_i[3]), 
         .Z(n26662)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n627_bdd_3_lut_24893.init = 16'hcaca;
    LUT4 mux_230_Mux_6_i542_3_lut (.A(n526_adj_2395), .B(n541), .C(index_q[4]), 
         .Z(n542_adj_2640)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_6_i542_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_0_i397_3_lut (.A(n27432), .B(n27387), .C(index_i[3]), 
         .Z(n397_adj_2641)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_0_i397_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_8_i653_3_lut_rep_409_3_lut_4_lut (.A(index_q[0]), .B(n27371), 
         .C(n27220), .D(index_q[3]), .Z(n27074)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(C+(D)))) */ ;
    defparam mux_230_Mux_8_i653_3_lut_rep_409_3_lut_4_lut.init = 16'h77f0;
    LUT4 n699_bdd_4_lut_24065_4_lut_4_lut (.A(index_q[0]), .B(n27371), .C(index_q[4]), 
         .D(index_q[3]), .Z(n25148)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (D))+!A (B (C (D)+!C !(D))+!B (D)))) */ ;
    defparam n699_bdd_4_lut_24065_4_lut_4_lut.init = 16'h0c73;
    LUT4 i20356_2_lut (.A(index_q[3]), .B(index_q[5]), .Z(n22730)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i20356_2_lut.init = 16'h8888;
    LUT4 i12736_2_lut_3_lut_4_lut (.A(n27123), .B(index_i[4]), .C(index_i[6]), 
         .D(index_i[5]), .Z(n15358)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12736_2_lut_3_lut_4_lut.init = 16'hfef0;
    PFUMX i21099 (.BLUT(n364_adj_2424), .ALUT(n379_adj_2345), .C0(index_q[4]), 
          .Z(n23473));
    LUT4 i19800_3_lut_3_lut_4_lut (.A(index_q[0]), .B(n27371), .C(n27219), 
         .D(index_q[3]), .Z(n22155)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(C+(D)))) */ ;
    defparam i19800_3_lut_3_lut_4_lut.init = 16'h77f0;
    LUT4 mux_229_Mux_10_i574_4_lut_4_lut (.A(n27123), .B(index_i[4]), .C(index_i[5]), 
         .D(n27108), .Z(n574_adj_2295)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_10_i574_4_lut_4_lut.init = 16'h1f1c;
    LUT4 mux_229_Mux_0_i188_3_lut (.A(n27442), .B(n931), .C(index_i[3]), 
         .Z(n188)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_0_i188_3_lut.init = 16'hcaca;
    LUT4 i11633_3_lut_4_lut (.A(index_q[0]), .B(n27371), .C(n27328), .D(index_q[5]), 
         .Z(n318_adj_2510)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (C (D))) */ ;
    defparam i11633_3_lut_4_lut.init = 16'hf800;
    LUT4 i19854_3_lut_3_lut_4_lut (.A(index_q[0]), .B(n27371), .C(index_q[3]), 
         .D(n27219), .Z(n22209)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A !(C+(D))) */ ;
    defparam i19854_3_lut_3_lut_4_lut.init = 16'h808f;
    PFUMX i20762 (.BLUT(n22091), .ALUT(n573_adj_2540), .C0(index_q[5]), 
          .Z(n23136));
    LUT4 index_i_5__bdd_4_lut_25624 (.A(n652), .B(index_i[2]), .C(index_i[3]), 
         .D(n27434), .Z(n26659)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (B+!(C (D))))) */ ;
    defparam index_i_5__bdd_4_lut_25624.init = 16'h3a0a;
    LUT4 mux_230_Mux_10_i574_4_lut_4_lut (.A(n27125), .B(index_q[4]), .C(index_q[5]), 
         .D(n27104), .Z(n574)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_10_i574_4_lut_4_lut.init = 16'h1f1c;
    LUT4 i12787_2_lut_3_lut_4_lut (.A(n27125), .B(index_q[4]), .C(index_q[6]), 
         .D(index_q[5]), .Z(n15412)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i12787_2_lut_3_lut_4_lut.init = 16'hfef0;
    PFUMX i20763 (.BLUT(n12091), .ALUT(n22094), .C0(index_q[5]), .Z(n23137));
    PFUMX i20764 (.BLUT(n669_adj_2642), .ALUT(n700_adj_2643), .C0(index_q[5]), 
          .Z(n23138));
    LUT4 mux_230_Mux_3_i251_3_lut_4_lut (.A(n27424), .B(index_q[1]), .C(index_q[3]), 
         .D(n27220), .Z(n15350)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_3_i251_3_lut_4_lut.init = 16'hfe0e;
    LUT4 mux_230_Mux_9_i364_3_lut_3_lut_4_lut (.A(n27424), .B(index_q[1]), 
         .C(index_q[3]), .D(n27220), .Z(n364_adj_2644)) /* synthesis lut_function=(!(A (C (D))+!A (B (C (D))+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_9_i364_3_lut_3_lut_4_lut.init = 16'h0efe;
    LUT4 i9560_4_lut_4_lut (.A(n27424), .B(index_q[1]), .C(index_q[3]), 
         .D(n21018), .Z(n12046)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A (B (C)+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i9560_4_lut_4_lut.init = 16'h0e3e;
    LUT4 n557_bdd_3_lut_23887_3_lut_4_lut (.A(n27424), .B(index_q[1]), .C(index_q[4]), 
         .D(index_q[3]), .Z(n25599)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam n557_bdd_3_lut_23887_3_lut_4_lut.init = 16'hf10f;
    LUT4 i21975_3_lut (.A(n26196), .B(n124_adj_2645), .C(index_i[4]), 
         .Z(n23496)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21975_3_lut.init = 16'hcaca;
    PFUMX i21100 (.BLUT(n397_adj_2646), .ALUT(n412_adj_2348), .C0(index_q[4]), 
          .Z(n23474));
    LUT4 mux_229_Mux_5_i731_3_lut (.A(n27393), .B(n27387), .C(index_i[3]), 
         .Z(n731_adj_2647)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_5_i731_3_lut.init = 16'hcaca;
    L6MUX21 i20765 (.D0(n22097), .D1(n763), .SD(index_q[5]), .Z(n23139));
    LUT4 n442_bdd_3_lut_24899 (.A(n27256), .B(n29956), .C(index_i[3]), 
         .Z(n26703)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n442_bdd_3_lut_24899.init = 16'hcaca;
    PFUMX i20767 (.BLUT(n860_adj_2648), .ALUT(n891_adj_2649), .C0(index_q[5]), 
          .Z(n23141));
    LUT4 i19984_3_lut_4_lut (.A(n27351), .B(index_i[2]), .C(index_i[3]), 
         .D(n29913), .Z(n22339)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19984_3_lut_4_lut.init = 16'hf606;
    L6MUX21 i24920 (.D0(n26728), .D1(n26725), .SD(index_i[5]), .Z(n26729));
    PFUMX i20768 (.BLUT(n924_adj_2650), .ALUT(n22100), .C0(index_q[5]), 
          .Z(n23142));
    PFUMX i24918 (.BLUT(n26727), .ALUT(n26726), .C0(index_i[4]), .Z(n26728));
    LUT4 i11602_2_lut_rep_399_3_lut_4_lut (.A(n27127), .B(index_q[4]), .C(index_q[6]), 
         .D(index_q[5]), .Z(n27064)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;
    defparam i11602_2_lut_rep_399_3_lut_4_lut.init = 16'hf080;
    LUT4 n269_bdd_3_lut_23798 (.A(n29948), .B(index_q[3]), .C(n27276), 
         .Z(n25515)) /* synthesis lut_function=(A (B+(C))+!A !(B+!(C))) */ ;
    defparam n269_bdd_3_lut_23798.init = 16'hb8b8;
    PFUMX i20769 (.BLUT(n22103), .ALUT(n1018_adj_2532), .C0(index_q[5]), 
          .Z(n23143));
    LUT4 mux_230_Mux_0_i572_3_lut_4_lut (.A(n27424), .B(index_q[1]), .C(index_q[3]), 
         .D(n27277), .Z(n572)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_0_i572_3_lut_4_lut.init = 16'hefe0;
    PFUMX i21101 (.BLUT(n428), .ALUT(n443), .C0(index_q[4]), .Z(n23475));
    LUT4 i19363_3_lut_4_lut (.A(n27351), .B(index_i[2]), .C(index_i[3]), 
         .D(n27387), .Z(n21718)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19363_3_lut_4_lut.init = 16'h6f60;
    PFUMX i19616 (.BLUT(n21969), .ALUT(n21970), .C0(index_q[5]), .Z(n21971));
    PFUMX mux_229_Mux_8_i574 (.BLUT(n542), .ALUT(n12127), .C0(index_i[5]), 
          .Z(n574_adj_2478)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 mux_229_Mux_3_i747_3_lut (.A(n27256), .B(n498), .C(index_i[3]), 
         .Z(n747_adj_2651)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_3_i747_3_lut.init = 16'hcaca;
    LUT4 i19608_4_lut_4_lut_3_lut_4_lut (.A(n27424), .B(index_q[1]), .C(index_q[4]), 
         .D(index_q[3]), .Z(n21963)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i19608_4_lut_4_lut_3_lut_4_lut.init = 16'h11ef;
    LUT4 i11575_2_lut_rep_422_3_lut_4_lut (.A(n27424), .B(index_q[1]), .C(index_q[4]), 
         .D(index_q[3]), .Z(n27087)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i11575_2_lut_rep_422_3_lut_4_lut.init = 16'hfef0;
    LUT4 mux_229_Mux_6_i285_3_lut_4_lut (.A(n27351), .B(index_i[2]), .C(index_i[3]), 
         .D(n27345), .Z(n285_adj_2489)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_6_i285_3_lut_4_lut.init = 16'hf606;
    L6MUX21 i21223 (.D0(n23595), .D1(n23596), .SD(index_i[5]), .Z(n23597));
    LUT4 mux_229_Mux_3_i460_3_lut_4_lut (.A(n27351), .B(index_i[2]), .C(index_i[3]), 
         .D(n29922), .Z(n460_adj_2488)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_3_i460_3_lut_4_lut.init = 16'h6f60;
    PFUMX i20787 (.BLUT(n158_adj_2652), .ALUT(n189_adj_2512), .C0(index_q[5]), 
          .Z(n23161));
    PFUMX i20039 (.BLUT(n22392), .ALUT(n22393), .C0(index_i[4]), .Z(n22394));
    L6MUX21 i23810 (.D0(n25525), .D1(n25522), .SD(index_q[5]), .Z(n25526));
    PFUMX i23808 (.BLUT(n25524), .ALUT(n475_adj_2653), .C0(index_q[4]), 
          .Z(n25525));
    PFUMX i20788 (.BLUT(n221_adj_2654), .ALUT(n22109), .C0(index_q[5]), 
          .Z(n23162));
    LUT4 mux_230_Mux_1_i924_3_lut (.A(n908_adj_2297), .B(n412_adj_2294), 
         .C(index_q[4]), .Z(n924_adj_2655)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_1_i924_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_8_i173_3_lut_3_lut_4_lut (.A(n27296), .B(index_q[2]), 
         .C(n954_adj_2285), .D(index_q[4]), .Z(n173_adj_2387)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_8_i173_3_lut_3_lut_4_lut.init = 16'hf077;
    PFUMX i20042 (.BLUT(n22395), .ALUT(n22396), .C0(index_i[4]), .Z(n22397));
    LUT4 n27628_bdd_3_lut (.A(n27628), .B(n27625), .C(index_i[4]), .Z(n27629)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n27628_bdd_3_lut.init = 16'hcaca;
    PFUMX i20789 (.BLUT(n286_adj_2656), .ALUT(n317_adj_2657), .C0(index_q[5]), 
          .Z(n23163));
    LUT4 i22309_3_lut (.A(n22233), .B(n22234), .C(index_q[4]), .Z(n22235)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22309_3_lut.init = 16'hcaca;
    LUT4 n285_bdd_3_lut_adj_82 (.A(n29948), .B(n27280), .C(index_q[3]), 
         .Z(n25518)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n285_bdd_3_lut_adj_82.init = 16'hacac;
    PFUMX i20790 (.BLUT(n349_adj_2658), .ALUT(n22115), .C0(index_q[5]), 
          .Z(n23164));
    LUT4 mux_230_Mux_8_i78_3_lut_4_lut (.A(n27296), .B(index_q[2]), .C(index_q[3]), 
         .D(n29936), .Z(n78_adj_2625)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_8_i78_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_230_Mux_1_i349_3_lut (.A(n506_adj_2304), .B(n348_adj_2659), 
         .C(index_q[4]), .Z(n349_adj_2660)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_1_i349_3_lut.init = 16'hcaca;
    LUT4 i20350_2_lut (.A(index_i[3]), .B(index_i[5]), .Z(n22724)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20350_2_lut.init = 16'h8888;
    LUT4 i22318_3_lut (.A(n22194), .B(n22195), .C(index_q[4]), .Z(n22196)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22318_3_lut.init = 16'hcaca;
    LUT4 i11484_3_lut (.A(index_i[3]), .B(index_i[1]), .C(index_i[0]), 
         .Z(n14081)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11484_3_lut.init = 16'hecec;
    PFUMX i20791 (.BLUT(n413_adj_2661), .ALUT(n22157), .C0(index_q[5]), 
          .Z(n23165));
    PFUMX mux_229_Mux_1_i636 (.BLUT(n620_adj_2551), .ALUT(n635), .C0(index_i[4]), 
          .Z(n636_adj_2662)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    PFUMX i24915 (.BLUT(n26724), .ALUT(n316_adj_2316), .C0(index_i[4]), 
          .Z(n26725));
    PFUMX i20792 (.BLUT(n22163), .ALUT(n507_adj_2663), .C0(index_q[5]), 
          .Z(n23166));
    LUT4 i19878_3_lut_3_lut_4_lut (.A(n27296), .B(index_q[2]), .C(n38), 
         .D(index_q[3]), .Z(n22233)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i19878_3_lut_3_lut_4_lut.init = 16'hf077;
    PFUMX i20793 (.BLUT(n22169), .ALUT(n573_adj_2538), .C0(index_q[5]), 
          .Z(n23167));
    LUT4 mux_230_Mux_1_i94_3_lut (.A(index_q[0]), .B(n93_adj_2664), .C(index_q[4]), 
         .Z(n94_adj_2665)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_1_i94_3_lut.init = 16'hcaca;
    LUT4 n22024_bdd_3_lut_24381 (.A(n27275), .B(n27277), .C(index_q[3]), 
         .Z(n25521)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n22024_bdd_3_lut_24381.init = 16'hcaca;
    PFUMX i21102 (.BLUT(n460_adj_2354), .ALUT(n475_adj_2400), .C0(index_q[4]), 
          .Z(n23476));
    LUT4 mux_229_Mux_3_i781_3_lut (.A(n27386), .B(n27383), .C(index_i[3]), 
         .Z(n781_adj_2568)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_3_i781_3_lut.init = 16'hcaca;
    PFUMX i20794 (.BLUT(n605_adj_2666), .ALUT(n22175), .C0(index_q[5]), 
          .Z(n23168));
    LUT4 n627_bdd_3_lut (.A(n27350), .B(n588), .C(index_i[3]), .Z(n26705)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n627_bdd_3_lut.init = 16'hacac;
    PFUMX i20795 (.BLUT(n669_adj_2667), .ALUT(n700_adj_2526), .C0(index_q[5]), 
          .Z(n23169));
    PFUMX i20796 (.BLUT(n732_adj_2668), .ALUT(n763_adj_2669), .C0(index_q[5]), 
          .Z(n23170));
    LUT4 mux_229_Mux_5_i124_3_lut (.A(n27385), .B(n27438), .C(index_i[3]), 
         .Z(n124_adj_2542)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_5_i124_3_lut.init = 16'hcaca;
    LUT4 i23063_2_lut_rep_419_3_lut_4_lut (.A(n27296), .B(index_q[2]), .C(index_q[5]), 
         .D(n27328), .Z(n27084)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i23063_2_lut_rep_419_3_lut_4_lut.init = 16'h0f7f;
    LUT4 i11871_2_lut_rep_401_3_lut_4_lut (.A(n27131), .B(index_i[4]), .C(index_i[6]), 
         .D(index_i[5]), .Z(n27066)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11871_2_lut_rep_401_3_lut_4_lut.init = 16'hf080;
    LUT4 mux_229_Mux_0_i525_3_lut_3_lut_rep_795 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29922)) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_0_i525_3_lut_3_lut_rep_795.init = 16'h6a6a;
    LUT4 i22347_3_lut (.A(n716_adj_2302), .B(n731_adj_2670), .C(index_q[4]), 
         .Z(n732_adj_2668)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22347_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_2_i669_3_lut (.A(n653_adj_2671), .B(n475_adj_2653), 
         .C(index_q[4]), .Z(n669_adj_2667)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_2_i669_3_lut.init = 16'hcaca;
    L6MUX21 i20798 (.D0(n860), .D1(n891), .SD(index_q[5]), .Z(n23172));
    PFUMX i20045 (.BLUT(n22398), .ALUT(n22399), .C0(index_i[4]), .Z(n22400));
    LUT4 mux_230_Mux_2_i605_3_lut (.A(n142_adj_2672), .B(n604_adj_2673), 
         .C(index_q[4]), .Z(n605_adj_2666)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_2_i605_3_lut.init = 16'hcaca;
    L6MUX21 i21230 (.D0(n23602), .D1(n23603), .SD(index_i[5]), .Z(n23604));
    LUT4 n316_bdd_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[3]), .C(index_i[1]), 
         .D(index_i[2]), .Z(n26724)) /* synthesis lut_function=(!(A (B+(C (D)+!C !(D)))+!A !(B+!((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n316_bdd_3_lut_3_lut_4_lut.init = 16'h4674;
    LUT4 i22352_3_lut (.A(n29959), .B(n22168), .C(index_q[4]), .Z(n22169)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22352_3_lut.init = 16'hcaca;
    LUT4 i22354_3_lut (.A(n22161), .B(n22162), .C(index_q[4]), .Z(n22163)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22354_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_2_i413_3_lut (.A(n397_adj_2674), .B(n954_adj_2285), 
         .C(index_q[4]), .Z(n413_adj_2661)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_2_i413_3_lut.init = 16'hcaca;
    L6MUX21 i21237 (.D0(n23609), .D1(n23610), .SD(index_i[5]), .Z(n23611));
    LUT4 i20041_3_lut (.A(n27435), .B(n851), .C(index_i[3]), .Z(n22396)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20041_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_2_i317_3_lut (.A(n668_adj_2412), .B(n316_adj_2675), 
         .C(index_q[4]), .Z(n317_adj_2657)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_2_i317_3_lut.init = 16'hcaca;
    PFUMX i21103 (.BLUT(n491_adj_2676), .ALUT(n11325), .C0(index_q[4]), 
          .Z(n23477));
    LUT4 mux_230_Mux_2_i286_3_lut (.A(n270_adj_2677), .B(n653_adj_2678), 
         .C(index_q[4]), .Z(n286_adj_2656)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_2_i286_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_2_i491_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n491_adj_2679)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A !(B (C)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_2_i491_3_lut_4_lut_4_lut.init = 16'h6a5a;
    L6MUX21 i24896 (.D0(n26706), .D1(n26704), .SD(index_i[5]), .Z(n26707));
    LUT4 i20040_3_lut (.A(n29914), .B(n27386), .C(index_i[3]), .Z(n22395)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20040_3_lut.init = 16'hcaca;
    LUT4 n308_bdd_3_lut_24384 (.A(n27289), .B(n27426), .C(index_q[3]), 
         .Z(n25524)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n308_bdd_3_lut_24384.init = 16'hacac;
    PFUMX i24894 (.BLUT(n572_adj_2680), .ALUT(n26705), .C0(index_i[4]), 
          .Z(n26706));
    LUT4 i22363_3_lut (.A(n142_adj_2301), .B(n14388), .C(index_q[4]), 
         .Z(n158_adj_2652)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22363_3_lut.init = 16'hcaca;
    LUT4 i20038_3_lut (.A(n29922), .B(n27342), .C(index_i[3]), .Z(n22393)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20038_3_lut.init = 16'hcaca;
    LUT4 n389_bdd_3_lut_24917 (.A(n27439), .B(n29956), .C(index_i[3]), 
         .Z(n26726)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n389_bdd_3_lut_24917.init = 16'hcaca;
    LUT4 i19615_3_lut (.A(n364), .B(n379), .C(index_q[4]), .Z(n21970)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19615_3_lut.init = 16'hcaca;
    LUT4 i19614_3_lut (.A(n333_adj_2681), .B(n348_adj_2601), .C(index_q[4]), 
         .Z(n21969)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19614_3_lut.init = 16'hcaca;
    LUT4 i22368_3_lut (.A(n22101), .B(n27470), .C(index_q[4]), .Z(n22103)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22368_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_3_i924_3_lut (.A(n908_adj_2682), .B(index_q[0]), .C(index_q[4]), 
         .Z(n924_adj_2650)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_3_i924_3_lut.init = 16'hcaca;
    PFUMX i23805 (.BLUT(n25521), .ALUT(n22024), .C0(index_q[4]), .Z(n25522));
    LUT4 mux_230_Mux_4_i900_3_lut_4_lut_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n900)) /* synthesis lut_function=(A ((C)+!B)+!A !(B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_4_i900_3_lut_4_lut_3_lut.init = 16'hb2b2;
    LUT4 mux_230_Mux_3_i891_3_lut (.A(n541), .B(n890_adj_2364), .C(index_q[4]), 
         .Z(n891_adj_2649)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_3_i891_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_0_i397_3_lut (.A(n29935), .B(n27280), .C(index_q[3]), 
         .Z(n397_adj_2646)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_0_i397_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_3_i669_3_lut (.A(n653_adj_2678), .B(n668_adj_2412), 
         .C(index_q[4]), .Z(n669_adj_2642)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_3_i669_3_lut.init = 16'hcaca;
    LUT4 i9605_4_lut (.A(n27371), .B(n27172), .C(index_q[3]), .D(index_q[4]), 
         .Z(n12091)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B ((D)+!C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i9605_4_lut.init = 16'h3afa;
    LUT4 i20032_3_lut (.A(n27435), .B(n27385), .C(index_i[3]), .Z(n22387)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20032_3_lut.init = 16'hcaca;
    LUT4 i20031_3_lut (.A(n27442), .B(n851), .C(index_i[3]), .Z(n22386)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20031_3_lut.init = 16'hcaca;
    PFUMX i20817 (.BLUT(n94_adj_2665), .ALUT(n22184), .C0(index_q[5]), 
          .Z(n23191));
    LUT4 mux_229_Mux_7_i173_3_lut (.A(n29914), .B(n27385), .C(index_i[3]), 
         .Z(n173_adj_2599)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_7_i173_3_lut.init = 16'hcaca;
    LUT4 i22377_3_lut (.A(n22089), .B(n22090), .C(index_q[4]), .Z(n22091)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22377_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_6_i653_3_lut (.A(n29929), .B(n619), .C(index_q[3]), 
         .Z(n653_adj_2633)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_6_i653_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_3_i476_3_lut (.A(n460_adj_2683), .B(n285_adj_2684), 
         .C(index_q[4]), .Z(n476_adj_2638)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_3_i476_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_5_i397_3_lut (.A(n29949), .B(n332), .C(index_q[3]), 
         .Z(n397_adj_2685)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_5_i397_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_5_i506_3_lut (.A(n29955), .B(n29940), .C(index_q[3]), 
         .Z(n506_adj_2686)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_5_i506_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_3_i413_3_lut (.A(n397_adj_2437), .B(n27310), .C(index_q[4]), 
         .Z(n413_adj_2636)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_3_i413_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_3_i286_4_lut (.A(n93_adj_2687), .B(index_q[2]), .C(index_q[4]), 
         .D(n15111), .Z(n286_adj_2627)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_3_i286_4_lut.init = 16'h3aca;
    LUT4 mux_230_Mux_5_i15_3_lut (.A(n29916), .B(n27425), .C(index_q[3]), 
         .Z(n15_adj_2464)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_5_i15_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_3_i158_3_lut (.A(n142_adj_2672), .B(n157_adj_2298), 
         .C(index_q[4]), .Z(n158_adj_2624)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_3_i158_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_5_i859_3_lut (.A(n308), .B(n29916), .C(index_q[3]), 
         .Z(n859_adj_2688)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_5_i859_3_lut.init = 16'hcaca;
    L6MUX21 i23803 (.D0(n25519), .D1(n25517), .SD(index_q[5]), .Z(n25520));
    L6MUX21 i20818 (.D0(n22187), .D1(n22193), .SD(index_q[5]), .Z(n23192));
    LUT4 mux_230_Mux_5_i875_3_lut (.A(n14_adj_2290), .B(n29934), .C(index_q[3]), 
         .Z(n875_adj_2689)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_5_i875_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_3_i125_3_lut (.A(n46_adj_2481), .B(n526_adj_2384), 
         .C(index_q[4]), .Z(n125_adj_2623)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_3_i125_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_8_i732_3_lut (.A(index_i[3]), .B(n15218), .C(index_i[5]), 
         .Z(n732_adj_2621)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_8_i732_3_lut.init = 16'h3a3a;
    LUT4 mux_230_Mux_4_i61_3_lut (.A(n27278), .B(n27311), .C(index_q[3]), 
         .Z(n61_adj_2467)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_4_i61_3_lut.init = 16'hcaca;
    PFUMX i23801 (.BLUT(n25518), .ALUT(n285_adj_2684), .C0(index_q[4]), 
          .Z(n25519));
    PFUMX i20820 (.BLUT(n22196), .ALUT(n317_adj_2690), .C0(index_q[5]), 
          .Z(n23194));
    PFUMX i24891 (.BLUT(n26703), .ALUT(n26702), .C0(index_i[4]), .Z(n26704));
    PFUMX i20821 (.BLUT(n349_adj_2660), .ALUT(n22202), .C0(index_q[5]), 
          .Z(n23195));
    L6MUX21 i20822 (.D0(n22205), .D1(n22211), .SD(index_q[5]), .Z(n23196));
    L6MUX21 i20823 (.D0(n22214), .D1(n22226), .SD(index_q[5]), .Z(n23197));
    LUT4 mux_229_Mux_2_i316_3_lut (.A(n29911), .B(n29922), .C(index_i[3]), 
         .Z(n316_adj_2451)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_2_i316_3_lut.init = 16'hcaca;
    LUT4 i20738_4_lut (.A(n27466), .B(n1002_adj_2691), .C(index_q[5]), 
         .D(index_q[4]), .Z(n23112)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;
    defparam i20738_4_lut.init = 16'hfaca;
    LUT4 n77_bdd_3_lut_24949 (.A(n27345), .B(n29923), .C(index_i[3]), 
         .Z(n26775)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n77_bdd_3_lut_24949.init = 16'hacac;
    PFUMX i20048 (.BLUT(n22401), .ALUT(n22402), .C0(index_i[4]), .Z(n22403));
    L6MUX21 i20825 (.D0(n22232), .D1(n636), .SD(index_q[5]), .Z(n23199));
    PFUMX i20826 (.BLUT(n22235), .ALUT(n700_adj_2389), .C0(index_q[5]), 
          .Z(n23200));
    LUT4 mux_230_Mux_4_i270_3_lut (.A(n29918), .B(n29955), .C(index_q[3]), 
         .Z(n270_adj_2692)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_4_i270_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_4_i15_3_lut (.A(n29940), .B(n14), .C(index_q[3]), 
         .Z(n15_adj_2469)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_4_i15_3_lut.init = 16'hcaca;
    PFUMX i23799 (.BLUT(n25516), .ALUT(n25515), .C0(index_q[4]), .Z(n25517));
    L6MUX21 i20828 (.D0(n22238), .D1(n22241), .SD(index_q[5]), .Z(n23202));
    LUT4 i19606_3_lut (.A(n491_adj_2693), .B(n506_adj_2304), .C(index_q[4]), 
         .Z(n21961)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19606_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_4_i348_3_lut (.A(n27291), .B(n29953), .C(index_q[3]), 
         .Z(n348)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_4_i348_3_lut.init = 16'hcaca;
    PFUMX i26899 (.BLUT(n29965), .ALUT(n29966), .C0(index_q[3]), .Z(n29967));
    LUT4 mux_229_Mux_0_i660_3_lut_rep_677 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27342)) /* synthesis lut_function=(A (B)+!A (B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_0_i660_3_lut_rep_677.init = 16'hc9c9;
    PFUMX i20830 (.BLUT(n924_adj_2655), .ALUT(n22247), .C0(index_q[5]), 
          .Z(n23204));
    LUT4 i21315_3_lut_4_lut_4_lut (.A(n27181), .B(index_q[5]), .C(index_q[4]), 
         .D(n27126), .Z(n23689)) /* synthesis lut_function=(A (B+(C (D)))+!A (B+((D)+!C))) */ ;
    defparam i21315_3_lut_4_lut_4_lut.init = 16'hfdcd;
    PFUMX i20831 (.BLUT(n987), .ALUT(n22250), .C0(index_q[5]), .Z(n23205));
    LUT4 i19605_3_lut (.A(n397_adj_2539), .B(n475_adj_2505), .C(index_q[4]), 
         .Z(n21960)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19605_3_lut.init = 16'hcaca;
    PFUMX mux_229_Mux_2_i891 (.BLUT(n875_adj_2314), .ALUT(n890_adj_2694), 
          .C0(index_i[4]), .Z(n891_adj_2695)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 mux_230_Mux_4_i860_3_lut (.A(n506_adj_2686), .B(n25710), .C(index_q[4]), 
         .Z(n860_adj_2611)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_4_i860_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_4_i684_3_lut (.A(n619), .B(n108), .C(index_q[3]), 
         .Z(n684_adj_2696)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_4_i684_3_lut.init = 16'hcaca;
    LUT4 i22397_3_lut (.A(n22071), .B(n22072), .C(index_q[4]), .Z(n22073)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22397_3_lut.init = 16'hcaca;
    LUT4 i22399_3_lut (.A(n22524), .B(n22525), .C(index_q[4]), .Z(n22526)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22399_3_lut.init = 16'hcaca;
    LUT4 i20017_3_lut (.A(n29944), .B(n27347), .C(index_i[3]), .Z(n22372)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20017_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_4_i700_3_lut (.A(n684_adj_2696), .B(index_q[1]), .C(index_q[4]), 
         .Z(n700_adj_2609)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_4_i700_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_4_i669_3_lut (.A(n653_adj_2317), .B(n668), .C(index_q[4]), 
         .Z(n669_adj_2608)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_4_i669_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_4_i542_3_lut (.A(n526_adj_2384), .B(n506_adj_2304), 
         .C(index_q[4]), .Z(n542_adj_2697)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_4_i542_3_lut.init = 16'hcaca;
    LUT4 i20732_4_lut (.A(n27181), .B(n27463), .C(index_q[5]), .D(index_q[4]), 
         .Z(n23106)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam i20732_4_lut.init = 16'hc5ca;
    LUT4 i19603_3_lut (.A(n251_adj_2342), .B(n443_adj_2344), .C(index_q[4]), 
         .Z(n21958)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19603_3_lut.init = 16'hcaca;
    LUT4 i19602_3_lut (.A(n397_adj_2539), .B(n15090), .C(index_q[4]), 
         .Z(n21957)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;
    defparam i19602_3_lut.init = 16'h3a3a;
    PFUMX mux_229_Mux_2_i860 (.BLUT(n844_adj_2320), .ALUT(n859_adj_2698), 
          .C0(index_i[4]), .Z(n860_adj_2699)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 mux_229_Mux_5_i939_3_lut_4_lut (.A(n27434), .B(index_i[2]), .C(index_i[4]), 
         .D(n954_adj_2331), .Z(n939_adj_2433)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C)) */ ;
    defparam mux_229_Mux_5_i939_3_lut_4_lut.init = 16'hf707;
    LUT4 i23088_2_lut (.A(index_i[5]), .B(index_i[4]), .Z(n22714)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i23088_2_lut.init = 16'heeee;
    LUT4 mux_230_Mux_4_i286_3_lut (.A(n270_adj_2692), .B(n15_adj_2469), 
         .C(index_q[4]), .Z(n286_adj_2606)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_4_i286_3_lut.init = 16'hcaca;
    LUT4 i20007_3_lut (.A(n29922), .B(n27393), .C(index_i[3]), .Z(n22362)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20007_3_lut.init = 16'hcaca;
    LUT4 i20034_3_lut_3_lut_4_lut (.A(n27434), .B(index_i[2]), .C(n1001), 
         .D(index_i[3]), .Z(n22389)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C+!(D))) */ ;
    defparam i20034_3_lut_3_lut_4_lut.init = 16'hf077;
    LUT4 i22614_3_lut (.A(n29963), .B(n27503), .C(index_q[5]), .Z(n21953)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22614_3_lut.init = 16'hcaca;
    LUT4 i19593_3_lut (.A(n78_adj_2625), .B(n93_adj_2590), .C(index_q[4]), 
         .Z(n21948)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19593_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_8_i78_3_lut_4_lut (.A(n27434), .B(index_i[2]), .C(index_i[3]), 
         .D(n27430), .Z(n78)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam mux_229_Mux_8_i78_3_lut_4_lut.init = 16'h8f80;
    LUT4 i19590_3_lut (.A(n15_adj_2700), .B(n526_adj_2384), .C(index_q[4]), 
         .Z(n21945)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19590_3_lut.init = 16'hcaca;
    PFUMX mux_229_Mux_3_i763 (.BLUT(n747_adj_2651), .ALUT(n762_adj_2303), 
          .C0(index_i[4]), .Z(n763_adj_2701)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 mux_230_Mux_4_i94_3_lut (.A(n61_adj_2467), .B(n27309), .C(index_q[4]), 
         .Z(n94_adj_2600)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_4_i94_3_lut.init = 16'hcaca;
    LUT4 i12490_3_lut_rep_831 (.A(index_q[2]), .B(index_q[1]), .C(index_q[0]), 
         .Z(n29958)) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i12490_3_lut_rep_831.init = 16'hc4c4;
    LUT4 i12504_3_lut (.A(index_q[3]), .B(index_q[1]), .C(index_q[0]), 
         .Z(n15111)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i12504_3_lut.init = 16'hc8c8;
    LUT4 i22419_3_lut (.A(n22386), .B(n22387), .C(index_i[4]), .Z(n22388)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i22419_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_3_i348_3_lut (.A(n27426), .B(n29919), .C(index_q[3]), 
         .Z(n348_adj_2702)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_3_i348_3_lut.init = 16'hcaca;
    LUT4 i23152_2_lut_rep_420_3_lut_4_lut (.A(n27434), .B(index_i[2]), .C(index_i[5]), 
         .D(n27335), .Z(n27085)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A (C (D)))) */ ;
    defparam i23152_2_lut_rep_420_3_lut_4_lut.init = 16'h0f7f;
    LUT4 i21953_3_lut (.A(n22356), .B(n22357), .C(index_i[4]), .Z(n22358)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21953_3_lut.init = 16'hcaca;
    LUT4 i22026_3_lut (.A(n27500), .B(n124_adj_2703), .C(index_q[4]), 
         .Z(n23465)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22026_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_3_i908_3_lut (.A(n27279), .B(n27311), .C(index_q[3]), 
         .Z(n908_adj_2682)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_3_i908_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_7_i333_3_lut (.A(n27297), .B(n14_adj_2290), .C(index_q[3]), 
         .Z(n333_adj_2681)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_7_i333_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_5_i891_3_lut (.A(n875_adj_2689), .B(n379), .C(index_q[4]), 
         .Z(n891_adj_2596)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_5_i891_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_2_i397_3_lut (.A(n29956), .B(n27386), .C(index_i[3]), 
         .Z(n397_adj_2449)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_2_i397_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_5_i860_3_lut (.A(n15_adj_2464), .B(n859_adj_2688), 
         .C(index_q[4]), .Z(n860_adj_2595)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_5_i860_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_7_i348_3_lut (.A(n29934), .B(n29935), .C(index_q[3]), 
         .Z(n348_adj_2601)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_7_i348_3_lut.init = 16'hcaca;
    LUT4 n557_bdd_2_lut_3_lut_4_lut (.A(n27434), .B(index_i[2]), .C(index_i[6]), 
         .D(index_i[3]), .Z(n25629)) /* synthesis lut_function=(A (B (C)+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D))) */ ;
    defparam n557_bdd_2_lut_3_lut_4_lut.init = 16'hf087;
    LUT4 mux_229_Mux_0_i963_3_lut_3_lut_rep_796 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29923)) /* synthesis lut_function=(!(A (B)+!A (B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_0_i963_3_lut_3_lut_rep_796.init = 16'h3636;
    LUT4 i1_3_lut_adj_83 (.A(index_i[0]), .B(index_i[4]), .C(index_i[2]), 
         .Z(n21014)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_3_lut_adj_83.init = 16'hfefe;
    PFUMX i20078 (.BLUT(n22431), .ALUT(n22432), .C0(index_i[4]), .Z(n22433));
    LUT4 mux_229_Mux_1_i317_3_lut (.A(n301), .B(n908_adj_2704), .C(index_i[4]), 
         .Z(n317_adj_2705)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_1_i317_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_2_i270_3_lut (.A(n29916), .B(n27427), .C(index_q[3]), 
         .Z(n270_adj_2677)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_2_i270_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_2_i316_3_lut (.A(n29947), .B(n27278), .C(index_q[3]), 
         .Z(n316_adj_2675)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_2_i316_3_lut.init = 16'hcaca;
    LUT4 i22429_3_lut (.A(n22044), .B(n22045), .C(index_q[4]), .Z(n22046)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22429_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_2_i397_3_lut (.A(n29958), .B(n29931), .C(index_q[3]), 
         .Z(n397_adj_2674)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_2_i397_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_5_i636_4_lut (.A(n157_adj_2374), .B(n27211), .C(index_q[4]), 
         .D(index_q[3]), .Z(n636_adj_2589)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_5_i636_4_lut.init = 16'h3aca;
    PFUMX mux_229_Mux_5_i732 (.BLUT(n11955), .ALUT(n731_adj_2647), .C0(index_i[4]), 
          .Z(n732_adj_2706)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 i9623_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n12109)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))+!A !(B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i9623_3_lut_4_lut_4_lut.init = 16'hb5b3;
    LUT4 i19989_3_lut (.A(n900_adj_2707), .B(n27342), .C(index_i[3]), 
         .Z(n22344)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19989_3_lut.init = 16'hcaca;
    LUT4 i22432_3_lut (.A(n18111), .B(n18112), .C(index_q[4]), .Z(n18113)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22432_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_5_i507_3_lut (.A(n491_adj_2519), .B(n506_adj_2686), 
         .C(index_q[4]), .Z(n507_adj_2585)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_5_i507_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_5_i573_3_lut_3_lut (.A(index_i[0]), .B(index_i[4]), 
         .C(n572_adj_2680), .Z(n573_adj_2708)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_5_i573_3_lut_3_lut.init = 16'hd1d1;
    LUT4 mux_230_Mux_5_i476_3_lut (.A(n460_adj_2709), .B(n475), .C(index_q[4]), 
         .Z(n476_adj_2584)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_5_i476_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_5_i413_3_lut (.A(n397_adj_2685), .B(n251_adj_2441), 
         .C(index_q[4]), .Z(n413_adj_2582)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_5_i413_3_lut.init = 16'hcaca;
    L6MUX21 i24851 (.D0(n26663), .D1(n26660), .SD(index_i[4]), .Z(n26664));
    LUT4 i21960_3_lut (.A(n27499), .B(n22339), .C(index_i[4]), .Z(n22340)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21960_3_lut.init = 16'hcaca;
    PFUMX i24849 (.BLUT(n26662), .ALUT(n26661), .C0(index_i[5]), .Z(n26663));
    LUT4 i15940_3_lut (.A(n18124), .B(n18125), .C(index_q[4]), .Z(n18126)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15940_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_5_i125_3_lut (.A(n109_adj_2408), .B(n124_adj_2393), 
         .C(index_q[4]), .Z(n125_adj_2581)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_5_i125_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_5_i94_3_lut (.A(n653_adj_2633), .B(n635_adj_2710), 
         .C(index_q[4]), .Z(n94_adj_2580)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_5_i94_3_lut.init = 16'hcaca;
    PFUMX i21123 (.BLUT(n142_adj_2711), .ALUT(n157_adj_2712), .C0(index_i[4]), 
          .Z(n23497));
    LUT4 mux_230_Mux_1_i986_3_lut (.A(n29934), .B(n27426), .C(index_q[3]), 
         .Z(n986_adj_2713)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_1_i986_3_lut.init = 16'hcaca;
    LUT4 i19974_3_lut (.A(n498), .B(n29952), .C(index_i[3]), .Z(n22329)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19974_3_lut.init = 16'hcaca;
    LUT4 i21985_3_lut (.A(n22329), .B(n22330), .C(index_i[4]), .Z(n22331)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21985_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_10_i637_3_lut_4_lut_4_lut (.A(n27183), .B(index_q[4]), 
         .C(index_q[5]), .D(n27125), .Z(n637_adj_2270)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_10_i637_3_lut_4_lut_4_lut.init = 16'h1f1c;
    LUT4 i20148_3_lut (.A(n526), .B(n541_adj_2392), .C(index_q[4]), .Z(n22503)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20148_3_lut.init = 16'hcaca;
    L6MUX21 i23352 (.D0(n24949), .D1(n24946), .SD(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2145[9]));
    LUT4 i9575_3_lut_4_lut_4_lut (.A(index_q[2]), .B(index_q[1]), .C(index_q[0]), 
         .D(n27328), .Z(n605_adj_2714)) /* synthesis lut_function=(A (B (C)+!B !(C+!(D)))+!A (B (C+!(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i9575_3_lut_4_lut_4_lut.init = 16'hc3c4;
    LUT4 i19966_3_lut (.A(n498), .B(n27358), .C(index_i[3]), .Z(n22321)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19966_3_lut.init = 16'hcaca;
    LUT4 i23708_then_3_lut (.A(index_q[0]), .B(index_q[4]), .C(index_q[3]), 
         .Z(n27523)) /* synthesis lut_function=(A (B)+!A (B (C)+!B !(C))) */ ;
    defparam i23708_then_3_lut.init = 16'hc9c9;
    LUT4 i22895_3_lut_4_lut (.A(n27182), .B(n20112), .C(index_q[8]), .D(n766), 
         .Z(n22138)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i22895_3_lut_4_lut.init = 16'hefe0;
    PFUMX i21124 (.BLUT(n173_adj_2547), .ALUT(n188), .C0(index_i[4]), 
          .Z(n23498));
    LUT4 i22629_3_lut (.A(n924_adj_2715), .B(n955), .C(index_q[5]), .Z(n23688)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22629_3_lut.init = 16'hcaca;
    LUT4 n803_bdd_3_lut_24122_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n25833)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A !(B (C+(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n803_bdd_3_lut_24122_4_lut_4_lut.init = 16'h9936;
    LUT4 i11925_3_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[3]), 
         .Z(n11265)) /* synthesis lut_function=(!((B (C))+!A)) */ ;
    defparam i11925_3_lut.init = 16'h2a2a;
    LUT4 i21991_3_lut (.A(n22317), .B(n22318), .C(index_i[4]), .Z(n22319)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21991_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_7_i956_3_lut_3_lut_4_lut (.A(n27185), .B(index_i[4]), 
         .C(n924_adj_2716), .D(index_i[5]), .Z(n956_adj_2717)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;
    defparam mux_229_Mux_7_i956_3_lut_3_lut_4_lut.init = 16'h11f0;
    LUT4 mux_230_Mux_6_i668_3_lut (.A(n108), .B(n29926), .C(index_q[3]), 
         .Z(n668_adj_2634)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_6_i668_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_6_i684_3_lut (.A(n14_adj_2290), .B(n29958), .C(index_q[3]), 
         .Z(n684_adj_2718)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_6_i684_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_10_i701_4_lut_4_lut (.A(n27185), .B(index_i[4]), .C(index_i[5]), 
         .D(n27124), .Z(n701_adj_2719)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B (C (D))+!B !(C)))) */ ;
    defparam mux_229_Mux_10_i701_4_lut_4_lut.init = 16'h3efe;
    LUT4 i19957_3_lut (.A(n27358), .B(n27438), .C(index_i[3]), .Z(n22312)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19957_3_lut.init = 16'hcaca;
    LUT4 i21993_3_lut (.A(n22311), .B(n22312), .C(index_i[4]), .Z(n22313)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21993_3_lut.init = 16'hcaca;
    LUT4 i23708_else_3_lut (.A(index_q[0]), .B(index_q[2]), .C(index_q[4]), 
         .D(index_q[3]), .Z(n27522)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C (D)+!C !(D))+!B !(C)))) */ ;
    defparam i23708_else_3_lut.init = 16'h1e58;
    PFUMX i21129 (.BLUT(n333), .ALUT(n348_adj_2720), .C0(index_i[4]), 
          .Z(n23503));
    LUT4 i22002_3_lut (.A(n22308), .B(n22309), .C(index_i[4]), .Z(n22310)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22002_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_6_i284_3_lut_4_lut_3_lut_rep_680 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27345)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_6_i284_3_lut_4_lut_3_lut_rep_680.init = 16'h6969;
    LUT4 i12105_2_lut_rep_797 (.A(index_i[1]), .B(index_i[2]), .C(index_i[0]), 
         .Z(n29924)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12105_2_lut_rep_797.init = 16'h7070;
    PFUMX i21130 (.BLUT(n364_adj_2721), .ALUT(n379_adj_2347), .C0(index_i[4]), 
          .Z(n23504));
    LUT4 index_i_7__bdd_4_lut_25344 (.A(index_i[7]), .B(n15194), .C(n25220), 
         .D(index_i[5]), .Z(n27060)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(B (C+(D))+!B !((D)+!C)))) */ ;
    defparam index_i_7__bdd_4_lut_25344.init = 16'h66f0;
    LUT4 i19779_3_lut_then_4_lut (.A(index_i[4]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n27526)) /* synthesis lut_function=(A (B (C)+!B !(C (D)+!C !(D)))+!A !(B (C)+!B !(C (D)+!C !(D)))) */ ;
    defparam i19779_3_lut_then_4_lut.init = 16'h96a5;
    LUT4 i19779_3_lut_else_4_lut (.A(index_i[4]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n27525)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C+!(D)))+!A !(B ((D)+!C)+!B (C (D)+!C !(D))))) */ ;
    defparam i19779_3_lut_else_4_lut.init = 16'h5685;
    L6MUX21 i21301 (.D0(n22010), .D1(n22013), .SD(index_q[5]), .Z(n23675));
    LUT4 i22855_3_lut_rep_403_4_lut (.A(n27178), .B(index_q[5]), .C(index_q[8]), 
         .D(n1021_adj_2722), .Z(n27068)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i22855_3_lut_rep_403_4_lut.init = 16'hf808;
    LUT4 n21795_bdd_3_lut (.A(n27069), .B(n701_adj_2719), .C(index_i[6]), 
         .Z(n26982)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n21795_bdd_3_lut.init = 16'hacac;
    PFUMX i25140 (.BLUT(n27449), .ALUT(n27450), .C0(index_i[1]), .Z(n27451));
    PFUMX i21131 (.BLUT(n397_adj_2641), .ALUT(n412), .C0(index_i[4]), 
          .Z(n23505));
    L6MUX21 i21305 (.D0(n22019), .D1(n18107), .SD(index_q[5]), .Z(n23679));
    L6MUX21 i21306 (.D0(n22022), .D1(n12055), .SD(index_q[5]), .Z(n23680));
    PFUMX i21308 (.BLUT(n542_adj_2640), .ALUT(n573_adj_2723), .C0(index_q[5]), 
          .Z(n23682));
    LUT4 mux_229_Mux_1_i732_3_lut (.A(n716_adj_2360), .B(n491_adj_2520), 
         .C(index_i[4]), .Z(n732_adj_2534)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_1_i732_3_lut.init = 16'hcaca;
    LUT4 i19780_3_lut_then_4_lut (.A(index_i[4]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n27529)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)+!C !(D)))+!A !(B (C+!(D))+!B (C (D)+!C !(D))))) */ ;
    defparam i19780_3_lut_then_4_lut.init = 16'h5a65;
    LUT4 i19780_3_lut_else_4_lut (.A(index_i[4]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n27528)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A !(B (C+!(D))+!B ((D)+!C)))) */ ;
    defparam i19780_3_lut_else_4_lut.init = 16'h59e5;
    PFUMX i21309 (.BLUT(n605_adj_2714), .ALUT(n636_adj_2724), .C0(index_q[5]), 
          .Z(n23683));
    PFUMX i21132 (.BLUT(n428_adj_2324), .ALUT(n443_adj_2312), .C0(index_i[4]), 
          .Z(n23506));
    LUT4 i19939_3_lut (.A(n356_adj_2398), .B(n27342), .C(index_i[3]), 
         .Z(n22294)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19939_3_lut.init = 16'hcaca;
    PFUMX i25253 (.BLUT(n27627), .ALUT(n27626), .C0(index_i[3]), .Z(n27628));
    LUT4 i22034_3_lut (.A(n22293), .B(n22294), .C(index_i[4]), .Z(n22295)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22034_3_lut.init = 16'hcaca;
    LUT4 i19936_3_lut (.A(n29911), .B(n27387), .C(index_i[3]), .Z(n22291)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19936_3_lut.init = 16'hcaca;
    LUT4 n26985_bdd_3_lut (.A(n28689), .B(n23583), .C(index_i[8]), .Z(n26986)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n26985_bdd_3_lut.init = 16'hcaca;
    PFUMX i19429 (.BLUT(n445_adj_2358), .ALUT(n508_adj_2513), .C0(index_q[6]), 
          .Z(n21784));
    LUT4 i22739_3_lut (.A(n22972), .B(n26707), .C(index_i[6]), .Z(n22981)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22739_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_9_i62_3_lut_4_lut_then_4_lut (.A(index_q[4]), .B(index_q[2]), 
         .C(index_q[1]), .D(index_q[0]), .Z(n27456)) /* synthesis lut_function=(!(A (B (C+(D)))+!A (B+(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_9_i62_3_lut_4_lut_then_4_lut.init = 16'h222b;
    LUT4 index_q_7__bdd_4_lut_25547 (.A(index_q[7]), .B(n15104), .C(n25198), 
         .D(index_q[5]), .Z(n27062)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(B (C+(D))+!B !((D)+!C)))) */ ;
    defparam index_q_7__bdd_4_lut_25547.init = 16'h66f0;
    PFUMX i21310 (.BLUT(n669_adj_2635), .ALUT(n700_adj_2725), .C0(index_q[5]), 
          .Z(n23684));
    PFUMX i21133 (.BLUT(n460), .ALUT(n475_adj_2378), .C0(index_i[4]), 
          .Z(n23507));
    PFUMX i21311 (.BLUT(n732_adj_2726), .ALUT(n22028), .C0(index_q[5]), 
          .Z(n23685));
    LUT4 mux_229_Mux_4_i158_3_lut (.A(n142), .B(n157_adj_2527), .C(index_i[4]), 
         .Z(n158_adj_2521)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_4_i158_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_3_i93_3_lut_4_lut (.A(n27429), .B(index_i[2]), .C(index_i[3]), 
         .D(n27430), .Z(n93_adj_2492)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam mux_229_Mux_3_i93_3_lut_4_lut.init = 16'hefe0;
    PFUMX i21312 (.BLUT(n797_adj_2630), .ALUT(n828_adj_2629), .C0(index_q[5]), 
          .Z(n23686));
    LUT4 mux_230_Mux_12_i254_4_lut (.A(n27084), .B(n20896), .C(index_q[6]), 
         .D(n27172), .Z(n254_adj_2727)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_12_i254_4_lut.init = 16'hca0a;
    LUT4 i22040_3_lut (.A(n22284), .B(n22285), .C(index_i[4]), .Z(n22286)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22040_3_lut.init = 16'hcaca;
    PFUMX i20892 (.BLUT(n956_adj_2717), .ALUT(n20714), .C0(index_i[6]), 
          .Z(n23266));
    LUT4 mux_229_Mux_12_i254_4_lut (.A(n27085), .B(n20888), .C(index_i[6]), 
         .D(n27229), .Z(n254_adj_2728)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_12_i254_4_lut.init = 16'hca0a;
    PFUMX i24847 (.BLUT(n26659), .ALUT(n26658), .C0(index_i[5]), .Z(n26660));
    PFUMX i21134 (.BLUT(n491), .ALUT(n11368), .C0(index_i[4]), .Z(n23508));
    LUT4 i22846_3_lut_rep_404_4_lut (.A(n27162), .B(index_i[5]), .C(index_i[8]), 
         .D(n1021), .Z(n27069)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i22846_3_lut_rep_404_4_lut.init = 16'hf808;
    LUT4 i19611_3_lut_4_lut_4_lut (.A(n27218), .B(index_q[4]), .C(index_q[3]), 
         .D(n27220), .Z(n21966)) /* synthesis lut_function=(A (B (C)+!B !(C+!(D)))+!A (B (C)+!B (C+(D)))) */ ;
    defparam i19611_3_lut_4_lut_4_lut.init = 16'hd3d0;
    LUT4 mux_229_Mux_0_i1002_3_lut_3_lut_4_lut (.A(n27429), .B(index_i[2]), 
         .C(n1001), .D(index_i[3]), .Z(n1002)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;
    defparam mux_229_Mux_0_i1002_3_lut_3_lut_4_lut.init = 16'hf011;
    PFUMX i21313 (.BLUT(n860_adj_2479), .ALUT(n891_adj_2626), .C0(index_q[5]), 
          .Z(n23687));
    LUT4 mux_230_Mux_7_i397_3_lut (.A(n29934), .B(n27297), .C(index_q[3]), 
         .Z(n397_adj_2594)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_7_i397_3_lut.init = 16'hcaca;
    LUT4 i22512_3_lut (.A(n29167), .B(n27451), .C(index_i[5]), .Z(n22910)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22512_3_lut.init = 16'hcaca;
    LUT4 i22519_3_lut (.A(n542_adj_2511), .B(n573_adj_2409), .C(index_i[5]), 
         .Z(n22904)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22519_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_0_i173_3_lut_4_lut (.A(n27424), .B(index_q[1]), .C(index_q[3]), 
         .D(n29953), .Z(n173_adj_2729)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_0_i173_3_lut_4_lut.init = 16'hdfd0;
    LUT4 i19921_3_lut (.A(n27393), .B(n27348), .C(index_i[3]), .Z(n22276)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19921_3_lut.init = 16'hcaca;
    LUT4 i19920_3_lut (.A(n29923), .B(n29913), .C(index_i[3]), .Z(n22275)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19920_3_lut.init = 16'hcaca;
    LUT4 i22049_3_lut (.A(n22275), .B(n22276), .C(index_i[4]), .Z(n22277)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22049_3_lut.init = 16'hcaca;
    LUT4 i19918_3_lut (.A(n29956), .B(n27436), .C(index_i[3]), .Z(n22273)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19918_3_lut.init = 16'hcaca;
    LUT4 i19917_3_lut (.A(n27440), .B(n652), .C(index_i[3]), .Z(n22272)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19917_3_lut.init = 16'hcaca;
    LUT4 i22051_3_lut (.A(n22272), .B(n22273), .C(index_i[4]), .Z(n22274)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22051_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_1_i620_3_lut_4_lut (.A(n27424), .B(index_q[1]), .C(index_q[3]), 
         .D(n29918), .Z(n620)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_1_i620_3_lut_4_lut.init = 16'hdfd0;
    LUT4 i19678_3_lut_4_lut (.A(n27424), .B(index_q[1]), .C(index_q[3]), 
         .D(n404), .Z(n22033)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i19678_3_lut_4_lut.init = 16'hdfd0;
    LUT4 mux_230_Mux_7_i956_3_lut_3_lut_4_lut (.A(n27195), .B(index_q[4]), 
         .C(n924_adj_2730), .D(index_q[5]), .Z(n956)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_7_i956_3_lut_3_lut_4_lut.init = 16'h11f0;
    LUT4 mux_229_Mux_7_i333_3_lut (.A(n27440), .B(n27385), .C(index_i[3]), 
         .Z(n333_adj_2572)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_7_i333_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_7_i348_3_lut (.A(n27435), .B(n27432), .C(index_i[3]), 
         .Z(n348_adj_2566)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_7_i348_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_8_i157_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n15_adj_2700)) /* synthesis lut_function=(A (B (C)+!B !(C (D)+!C !(D)))+!A !(B ((D)+!C)+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_8_i157_3_lut_4_lut_4_lut.init = 16'h83e0;
    PFUMX i20090 (.BLUT(n22443), .ALUT(n22444), .C0(index_i[4]), .Z(n22445));
    LUT4 mux_229_Mux_7_i397_3_lut (.A(n27435), .B(n27440), .C(index_i[3]), 
         .Z(n397_adj_2565)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_7_i397_3_lut.init = 16'hcaca;
    LUT4 i22545_3_lut (.A(n924_adj_2731), .B(n955_adj_2732), .C(index_i[5]), 
         .Z(n22833)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22545_3_lut.init = 16'hcaca;
    LUT4 i19846_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n22201)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(D))+!A (B (D)+!B ((D)+!C))) */ ;
    defparam i19846_3_lut_4_lut_4_lut.init = 16'hd52b;
    LUT4 mux_230_Mux_4_i205_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n205_adj_2733)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_4_i205_3_lut_4_lut_4_lut.init = 16'h5a2a;
    LUT4 mux_230_Mux_0_i684_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n684_adj_2399)) /* synthesis lut_function=(!(A ((D)+!B)+!A !(B (D)+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_0_i684_3_lut_4_lut_4_lut.init = 16'h5498;
    LUT4 i22834_3_lut (.A(n25840), .B(n26455), .C(index_i[6]), .Z(n22836)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22834_3_lut.init = 16'hcaca;
    LUT4 i20412_3_lut_3_lut_4_lut (.A(n27195), .B(index_q[4]), .C(n252), 
         .D(index_q[5]), .Z(n22786)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i20412_3_lut_3_lut_4_lut.init = 16'hf011;
    PFUMX i23350 (.BLUT(n24948), .ALUT(n24947), .C0(index_i[8]), .Z(n24949));
    LUT4 mux_229_Mux_6_i732_3_lut_4_lut (.A(n27440), .B(index_i[3]), .C(index_i[4]), 
         .D(n781_adj_2568), .Z(n732_adj_2734)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_6_i732_3_lut_4_lut.init = 16'hf909;
    LUT4 mux_230_Mux_10_i701_4_lut_4_lut (.A(n27195), .B(index_q[4]), .C(index_q[5]), 
         .D(n27126), .Z(n701)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B (C (D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_10_i701_4_lut_4_lut.init = 16'h3efe;
    LUT4 mux_229_Mux_6_i700_3_lut_4_lut (.A(n27440), .B(index_i[3]), .C(index_i[4]), 
         .D(n684_adj_2735), .Z(n700_adj_2736)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_6_i700_3_lut_4_lut.init = 16'h9f90;
    LUT4 i1_4_lut (.A(index_q[6]), .B(n27166), .C(index_q[5]), .D(index_q[4]), 
         .Z(n20711)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i1_4_lut.init = 16'hfffe;
    LUT4 i17974_4_lut (.A(n27323), .B(n892_adj_2476), .C(index_q[6]), 
         .D(index_q[5]), .Z(n20187)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D))))) */ ;
    defparam i17974_4_lut.init = 16'h3a35;
    LUT4 i22836_3_lut (.A(n20187), .B(n20711), .C(index_q[7]), .Z(n23785)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22836_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_6_i653_3_lut (.A(n27436), .B(n652), .C(index_i[3]), 
         .Z(n653_adj_2544)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_6_i653_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_6_i668_3_lut (.A(n660), .B(n27442), .C(index_i[3]), 
         .Z(n668_adj_2558)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_6_i668_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_6_i684_3_lut (.A(n27385), .B(n29956), .C(index_i[3]), 
         .Z(n684_adj_2735)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_6_i684_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_0_i1017_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .D(index_i[3]), .Z(n1017)) /* synthesis lut_function=(A (B (D)+!B !((D)+!C))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_0_i1017_4_lut_4_lut_4_lut.init = 16'hdd70;
    LUT4 mux_230_Mux_6_i732_3_lut_4_lut (.A(n27297), .B(index_q[3]), .C(index_q[4]), 
         .D(n731_adj_2603), .Z(n732_adj_2726)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_6_i732_3_lut_4_lut.init = 16'hf909;
    LUT4 mux_230_Mux_9_i62_3_lut_4_lut_else_4_lut (.A(index_q[4]), .B(index_q[2]), 
         .C(index_q[1]), .D(index_q[0]), .Z(n27455)) /* synthesis lut_function=((B+(C (D)))+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_9_i62_3_lut_4_lut_else_4_lut.init = 16'hfddd;
    LUT4 mux_230_Mux_6_i700_3_lut_4_lut (.A(n27297), .B(index_q[3]), .C(index_q[4]), 
         .D(n684_adj_2718), .Z(n700_adj_2725)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_6_i700_3_lut_4_lut.init = 16'h9f90;
    LUT4 mux_229_Mux_0_i220_3_lut (.A(n27383), .B(n27389), .C(index_i[3]), 
         .Z(n220_adj_2575)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_0_i220_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_1_i986_3_lut (.A(n27435), .B(n27389), .C(index_i[3]), 
         .Z(n986_adj_2737)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_1_i986_3_lut.init = 16'hcaca;
    PFUMX i20925 (.BLUT(n23295), .ALUT(n23296), .C0(index_q[5]), .Z(n23299));
    PFUMX i21151 (.BLUT(n557_adj_2310), .ALUT(n572_adj_2620), .C0(index_i[4]), 
          .Z(n23525));
    LUT4 i19711_3_lut_3_lut (.A(n27297), .B(index_q[3]), .C(n38), .Z(n22066)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam i19711_3_lut_3_lut.init = 16'h7474;
    LUT4 i22851_3_lut (.A(n23676), .B(n26221), .C(index_q[6]), .Z(n23691)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22851_3_lut.init = 16'hcaca;
    PFUMX i21152 (.BLUT(n589_adj_2617), .ALUT(n604_adj_2356), .C0(index_i[4]), 
          .Z(n23526));
    LUT4 i22636_3_lut (.A(n26486), .B(n22219), .C(index_i[5]), .Z(n22220)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22636_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_3_i349_3_lut_3_lut (.A(index_q[1]), .B(index_q[4]), 
         .C(n348_adj_2702), .Z(n349_adj_2631)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_3_i349_3_lut_3_lut.init = 16'hd1d1;
    PFUMX i21153 (.BLUT(n620_adj_2614), .ALUT(n635_adj_2738), .C0(index_i[4]), 
          .Z(n23527));
    PFUMX i20926 (.BLUT(n23297), .ALUT(n23298), .C0(index_q[5]), .Z(n23300));
    LUT4 i23080_2_lut (.A(index_i[3]), .B(index_i[2]), .Z(n22740)) /* synthesis lut_function=(A+!(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i23080_2_lut.init = 16'hbbbb;
    LUT4 i19848_3_lut (.A(n27278), .B(n29938), .C(index_q[3]), .Z(n22203)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19848_3_lut.init = 16'hcaca;
    LUT4 i19737_3_lut_3_lut_4_lut (.A(n27293), .B(index_q[2]), .C(n14_adj_2290), 
         .D(index_q[3]), .Z(n22092)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (B (C (D))+!B (C+!(D)))) */ ;
    defparam i19737_3_lut_3_lut_4_lut.init = 16'hf099;
    LUT4 i17997_4_lut (.A(n27321), .B(n892_adj_2439), .C(index_i[6]), 
         .D(index_i[5]), .Z(n20213)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D))))) */ ;
    defparam i17997_4_lut.init = 16'h3a35;
    LUT4 i22859_3_lut (.A(n20213), .B(n20603), .C(index_i[7]), .Z(n23255)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22859_3_lut.init = 16'hcaca;
    LUT4 n476_bdd_3_lut_23668_3_lut_4_lut (.A(n27293), .B(index_q[2]), .C(n491_adj_2739), 
         .D(index_q[4]), .Z(n25353)) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))+!A !(B ((D)+!C)+!B !(C+(D)))) */ ;
    defparam n476_bdd_3_lut_23668_3_lut_4_lut.init = 16'h99f0;
    LUT4 i19671_3_lut_3_lut_4_lut (.A(n27293), .B(index_q[2]), .C(n29931), 
         .D(index_q[3]), .Z(n22026)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (B (C (D))+!B (C+!(D)))) */ ;
    defparam i19671_3_lut_3_lut_4_lut.init = 16'hf099;
    PFUMX i21154 (.BLUT(n653_adj_2613), .ALUT(n668_adj_2583), .C0(index_i[4]), 
          .Z(n23528));
    LUT4 i22316_3_lut (.A(n22200), .B(n22201), .C(index_q[4]), .Z(n22202)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22316_3_lut.init = 16'hcaca;
    LUT4 i22408_3_lut (.A(n22056), .B(n22057), .C(index_q[4]), .Z(n22058)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22408_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_0_i716_3_lut (.A(n29946), .B(n27311), .C(index_q[3]), 
         .Z(n716_adj_2406)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_0_i716_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_6_i636_4_lut_4_lut (.A(index_q[1]), .B(index_q[4]), 
         .C(n635_adj_2710), .D(n14725), .Z(n636_adj_2724)) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_6_i636_4_lut_4_lut.init = 16'hf3d1;
    PFUMX i20932 (.BLUT(n23302), .ALUT(n23303), .C0(index_q[5]), .Z(n23306));
    LUT4 mux_230_Mux_1_i732_3_lut (.A(n716_adj_2357), .B(n491_adj_2519), 
         .C(index_q[4]), .Z(n732_adj_2402)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_1_i732_3_lut.init = 16'hcaca;
    PFUMX i21155 (.BLUT(n684_adj_2463), .ALUT(n699_adj_2336), .C0(index_i[4]), 
          .Z(n23529));
    PFUMX i20933 (.BLUT(n23304), .ALUT(n23305), .C0(index_q[5]), .Z(n23307));
    LUT4 mux_230_Mux_5_i731_3_lut (.A(n29938), .B(n27280), .C(index_q[3]), 
         .Z(n731)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_5_i731_3_lut.init = 16'hcaca;
    PFUMX i21156 (.BLUT(n716_adj_2612), .ALUT(n731_adj_2440), .C0(index_i[4]), 
          .Z(n23530));
    LUT4 i22795_3_lut (.A(n23173), .B(n26132), .C(index_q[6]), .Z(n23182)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22795_3_lut.init = 16'hcaca;
    PFUMX i21157 (.BLUT(n747_adj_2330), .ALUT(n762_adj_2740), .C0(index_i[4]), 
          .Z(n23531));
    LUT4 mux_229_Mux_4_i828_3_lut_4_lut (.A(index_i[4]), .B(index_i[3]), 
         .C(n812), .D(n29951), .Z(n828_adj_2741)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_4_i828_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i19782_3_lut (.A(n25203), .B(n21785), .C(index_q[8]), .Z(n22137)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19782_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_5_i797_3_lut_4_lut (.A(index_i[4]), .B(index_i[3]), 
         .C(n27476), .D(n27256), .Z(n797_adj_2742)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_5_i797_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i20946 (.BLUT(n23316), .ALUT(n23317), .C0(index_i[5]), .Z(n23320));
    LUT4 mux_230_Mux_0_i653_3_lut (.A(n14_adj_2290), .B(n29955), .C(index_q[3]), 
         .Z(n653_adj_2396)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_0_i653_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_1_i763_3_lut_4_lut (.A(index_i[4]), .B(index_i[3]), 
         .C(n27542), .D(n27256), .Z(n763_adj_2535)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_1_i763_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12406_2_lut_rep_598 (.A(index_i[2]), .B(index_i[0]), .Z(n27263)) /* synthesis lut_function=(A (B)) */ ;
    defparam i12406_2_lut_rep_598.init = 16'h8888;
    PFUMX i21158 (.BLUT(n781_adj_2322), .ALUT(n796_adj_2473), .C0(index_i[4]), 
          .Z(n23532));
    PFUMX i20947 (.BLUT(n23318), .ALUT(n23319), .C0(index_i[5]), .Z(n23321));
    LUT4 mux_230_Mux_3_i860_3_lut_4_lut (.A(n27293), .B(index_q[2]), .C(index_q[4]), 
         .D(n859_adj_2381), .Z(n860_adj_2648)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam mux_230_Mux_3_i860_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_230_Mux_7_i443_3_lut_4_lut (.A(n27293), .B(index_q[2]), .C(index_q[3]), 
         .D(n29931), .Z(n443_adj_2602)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;
    defparam mux_230_Mux_7_i443_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_229_Mux_0_i124_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n124_adj_2645)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A !(B (D)+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_0_i124_3_lut_4_lut_4_lut.init = 16'h6c99;
    LUT4 i19938_3_lut_4_lut_4_lut (.A(index_i[0]), .B(n27394), .C(index_i[3]), 
         .D(n27322), .Z(n22293)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19938_3_lut_4_lut_4_lut.init = 16'hc5c0;
    PFUMX i21159 (.BLUT(n812_adj_2743), .ALUT(n11924), .C0(index_i[4]), 
          .Z(n23533));
    LUT4 mux_229_Mux_3_i796_3_lut_3_lut (.A(index_i[4]), .B(n781_adj_2568), 
         .C(index_i[2]), .Z(n796_adj_2744)) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam mux_229_Mux_3_i796_3_lut_3_lut.init = 16'he4e4;
    LUT4 i9638_4_lut_4_lut (.A(index_i[4]), .B(n22724), .C(n27506), .D(n27430), 
         .Z(n12124)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam i9638_4_lut_4_lut.init = 16'hf4b0;
    LUT4 i20598_4_lut_4_lut (.A(index_i[4]), .B(index_i[5]), .C(n27509), 
         .D(n908_adj_2704), .Z(n22972)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam i20598_4_lut_4_lut.init = 16'hd1c0;
    LUT4 mux_229_Mux_3_i94_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[4]), .D(n93_adj_2492), .Z(n94_adj_2745)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_3_i94_3_lut_4_lut.init = 16'hf606;
    PFUMX i21161 (.BLUT(n875_adj_2746), .ALUT(n890_adj_2355), .C0(index_i[4]), 
          .Z(n23535));
    LUT4 i20639_3_lut (.A(n23005), .B(n23006), .C(index_i[7]), .Z(n23013)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20639_3_lut.init = 16'hcaca;
    LUT4 i20632_3_lut (.A(n22991), .B(n26780), .C(index_i[6]), .Z(n23006)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20632_3_lut.init = 16'hcaca;
    LUT4 i20641_3_lut (.A(n23009), .B(n23010), .C(index_i[7]), .Z(n23015)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20641_3_lut.init = 16'hcaca;
    LUT4 i20635_3_lut (.A(n22997), .B(n22998), .C(index_i[6]), .Z(n23009)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20635_3_lut.init = 16'hcaca;
    PFUMX i21162 (.BLUT(n908_adj_2500), .ALUT(n923_adj_2607), .C0(index_i[4]), 
          .Z(n23536));
    LUT4 mux_229_Mux_3_i62_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[4]), .D(n812_adj_2554), .Z(n62_adj_2747)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_3_i62_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_229_Mux_3_i700_3_lut_4_lut (.A(index_i[4]), .B(index_i[3]), 
         .C(n684_adj_2482), .D(n29951), .Z(n700_adj_2748)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_3_i700_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i1_4_lut_adj_84 (.A(index_i[7]), .B(n27070), .C(index_i[6]), 
         .D(index_i[8]), .Z(n20675)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_4_lut_adj_84.init = 16'hfffe;
    LUT4 i23135_2_lut_rep_599 (.A(index_i[4]), .B(index_i[3]), .Z(n27264)) /* synthesis lut_function=((B)+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i23135_2_lut_rep_599.init = 16'hdddd;
    LUT4 mux_229_Mux_3_i797_3_lut_4_lut (.A(index_i[4]), .B(index_i[3]), 
         .C(n796_adj_2744), .D(n27430), .Z(n797_adj_2495)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_3_i797_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i25176 (.BLUT(n27507), .ALUT(n27508), .C0(index_i[0]), .Z(n27509));
    LUT4 i11768_3_lut_3_lut_rep_760 (.A(index_q[1]), .B(index_q[0]), .C(index_q[2]), 
         .Z(n27425)) /* synthesis lut_function=(!(A+!((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i11768_3_lut_3_lut_rep_760.init = 16'h5151;
    PFUMX i19697 (.BLUT(n22050), .ALUT(n22051), .C0(index_q[5]), .Z(n22052));
    PFUMX i23710 (.BLUT(n25416), .ALUT(n25412), .C0(index_q[6]), .Z(n25417));
    LUT4 n21809_bdd_3_lut_23390 (.A(n23301), .B(n23308), .C(index_q[7]), 
         .Z(n24992)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n21809_bdd_3_lut_23390.init = 16'hcaca;
    LUT4 mux_230_Mux_6_i452_3_lut_4_lut_3_lut_rep_761 (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[0]), .Z(n27426)) /* synthesis lut_function=(A (B (C))+!A !(B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_6_i452_3_lut_4_lut_3_lut_rep_761.init = 16'h9595;
    L6MUX21 i24731 (.D0(n26534), .D1(n26532), .SD(index_q[5]), .Z(n26535));
    PFUMX i19438 (.BLUT(n445), .ALUT(n508), .C0(index_i[6]), .Z(n21793));
    PFUMX i23347 (.BLUT(n24945), .ALUT(n23255), .C0(index_i[8]), .Z(n24946));
    PFUMX i24729 (.BLUT(n26533), .ALUT(n14_adj_2290), .C0(index_q[3]), 
          .Z(n26534));
    LUT4 mux_230_Mux_7_i45_3_lut_4_lut_3_lut_rep_762 (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[0]), .Z(n27427)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_7_i45_3_lut_4_lut_3_lut_rep_762.init = 16'h6565;
    PFUMX mux_230_Mux_1_i891 (.BLUT(n882), .ALUT(n890_adj_2749), .C0(n27268), 
          .Z(n891_adj_2405)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 n22912_bdd_3_lut_23405 (.A(n22914), .B(n22915), .C(index_i[7]), 
         .Z(n25008)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n22912_bdd_3_lut_23405.init = 16'hcaca;
    PFUMX i24727 (.BLUT(n26531), .ALUT(n22003), .C0(index_q[4]), .Z(n26532));
    LUT4 mux_230_Mux_7_i620_3_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[0]), .D(index_q[3]), .Z(n620_adj_2750)) /* synthesis lut_function=(A (B (C+!(D)))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_7_i620_3_lut_4_lut_4_lut.init = 16'h9199;
    LUT4 i12501_2_lut_rep_602 (.A(index_q[2]), .B(index_q[0]), .Z(n27267)) /* synthesis lut_function=(A (B)) */ ;
    defparam i12501_2_lut_rep_602.init = 16'h8888;
    PFUMX i19757 (.BLUT(n22110), .ALUT(n22111), .C0(index_q[5]), .Z(n22112));
    PFUMX i19763 (.BLUT(n22116), .ALUT(n22117), .C0(index_q[5]), .Z(n22118));
    LUT4 mux_230_Mux_8_i93_3_lut_3_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[0]), .D(index_q[3]), .Z(n93_adj_2590)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(D))+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_8_i93_3_lut_3_lut_4_lut.init = 16'h3391;
    PFUMX i19766 (.BLUT(n22119), .ALUT(n22120), .C0(index_q[5]), .Z(n22121));
    LUT4 mux_230_Mux_2_i890_3_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[0]), .D(index_q[3]), .Z(n890)) /* synthesis lut_function=(A (B (C (D))+!B (C (D)+!C !(D)))+!A !(B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_2_i890_3_lut_4_lut_4_lut.init = 16'ha546;
    LUT4 i22696_3_lut (.A(n28767), .B(n27570), .C(index_q[5]), .Z(n23111)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22696_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_0_i620_3_lut (.A(n29934), .B(n29918), .C(index_q[3]), 
         .Z(n620_adj_2390)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_0_i620_3_lut.init = 16'hcaca;
    LUT4 i20799_4_lut_4_lut (.A(index_q[4]), .B(index_q[5]), .C(n27473), 
         .D(n908_adj_2751), .Z(n23173)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam i20799_4_lut_4_lut.init = 16'hd1c0;
    LUT4 i9557_4_lut_4_lut (.A(index_q[4]), .B(n22730), .C(n29967), .D(n29936), 
         .Z(n12043)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam i9557_4_lut_4_lut.init = 16'hf4b0;
    PFUMX i19769 (.BLUT(n22122), .ALUT(n22123), .C0(index_q[5]), .Z(n22124));
    LUT4 i23101_2_lut_rep_603 (.A(index_q[4]), .B(index_q[3]), .Z(n27268)) /* synthesis lut_function=((B)+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i23101_2_lut_rep_603.init = 16'hdddd;
    LUT4 mux_229_Mux_6_i363_3_lut_4_lut_3_lut_rep_681 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27346)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_6_i363_3_lut_4_lut_3_lut_rep_681.init = 16'h9292;
    PFUMX i19775 (.BLUT(n22128), .ALUT(n22129), .C0(index_i[5]), .Z(n22130));
    LUT4 mux_230_Mux_3_i797_3_lut_4_lut (.A(index_q[4]), .B(index_q[3]), 
         .C(n796_adj_2619), .D(n29936), .Z(n797)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_3_i797_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i19778 (.BLUT(n22131), .ALUT(n22132), .C0(index_i[5]), .Z(n22133));
    LUT4 i11777_2_lut_rep_604 (.A(index_q[0]), .B(index_q[1]), .Z(n27269)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i11777_2_lut_rep_604.init = 16'h4444;
    LUT4 i20780_3_lut (.A(n23148), .B(n23149), .C(index_q[7]), .Z(n23154)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20780_3_lut.init = 16'hcaca;
    LUT4 i22701_3_lut (.A(n542_adj_2697), .B(n573_adj_2537), .C(index_q[5]), 
         .Z(n23105)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22701_3_lut.init = 16'hcaca;
    LUT4 i20775_3_lut (.A(n23138), .B(n23139), .C(index_q[6]), .Z(n23149)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20775_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_0_i589_3_lut (.A(n29935), .B(n14), .C(index_q[3]), 
         .Z(n589)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_0_i589_3_lut.init = 16'hcaca;
    LUT4 i21022_3_lut (.A(n308), .B(n27238), .C(index_q[3]), .Z(n23396)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21022_3_lut.init = 16'hcaca;
    LUT4 i21021_3_lut (.A(n619), .B(n29934), .C(index_q[3]), .Z(n23395)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21021_3_lut.init = 16'hcaca;
    LUT4 i22417_3_lut (.A(n22053), .B(n22054), .C(index_q[4]), .Z(n22055)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22417_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_2_i604_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[0]), .D(index_q[3]), .Z(n604_adj_2673)) /* synthesis lut_function=(!(A (B (D)+!B !(C+!(D)))+!A !(B (D)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_2_i604_3_lut_4_lut_4_lut_4_lut.init = 16'h65bb;
    LUT4 i22708_3_lut (.A(n286_adj_2564), .B(n317_adj_2752), .C(index_i[5]), 
         .Z(n23577)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22708_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_5_i781_3_lut_4_lut_4_lut_then_4_lut (.A(index_q[3]), 
         .B(index_q[0]), .C(index_q[4]), .D(index_q[2]), .Z(n27459)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_5_i781_3_lut_4_lut_4_lut_then_4_lut.init = 16'hece0;
    LUT4 n811_bdd_4_lut_then_4_lut (.A(index_i[3]), .B(index_i[4]), .C(index_i[1]), 
         .D(index_i[2]), .Z(n27541)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B+(C (D)+!C !(D)))) */ ;
    defparam n811_bdd_4_lut_then_4_lut.init = 16'hf44f;
    LUT4 i19876_3_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[2]), .C(index_q[0]), 
         .D(index_q[3]), .Z(n22231)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A (B (C)+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i19876_3_lut_4_lut_4_lut.init = 16'h3c9d;
    LUT4 mux_230_Mux_5_i781_3_lut_4_lut_4_lut_else_4_lut (.A(index_q[3]), 
         .B(index_q[0]), .C(index_q[4]), .Z(n27458)) /* synthesis lut_function=(!(A (C)+!A (B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_5_i781_3_lut_4_lut_4_lut_else_4_lut.init = 16'h1f1f;
    LUT4 n811_bdd_4_lut_else_4_lut (.A(index_i[3]), .B(index_i[4]), .C(index_i[1]), 
         .D(index_i[2]), .Z(n27540)) /* synthesis lut_function=(!(A (B (D)+!B ((D)+!C))+!A !(B+!((D)+!C)))) */ ;
    defparam n811_bdd_4_lut_else_4_lut.init = 16'h44fc;
    LUT4 mux_230_Mux_0_i954_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n954_adj_2428)) /* synthesis lut_function=(A (D)+!A !(B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_0_i954_3_lut_4_lut_4_lut.init = 16'haf40;
    LUT4 mux_229_Mux_2_i349_3_lut_3_lut (.A(index_i[0]), .B(index_i[4]), 
         .C(n348_adj_2753), .Z(n349_adj_2754)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_2_i349_3_lut_3_lut.init = 16'hd1d1;
    LUT4 i21020_3_lut (.A(n27425), .B(n27297), .C(index_q[3]), .Z(n23394)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21020_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_6_i347_3_lut_4_lut_3_lut_rep_606 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n27271)) /* synthesis lut_function=(!(A (B+!(C))+!A ((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_6_i347_3_lut_4_lut_3_lut_rep_606.init = 16'h2424;
    LUT4 mux_229_Mux_2_i859_3_lut_4_lut_4_lut (.A(index_i[0]), .B(n29952), 
         .C(index_i[3]), .D(n27322), .Z(n859_adj_2698)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B ((D)+!C)+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_2_i859_3_lut_4_lut_4_lut.init = 16'h5c0c;
    LUT4 mux_230_Mux_0_i491_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n491_adj_2676)) /* synthesis lut_function=(!(A (B (D)+!B !(C+!(D)))+!A ((C+!(D))+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_0_i491_3_lut_4_lut.init = 16'h24aa;
    PFUMX i19790 (.BLUT(n22143), .ALUT(n22144), .C0(index_i[5]), .Z(n22145));
    LUT4 i21019_3_lut (.A(n27238), .B(n29935), .C(index_q[3]), .Z(n23393)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21019_3_lut.init = 16'hcaca;
    LUT4 i12247_2_lut (.A(index_i[1]), .B(index_i[3]), .Z(n541_adj_2377)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i12247_2_lut.init = 16'h1111;
    LUT4 n572_bdd_3_lut_24963_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n26170)) /* synthesis lut_function=(A (B (C+(D)))+!A (B ((D)+!C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam n572_bdd_3_lut_24963_4_lut.init = 16'hcc94;
    L6MUX21 i21004 (.D0(n23376), .D1(n23377), .SD(index_q[5]), .Z(n23378));
    LUT4 mux_229_Mux_2_i507_3_lut_3_lut (.A(index_i[0]), .B(index_i[4]), 
         .C(n491_adj_2679), .Z(n507_adj_2755)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_2_i507_3_lut_3_lut.init = 16'h7474;
    PFUMX i19793 (.BLUT(n22146), .ALUT(n22147), .C0(index_i[5]), .Z(n22148));
    LUT4 i19680_3_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[2]), .C(index_q[0]), 
         .D(index_q[3]), .Z(n22035)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C+(D)))+!A !(B (C (D)+!C !(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i19680_3_lut_4_lut_4_lut.init = 16'h955a;
    LUT4 mux_230_Mux_2_i653_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n653_adj_2671)) /* synthesis lut_function=(A (B (C+!(D))+!B !(D))+!A !(B (C+!(D))+!B !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_2_i653_3_lut_4_lut.init = 16'h94aa;
    LUT4 mux_229_Mux_0_i526_3_lut (.A(n27346), .B(n29922), .C(index_i[3]), 
         .Z(n526_adj_2376)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_0_i526_3_lut.init = 16'hcaca;
    PFUMX i19796 (.BLUT(n22149), .ALUT(n22150), .C0(index_i[5]), .Z(n22151));
    LUT4 i9676_3_lut_4_lut_3_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[4]), 
         .Z(n12165)) /* synthesis lut_function=(!(A (B)+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i9676_3_lut_4_lut_3_lut.init = 16'h6262;
    PFUMX i19799 (.BLUT(n22152), .ALUT(n22153), .C0(index_i[5]), .Z(n22154));
    LUT4 i19881_3_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[2]), .C(index_q[0]), 
         .D(index_q[3]), .Z(n22236)) /* synthesis lut_function=(A (B (C)+!B !(C+!(D)))+!A (B (C (D)+!C !(D))+!B !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i19881_3_lut_4_lut_4_lut.init = 16'hc395;
    LUT4 mux_229_Mux_4_i221_3_lut_3_lut (.A(index_i[0]), .B(index_i[4]), 
         .C(n205_adj_2756), .Z(n221_adj_2757)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_4_i221_3_lut_3_lut.init = 16'h7474;
    LUT4 mux_230_Mux_4_i14_3_lut_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n14)) /* synthesis lut_function=(!(A (B+(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_4_i14_3_lut_3_lut.init = 16'h5656;
    LUT4 mux_230_Mux_2_i908_3_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[0]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n908_adj_2751)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C)+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_2_i908_3_lut_4_lut_4_lut.init = 16'h5a51;
    LUT4 mux_230_Mux_5_i828_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[4]), .D(n27307), .Z(n828_adj_2593)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_5_i828_4_lut_4_lut.init = 16'hc66c;
    LUT4 mux_230_Mux_7_i108_3_lut_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n108)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_7_i108_3_lut_3_lut.init = 16'hc6c6;
    PFUMX i24686 (.BLUT(n26485), .ALUT(n26484), .C0(index_i[4]), .Z(n26486));
    LUT4 mux_230_Mux_3_i507_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[4]), .D(n491_adj_2401), .Z(n507_adj_2639)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_3_i507_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_230_Mux_1_i882_3_lut_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n882)) /* synthesis lut_function=(A ((C)+!B)+!A !((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_1_i882_3_lut_3_lut.init = 16'ha6a6;
    LUT4 mux_229_Mux_6_i396_3_lut_4_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[1]), .Z(n356_adj_2398)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_6_i396_3_lut_4_lut_4_lut_3_lut.init = 16'h7979;
    LUT4 mux_229_Mux_6_i134_3_lut_4_lut_3_lut_rep_682 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27347)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_6_i134_3_lut_4_lut_3_lut_rep_682.init = 16'h9696;
    LUT4 mux_230_Mux_6_i442_rep_609 (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .Z(n27274)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_6_i442_rep_609.init = 16'h6464;
    LUT4 mux_230_Mux_6_i483_3_lut_3_lut_rep_610 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n27275)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_6_i483_3_lut_3_lut_rep_610.init = 16'h6c6c;
    LUT4 mux_230_Mux_6_i134_3_lut_4_lut_3_lut_rep_611 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n27276)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_6_i134_3_lut_4_lut_3_lut_rep_611.init = 16'h9696;
    PFUMX i19805 (.BLUT(n22158), .ALUT(n22159), .C0(index_i[5]), .Z(n22160));
    LUT4 i19365_3_lut_4_lut_4_lut (.A(index_i[0]), .B(n29922), .C(index_i[3]), 
         .D(n27381), .Z(n21720)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19365_3_lut_4_lut_4_lut.init = 16'hcfc5;
    LUT4 mux_229_Mux_2_i763_4_lut_4_lut (.A(index_i[0]), .B(n11969), .C(index_i[4]), 
         .D(n157_adj_2299), .Z(n763_adj_2758)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_2_i763_4_lut_4_lut.init = 16'hdfd0;
    CCU2D add_417_15 (.A0(quarter_wave_sample_register_i[14]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(\quarter_wave_sample_register_q[15] ), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17900), .S0(o_val_pipeline_i_0__15__N_2176[14]), 
          .S1(o_val_pipeline_i_0__15__N_2176[15]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam add_417_15.INIT0 = 16'hf555;
    defparam add_417_15.INIT1 = 16'hf555;
    defparam add_417_15.INJECT1_0 = "NO";
    defparam add_417_15.INJECT1_1 = "NO";
    LUT4 mux_230_Mux_6_i490_3_lut_3_lut_rep_612 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n27277)) /* synthesis lut_function=(!(A (B)+!A (B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_6_i490_3_lut_3_lut_rep_612.init = 16'h3636;
    LUT4 i12146_2_lut_3_lut_3_lut (.A(index_i[0]), .B(index_i[3]), .C(index_i[2]), 
         .Z(n14744)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12146_2_lut_3_lut_3_lut.init = 16'h4040;
    LUT4 mux_229_Mux_0_i652_3_lut_4_lut_3_lut_rep_683 (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[1]), .Z(n27348)) /* synthesis lut_function=(!(A (B+(C))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_0_i652_3_lut_4_lut_3_lut_rep_683.init = 16'h4646;
    LUT4 mux_229_Mux_2_i773_3_lut_rep_685 (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[1]), .Z(n27350)) /* synthesis lut_function=(A ((C)+!B)+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_2_i773_3_lut_rep_685.init = 16'he6e6;
    LUT4 i11400_2_lut_rep_686 (.A(index_i[0]), .B(index_i[1]), .Z(n27351)) /* synthesis lut_function=((B)+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11400_2_lut_rep_686.init = 16'hdddd;
    LUT4 mux_230_Mux_5_i581_3_lut_3_lut_rep_613 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n27278)) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_5_i581_3_lut_3_lut_rep_613.init = 16'h6a6a;
    LUT4 i19875_3_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[0]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n22230)) /* synthesis lut_function=(!(A ((D)+!C)+!A !(B (C (D))+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i19875_3_lut_4_lut_4_lut.init = 16'h51a0;
    LUT4 i11471_2_lut_rep_764 (.A(index_i[0]), .B(index_i[1]), .Z(n27429)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11471_2_lut_rep_764.init = 16'h8888;
    LUT4 mux_230_Mux_5_i459_3_lut_4_lut_3_lut_rep_614 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n27279)) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_5_i459_3_lut_4_lut_3_lut_rep_614.init = 16'h6b6b;
    LUT4 mux_229_Mux_4_i77_3_lut_4_lut_3_lut_rep_687 (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[1]), .Z(n27352)) /* synthesis lut_function=(A (B (C))+!A !(B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_4_i77_3_lut_4_lut_3_lut_rep_687.init = 16'h9595;
    LUT4 mux_230_Mux_6_i262_3_lut_4_lut_3_lut_rep_615 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n27280)) /* synthesis lut_function=(A ((C)+!B)+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_6_i262_3_lut_4_lut_3_lut_rep_615.init = 16'hb6b6;
    LUT4 mux_229_Mux_6_i60_3_lut_4_lut_4_lut_3_lut_rep_688 (.A(index_i[0]), 
         .B(index_i[2]), .C(index_i[1]), .Z(n27353)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_6_i60_3_lut_4_lut_4_lut_3_lut_rep_688.init = 16'hd6d6;
    LUT4 mux_230_Mux_1_i301_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n301_adj_2759)) /* synthesis lut_function=(A (B (C+(D))+!B !(D))+!A !(B (C+(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_1_i301_3_lut_4_lut_4_lut.init = 16'h99b6;
    LUT4 i12516_2_lut (.A(index_q[1]), .B(index_q[3]), .Z(n541_adj_2371)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i12516_2_lut.init = 16'h1111;
    LUT4 mux_230_Mux_0_i526_3_lut (.A(n29953), .B(n27278), .C(index_q[3]), 
         .Z(n526_adj_2370)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_0_i526_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_5_i460_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n460_adj_2709)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A !(B (C)+!B !(C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_5_i460_3_lut_4_lut_4_lut.init = 16'h6b5a;
    LUT4 n15000_bdd_3_lut_24607_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n26385)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+!(D)))+!A (B (D)+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n15000_bdd_3_lut_24607_4_lut_4_lut_4_lut.init = 16'h30f7;
    LUT4 i9593_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n12079)) /* synthesis lut_function=(!(A (B (D)+!B (C+!(D)))+!A !(B (D)+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i9593_3_lut_4_lut_4_lut.init = 16'h4699;
    LUT4 mux_229_Mux_6_i459_rep_693 (.A(index_i[0]), .B(index_i[2]), .C(index_i[1]), 
         .Z(n27358)) /* synthesis lut_function=(!(A (B+!(C))+!A !((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_6_i459_rep_693.init = 16'h7171;
    PFUMX i19817 (.BLUT(n22170), .ALUT(n22171), .C0(index_i[5]), .Z(n22172));
    LUT4 mux_229_Mux_3_i653_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[1]), .D(index_i[3]), .Z(n653_adj_2454)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C))+!A !(B (C (D)+!C !(D))+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_3_i653_3_lut_4_lut_4_lut.init = 16'h71a5;
    PFUMX i19826 (.BLUT(n22179), .ALUT(n22180), .C0(index_i[5]), .Z(n22181));
    LUT4 mux_230_Mux_2_i491_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n491_adj_2760)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A !(B (C)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_2_i491_3_lut_4_lut_4_lut.init = 16'h6a5a;
    LUT4 n172_bdd_3_lut_4_lut_4_lut_4_lut_adj_85 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n26485)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)+!C !(D)))+!A (B (C+!(D))+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n172_bdd_3_lut_4_lut_4_lut_4_lut_adj_85.init = 16'h0f38;
    LUT4 i22722_3_lut (.A(n26360), .B(n22126), .C(index_q[5]), .Z(n22127)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22722_3_lut.init = 16'hcaca;
    LUT4 i19998_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[2]), .C(index_i[1]), 
         .D(index_i[3]), .Z(n22353)) /* synthesis lut_function=(!(A (B (D)+!B !(C+(D)))+!A !(B (D)+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19998_3_lut_4_lut_4_lut.init = 16'h66b9;
    LUT4 n123_bdd_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[2]), .C(index_i[1]), 
         .D(index_i[3]), .Z(n25814)) /* synthesis lut_function=(A (B+!((D)+!C))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n123_bdd_3_lut_4_lut_4_lut.init = 16'h99b9;
    LUT4 i20016_3_lut_4_lut (.A(index_i[0]), .B(index_i[2]), .C(index_i[1]), 
         .D(index_i[3]), .Z(n22371)) /* synthesis lut_function=(A (B (D)+!B (C+(D)))+!A !(B (D)+!B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20016_3_lut_4_lut.init = 16'haa65;
    LUT4 mux_229_Mux_3_i444_3_lut_4_lut (.A(index_i[0]), .B(index_i[3]), 
         .C(n27381), .D(index_i[4]), .Z(n444_adj_2761)) /* synthesis lut_function=(!(A (B (D)+!B (C (D)))+!A !(B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_3_i444_3_lut_4_lut.init = 16'h46aa;
    LUT4 mux_229_Mux_3_i1002_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n20166)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (D))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_3_i1002_3_lut_3_lut_4_lut.init = 16'hf708;
    LUT4 mux_229_Mux_6_i572_3_lut_4_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[1]), .D(index_i[3]), .Z(n572_adj_2615)) /* synthesis lut_function=(A (C)+!A (B (C+!(D))+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_6_i572_3_lut_4_lut.init = 16'hf0e5;
    LUT4 mux_230_Mux_6_i475_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n475_adj_2653)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A !(B (C+(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_6_i475_3_lut_4_lut_4_lut.init = 16'h9936;
    LUT4 n284_bdd_3_lut_24447_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n26172)) /* synthesis lut_function=(A (B (C+(D))+!B ((D)+!C))+!A !(B (C+(D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam n284_bdd_3_lut_24447_4_lut.init = 16'haa96;
    LUT4 i19366_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[2]), .C(index_i[1]), 
         .D(index_i[3]), .Z(n21721)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+!(D)))+!A (B (D)+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19366_3_lut_4_lut_4_lut.init = 16'hd699;
    LUT4 mux_229_Mux_6_i15_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[1]), .D(index_i[3]), .Z(n15_adj_2503)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !((D)+!C))+!A !(B+!((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_6_i15_3_lut_4_lut_4_lut.init = 16'h66d6;
    LUT4 mux_229_Mux_9_i316_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n316_adj_2487)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C+(D)))+!A (B (C (D)+!C !(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_9_i316_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h3ff8;
    LUT4 mux_229_Mux_5_i572_3_lut_4_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[1]), .D(index_i[3]), .Z(n572_adj_2680)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A !(B (C+(D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_5_i572_3_lut_4_lut.init = 16'haa95;
    LUT4 mux_230_Mux_0_i124_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n124_adj_2703)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A !(B (D)+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_0_i124_3_lut_4_lut_4_lut.init = 16'h6c99;
    LUT4 i20169_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n22524)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i20169_3_lut_4_lut.init = 16'h64cc;
    PFUMX i23671 (.BLUT(n25357), .ALUT(n25354), .C0(index_q[6]), .Z(n23116));
    LUT4 mux_229_Mux_1_i93_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[1]), .D(index_i[3]), .Z(n93_adj_2426)) /* synthesis lut_function=(A (B (C (D))+!B !(D))+!A !(B (C (D))+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_1_i93_3_lut_4_lut_4_lut.init = 16'h9566;
    LUT4 mux_229_Mux_5_i475_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[1]), .D(index_i[3]), .Z(n475_adj_2530)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (D)+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_5_i475_3_lut_4_lut_4_lut.init = 16'hd499;
    LUT4 mux_229_Mux_0_i157_3_lut_4_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[1]), .D(index_i[3]), .Z(n157_adj_2712)) /* synthesis lut_function=(A (B (C+!(D))+!B !(D))+!A (B (D)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_0_i157_3_lut_4_lut.init = 16'hd4aa;
    LUT4 mux_229_Mux_0_i635_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n635_adj_2738)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_0_i635_3_lut_4_lut_4_lut.init = 16'hfd0a;
    LUT4 i22900_3_lut (.A(n23744), .B(n23745), .C(index_q[8]), .Z(n23748)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22900_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_520_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n27185)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_2_lut_rep_520_3_lut_4_lut.init = 16'h8000;
    LUT4 i20088_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n22443)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (D))+!A !(D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20088_3_lut_4_lut_4_lut_4_lut.init = 16'ha25d;
    LUT4 mux_229_Mux_8_i635_3_lut_4_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n635_adj_2365)) /* synthesis lut_function=(!(A (B (C (D))+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_8_i635_3_lut_4_lut_3_lut_4_lut.init = 16'h0ff8;
    LUT4 i19395_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[2]), .C(index_i[1]), 
         .D(index_i[3]), .Z(n21750)) /* synthesis lut_function=(A ((C (D))+!B)+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19395_3_lut_4_lut_4_lut.init = 16'he666;
    LUT4 mux_229_Mux_4_i252_4_lut_4_lut (.A(index_i[0]), .B(index_i[3]), 
         .C(n27322), .D(index_i[4]), .Z(n252_adj_2762)) /* synthesis lut_function=(!(A (B (D)+!B !(D))+!A !(B ((D)+!C)+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_4_i252_4_lut_4_lut.init = 16'h669d;
    LUT4 mux_229_Mux_2_i348_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[1]), .D(index_i[3]), .Z(n348_adj_2753)) /* synthesis lut_function=(!(A (B (D)+!B (C+!(D)))+!A !(B (D)+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_2_i348_3_lut_4_lut_4_lut.init = 16'h4699;
    LUT4 i21015_3_lut (.A(n27427), .B(n29935), .C(index_q[3]), .Z(n23389)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21015_3_lut.init = 16'hcaca;
    LUT4 i21014_3_lut (.A(n27425), .B(n108), .C(index_q[3]), .Z(n23388)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21014_3_lut.init = 16'hcaca;
    PFUMX i24654 (.BLUT(n26453), .ALUT(n26452), .C0(index_i[5]), .Z(n26454));
    LUT4 i20076_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[2]), .C(index_i[1]), 
         .D(index_i[3]), .Z(n22431)) /* synthesis lut_function=(!(A (B+!((D)+!C))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20076_3_lut_4_lut_4_lut.init = 16'h6646;
    LUT4 mux_229_Mux_4_i205_3_lut_4_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[1]), .D(index_i[3]), .Z(n205_adj_2756)) /* synthesis lut_function=(!(A (B (D)+!B (C (D)))+!A !(B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_4_i205_3_lut_4_lut.init = 16'h46aa;
    LUT4 n15000_bdd_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n26388)) /* synthesis lut_function=(A (B (C+!(D))+!B ((D)+!C))+!A (B (C (D)+!C !(D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n15000_bdd_3_lut_4_lut_4_lut_4_lut.init = 16'hf38f;
    LUT4 mux_229_Mux_1_i62_3_lut_4_lut (.A(index_i[0]), .B(index_i[3]), 
         .C(index_i[2]), .D(index_i[4]), .Z(n62_adj_2763)) /* synthesis lut_function=(A (B (D)+!B ((D)+!C))+!A !(B (D)+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_1_i62_3_lut_4_lut.init = 16'haa56;
    LUT4 i20019_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n22374)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A (B (C)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20019_3_lut_4_lut_4_lut.init = 16'h3c8c;
    PFUMX i19835 (.BLUT(n22188), .ALUT(n22189), .C0(index_i[5]), .Z(n22190));
    LUT4 index_q_1__bdd_4_lut_26068 (.A(index_q[1]), .B(index_q[0]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n27480)) /* synthesis lut_function=(!(A (B (D)+!B (C+!(D)))+!A !(B (C (D)+!C !(D))+!B !((D)+!C)))) */ ;
    defparam index_q_1__bdd_4_lut_26068.init = 16'h429c;
    LUT4 i7273_2_lut_rep_663 (.A(index_q[3]), .B(index_q[4]), .Z(n27328)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i7273_2_lut_rep_663.init = 16'heeee;
    L6MUX21 i20446 (.D0(n22433), .D1(n22445), .SD(index_i[5]), .Z(n22820));
    L6MUX21 i21011 (.D0(n23383), .D1(n23384), .SD(index_q[5]), .Z(n23385));
    L6MUX21 i21018 (.D0(n23390), .D1(n23391), .SD(index_q[5]), .Z(n23392));
    L6MUX21 i20450 (.D0(n21695), .D1(n18090), .SD(index_i[5]), .Z(n22824));
    L6MUX21 i20451 (.D0(n21698), .D1(n11931), .SD(index_i[5]), .Z(n22825));
    LUT4 n23315_bdd_3_lut_23503 (.A(n23315), .B(n21815), .C(index_q[7]), 
         .Z(n24990)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n23315_bdd_3_lut_23503.init = 16'hcaca;
    L6MUX21 i21025 (.D0(n23397), .D1(n23398), .SD(index_q[5]), .Z(n23399));
    LUT4 i21013_3_lut (.A(n619), .B(n27297), .C(index_q[3]), .Z(n23387)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21013_3_lut.init = 16'hcaca;
    LUT4 i21012_3_lut (.A(n14_adj_2290), .B(n29916), .C(index_q[3]), .Z(n23386)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21012_3_lut.init = 16'hcaca;
    PFUMX i20453 (.BLUT(n542_adj_2561), .ALUT(n573_adj_2616), .C0(index_i[5]), 
          .Z(n22827));
    LUT4 i19715_then_4_lut (.A(index_q[2]), .B(index_q[1]), .C(index_q[4]), 
         .D(index_q[3]), .Z(n27462)) /* synthesis lut_function=(A (B (C+(D))+!B !(C))+!A !(B (C+(D))+!B !(C+!(D)))) */ ;
    defparam i19715_then_4_lut.init = 16'h9a97;
    PFUMX i20454 (.BLUT(n605_adj_2764), .ALUT(n636_adj_2765), .C0(index_i[5]), 
          .Z(n22828));
    LUT4 i11564_2_lut_3_lut_4_lut (.A(n27220), .B(n27328), .C(index_q[6]), 
         .D(index_q[5]), .Z(n254)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i11564_2_lut_3_lut_4_lut.init = 16'hfef0;
    L6MUX21 i23335 (.D0(n24932), .D1(n24929), .SD(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_2160[4]));
    LUT4 i19715_else_4_lut (.A(index_q[2]), .B(index_q[1]), .C(index_q[4]), 
         .D(index_q[3]), .Z(n27461)) /* synthesis lut_function=(!(A (B (C)+!B (C+(D)))+!A !(B (C (D)+!C !(D))+!B (C+!(D))))) */ ;
    defparam i19715_else_4_lut.init = 16'h581f;
    PFUMX i20455 (.BLUT(n669_adj_2559), .ALUT(n700_adj_2736), .C0(index_i[5]), 
          .Z(n22829));
    LUT4 i11776_2_lut_rep_620 (.A(index_q[0]), .B(index_q[1]), .Z(n27285)) /* synthesis lut_function=((B)+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i11776_2_lut_rep_620.init = 16'hdddd;
    PFUMX i20456 (.BLUT(n732_adj_2734), .ALUT(n21704), .C0(index_i[5]), 
          .Z(n22830));
    PFUMX i26394 (.BLUT(n29231), .ALUT(n173_adj_2729), .C0(index_q[5]), 
          .Z(n29232));
    LUT4 mux_230_Mux_6_i285_3_lut_4_lut (.A(n27285), .B(index_q[2]), .C(index_q[3]), 
         .D(n29945), .Z(n285_adj_2684)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_6_i285_3_lut_4_lut.init = 16'hf606;
    PFUMX i26392 (.BLUT(n29229), .ALUT(n29228), .C0(index_q[3]), .Z(n29230));
    PFUMX i20457 (.BLUT(n797_adj_2557), .ALUT(n828_adj_2555), .C0(index_i[5]), 
          .Z(n22831));
    LUT4 mux_230_Mux_6_i325_3_lut_4_lut_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n356)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_6_i325_3_lut_4_lut_3_lut.init = 16'h6d6d;
    L6MUX21 i26396 (.D0(n29232), .D1(n29230), .SD(index_q[4]), .Z(n29233));
    PFUMX i20458 (.BLUT(n860_adj_2766), .ALUT(n891_adj_2553), .C0(index_i[5]), 
          .Z(n22832));
    LUT4 mux_230_Mux_0_i635_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n635_adj_2391)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_0_i635_3_lut_4_lut_4_lut.init = 16'hfd0a;
    PFUMX i19844 (.BLUT(n22197), .ALUT(n22198), .C0(index_i[5]), .Z(n22199));
    LUT4 i19828_3_lut_4_lut (.A(n27285), .B(index_q[2]), .C(index_q[3]), 
         .D(n29949), .Z(n22183)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i19828_3_lut_4_lut.init = 16'hf606;
    LUT4 i21008_3_lut (.A(n29935), .B(n29926), .C(index_q[3]), .Z(n23382)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21008_3_lut.init = 16'hcaca;
    LUT4 i21007_3_lut (.A(n38), .B(n27427), .C(index_q[3]), .Z(n23381)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21007_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_6_i564_3_lut_4_lut_3_lut_rep_623 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n27288)) /* synthesis lut_function=(A (B)+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_6_i564_3_lut_4_lut_3_lut_rep_623.init = 16'hd9d9;
    LUT4 mux_229_Mux_7_i526_3_lut_3_lut_4_lut_4_lut_3_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n526_adj_2562)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(D))+!A !(D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_7_i526_3_lut_3_lut_4_lut_4_lut_3_lut_4_lut.init = 16'h887f;
    PFUMX i19853 (.BLUT(n22206), .ALUT(n22207), .C0(index_i[5]), .Z(n22208));
    PFUMX i19862 (.BLUT(n22215), .ALUT(n22216), .C0(index_i[5]), .Z(n22217));
    LUT4 mux_230_Mux_3_i652_rep_624 (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .Z(n27289)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_3_i652_rep_624.init = 16'h4d4d;
    LUT4 i20606_3_lut (.A(n26664), .B(n22971), .C(index_i[6]), .Z(n22980)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20606_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_8_i93_3_lut_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n93_adj_2550)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (D))+!A (B ((D)+!C)+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_8_i93_3_lut_3_lut_4_lut_4_lut.init = 16'h08f3;
    LUT4 mux_230_Mux_6_i300_3_lut_rep_626 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n27291)) /* synthesis lut_function=(A (B+!(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_6_i300_3_lut_rep_626.init = 16'hdada;
    LUT4 i19813_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n22168)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D))+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i19813_3_lut_4_lut.init = 16'hccdb;
    LUT4 i19719_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n22074)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i19719_3_lut_4_lut_4_lut.init = 16'hda5a;
    LUT4 i9567_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n12053)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A (B (C+!(D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i9567_3_lut_4_lut_4_lut.init = 16'hd966;
    LUT4 i19839_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n22194)) /* synthesis lut_function=(!(A (B (C (D))+!B (C (D)+!C !(D)))+!A !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i19839_3_lut_4_lut_4_lut.init = 16'h5aad;
    LUT4 mux_230_Mux_3_i653_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n653_adj_2678)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A !(B (D)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_3_i653_3_lut_4_lut_4_lut.init = 16'h4d99;
    LUT4 mux_230_Mux_6_i572_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n572_adj_2767)) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_6_i572_3_lut_4_lut.init = 16'hccd9;
    LUT4 i19738_3_lut_4_lut_4_lut (.A(index_q[2]), .B(index_q[1]), .C(index_q[0]), 
         .D(index_q[3]), .Z(n22093)) /* synthesis lut_function=(A (B (C)+!B !(C+!(D)))+!A (B (C+!(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i19738_3_lut_4_lut_4_lut.init = 16'hc3c4;
    LUT4 i19692_3_lut (.A(n27274), .B(n29938), .C(index_q[3]), .Z(n22047)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19692_3_lut.init = 16'hcaca;
    LUT4 n21642_bdd_3_lut_24366_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n25710)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C))+!A !(B (C+!(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam n21642_bdd_3_lut_24366_4_lut_4_lut.init = 16'h5ad6;
    LUT4 mux_230_Mux_4_i812_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[2]), 
         .C(index_q[4]), .D(index_q[3]), .Z(n812_adj_2768)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A !(B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_4_i812_3_lut_4_lut_4_lut.init = 16'ha595;
    LUT4 i20026_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n22381)) /* synthesis lut_function=(A (B (C+(D))+!B ((D)+!C))+!A !(B (C+(D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20026_3_lut_4_lut.init = 16'haa96;
    LUT4 mux_229_Mux_6_i812_3_lut_4_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n812_adj_2554)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(D))+!A !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_6_i812_3_lut_4_lut_3_lut_4_lut.init = 16'h7780;
    LUT4 n18312_bdd_4_lut_then_4_lut (.A(index_q[3]), .B(index_q[4]), .C(index_q[1]), 
         .D(index_q[2]), .Z(n27550)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B+(C (D)+!C !(D)))) */ ;
    defparam n18312_bdd_4_lut_then_4_lut.init = 16'hf44f;
    LUT4 mux_230_Mux_4_i827_3_lut_rep_528_3_lut (.A(index_q[0]), .B(index_q[2]), 
         .C(index_q[3]), .Z(n27193)) /* synthesis lut_function=(A (B+(C))+!A !(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_4_i827_3_lut_rep_528_3_lut.init = 16'ha9a9;
    LUT4 mux_229_Mux_4_i1002_3_lut_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n1002_adj_2499)) /* synthesis lut_function=(A (B (C (D))+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_4_i1002_3_lut_3_lut_3_lut_4_lut.init = 16'hf007;
    LUT4 i12452_2_lut_rep_628 (.A(index_q[0]), .B(index_q[1]), .Z(n27293)) /* synthesis lut_function=(A (B)) */ ;
    defparam i12452_2_lut_rep_628.init = 16'h8888;
    LUT4 mux_230_Mux_8_i860_3_lut_4_lut (.A(n27219), .B(index_q[3]), .C(index_q[4]), 
         .D(n27166), .Z(n860_adj_2501)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_8_i860_3_lut_4_lut.init = 16'h08f8;
    LUT4 i20924_3_lut_4_lut (.A(n27219), .B(index_q[3]), .C(index_q[4]), 
         .D(n364_adj_2644), .Z(n23298)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i20924_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_230_Mux_3_i1002_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n20198)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (D))+!A (D)) */ ;
    defparam mux_230_Mux_3_i1002_3_lut_3_lut_4_lut.init = 16'hf708;
    PFUMX i20492 (.BLUT(n94_adj_2545), .ALUT(n125_adj_2543), .C0(index_i[5]), 
          .Z(n22866));
    LUT4 mux_230_Mux_7_i491_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n491_adj_2769)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(D))+!A (B (C+!(D))+!B !(D)))) */ ;
    defparam mux_230_Mux_7_i491_3_lut_4_lut_4_lut_4_lut.init = 16'h3780;
    PFUMX i20493 (.BLUT(n18119), .ALUT(n14743), .C0(index_i[5]), .Z(n22867));
    LUT4 mux_230_Mux_1_i348_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n348_adj_2659)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A (B (C+!(D))+!B !(D)))) */ ;
    defparam mux_230_Mux_1_i348_3_lut_4_lut_4_lut.init = 16'h3f80;
    L6MUX21 i24611 (.D0(n26389), .D1(n26386), .SD(index_i[5]), .Z(n26390));
    LUT4 i19869_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n22224)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A (B (C)+!B !(C (D))))) */ ;
    defparam i19869_3_lut_4_lut_4_lut.init = 16'h3c8c;
    LUT4 i11632_2_lut_rep_453_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[4]), .D(n27317), .Z(n27118)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;
    defparam i11632_2_lut_rep_453_3_lut_4_lut.init = 16'hf8f0;
    LUT4 i22131_3_lut (.A(n620_adj_2770), .B(n14788), .C(index_i[4]), 
         .Z(n22198)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22131_3_lut.init = 16'hcaca;
    PFUMX i24609 (.BLUT(n26388), .ALUT(n26387), .C0(index_i[4]), .Z(n26389));
    LUT4 i11631_2_lut_rep_507_3_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .Z(n27172)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam i11631_2_lut_rep_507_3_lut.init = 16'hf8f8;
    L6MUX21 i20495 (.D0(n21710), .D1(n21713), .SD(index_i[5]), .Z(n22869));
    L6MUX21 i20496 (.D0(n21716), .D1(n21719), .SD(index_i[5]), .Z(n22870));
    LUT4 i7987_2_lut_rep_706 (.A(index_q[1]), .B(index_q[2]), .Z(n27371)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i7987_2_lut_rep_706.init = 16'h8888;
    LUT4 i9609_2_lut_3_lut (.A(index_q[1]), .B(index_q[2]), .C(index_q[3]), 
         .Z(n12095)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i9609_2_lut_3_lut.init = 16'h8080;
    LUT4 mux_230_Mux_5_i700_3_lut (.A(n460_adj_2709), .B(n29945), .C(index_q[4]), 
         .Z(n700_adj_2591)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_5_i700_3_lut.init = 16'hcaca;
    LUT4 n18312_bdd_4_lut_else_4_lut (.A(index_q[3]), .B(index_q[4]), .C(index_q[1]), 
         .D(index_q[2]), .Z(n27549)) /* synthesis lut_function=(!(A (B (D)+!B ((D)+!C))+!A !(B+!((D)+!C)))) */ ;
    defparam n18312_bdd_4_lut_else_4_lut.init = 16'h44fc;
    L6MUX21 i21431 (.D0(n23789), .D1(n23790), .SD(index_q[5]), .Z(n23805));
    LUT4 i19687_3_lut_4_lut (.A(n27285), .B(index_q[2]), .C(index_q[3]), 
         .D(n27280), .Z(n22042)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i19687_3_lut_4_lut.init = 16'h6f60;
    L6MUX21 i21432 (.D0(n23791), .D1(n23792), .SD(index_q[5]), .Z(n23806));
    L6MUX21 i21433 (.D0(n23793), .D1(n23794), .SD(index_q[5]), .Z(n23807));
    LUT4 i15925_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .D(index_q[0]), .Z(n18111)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C (D)+!C !(D)))+!A !(B (D)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i15925_3_lut_4_lut_4_lut_4_lut.init = 16'h83fc;
    LUT4 index_q_6__bdd_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[6]), .D(n27307), .Z(n25777)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)+!C !(D)))+!A (B (C (D))+!B (C (D)+!C !(D))))) */ ;
    defparam index_q_6__bdd_4_lut_4_lut_4_lut.init = 16'h0f7c;
    PFUMX i24605 (.BLUT(n78), .ALUT(n26385), .C0(index_i[4]), .Z(n26386));
    LUT4 i11656_2_lut_rep_516_3_lut (.A(index_q[1]), .B(index_q[2]), .C(index_q[3]), 
         .Z(n27181)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i11656_2_lut_rep_516_3_lut.init = 16'hf8f8;
    PFUMX i20497 (.BLUT(n413_adj_2533), .ALUT(n444_adj_2435), .C0(index_i[5]), 
          .Z(n22871));
    LUT4 mux_230_Mux_1_i317_3_lut (.A(n301_adj_2759), .B(n908_adj_2751), 
         .C(index_q[4]), .Z(n317_adj_2690)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_1_i317_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_3_i93_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n93_adj_2687)) /* synthesis lut_function=(A (B (C+!(D))+!B (D))+!A (B ((D)+!C)+!B (D))) */ ;
    defparam mux_230_Mux_3_i93_3_lut_4_lut_4_lut_4_lut.init = 16'hf78c;
    LUT4 mux_230_Mux_8_i412_3_lut_4_lut_3_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .Z(n15090)) /* synthesis lut_function=(A (B+!(C))+!A !((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_8_i412_3_lut_4_lut_3_lut.init = 16'h8e8e;
    LUT4 mux_230_Mux_9_i412_3_lut_3_lut_4_lut_3_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .Z(n412_adj_2294)) /* synthesis lut_function=(!(A (B (C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_9_i412_3_lut_3_lut_4_lut_3_lut.init = 16'h7e7e;
    PFUMX i20498 (.BLUT(n476_adj_2531), .ALUT(n507), .C0(index_i[5]), 
          .Z(n22872));
    LUT4 n347_bdd_3_lut_25118_4_lut (.A(n27384), .B(index_i[2]), .C(index_i[3]), 
         .D(n27350), .Z(n25825)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n347_bdd_3_lut_25118_4_lut.init = 16'hf606;
    LUT4 mux_230_Mux_3_i460_3_lut_4_lut (.A(n27285), .B(index_q[2]), .C(index_q[3]), 
         .D(n27278), .Z(n460_adj_2683)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_3_i460_3_lut_4_lut.init = 16'h6f60;
    PFUMX i20499 (.BLUT(n18093), .ALUT(n573_adj_2708), .C0(index_i[5]), 
          .Z(n22873));
    PFUMX i20500 (.BLUT(n605), .ALUT(n636_adj_2528), .C0(index_i[5]), 
          .Z(n22874));
    LUT4 mux_230_Mux_9_i30_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[0]), .D(index_q[3]), .Z(n30_adj_2546)) /* synthesis lut_function=(A (B (C (D))+!B !(D))+!A !(B+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_9_i30_3_lut_4_lut_4_lut_4_lut.init = 16'h8033;
    LUT4 mux_230_Mux_8_i526_3_lut_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n526_adj_2367)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D)))) */ ;
    defparam mux_230_Mux_8_i526_3_lut_3_lut_3_lut_4_lut.init = 16'h0f70;
    L6MUX21 i21434 (.D0(n23795), .D1(n23796), .SD(index_q[5]), .Z(n23808));
    LUT4 i11994_2_lut_rep_543_3_lut (.A(index_q[1]), .B(index_q[2]), .C(index_q[0]), 
         .Z(n27208)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i11994_2_lut_rep_543_3_lut.init = 16'h7070;
    LUT4 mux_230_Mux_4_i93_3_lut_4_lut_3_lut_rep_644_4_lut (.A(index_q[1]), 
         .B(index_q[2]), .C(index_q[3]), .D(index_q[0]), .Z(n27309)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_4_i93_3_lut_4_lut_3_lut_rep_644_4_lut.init = 16'h07f0;
    LUT4 i12124_2_lut_rep_546_3_lut (.A(index_q[1]), .B(index_q[2]), .C(index_q[0]), 
         .Z(n27211)) /* synthesis lut_function=(A (B+!(C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i12124_2_lut_rep_546_3_lut.init = 16'h8f8f;
    PFUMX i20501 (.BLUT(n21722), .ALUT(n700_adj_2771), .C0(index_i[5]), 
          .Z(n22875));
    LUT4 i22751_3_lut (.A(n12129), .B(n892_adj_2598), .C(index_i[6]), 
         .Z(n22856)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22751_3_lut.init = 16'hcaca;
    LUT4 i19699_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .D(index_q[0]), .Z(n22054)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C (D)+!C !(D)))+!A !(B (D)+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i19699_3_lut_4_lut_4_lut_4_lut.init = 16'h7c03;
    LUT4 i19717_3_lut_3_lut_4_lut (.A(index_q[1]), .B(index_q[2]), .C(index_q[3]), 
         .D(index_q[0]), .Z(n22072)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i19717_3_lut_3_lut_4_lut.init = 16'hf80f;
    LUT4 i12580_2_lut_rep_553_3_lut (.A(index_q[1]), .B(index_q[2]), .C(index_q[0]), 
         .Z(n27218)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i12580_2_lut_rep_553_3_lut.init = 16'h8080;
    LUT4 i1_3_lut_rep_513_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(n27328), .Z(n27178)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;
    defparam i1_3_lut_rep_513_4_lut.init = 16'hfff8;
    LUT4 mux_229_Mux_0_i348_3_lut_4_lut (.A(n27384), .B(index_i[2]), .C(index_i[3]), 
         .D(n27388), .Z(n348_adj_2720)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_0_i348_3_lut_4_lut.init = 16'h6f60;
    LUT4 i11888_4_lut (.A(n15358), .B(index_i[8]), .C(n765_adj_2772), 
         .D(index_i[7]), .Z(n1022)) /* synthesis lut_function=(A (B+(C (D)))+!A (B+(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11888_4_lut.init = 16'hfcdd;
    LUT4 mux_230_Mux_3_i142_3_lut_3_lut_3_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .Z(n142_adj_2672)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_3_i142_3_lut_3_lut_3_lut.init = 16'h3838;
    L6MUX21 i20502 (.D0(n732_adj_2706), .D1(n21725), .SD(index_i[5]), 
            .Z(n22876));
    PFUMX i20503 (.BLUT(n797_adj_2742), .ALUT(n828_adj_2773), .C0(index_i[5]), 
          .Z(n22877));
    LUT4 i9591_3_lut_3_lut_4_lut (.A(index_q[3]), .B(index_q[4]), .C(n27278), 
         .D(index_q[0]), .Z(n605_adj_2588)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i9591_3_lut_3_lut_4_lut.init = 16'h10fe;
    LUT4 i1_3_lut_4_lut_adj_86 (.A(index_q[3]), .B(index_q[4]), .C(index_q[5]), 
         .D(n27371), .Z(n20671)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i1_3_lut_4_lut_adj_86.init = 16'hfffe;
    LUT4 i11623_2_lut_rep_461_3_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .D(index_q[0]), .Z(n27126)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i11623_2_lut_rep_461_3_lut_4_lut.init = 16'hf8f0;
    LUT4 i12497_2_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(n27323), 
         .D(index_q[2]), .Z(n15104)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;
    defparam i12497_2_lut_3_lut_4_lut.init = 16'hf080;
    LUT4 mux_230_Mux_7_i315_3_lut_rep_573_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n27238)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B+!(C)))) */ ;
    defparam mux_230_Mux_7_i315_3_lut_rep_573_3_lut.init = 16'h3838;
    LUT4 i11625_4_lut (.A(n15412), .B(index_q[8]), .C(n765), .D(index_q[7]), 
         .Z(n1022_adj_2774)) /* synthesis lut_function=(A (B+(C (D)))+!A (B+(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i11625_4_lut.init = 16'hfcdd;
    PFUMX i20504 (.BLUT(n860_adj_2525), .ALUT(n891_adj_2524), .C0(index_i[5]), 
          .Z(n22878));
    LUT4 mux_230_Mux_8_i491_3_lut_3_lut_3_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .D(index_q[0]), .Z(n491_adj_2693)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_8_i491_3_lut_3_lut_3_lut_4_lut.init = 16'h7870;
    LUT4 i19801_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[0]), .D(index_q[3]), .Z(n22156)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(D))+!A (B+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i19801_3_lut_4_lut_4_lut_4_lut.init = 16'h3380;
    LUT4 index_q_6__bdd_3_lut_24247_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(n27317), .D(index_q[6]), .Z(n25778)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (C+!(D))) */ ;
    defparam index_q_6__bdd_3_lut_24247_4_lut.init = 16'hf07f;
    PFUMX i25174 (.BLUT(n27504), .ALUT(n27505), .C0(index_i[3]), .Z(n27506));
    LUT4 i19830_3_lut (.A(n900), .B(n29919), .C(index_q[3]), .Z(n22185)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19830_3_lut.init = 16'hcaca;
    PFUMX mux_230_Mux_7_i190 (.BLUT(n22001), .ALUT(n173_adj_2292), .C0(index_q[5]), 
          .Z(n190)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 i2685_2_lut_rep_582 (.A(index_i[0]), .B(index_i[1]), .Z(n27247)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i2685_2_lut_rep_582.init = 16'h6666;
    L6MUX21 i21435 (.D0(n23797), .D1(n23798), .SD(index_q[5]), .Z(n23809));
    PFUMX mux_230_Mux_8_i764 (.BLUT(n716_adj_2271), .ALUT(n732_adj_2522), 
          .C0(n22671), .Z(n764)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 mux_229_Mux_3_i507_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[4]), .D(n491_adj_2379), .Z(n507_adj_2775)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_3_i507_3_lut_4_lut.init = 16'h6f60;
    PFUMX mux_230_Mux_8_i574 (.BLUT(n542_adj_2368), .ALUT(n12046), .C0(index_q[5]), 
          .Z(n574_adj_2430)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 i19727_then_4_lut (.A(index_q[0]), .B(index_q[4]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n27465)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C))+!A (B (C)+!B !(C+!(D)))) */ ;
    defparam i19727_then_4_lut.init = 16'hc34a;
    LUT4 i11721_2_lut_rep_439_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n27104)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;
    defparam i11721_2_lut_rep_439_3_lut_4_lut.init = 16'hf080;
    L6MUX21 i21436 (.D0(n23799), .D1(n23800), .SD(index_q[5]), .Z(n23810));
    LUT4 mux_230_Mux_4_i1002_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n1002_adj_2691)) /* synthesis lut_function=(A (B (C (D))+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D))) */ ;
    defparam mux_230_Mux_4_i1002_3_lut_3_lut_4_lut.init = 16'hf007;
    LUT4 i21005_3_lut (.A(n29926), .B(n14_adj_2290), .C(index_q[3]), .Z(n23379)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21005_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_6_i812_3_lut_4_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n812_adj_2628)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(D))+!A !(D))) */ ;
    defparam mux_230_Mux_6_i812_3_lut_4_lut_3_lut_4_lut.init = 16'h7780;
    PFUMX i24590 (.BLUT(n26359), .ALUT(n26358), .C0(index_q[4]), .Z(n26360));
    L6MUX21 i21437 (.D0(n23801), .D1(n23802), .SD(index_q[5]), .Z(n23811));
    PFUMX i20523 (.BLUT(n94_adj_2518), .ALUT(n21728), .C0(index_i[5]), 
          .Z(n22897));
    LUT4 i19390_3_lut (.A(n900_adj_2707), .B(n356_adj_2398), .C(index_i[3]), 
         .Z(n21745)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19390_3_lut.init = 16'hcaca;
    L6MUX21 i21438 (.D0(n23803), .D1(n23804), .SD(index_q[5]), .Z(n23812));
    LUT4 mux_230_Mux_5_i30_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n30_adj_2465)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A (B+!(C+(D)))) */ ;
    defparam mux_230_Mux_5_i30_3_lut_4_lut.init = 16'hcc67;
    LUT4 n12162_bdd_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[4]), 
         .D(index_q[2]), .Z(n26533)) /* synthesis lut_function=(A (B)+!A !(B (D)+!B !(C (D)))) */ ;
    defparam n12162_bdd_3_lut_4_lut.init = 16'h98cc;
    LUT4 i19806_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n22161)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+(D)))+!A !(B (D)+!B !((D)+!C))) */ ;
    defparam i19806_3_lut_4_lut_4_lut.init = 16'h99c7;
    LUT4 i19727_else_4_lut (.A(index_q[0]), .B(index_q[4]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n27464)) /* synthesis lut_function=(A (C)+!A !(B ((D)+!C)+!B !(C))) */ ;
    defparam i19727_else_4_lut.init = 16'hb0f0;
    LUT4 i12548_2_lut_rep_631 (.A(index_q[0]), .B(index_q[1]), .Z(n27296)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i12548_2_lut_rep_631.init = 16'heeee;
    LUT4 i22324_3_lut (.A(n27480), .B(n22183), .C(index_q[4]), .Z(n22184)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22324_3_lut.init = 16'hcaca;
    PFUMX i20525 (.BLUT(n221_adj_2757), .ALUT(n252_adj_2762), .C0(index_i[5]), 
          .Z(n22899));
    LUT4 mux_229_Mux_3_i890_3_lut_4_lut (.A(n27384), .B(index_i[2]), .C(index_i[3]), 
         .D(n356_adj_2398), .Z(n890_adj_2484)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_3_i890_3_lut_4_lut.init = 16'h6f60;
    PFUMX i23333 (.BLUT(n24931), .ALUT(n24930), .C0(index_q[8]), .Z(n24932));
    PFUMX i20526 (.BLUT(n286_adj_2515), .ALUT(n21731), .C0(index_i[5]), 
          .Z(n22900));
    LUT4 i11917_4_lut (.A(n15146), .B(index_i[7]), .C(n892_adj_2439), 
         .D(index_i[6]), .Z(n1021)) /* synthesis lut_function=(A (B+(C (D)))+!A (B+(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11917_4_lut.init = 16'hfcdd;
    LUT4 mux_230_Mux_7_i572_3_lut_rep_410_3_lut_3_lut_4_lut (.A(index_q[0]), 
         .B(index_q[1]), .C(index_q[3]), .D(index_q[2]), .Z(n27075)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)+!C !(D)))) */ ;
    defparam mux_230_Mux_7_i572_3_lut_rep_410_3_lut_3_lut_4_lut.init = 16'hfe01;
    LUT4 i11820_2_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n635_adj_2275)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A (B (C+!(D))+!B (C+(D)))) */ ;
    defparam i11820_2_lut_4_lut_4_lut.init = 16'hf1fc;
    PFUMX i20527 (.BLUT(n349_adj_2276), .ALUT(n21734), .C0(index_i[5]), 
          .Z(n22901));
    LUT4 mux_229_Mux_4_i653_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n653_adj_2459)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A (B (C (D)+!C !(D))+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_4_i653_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hc837;
    LUT4 i22154_3_lut (.A(n491_adj_2776), .B(n506_adj_2777), .C(index_i[4]), 
         .Z(n22180)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22154_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_0_i333_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n333_adj_2632)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B (D))) */ ;
    defparam mux_230_Mux_0_i333_3_lut_3_lut_4_lut.init = 16'hf10e;
    LUT4 i20077_3_lut_4_lut (.A(n27384), .B(index_i[2]), .C(index_i[3]), 
         .D(n27345), .Z(n22432)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20077_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_230_Mux_3_i30_3_lut_3_lut_4_lut_3_lut_4_lut (.A(index_q[0]), 
         .B(index_q[1]), .C(index_q[3]), .D(index_q[2]), .Z(n30_adj_2471)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C+!(D)))) */ ;
    defparam mux_230_Mux_3_i30_3_lut_3_lut_4_lut_3_lut_4_lut.init = 16'hfe11;
    LUT4 i19818_3_lut (.A(n404), .B(n29948), .C(index_q[3]), .Z(n22173)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19818_3_lut.init = 16'hcaca;
    LUT4 i12444_1_lut_rep_416_2_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n27081)) /* synthesis lut_function=(!(A (C+(D))+!A (B (C+(D))+!B (C)))) */ ;
    defparam i12444_1_lut_rep_416_2_lut_3_lut_4_lut.init = 16'h010f;
    LUT4 i11660_2_lut_rep_462_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n27127)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i11660_2_lut_rep_462_3_lut_4_lut.init = 16'hfef0;
    LUT4 i22350_3_lut (.A(n22173), .B(n22174), .C(index_q[4]), .Z(n22175)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22350_3_lut.init = 16'hcaca;
    LUT4 i22768_3_lut (.A(n12048), .B(n892_adj_2502), .C(index_q[6]), 
         .Z(n23742)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22768_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_8_i397_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n397_adj_2539)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B ((D)+!C))) */ ;
    defparam mux_230_Mux_8_i397_3_lut_3_lut_4_lut.init = 16'hf10f;
    LUT4 n21809_bdd_3_lut_23506 (.A(n21809), .B(n27675), .C(index_q[7]), 
         .Z(n24993)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n21809_bdd_3_lut_23506.init = 16'hcaca;
    LUT4 i19383_3_lut (.A(n29956), .B(n27388), .C(index_i[3]), .Z(n21738)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19383_3_lut.init = 16'hcaca;
    PFUMX i20532 (.BLUT(n669_adj_2509), .ALUT(n700_adj_2507), .C0(index_i[5]), 
          .Z(n22906));
    LUT4 n168_bdd_3_lut_24457_4_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[3]), 
         .C(index_i[1]), .Z(n25837)) /* synthesis lut_function=(A (C)+!A (B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n168_bdd_3_lut_24457_4_lut_4_lut_3_lut.init = 16'he5e5;
    LUT4 mux_230_Mux_8_i46_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n46_adj_2481)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (B (C)+!B !(C (D)+!C !(D)))) */ ;
    defparam mux_230_Mux_8_i46_3_lut_4_lut_4_lut_4_lut.init = 16'hc1f0;
    LUT4 mux_229_Mux_0_i812_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n812_adj_2743)) /* synthesis lut_function=(A (B (C+(D))+!B !(C))+!A (B (D)+!B !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_0_i812_3_lut_4_lut_4_lut_4_lut.init = 16'hcf92;
    LUT4 mux_230_Mux_7_i924_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[4]), .D(n27317), .Z(n924_adj_2730)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B ((D)+!C))) */ ;
    defparam mux_230_Mux_7_i924_3_lut_3_lut_4_lut.init = 16'hf10f;
    LUT4 mux_230_Mux_3_i157_3_lut_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n157_adj_2298)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B !(C+(D))))) */ ;
    defparam mux_230_Mux_3_i157_3_lut_3_lut_3_lut_4_lut.init = 16'h1ff0;
    PFUMX i20533 (.BLUT(n21746), .ALUT(n763_adj_2438), .C0(index_i[5]), 
          .Z(n22907));
    LUT4 i19807_3_lut (.A(n404), .B(n27289), .C(index_q[3]), .Z(n22162)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19807_3_lut.init = 16'hcaca;
    PFUMX i20534 (.BLUT(n21749), .ALUT(n828_adj_2741), .C0(index_i[5]), 
          .Z(n22908));
    L6MUX21 i26153 (.D0(n28897), .D1(n28894), .SD(index_q[4]), .Z(n28898));
    PFUMX i26151 (.BLUT(n28896), .ALUT(n28895), .C0(index_q[5]), .Z(n28897));
    PFUMX i20535 (.BLUT(n860_adj_2504), .ALUT(n21752), .C0(index_i[5]), 
          .Z(n22909));
    LUT4 mux_229_Mux_0_i931_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n588)) /* synthesis lut_function=(!(A (B+(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_0_i931_3_lut_3_lut.init = 16'h5656;
    LUT4 mux_229_Mux_9_i62_3_lut_4_lut_then_4_lut (.A(index_i[4]), .B(index_i[2]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n27468)) /* synthesis lut_function=(!(A (B (C+(D)))+!A (B+(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_9_i62_3_lut_4_lut_then_4_lut.init = 16'h222b;
    PFUMX i26147 (.BLUT(n28893), .ALUT(n28892), .C0(index_q[3]), .Z(n28894));
    LUT4 i19849_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n22204)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B ((D)+!C)+!B (C))) */ ;
    defparam i19849_3_lut_4_lut_4_lut.init = 16'hfc1c;
    PFUMX i20554 (.BLUT(n94_adj_2745), .ALUT(n125_adj_2497), .C0(index_i[5]), 
          .Z(n22928));
    PFUMX i20555 (.BLUT(n158_adj_2494), .ALUT(n189_adj_2778), .C0(index_i[5]), 
          .Z(n22929));
    PFUMX i25172 (.BLUT(n27501), .ALUT(n27502), .C0(index_q[1]), .Z(n27503));
    LUT4 i11599_2_lut_rep_555_3_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .Z(n27220)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i11599_2_lut_rep_555_3_lut.init = 16'he0e0;
    PFUMX i20556 (.BLUT(n221_adj_2577), .ALUT(n252_adj_2779), .C0(index_i[5]), 
          .Z(n22930));
    LUT4 i11663_2_lut_rep_448_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[4]), .D(n27317), .Z(n27113)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i11663_2_lut_rep_448_3_lut_4_lut.init = 16'hfef0;
    LUT4 mux_229_Mux_1_i882_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n882_adj_2780)) /* synthesis lut_function=(A ((C)+!B)+!A !((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_1_i882_3_lut_3_lut.init = 16'ha6a6;
    PFUMX i20557 (.BLUT(n286_adj_2493), .ALUT(n22274), .C0(index_i[5]), 
          .Z(n22931));
    LUT4 mux_230_Mux_7_i141_3_lut_4_lut_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n308)) /* synthesis lut_function=(A ((C)+!B)+!A (B+!(C))) */ ;
    defparam mux_230_Mux_7_i141_3_lut_4_lut_3_lut.init = 16'he7e7;
    PFUMX i20558 (.BLUT(n349_adj_2781), .ALUT(n22277), .C0(index_i[5]), 
          .Z(n22932));
    LUT4 i11674_4_lut (.A(n27182), .B(index_q[7]), .C(n892_adj_2476), 
         .D(index_q[6]), .Z(n1021_adj_2722)) /* synthesis lut_function=(A (B+(C (D)))+!A (B+(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i11674_4_lut.init = 16'hfcdd;
    LUT4 mux_229_Mux_9_i62_3_lut_4_lut_else_4_lut (.A(index_i[4]), .B(index_i[2]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n27467)) /* synthesis lut_function=((B+(C (D)))+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_9_i62_3_lut_4_lut_else_4_lut.init = 16'hfddd;
    PFUMX i20559 (.BLUT(n413_adj_2491), .ALUT(n444_adj_2761), .C0(index_i[5]), 
          .Z(n22933));
    LUT4 n27296_bdd_4_lut (.A(n27296), .B(index_q[6]), .C(index_q[2]), 
         .D(index_q[5]), .Z(n27673)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A !(B (C+(D))+!B (D)))) */ ;
    defparam n27296_bdd_4_lut.init = 16'h5fe0;
    LUT4 i19752_3_lut_3_lut_4_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n22107)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B !((D)+!C)))) */ ;
    defparam i19752_3_lut_3_lut_4_lut_3_lut_4_lut.init = 16'h11ef;
    LUT4 n348_bdd_3_lut_24996_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n26116)) /* synthesis lut_function=(A (B (D)+!B (C+(D)))+!A (B (D)+!B !(C (D)+!C !(D)))) */ ;
    defparam n348_bdd_3_lut_24996_4_lut_4_lut.init = 16'hef30;
    PFUMX i20560 (.BLUT(n476_adj_2490), .ALUT(n507_adj_2775), .C0(index_i[5]), 
          .Z(n22934));
    LUT4 i19836_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n22191)) /* synthesis lut_function=(A (B (D)+!B ((D)+!C))+!A (B (D)+!B (C+!(D)))) */ ;
    defparam i19836_3_lut_4_lut_4_lut_4_lut.init = 16'hfe13;
    LUT4 mux_230_Mux_7_i29_3_lut_rep_632 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n27297)) /* synthesis lut_function=(A (B+!(C))+!A !((C)+!B)) */ ;
    defparam mux_230_Mux_7_i29_3_lut_rep_632.init = 16'h8e8e;
    LUT4 i19378_3_lut (.A(n27346), .B(n27256), .C(index_i[3]), .Z(n21733)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19378_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_5_i53_3_lut_4_lut_3_lut_rep_634 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n27299)) /* synthesis lut_function=(A ((C)+!B)+!A (B)) */ ;
    defparam mux_230_Mux_5_i53_3_lut_4_lut_3_lut_rep_634.init = 16'he6e6;
    LUT4 mux_230_Mux_6_i635_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n635_adj_2710)) /* synthesis lut_function=(A (B (C+(D))+!B !(D))+!A (B)) */ ;
    defparam mux_230_Mux_6_i635_3_lut_4_lut.init = 16'hcce6;
    LUT4 i20814_3_lut (.A(n23185), .B(n23186), .C(index_q[8]), .Z(n23188)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20814_3_lut.init = 16'hcaca;
    LUT4 i20813_3_lut (.A(n23183), .B(n23184), .C(index_q[8]), .Z(n23187)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20813_3_lut.init = 16'hcaca;
    LUT4 i19831_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n22186)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A (B (D)+!B !(C (D))))) */ ;
    defparam i19831_3_lut_4_lut.init = 16'h18cc;
    LUT4 i19734_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n22089)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)))+!A !(B (C+!(D))+!B (D)))) */ ;
    defparam i19734_3_lut_3_lut_4_lut.init = 16'h71cc;
    PFUMX i20561 (.BLUT(n22283), .ALUT(n573_adj_2411), .C0(index_i[5]), 
          .Z(n22935));
    LUT4 mux_230_Mux_0_i557_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n557_adj_2386)) /* synthesis lut_function=(A ((D)+!C)+!A !((D)+!B)) */ ;
    defparam mux_230_Mux_0_i557_3_lut_4_lut.init = 16'haa4e;
    LUT4 mux_230_Mux_3_i700_3_lut_4_lut (.A(index_q[4]), .B(index_q[3]), 
         .C(n684_adj_2477), .D(n29950), .Z(n700_adj_2643)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_3_i700_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i19377_3_lut (.A(n29952), .B(n356_adj_2398), .C(index_i[3]), 
         .Z(n21732)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19377_3_lut.init = 16'hcaca;
    LUT4 i22080_3_lut (.A(n21732), .B(n21733), .C(index_i[4]), .Z(n21734)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22080_3_lut.init = 16'hcaca;
    LUT4 i11494_2_lut_rep_716 (.A(index_i[1]), .B(index_i[2]), .Z(n27381)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11494_2_lut_rep_716.init = 16'h8888;
    LUT4 mux_229_Mux_7_i491_3_lut_4_lut_4_lut_4_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[2]), .D(index_i[3]), .Z(n491_adj_2776)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A (B ((D)+!C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_7_i491_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'h3870;
    PFUMX i20562 (.BLUT(n11965), .ALUT(n22286), .C0(index_i[5]), .Z(n22936));
    LUT4 mux_229_Mux_8_i491_3_lut_3_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n491_adj_2574)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_8_i491_3_lut_3_lut_3_lut_4_lut.init = 16'h7870;
    PFUMX i20563 (.BLUT(n669_adj_2486), .ALUT(n700_adj_2748), .C0(index_i[5]), 
          .Z(n22937));
    LUT4 i11862_2_lut_3_lut_4_lut (.A(n27224), .B(n27335), .C(index_i[6]), 
         .D(index_i[5]), .Z(n254_adj_2429)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i11862_2_lut_3_lut_4_lut.init = 16'hfef0;
    L6MUX21 i20564 (.D0(n22292), .D1(n763_adj_2701), .SD(index_i[5]), 
            .Z(n22938));
    LUT4 i22356_3_lut (.A(n22155), .B(n22156), .C(index_q[4]), .Z(n22157)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22356_3_lut.init = 16'hcaca;
    LUT4 n77_bdd_3_lut_3_lut_4_lut_4_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n26776)) /* synthesis lut_function=(A (B (C)+!B !(D))+!A !(D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n77_bdd_3_lut_3_lut_4_lut_4_lut_3_lut_4_lut.init = 16'h80f7;
    LUT4 i11489_2_lut_rep_487_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[3]), 
         .Z(n27152)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11489_2_lut_rep_487_3_lut.init = 16'hf8f8;
    PFUMX i20566 (.BLUT(n860_adj_2569), .ALUT(n891_adj_2485), .C0(index_i[5]), 
          .Z(n22940));
    LUT4 mux_229_Mux_5_i828_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[4]), .D(n27302), .Z(n828_adj_2773)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_5_i828_4_lut_4_lut.init = 16'hc66c;
    LUT4 i11778_2_lut_3_lut_3_lut (.A(index_q[3]), .B(index_q[1]), .C(index_q[0]), 
         .Z(n14376)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i11778_2_lut_3_lut_3_lut.init = 16'h4040;
    LUT4 i11845_4_lut_4_lut (.A(index_q[3]), .B(index_q[2]), .C(index_q[0]), 
         .D(index_q[1]), .Z(n875_adj_2425)) /* synthesis lut_function=((B (C)+!B (D))+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i11845_4_lut_4_lut.init = 16'hf7d5;
    PFUMX i20567 (.BLUT(n924_adj_2483), .ALUT(n22295), .C0(index_i[5]), 
          .Z(n22941));
    LUT4 i11832_2_lut_4_lut_4_lut_4_lut (.A(index_q[3]), .B(index_q[2]), 
         .C(index_q[1]), .D(index_q[0]), .Z(n668_adj_2397)) /* synthesis lut_function=(!(A+!(B (C)+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i11832_2_lut_4_lut_4_lut_4_lut.init = 16'h5041;
    LUT4 i20929_3_lut_4_lut_3_lut (.A(index_q[3]), .B(index_q[4]), .C(n27172), 
         .Z(n23303)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i20929_3_lut_4_lut_3_lut.init = 16'h6464;
    PFUMX i20568 (.BLUT(n22301), .ALUT(n1018), .C0(index_i[5]), .Z(n22942));
    PFUMX mux_229_Mux_1_i891 (.BLUT(n882_adj_2780), .ALUT(n890_adj_2587), 
          .C0(n27264), .Z(n891_adj_2536)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 i19771_4_lut_3_lut (.A(index_q[3]), .B(index_q[4]), .C(n27218), 
         .Z(n22126)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i19771_4_lut_3_lut.init = 16'h6565;
    LUT4 i8881_4_lut_4_lut (.A(index_q[3]), .B(index_q[0]), .C(index_q[1]), 
         .D(index_q[2]), .Z(n11325)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (D)+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i8881_4_lut_4_lut.init = 16'h0bf4;
    LUT4 i12143_2_lut_rep_547_2_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .Z(n27212)) /* synthesis lut_function=(A (B+!(C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12143_2_lut_rep_547_2_lut_3_lut.init = 16'h8f8f;
    LUT4 mux_229_Mux_8_i412_3_lut_4_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .Z(n15204)) /* synthesis lut_function=(A (B+!(C))+!A !((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_8_i412_3_lut_4_lut_3_lut.init = 16'h8e8e;
    LUT4 mux_230_Mux_1_i987_3_lut_4_lut_4_lut (.A(index_q[3]), .B(n986_adj_2713), 
         .C(index_q[4]), .D(n27238), .Z(n987)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_1_i987_3_lut_4_lut_4_lut.init = 16'hc5c0;
    LUT4 i9483_2_lut_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[3]), 
         .Z(n11969)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9483_2_lut_3_lut.init = 16'h8080;
    LUT4 i19963_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .D(index_i[3]), .Z(n22318)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(D))+!A (B+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19963_3_lut_4_lut_4_lut_4_lut.init = 16'h3380;
    L6MUX21 i23589 (.D0(n25265), .D1(n25263), .SD(index_i[6]), .Z(n25266));
    LUT4 i9677_3_lut_4_lut_4_lut_4_lut (.A(index_q[3]), .B(index_q[2]), 
         .C(index_q[1]), .D(index_q[0]), .Z(n12166)) /* synthesis lut_function=(!(A ((D)+!C)+!A !(B (C+!(D))+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i9677_3_lut_4_lut_4_lut_4_lut.init = 16'h51e5;
    LUT4 i11819_2_lut_rep_442_4_lut_4_lut_4_lut (.A(index_q[3]), .B(index_q[2]), 
         .C(index_q[1]), .D(index_q[0]), .Z(n27107)) /* synthesis lut_function=(!(A+(B (C)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i11819_2_lut_rep_442_4_lut_4_lut_4_lut.init = 16'h1404;
    LUT4 mux_230_Mux_2_i221_4_lut_4_lut (.A(index_q[3]), .B(index_q[4]), 
         .C(n27218), .D(n27104), .Z(n221_adj_2654)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (B+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_2_i221_4_lut_4_lut.init = 16'hf7c4;
    PFUMX i21104 (.BLUT(n23462), .ALUT(n23463), .C0(index_q[5]), .Z(n23478));
    LUT4 i9562_3_lut_3_lut (.A(index_q[3]), .B(index_q[4]), .C(n12047), 
         .Z(n12048)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i9562_3_lut_3_lut.init = 16'h7474;
    PFUMX i21105 (.BLUT(n23464), .ALUT(n23465), .C0(index_q[5]), .Z(n23479));
    LUT4 mux_229_Mux_9_i30_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .D(index_i[3]), .Z(n30_adj_2579)) /* synthesis lut_function=(A (B (C (D))+!B !(D))+!A !(B+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_9_i30_3_lut_4_lut_4_lut_4_lut.init = 16'h8033;
    LUT4 i19393_3_lut_4_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n21748)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19393_3_lut_4_lut_3_lut_4_lut.init = 16'hf80f;
    LUT4 i22961_2_lut_rep_636 (.A(index_i[1]), .B(index_i[2]), .Z(n27301)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i22961_2_lut_rep_636.init = 16'h9999;
    LUT4 n442_bdd_2_lut_24898_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[3]), 
         .Z(n26702)) /* synthesis lut_function=(A (B+(C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n442_bdd_2_lut_24898_3_lut.init = 16'hf9f9;
    LUT4 mux_229_Mux_4_i93_3_lut_4_lut_3_lut_rep_690_4_lut (.A(index_i[1]), 
         .B(index_i[2]), .C(index_i[3]), .D(index_i[0]), .Z(n27355)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_4_i93_3_lut_4_lut_3_lut_rep_690_4_lut.init = 16'h07f0;
    LUT4 mux_230_Mux_3_i747_3_lut (.A(n27274), .B(n404), .C(index_q[3]), 
         .Z(n747_adj_2296)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_3_i747_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_0_i93_3_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .Z(n93_adj_2578)) /* synthesis lut_function=(A (B)+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_0_i93_3_lut_3_lut.init = 16'h9c9c;
    LUT4 i11941_2_lut_rep_548_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[0]), 
         .Z(n27213)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11941_2_lut_rep_548_3_lut.init = 16'h8080;
    LUT4 i11478_2_lut_rep_459_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n27124)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11478_2_lut_rep_459_3_lut_4_lut.init = 16'hf8f0;
    LUT4 i19372_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n21727)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C (D)+!C !(D)))+!A !(B (D)+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19372_3_lut_4_lut_4_lut_4_lut.init = 16'h7c03;
    LUT4 mux_229_Mux_3_i142_3_lut_3_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .Z(n142_adj_2444)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_3_i142_3_lut_3_lut_3_lut.init = 16'h3838;
    LUT4 i19375_3_lut (.A(n27353), .B(n27348), .C(index_i[3]), .Z(n21730)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19375_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_1_i923_3_lut_3_lut_4_lut_3_lut_rep_717 (.A(index_i[1]), 
         .B(index_i[2]), .C(index_i[3]), .Z(n27382)) /* synthesis lut_function=(!(A (B (C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_1_i923_3_lut_3_lut_4_lut_3_lut_rep_717.init = 16'h7e7e;
    LUT4 mux_229_Mux_4_i491_3_lut_4_lut_4_lut (.A(index_i[2]), .B(n27435), 
         .C(index_i[3]), .D(n27429), .Z(n491_adj_2570)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_4_i491_3_lut_4_lut_4_lut.init = 16'hfc5c;
    LUT4 n890_bdd_3_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[3]), 
         .D(index_i[5]), .Z(n25626)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A (B (C (D))+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n890_bdd_3_lut_3_lut_4_lut.init = 16'h0f7e;
    LUT4 mux_229_Mux_4_i900_3_lut_4_lut_4_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .Z(n900_adj_2707)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_4_i900_3_lut_4_lut_4_lut_3_lut.init = 16'hd4d4;
    LUT4 mux_229_Mux_3_i349_3_lut_3_lut (.A(index_i[1]), .B(index_i[4]), 
         .C(n348_adj_2291), .Z(n349_adj_2781)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_3_i349_3_lut_3_lut.init = 16'hd1d1;
    LUT4 i22082_3_lut (.A(n21729), .B(n21730), .C(index_i[4]), .Z(n21731)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22082_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_5_i109_3_lut_4_lut_3_lut (.A(index_i[1]), .B(index_i[3]), 
         .C(index_i[0]), .Z(n109_adj_2541)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_5_i109_3_lut_4_lut_3_lut.init = 16'h6565;
    LUT4 i12145_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[4]), 
         .C(n27316), .D(index_i[0]), .Z(n14743)) /* synthesis lut_function=(!(A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12145_3_lut_4_lut_4_lut_4_lut.init = 16'h55d5;
    LUT4 i20095_3_lut_4_lut_3_lut (.A(index_i[1]), .B(index_i[3]), .C(index_i[2]), 
         .Z(n22450)) /* synthesis lut_function=(A (B)+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20095_3_lut_4_lut_3_lut.init = 16'hd9d9;
    PFUMX i21107 (.BLUT(n23468), .ALUT(n23469), .C0(index_q[5]), .Z(n23481));
    LUT4 mux_229_Mux_6_i660_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n660)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_6_i660_3_lut_3_lut.init = 16'hc6c6;
    LUT4 mux_229_Mux_1_i348_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n348_adj_2421)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A (B ((D)+!C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_1_i348_3_lut_4_lut_4_lut_4_lut.init = 16'h38f0;
    LUT4 i19956_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n22311)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C))+!A !(B ((D)+!C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19956_3_lut_4_lut_4_lut.init = 16'h925a;
    LUT4 n476_bdd_3_lut_25057_3_lut (.A(index_i[1]), .B(index_i[4]), .C(n124_adj_2542), 
         .Z(n25978)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n476_bdd_3_lut_25057_3_lut.init = 16'hd1d1;
    LUT4 mux_229_Mux_6_i498_3_lut_4_lut_4_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .Z(n498)) /* synthesis lut_function=(A (C)+!A !(B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_6_i498_3_lut_4_lut_4_lut_3_lut.init = 16'hb5b5;
    PFUMX i23587 (.BLUT(n924_adj_2782), .ALUT(n25264), .C0(index_i[5]), 
          .Z(n25265));
    LUT4 mux_229_Mux_5_i924_4_lut_3_lut (.A(index_i[2]), .B(n14081), .C(index_i[4]), 
         .Z(n924_adj_2782)) /* synthesis lut_function=(!(A (B+(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_5_i924_4_lut_3_lut.init = 16'h5656;
    LUT4 i11902_2_lut_rep_637 (.A(index_i[2]), .B(index_i[3]), .Z(n27302)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11902_2_lut_rep_637.init = 16'heeee;
    L6MUX21 i26016 (.D0(n28688), .D1(n28685), .SD(index_i[7]), .Z(n28689));
    LUT4 i11482_3_lut_3_lut_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[0]), 
         .Z(n652)) /* synthesis lut_function=(!(A ((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11482_3_lut_3_lut_3_lut.init = 16'h5d5d;
    PFUMX i26014 (.BLUT(n28687), .ALUT(n28686), .C0(index_i[5]), .Z(n28688));
    LUT4 i9447_3_lut_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), .C(index_i[1]), 
         .D(index_i[0]), .Z(n526_adj_2560)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9447_3_lut_3_lut_4_lut.init = 16'h1ef0;
    LUT4 i24257_then_3_lut (.A(index_i[0]), .B(index_i[4]), .C(index_i[3]), 
         .Z(n27559)) /* synthesis lut_function=(A (B)+!A (B (C)+!B !(C))) */ ;
    defparam i24257_then_3_lut.init = 16'hc9c9;
    LUT4 i22087_3_lut (.A(n21726), .B(n21727), .C(index_i[4]), .Z(n21728)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22087_3_lut.init = 16'hcaca;
    PFUMX i26012 (.BLUT(n23586), .ALUT(n28684), .C0(index_i[6]), .Z(n28685));
    LUT4 i12572_2_lut_rep_500_3_lut (.A(index_i[2]), .B(index_i[3]), .C(index_i[1]), 
         .Z(n27165)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12572_2_lut_rep_500_3_lut.init = 16'hfefe;
    L6MUX21 i21109 (.D0(n23472), .D1(n23473), .SD(index_q[5]), .Z(n23483));
    LUT4 i19368_3_lut (.A(n27256), .B(n27393), .C(index_i[3]), .Z(n21723)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19368_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_2_i731_3_lut_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n731_adj_2442)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(B (C)+!B !(C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_2_i731_3_lut_3_lut_4_lut.init = 16'h69f0;
    LUT4 index_q_4__bdd_3_lut_23545_4_lut (.A(n27219), .B(index_q[3]), .C(index_q[5]), 
         .D(index_q[4]), .Z(n25201)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam index_q_4__bdd_3_lut_23545_4_lut.init = 16'hf080;
    LUT4 i20719_3_lut (.A(n23088), .B(n25152), .C(index_q[7]), .Z(n23093)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20719_3_lut.init = 16'hcaca;
    LUT4 i20807_3_lut (.A(n26121), .B(n23172), .C(index_q[6]), .Z(n23181)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20807_3_lut.init = 16'hcaca;
    PFUMX i20586 (.BLUT(n158_adj_2474), .ALUT(n189_adj_2418), .C0(index_i[5]), 
          .Z(n22960));
    L6MUX21 i21110 (.D0(n23474), .D1(n23475), .SD(index_q[5]), .Z(n23484));
    LUT4 mux_229_Mux_6_i924_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[4]), .D(n908_adj_2549), .Z(n924_adj_2731)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_6_i924_3_lut_4_lut.init = 16'h6f60;
    L6MUX21 i21111 (.D0(n23476), .D1(n23477), .SD(index_q[5]), .Z(n23485));
    LUT4 i24257_else_3_lut (.A(index_i[2]), .B(index_i[0]), .C(index_i[4]), 
         .D(index_i[3]), .Z(n27558)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)+!C !(D)))+!A (B (C+!(D))+!B !(C)))) */ ;
    defparam i24257_else_3_lut.init = 16'h1e38;
    PFUMX i20816 (.BLUT(n12104), .ALUT(n62_adj_2783), .C0(index_q[5]), 
          .Z(n23190));
    LUT4 i20718_3_lut (.A(n23086), .B(n23087), .C(index_q[7]), .Z(n23092)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20718_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_5_i700_3_lut (.A(n460_adj_2529), .B(n27345), .C(index_i[4]), 
         .Z(n700_adj_2771)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_5_i700_3_lut.init = 16'hcaca;
    LUT4 i22936_3_lut (.A(n23092), .B(n23093), .C(index_q[8]), .Z(n23095)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22936_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_0_i236_3_lut_3_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[3]), .Z(n236)) /* synthesis lut_function=(A (B+(C))+!A !(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_0_i236_3_lut_3_lut.init = 16'ha9a9;
    LUT4 i22975_2_lut_rep_640 (.A(index_q[1]), .B(index_q[2]), .Z(n27305)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i22975_2_lut_rep_640.init = 16'h9999;
    PFUMX i20754 (.BLUT(n31_adj_2472), .ALUT(n62_adj_2784), .C0(index_q[5]), 
          .Z(n23128));
    LUT4 mux_230_Mux_0_i93_3_lut_3_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .Z(n93_adj_2372)) /* synthesis lut_function=(A (B)+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_0_i93_3_lut_3_lut.init = 16'h9c9c;
    LUT4 n442_bdd_2_lut_24408_3_lut (.A(index_q[1]), .B(index_q[2]), .C(index_q[3]), 
         .Z(n26127)) /* synthesis lut_function=(A (B+(C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam n442_bdd_2_lut_24408_3_lut.init = 16'hf9f9;
    PFUMX i20723 (.BLUT(n31_adj_2470), .ALUT(n62_adj_2468), .C0(index_q[5]), 
          .Z(n23097));
    PFUMX i20692 (.BLUT(n31_adj_2466), .ALUT(n22031), .C0(index_q[5]), 
          .Z(n23066));
    LUT4 i9683_3_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[4]), 
         .Z(n12172)) /* synthesis lut_function=(A (B)+!A !(B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9683_3_lut_4_lut_3_lut.init = 16'h9898;
    LUT4 n27296_bdd_3_lut_25595 (.A(n27218), .B(index_q[6]), .C(index_q[5]), 
         .Z(n27672)) /* synthesis lut_function=(!(A (B)+!A (C))) */ ;
    defparam n27296_bdd_3_lut_25595.init = 16'h2727;
    LUT4 i20011_3_lut_4_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n22366)) /* synthesis lut_function=(!(A (B (D)+!B !((D)+!C))+!A (B (C+(D))+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20011_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'h338f;
    LUT4 index_q_8__bdd_3_lut_then_4_lut (.A(index_q[4]), .B(index_q[6]), 
         .C(index_q[5]), .D(n27127), .Z(n27562)) /* synthesis lut_function=(!(A (B (C+(D)))+!A (B (C)))) */ ;
    defparam index_q_8__bdd_3_lut_then_4_lut.init = 16'h373f;
    PFUMX i23585 (.BLUT(n25262), .ALUT(n27162), .C0(index_i[5]), .Z(n25263));
    LUT4 i19401_3_lut (.A(n25225), .B(n21794), .C(index_i[8]), .Z(n21756)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19401_3_lut.init = 16'hcaca;
    LUT4 i19975_3_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[3]), .C(index_i[2]), 
         .D(index_i[0]), .Z(n22330)) /* synthesis lut_function=(A (B (D)+!B (C (D)+!C !(D)))+!A (B (D)+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19975_3_lut_4_lut_4_lut.init = 16'hfc13;
    PFUMX i20615 (.BLUT(n11978), .ALUT(n62_adj_2763), .C0(index_i[5]), 
          .Z(n22989));
    LUT4 i22174_3_lut (.A(n109), .B(n124_adj_2498), .C(index_i[4]), .Z(n22132)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22174_3_lut.init = 16'hcaca;
    PFUMX i20587 (.BLUT(n221_adj_2785), .ALUT(n22310), .C0(index_i[5]), 
          .Z(n22961));
    LUT4 i8920_4_lut_4_lut (.A(index_i[3]), .B(index_i[0]), .C(index_i[1]), 
         .D(index_i[2]), .Z(n11368)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (D)+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i8920_4_lut_4_lut.init = 16'h0bf4;
    LUT4 mux_229_Mux_2_i221_4_lut_4_lut (.A(index_i[3]), .B(index_i[4]), 
         .C(n27213), .D(n27108), .Z(n221_adj_2785)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (B+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_2_i221_4_lut_4_lut.init = 16'hf7c4;
    LUT4 n22303_bdd_3_lut_3_lut (.A(index_i[1]), .B(n526_adj_2560), .C(index_i[4]), 
         .Z(n25980)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n22303_bdd_3_lut_3_lut.init = 16'h5c5c;
    LUT4 i12399_2_lut_rep_564_3_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .Z(n27229)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12399_2_lut_rep_564_3_lut.init = 16'hf8f8;
    LUT4 index_q_8__bdd_3_lut_else_4_lut (.A(n27179), .B(index_q[4]), .C(index_q[6]), 
         .D(index_q[5]), .Z(n27561)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;
    defparam index_q_8__bdd_3_lut_else_4_lut.init = 16'hf080;
    LUT4 index_q_0__bdd_4_lut_25171 (.A(index_q[0]), .B(index_q[3]), .C(index_q[1]), 
         .D(index_q[2]), .Z(n27470)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C))+!A (B (C (D)+!C !(D))+!B !(C+!(D))))) */ ;
    defparam index_q_0__bdd_4_lut_25171.init = 16'h16d3;
    LUT4 mux_229_Mux_1_i573_3_lut_4_lut_4_lut (.A(index_i[3]), .B(n557), 
         .C(index_i[4]), .D(n27383), .Z(n573_adj_2786)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B ((D)+!C)+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_1_i573_3_lut_4_lut_4_lut.init = 16'h5c0c;
    CCU2D add_417_13 (.A0(quarter_wave_sample_register_i[12]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[13]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17899), .COUT(n17900), 
          .S0(o_val_pipeline_i_0__15__N_2176[12]), .S1(o_val_pipeline_i_0__15__N_2176[13]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam add_417_13.INIT0 = 16'hf555;
    defparam add_417_13.INIT1 = 16'hf555;
    defparam add_417_13.INJECT1_0 = "NO";
    defparam add_417_13.INJECT1_1 = "NO";
    LUT4 i11408_4_lut_4_lut (.A(index_i[3]), .B(index_i[2]), .C(index_i[0]), 
         .D(index_i[1]), .Z(n875_adj_2746)) /* synthesis lut_function=((B (C)+!B (D))+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11408_4_lut_4_lut.init = 16'hf7d5;
    LUT4 i19362_3_lut (.A(n356_adj_2398), .B(n27393), .C(index_i[3]), 
         .Z(n21717)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19362_3_lut.init = 16'hcaca;
    LUT4 i19864_4_lut_3_lut (.A(index_i[3]), .B(index_i[4]), .C(n27213), 
         .Z(n22219)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19864_4_lut_3_lut.init = 16'h6565;
    PFUMX i20553 (.BLUT(n31_adj_2461), .ALUT(n62_adj_2747), .C0(index_i[5]), 
          .Z(n22927));
    LUT4 mux_229_Mux_6_i730_3_lut_rep_718_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27383)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_6_i730_3_lut_rep_718_3_lut.init = 16'h3838;
    LUT4 mux_229_Mux_1_i987_3_lut_4_lut_4_lut (.A(index_i[3]), .B(n986_adj_2737), 
         .C(index_i[4]), .D(n27383), .Z(n987_adj_2787)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_1_i987_3_lut_4_lut_4_lut.init = 16'hc5c0;
    LUT4 i9643_3_lut_3_lut (.A(index_i[3]), .B(index_i[4]), .C(n12128), 
         .Z(n12129)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9643_3_lut_3_lut.init = 16'h7474;
    LUT4 i11654_2_lut_rep_642 (.A(index_q[2]), .B(index_q[3]), .Z(n27307)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i11654_2_lut_rep_642.init = 16'heeee;
    LUT4 n557_bdd_2_lut_24052_3_lut (.A(index_q[2]), .B(index_q[3]), .C(index_q[4]), 
         .Z(n25717)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam n557_bdd_2_lut_24052_3_lut.init = 16'he0e0;
    PFUMX i20522 (.BLUT(n31_adj_2458), .ALUT(n62_adj_2457), .C0(index_i[5]), 
          .Z(n22896));
    LUT4 i22182_3_lut (.A(n620_adj_2750), .B(n14372), .C(index_q[4]), 
         .Z(n22117)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22182_3_lut.init = 16'hcaca;
    LUT4 i19759_3_lut (.A(n27289), .B(n27299), .C(index_q[3]), .Z(n22114)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19759_3_lut.init = 16'hcaca;
    LUT4 n21642_bdd_3_lut_23998 (.A(n29950), .B(n29945), .C(index_q[3]), 
         .Z(n25709)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n21642_bdd_3_lut_23998.init = 16'hcaca;
    PFUMX i20491 (.BLUT(n31), .ALUT(n21707), .C0(index_i[5]), .Z(n22865));
    LUT4 i23095_2_lut_rep_482_3_lut_4_lut (.A(index_q[2]), .B(index_q[3]), 
         .C(index_q[1]), .D(index_q[0]), .Z(n27147)) /* synthesis lut_function=(!(A+(B+(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i23095_2_lut_rep_482_3_lut_4_lut.init = 16'h0111;
    LUT4 i11999_2_lut_rep_514_3_lut (.A(index_q[2]), .B(index_q[3]), .C(index_q[1]), 
         .Z(n27179)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i11999_2_lut_rep_514_3_lut.init = 16'hfefe;
    LUT4 i24206_then_4_lut (.A(index_i[0]), .B(index_i[4]), .C(index_i[1]), 
         .D(index_i[3]), .Z(n27566)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam i24206_then_4_lut.init = 16'h3c69;
    LUT4 i9571_3_lut_3_lut_4_lut (.A(index_q[2]), .B(index_q[3]), .C(index_q[1]), 
         .D(index_q[0]), .Z(n526_adj_2395)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i9571_3_lut_3_lut_4_lut.init = 16'h1ef0;
    PFUMX i20588 (.BLUT(n286_adj_2455), .ALUT(n317_adj_2452), .C0(index_i[5]), 
          .Z(n22962));
    LUT4 n526_bdd_2_lut_24009_3_lut_4_lut (.A(index_q[2]), .B(index_q[3]), 
         .C(index_q[4]), .D(index_q[1]), .Z(n25714)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam n526_bdd_2_lut_24009_3_lut_4_lut.init = 16'h0f1f;
    LUT4 i22358_3_lut (.A(n22113), .B(n22114), .C(index_q[4]), .Z(n22115)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22358_3_lut.init = 16'hcaca;
    PFUMX i24497 (.BLUT(n26220), .ALUT(n26219), .C0(index_q[5]), .Z(n26221));
    PFUMX i20589 (.BLUT(n349_adj_2754), .ALUT(n22313), .C0(index_i[5]), 
          .Z(n22963));
    CCU2D add_417_11 (.A0(quarter_wave_sample_register_i[10]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[11]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17898), .COUT(n17899), 
          .S0(o_val_pipeline_i_0__15__N_2176[10]), .S1(o_val_pipeline_i_0__15__N_2176[11]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam add_417_11.INIT0 = 16'hf555;
    defparam add_417_11.INIT1 = 16'hf555;
    defparam add_417_11.INJECT1_0 = "NO";
    defparam add_417_11.INJECT1_1 = "NO";
    LUT4 mux_229_Mux_6_i204_3_lut_4_lut_3_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .Z(n204)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_6_i204_3_lut_4_lut_3_lut_3_lut.init = 16'h3d3d;
    LUT4 i9612_3_lut_4_lut_3_lut_4_lut (.A(index_q[2]), .B(index_q[3]), 
         .C(index_q[1]), .D(index_q[0]), .Z(n844_adj_2283)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i9612_3_lut_4_lut_3_lut_4_lut.init = 16'hf00e;
    LUT4 mux_230_Mux_2_i955_then_4_lut (.A(index_q[4]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n27472)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B (C+!(D))+!B !(C (D)))) */ ;
    defparam mux_230_Mux_2_i955_then_4_lut.init = 16'he95d;
    PFUMX i20590 (.BLUT(n413_adj_2450), .ALUT(n22319), .C0(index_i[5]), 
          .Z(n22964));
    LUT4 i24206_else_4_lut (.A(index_i[0]), .B(index_i[4]), .C(index_i[1]), 
         .D(index_i[3]), .Z(n27565)) /* synthesis lut_function=(!(A (B (C)+!B !(C (D)+!C !(D)))+!A (B ((D)+!C)+!B !((D)+!C)))) */ ;
    defparam i24206_else_4_lut.init = 16'h394b;
    PFUMX i20591 (.BLUT(n22322), .ALUT(n507_adj_2755), .C0(index_i[5]), 
          .Z(n22965));
    LUT4 mux_229_Mux_8_i860_3_lut_4_lut (.A(n27214), .B(index_i[3]), .C(index_i[4]), 
         .D(n27159), .Z(n860_adj_2597)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_8_i860_3_lut_4_lut.init = 16'h08f8;
    PFUMX i20592 (.BLUT(n22328), .ALUT(n573), .C0(index_i[5]), .Z(n22966));
    LUT4 mux_230_Mux_2_i955_else_4_lut (.A(index_q[4]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n27471)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+(D)))+!A !(B (C+!(D))+!B !(C+!(D))))) */ ;
    defparam mux_230_Mux_2_i955_else_4_lut.init = 16'h49c6;
    PFUMX i20593 (.BLUT(n605_adj_2446), .ALUT(n22331), .C0(index_i[5]), 
          .Z(n22967));
    LUT4 i11550_2_lut_rep_583 (.A(index_i[0]), .B(index_i[1]), .Z(n27248)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11550_2_lut_rep_583.init = 16'h2222;
    PFUMX i20594 (.BLUT(n669), .ALUT(n700_adj_2448), .C0(index_i[5]), 
          .Z(n22968));
    LUT4 mux_229_Mux_6_i636_4_lut_4_lut (.A(index_i[1]), .B(index_i[4]), 
         .C(n635_adj_2318), .D(n14744), .Z(n636_adj_2765)) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_6_i636_4_lut_4_lut.init = 16'hf3d1;
    LUT4 i11473_2_lut_2_lut_3_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .Z(n14070)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11473_2_lut_2_lut_3_lut.init = 16'h0808;
    PFUMX i20595 (.BLUT(n732_adj_2443), .ALUT(n763_adj_2758), .C0(index_i[5]), 
          .Z(n22969));
    LUT4 n22923_bdd_3_lut (.A(n22916), .B(n22917), .C(index_i[7]), .Z(n25006)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n22923_bdd_3_lut.init = 16'hcaca;
    LUT4 i15920_3_lut (.A(n27271), .B(n29949), .C(index_q[3]), .Z(n18106)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15920_3_lut.init = 16'hcaca;
    LUT4 i11551_2_lut_rep_719 (.A(index_i[1]), .B(index_i[0]), .Z(n27384)) /* synthesis lut_function=((B)+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11551_2_lut_rep_719.init = 16'hdddd;
    LUT4 mux_229_Mux_5_i867_3_lut_4_lut_3_lut_rep_720 (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .Z(n27385)) /* synthesis lut_function=(!(A ((C)+!B)+!A !((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_5_i867_3_lut_4_lut_3_lut_rep_720.init = 16'h5959;
    L6MUX21 i20597 (.D0(n860_adj_2699), .D1(n891_adj_2695), .SD(index_i[5]), 
            .Z(n22971));
    LUT4 mux_229_Mux_5_i347_3_lut_4_lut_4_lut_3_lut_rep_722 (.A(index_i[1]), 
         .B(index_i[2]), .C(index_i[0]), .Z(n27387)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_5_i347_3_lut_4_lut_4_lut_3_lut_rep_722.init = 16'hd6d6;
    LUT4 i12190_3_lut_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n14788)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (D))+!A (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12190_3_lut_3_lut_3_lut_4_lut.init = 16'h00f7;
    LUT4 i11487_3_lut_3_lut_3_lut_rep_723 (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .Z(n27388)) /* synthesis lut_function=(!(A+!(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11487_3_lut_3_lut_3_lut_rep_723.init = 16'h4545;
    LUT4 mux_229_Mux_5_i300_3_lut_4_lut_3_lut_rep_724 (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .Z(n27389)) /* synthesis lut_function=(A (B (C))+!A !(B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_5_i300_3_lut_4_lut_3_lut_rep_724.init = 16'h9595;
    LUT4 i15919_3_lut (.A(n29949), .B(n29953), .C(index_q[3]), .Z(n18105)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15919_3_lut.init = 16'hcaca;
    LUT4 i21148_3_lut (.A(n23519), .B(n23520), .C(index_i[7]), .Z(n23522)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21148_3_lut.init = 16'hcaca;
    PFUMX i23330 (.BLUT(n24928), .ALUT(n23124), .C0(index_q[8]), .Z(n24929));
    LUT4 mux_229_Mux_2_i269_3_lut_4_lut_3_lut_rep_727 (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .Z(n27392)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_2_i269_3_lut_4_lut_3_lut_rep_727.init = 16'h6565;
    LUT4 mux_229_Mux_6_i420_3_lut_4_lut_4_lut_3_lut_rep_728 (.A(index_i[1]), 
         .B(index_i[2]), .C(index_i[0]), .Z(n27393)) /* synthesis lut_function=(A (B+(C))+!A !(B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_6_i420_3_lut_4_lut_4_lut_3_lut_rep_728.init = 16'hbdbd;
    LUT4 i21147_3_lut (.A(n23517), .B(n23518), .C(index_i[7]), .Z(n23521)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21147_3_lut.init = 16'hcaca;
    PFUMX i21135 (.BLUT(n23493), .ALUT(n23494), .C0(index_i[5]), .Z(n23509));
    LUT4 mux_229_Mux_5_i459_3_lut_4_lut_4_lut_3_lut_rep_729 (.A(index_i[1]), 
         .B(index_i[2]), .C(index_i[0]), .Z(n27394)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_5_i459_3_lut_4_lut_4_lut_3_lut_rep_729.init = 16'h7979;
    LUT4 i21117_3_lut (.A(n23488), .B(n23489), .C(index_q[7]), .Z(n23491)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21117_3_lut.init = 16'hcaca;
    LUT4 i21116_3_lut (.A(n23486), .B(n23487), .C(index_q[7]), .Z(n23490)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21116_3_lut.init = 16'hcaca;
    PFUMX i21136 (.BLUT(n23495), .ALUT(n23496), .C0(index_i[5]), .Z(n23510));
    LUT4 mux_229_Mux_5_i460_3_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .D(index_i[3]), .Z(n460_adj_2529)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B (C (D)+!C !(D))+!B (C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_5_i460_3_lut_4_lut_4_lut.init = 16'h793c;
    LUT4 i22184_3_lut (.A(n491_adj_2769), .B(n506_adj_2788), .C(index_q[4]), 
         .Z(n22111)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22184_3_lut.init = 16'hcaca;
    L6MUX21 i21137 (.D0(n23497), .D1(n23498), .SD(index_i[5]), .Z(n23511));
    PFUMX i21138 (.BLUT(n23499), .ALUT(n23500), .C0(index_i[5]), .Z(n23512));
    LUT4 i19686_3_lut (.A(n356), .B(n29938), .C(index_q[3]), .Z(n22041)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19686_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_0_i364_3_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .D(index_i[3]), .Z(n364_adj_2721)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !(B (C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_0_i364_3_lut_3_lut_4_lut.init = 16'hbd0f;
    LUT4 mux_229_Mux_7_i620_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n620_adj_2770)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A !(B (C+!(D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_7_i620_3_lut_4_lut_4_lut_4_lut.init = 16'h8c33;
    LUT4 n557_bdd_3_lut_24051_4_lut (.A(n27219), .B(index_q[3]), .C(index_q[4]), 
         .D(n27166), .Z(n25716)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam n557_bdd_3_lut_24051_4_lut.init = 16'hf707;
    LUT4 i19972_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[0]), 
         .D(index_i[3]), .Z(n22327)) /* synthesis lut_function=(A (B+(C+(D)))+!A !(B (C+(D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19972_3_lut_4_lut.init = 16'haabd;
    L6MUX21 i21140 (.D0(n23503), .D1(n23504), .SD(index_i[5]), .Z(n23514));
    LUT4 i9663_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .D(index_i[3]), .Z(n12152)) /* synthesis lut_function=(!(A (B (C (D))+!B (C (D)+!C !(D)))+!A (B (C+(D))+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9663_3_lut_4_lut_4_lut_4_lut.init = 16'h0abd;
    LUT4 i22361_3_lut (.A(n22107), .B(n22108), .C(index_q[4]), .Z(n22109)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22361_3_lut.init = 16'hcaca;
    LUT4 i20549_3_lut (.A(n22918), .B(n22919), .C(index_i[7]), .Z(n22923)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20549_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_6_i483_3_lut_3_lut_rep_798 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29925)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_6_i483_3_lut_3_lut_rep_798.init = 16'h6c6c;
    LUT4 i9662_3_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[4]), 
         .Z(n12151)) /* synthesis lut_function=(!(A (B)+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9662_3_lut_4_lut_3_lut.init = 16'h6262;
    L6MUX21 i21141 (.D0(n23505), .D1(n23506), .SD(index_i[5]), .Z(n23515));
    LUT4 mux_229_Mux_2_i604_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .D(index_i[3]), .Z(n604_adj_2445)) /* synthesis lut_function=(!(A (B (D)+!B !(C+!(D)))+!A !(B (D)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_2_i604_3_lut_4_lut_4_lut_4_lut.init = 16'h65bb;
    L6MUX21 i21142 (.D0(n23507), .D1(n23508), .SD(index_i[5]), .Z(n23516));
    LUT4 mux_230_Mux_2_i507_3_lut_3_lut (.A(index_q[0]), .B(index_q[4]), 
         .C(n491_adj_2760), .Z(n507_adj_2663)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_2_i507_3_lut_3_lut.init = 16'h7474;
    LUT4 mux_229_Mux_2_i890_3_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .D(index_i[3]), .Z(n890_adj_2694)) /* synthesis lut_function=(A (B (C (D))+!B (C (D)+!C !(D)))+!A !(B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_2_i890_3_lut_4_lut_4_lut.init = 16'ha546;
    LUT4 mux_230_Mux_2_i349_3_lut_3_lut (.A(index_q[0]), .B(index_q[4]), 
         .C(n348_adj_2573), .Z(n349_adj_2658)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_2_i349_3_lut_3_lut.init = 16'hd1d1;
    LUT4 mux_230_Mux_2_i763_4_lut_4_lut (.A(index_q[0]), .B(n12095), .C(index_q[4]), 
         .D(n157_adj_2516), .Z(n763_adj_2669)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_2_i763_4_lut_4_lut.init = 16'hdfd0;
    LUT4 i19374_3_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[0]), 
         .D(index_i[3]), .Z(n21729)) /* synthesis lut_function=(A (B (C (D))+!B !(C (D)+!C !(D)))+!A (B (C)+!B !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19374_3_lut_4_lut_4_lut.init = 16'hc371;
    LUT4 i19356_3_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[0]), 
         .D(index_i[3]), .Z(n21711)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C+(D)))+!A !(B (C (D)+!C !(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19356_3_lut_4_lut_4_lut.init = 16'h955a;
    LUT4 i20037_3_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[0]), 
         .D(index_i[3]), .Z(n22392)) /* synthesis lut_function=(A (B (C)+!B !(C+!(D)))+!A (B (C (D)+!C !(D))+!B !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20037_3_lut_4_lut_4_lut.init = 16'hc395;
    LUT4 mux_229_Mux_2_i908_3_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .D(index_i[3]), .Z(n908_adj_2704)) /* synthesis lut_function=(!(A (B+!(D))+!A !(B+!(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_2_i908_3_lut_4_lut_4_lut.init = 16'h6645;
    LUT4 mux_229_Mux_6_i860_3_lut_3_lut (.A(n27096), .B(index_i[4]), .C(n844_adj_2556), 
         .Z(n860_adj_2766)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam mux_229_Mux_6_i860_3_lut_3_lut.init = 16'h7474;
    LUT4 i19360_3_lut (.A(n29913), .B(n27387), .C(index_i[3]), .Z(n21715)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19360_3_lut.init = 16'hcaca;
    PFUMX i24472 (.BLUT(n26195), .ALUT(n29956), .C0(index_i[3]), .Z(n26196));
    LUT4 i20028_3_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[0]), 
         .D(index_i[3]), .Z(n22383)) /* synthesis lut_function=(!(A ((D)+!B)+!A !(B (D)+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20028_3_lut_4_lut_4_lut.init = 16'h4588;
    LUT4 mux_229_Mux_1_i301_3_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .D(index_i[3]), .Z(n301)) /* synthesis lut_function=(A (B (C)+!B (C (D)+!C !(D)))+!A !(B (C (D))+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_1_i301_3_lut_4_lut_4_lut.init = 16'ha5d6;
    LUT4 i19359_3_lut (.A(n27342), .B(n29923), .C(index_i[3]), .Z(n21714)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19359_3_lut.init = 16'hcaca;
    LUT4 i9684_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[0]), 
         .D(index_i[3]), .Z(n12173)) /* synthesis lut_function=(!(A (B (C (D))+!B (D))+!A !(B (C (D))+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9684_3_lut_4_lut.init = 16'h59aa;
    L6MUX21 i23559 (.D0(n25224), .D1(n27060), .SD(index_i[6]), .Z(n25225));
    LUT4 mux_230_Mux_5_i573_3_lut_3_lut (.A(index_q[0]), .B(index_q[4]), 
         .C(n572_adj_2789), .Z(n573_adj_2586)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_5_i573_3_lut_3_lut.init = 16'hd1d1;
    CCU2D add_417_9 (.A0(quarter_wave_sample_register_i[8]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[9]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17897), .COUT(n17898), 
          .S0(o_val_pipeline_i_0__15__N_2176[8]), .S1(o_val_pipeline_i_0__15__N_2176[9]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam add_417_9.INIT0 = 16'hf555;
    defparam add_417_9.INIT1 = 16'hf555;
    defparam add_417_9.INJECT1_0 = "NO";
    defparam add_417_9.INJECT1_1 = "NO";
    LUT4 index_i_5__bdd_4_lut_24846_4_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n26453)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B (C)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam index_i_5__bdd_4_lut_24846_4_lut_4_lut.init = 16'h3d2d;
    LUT4 i21444_3_lut (.A(n23815), .B(n23816), .C(index_q[7]), .Z(n23818)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21444_3_lut.init = 16'hcaca;
    LUT4 i20029_3_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[0]), 
         .D(index_i[3]), .Z(n22384)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A (B (C)+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20029_3_lut_4_lut_4_lut.init = 16'h3c9d;
    LUT4 mux_230_Mux_4_i221_3_lut_3_lut (.A(index_q[0]), .B(index_q[4]), 
         .C(n205_adj_2733), .Z(n221_adj_2604)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_4_i221_3_lut_3_lut.init = 16'h7474;
    LUT4 i23458_then_4_lut (.A(index_q[0]), .B(index_q[4]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n27569)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)+!C !(D))+!B (C (D)))) */ ;
    defparam i23458_then_4_lut.init = 16'hda0e;
    LUT4 i21443_3_lut (.A(n23813), .B(n23814), .C(index_q[7]), .Z(n23817)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21443_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_4_i142_3_lut_4_lut_3_lut (.A(index_q[0]), .B(index_q[3]), 
         .C(index_q[2]), .Z(n142_adj_2373)) /* synthesis lut_function=(A (B (C))+!A !(B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_4_i142_3_lut_4_lut_3_lut.init = 16'h9595;
    LUT4 mux_230_Mux_0_i985_3_lut_4_lut_3_lut (.A(index_q[0]), .B(index_q[2]), 
         .C(index_q[1]), .Z(n985_adj_2277)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_0_i985_3_lut_4_lut_3_lut.init = 16'h1919;
    LUT4 mux_230_Mux_1_i890_4_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[4]), 
         .C(n14_adj_2290), .D(index_q[3]), .Z(n890_adj_2749)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A !(B+(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_1_i890_4_lut_4_lut_4_lut_4_lut.init = 16'h7477;
    PFUMX i23557 (.BLUT(n27070), .ALUT(n27085), .C0(index_i[7]), .Z(n25224));
    PFUMX i20616 (.BLUT(n94), .ALUT(n22340), .C0(index_i[5]), .Z(n22990));
    LUT4 mux_230_Mux_5_i564_3_lut_4_lut_3_lut_rep_646 (.A(index_q[0]), .B(index_q[2]), 
         .C(index_q[1]), .Z(n27311)) /* synthesis lut_function=(A (B (C))+!A !(B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_5_i564_3_lut_4_lut_3_lut_rep_646.init = 16'h9595;
    LUT4 mux_230_Mux_5_i572_3_lut_4_lut (.A(index_q[0]), .B(index_q[2]), 
         .C(index_q[1]), .D(index_q[3]), .Z(n572_adj_2789)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A !(B (C+(D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_5_i572_3_lut_4_lut.init = 16'haa95;
    LUT4 mux_230_Mux_1_i93_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[2]), 
         .C(index_q[1]), .D(index_q[3]), .Z(n93_adj_2664)) /* synthesis lut_function=(A (B (C (D))+!B !(D))+!A !(B (C (D))+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_1_i93_3_lut_4_lut_4_lut.init = 16'h9566;
    LUT4 mux_230_Mux_4_i252_4_lut_4_lut (.A(index_q[0]), .B(index_q[3]), 
         .C(n27334), .D(index_q[4]), .Z(n252_adj_2605)) /* synthesis lut_function=(!(A (B (D)+!B !(D))+!A !(B ((D)+!C)+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_4_i252_4_lut_4_lut.init = 16'h669d;
    L6MUX21 i20617 (.D0(n22346), .D1(n22349), .SD(index_i[5]), .Z(n22991));
    LUT4 mux_230_Mux_3_i444_3_lut_4_lut (.A(index_q[0]), .B(index_q[3]), 
         .C(n27371), .D(index_q[4]), .Z(n444_adj_2637)) /* synthesis lut_function=(!(A (B (D)+!B (C (D)))+!A !(B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_3_i444_3_lut_4_lut.init = 16'h46aa;
    LUT4 i19857_3_lut_4_lut (.A(index_q[0]), .B(index_q[2]), .C(index_q[1]), 
         .D(index_q[3]), .Z(n22212)) /* synthesis lut_function=(A (B (D)+!B (C+(D)))+!A !(B (D)+!B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i19857_3_lut_4_lut.init = 16'haa65;
    PFUMX i20619 (.BLUT(n22355), .ALUT(n317_adj_2705), .C0(index_i[5]), 
          .Z(n22993));
    LUT4 mux_230_Mux_1_i62_3_lut_4_lut (.A(index_q[0]), .B(index_q[3]), 
         .C(index_q[2]), .D(index_q[4]), .Z(n62_adj_2783)) /* synthesis lut_function=(A (B (D)+!B ((D)+!C))+!A !(B (D)+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_1_i62_3_lut_4_lut.init = 16'haa56;
    PFUMX i20620 (.BLUT(n349_adj_2422), .ALUT(n22358), .C0(index_i[5]), 
          .Z(n22994));
    LUT4 i19744_3_lut (.A(n356), .B(n29919), .C(index_q[3]), .Z(n22099)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19744_3_lut.init = 16'hcaca;
    L6MUX21 i20621 (.D0(n22364), .D1(n22367), .SD(index_i[5]), .Z(n22995));
    L6MUX21 i20622 (.D0(n22373), .D1(n22376), .SD(index_i[5]), .Z(n22996));
    PFUMX i20623 (.BLUT(n22382), .ALUT(n573_adj_2786), .C0(index_i[5]), 
          .Z(n22997));
    LUT4 i21181_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n23555)) /* synthesis lut_function=(A (B (C)+!B !(C (D)+!C !(D)))+!A !(B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21181_3_lut_4_lut_4_lut_4_lut.init = 16'h83f0;
    LUT4 i22370_3_lut (.A(n22098), .B(n22099), .C(index_q[4]), .Z(n22100)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22370_3_lut.init = 16'hcaca;
    LUT4 i19753_3_lut_4_lut_4_lut (.A(index_q[2]), .B(n308), .C(index_q[3]), 
         .D(n27296), .Z(n22108)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i19753_3_lut_4_lut_4_lut.init = 16'hc5c0;
    L6MUX21 i24450 (.D0(n26174), .D1(n26171), .SD(index_q[5]), .Z(n26175));
    LUT4 i20485_3_lut (.A(n22852), .B(n22853), .C(index_i[7]), .Z(n22859)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20485_3_lut.init = 16'hcaca;
    PFUMX i24448 (.BLUT(n26173), .ALUT(n26172), .C0(index_q[4]), .Z(n26174));
    L6MUX21 i20624 (.D0(n22385), .D1(n636_adj_2662), .SD(index_i[5]), 
            .Z(n22998));
    L6MUX21 i21166 (.D0(n23524), .D1(n23525), .SD(index_i[5]), .Z(n23540));
    PFUMX i20625 (.BLUT(n22391), .ALUT(n700), .C0(index_i[5]), .Z(n22999));
    LUT4 i23458_else_4_lut (.A(index_q[0]), .B(index_q[4]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n27568)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C))+!A (B (C)+!B (C+(D)))) */ ;
    defparam i23458_else_4_lut.init = 16'hf178;
    LUT4 mux_230_Mux_7_i506_3_lut_4_lut_4_lut (.A(index_q[2]), .B(n29934), 
         .C(index_q[3]), .D(n27296), .Z(n506_adj_2788)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B ((D)+!C)+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_7_i506_3_lut_4_lut_4_lut.init = 16'h5c0c;
    L6MUX21 i20627 (.D0(n22394), .D1(n22400), .SD(index_i[5]), .Z(n23001));
    L6MUX21 i21167 (.D0(n23526), .D1(n23527), .SD(index_i[5]), .Z(n23541));
    L6MUX21 i21168 (.D0(n23528), .D1(n23529), .SD(index_i[5]), .Z(n23542));
    LUT4 i19357_3_lut (.A(n27358), .B(n29923), .C(index_i[3]), .Z(n21712)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19357_3_lut.init = 16'hcaca;
    L6MUX21 i21169 (.D0(n23530), .D1(n23531), .SD(index_i[5]), .Z(n23543));
    LUT4 mux_229_Mux_5_i781_3_lut_4_lut_4_lut_then_4_lut (.A(index_i[3]), 
         .B(index_i[0]), .C(index_i[4]), .D(index_i[2]), .Z(n27475)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_5_i781_3_lut_4_lut_4_lut_then_4_lut.init = 16'hece0;
    L6MUX21 i21170 (.D0(n23532), .D1(n23533), .SD(index_i[5]), .Z(n23544));
    LUT4 i20484_3_lut (.A(n22850), .B(n22851), .C(index_i[7]), .Z(n22858)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20484_3_lut.init = 16'hcaca;
    PFUMX i20629 (.BLUT(n924), .ALUT(n22448), .C0(index_i[5]), .Z(n23003));
    LUT4 i20489_3_lut (.A(n22860), .B(n22861), .C(index_i[8]), .Z(n22863)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20489_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_8_i526_3_lut_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n526_adj_2366)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_8_i526_3_lut_3_lut_3_lut_4_lut.init = 16'h0f70;
    LUT4 n300_bdd_3_lut_24390_4_lut_4_lut (.A(index_q[2]), .B(n619), .C(index_q[3]), 
         .D(n27296), .Z(n26118)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B ((D)+!C)+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam n300_bdd_3_lut_24390_4_lut_4_lut.init = 16'h5c0c;
    PFUMX i24445 (.BLUT(n26170), .ALUT(n27107), .C0(index_q[4]), .Z(n26171));
    LUT4 i19741_3_lut (.A(n29947), .B(n27280), .C(index_q[3]), .Z(n22096)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19741_3_lut.init = 16'hcaca;
    PFUMX i20630 (.BLUT(n987_adj_2787), .ALUT(n22451), .C0(index_i[5]), 
          .Z(n23004));
    LUT4 i20472_3_lut (.A(n22841), .B(n22842), .C(index_i[7]), .Z(n22846)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20472_3_lut.init = 16'hcaca;
    LUT4 i23148_2_lut_rep_490_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n27155)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i23148_2_lut_rep_490_3_lut_4_lut.init = 16'h0007;
    LUT4 i20464_3_lut (.A(n22825), .B(n25836), .C(index_i[6]), .Z(n22838)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20464_3_lut.init = 16'hcaca;
    LUT4 i20463_3_lut (.A(n25829), .B(n22824), .C(index_i[6]), .Z(n22837)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20463_3_lut.init = 16'hcaca;
    L6MUX21 i21171 (.D0(n23534), .D1(n23535), .SD(index_i[5]), .Z(n23545));
    LUT4 mux_230_Mux_6_i573_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[4]), .D(n572_adj_2767), .Z(n573_adj_2723)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_6_i573_3_lut_4_lut.init = 16'hf909;
    L6MUX21 i24443 (.D0(n26168), .D1(n26166), .SD(index_q[4]), .Z(n26169));
    PFUMX i24441 (.BLUT(n27104), .ALUT(n26167), .C0(index_q[5]), .Z(n26168));
    L6MUX21 i21172 (.D0(n23536), .D1(n23537), .SD(index_i[5]), .Z(n23546));
    L6MUX21 i21173 (.D0(n23538), .D1(n23539), .SD(index_i[5]), .Z(n23547));
    L6MUX21 i23543 (.D0(n25202), .D1(n27062), .SD(index_q[6]), .Z(n25203));
    LUT4 mux_229_Mux_7_i747_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n747_adj_2548)) /* synthesis lut_function=(A (B (C)+!B (C (D)+!C !(D)))+!A (B (C+!(D))+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_7_i747_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hf0c7;
    PFUMX i24439 (.BLUT(n26165), .ALUT(n26164), .C0(index_q[5]), .Z(n26166));
    PFUMX i23541 (.BLUT(n25201), .ALUT(n27084), .C0(index_q[7]), .Z(n25202));
    LUT4 i11774_3_lut_3_lut_4_lut_4_lut (.A(index_q[2]), .B(index_q[3]), 
         .C(index_q[1]), .D(index_q[0]), .Z(n14372)) /* synthesis lut_function=(!(A+!(B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i11774_3_lut_3_lut_4_lut_4_lut.init = 16'h4555;
    LUT4 mux_230_Mux_4_i491_3_lut_4_lut_4_lut (.A(index_q[2]), .B(n29934), 
         .C(index_q[3]), .D(n27293), .Z(n491_adj_2739)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_4_i491_3_lut_4_lut_4_lut.init = 16'hfc5c;
    LUT4 n22912_bdd_3_lut (.A(n22912), .B(n22913), .C(index_i[7]), .Z(n25009)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n22912_bdd_3_lut.init = 16'hcaca;
    LUT4 i22375_3_lut (.A(n22092), .B(n22093), .C(index_q[4]), .Z(n22094)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22375_3_lut.init = 16'hcaca;
    LUT4 i11391_2_lut_rep_443_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n27108)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11391_2_lut_rep_443_3_lut_4_lut.init = 16'hf080;
    LUT4 i20461_3_lut (.A(n25819), .B(n22820), .C(index_i[6]), .Z(n22835)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20461_3_lut.init = 16'hcaca;
    LUT4 index_q_5__bdd_3_lut_25454 (.A(index_q[5]), .B(n27670), .C(index_q[3]), 
         .Z(n27671)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam index_q_5__bdd_3_lut_25454.init = 16'hcaca;
    L6MUX21 i24406 (.D0(n26131), .D1(n26129), .SD(index_q[5]), .Z(n26132));
    PFUMX i24404 (.BLUT(n572_adj_2789), .ALUT(n26130), .C0(index_q[4]), 
          .Z(n26131));
    LUT4 i11790_3_lut_3_lut_4_lut_4_lut (.A(index_q[2]), .B(index_q[3]), 
         .C(index_q[1]), .D(index_q[0]), .Z(n14388)) /* synthesis lut_function=(!(A ((C+(D))+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i11790_3_lut_3_lut_4_lut_4_lut.init = 16'h555d;
    LUT4 mux_230_Mux_5_i924_4_lut_3_lut (.A(index_q[2]), .B(n15103), .C(index_q[4]), 
         .Z(n924_adj_2790)) /* synthesis lut_function=(!(A (B+(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_5_i924_4_lut_3_lut.init = 16'h5656;
    LUT4 i19684_3_lut (.A(n29949), .B(n27280), .C(index_q[3]), .Z(n22039)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19684_3_lut.init = 16'hcaca;
    CCU2D add_417_7 (.A0(quarter_wave_sample_register_i[6]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[7]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17896), .COUT(n17897), 
          .S1(o_val_pipeline_i_0__15__N_2176[7]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam add_417_7.INIT0 = 16'hf555;
    defparam add_417_7.INIT1 = 16'hf555;
    defparam add_417_7.INJECT1_0 = "NO";
    defparam add_417_7.INJECT1_1 = "NO";
    LUT4 index_i_6__bdd_4_lut_24140_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[6]), .D(n27302), .Z(n25795)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)+!C !(D)))+!A (B (C (D))+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam index_i_6__bdd_4_lut_24140_4_lut_4_lut.init = 16'h0f7c;
    LUT4 index_i_8__bdd_3_lut_23364_then_4_lut (.A(index_i[4]), .B(index_i[6]), 
         .C(index_i[5]), .D(n27131), .Z(n27575)) /* synthesis lut_function=(!(A (B (C+(D)))+!A (B (C)))) */ ;
    defparam index_i_8__bdd_3_lut_23364_then_4_lut.init = 16'h373f;
    LUT4 index_i_8__bdd_3_lut_23364_else_4_lut (.A(n27165), .B(index_i[4]), 
         .C(index_i[6]), .D(index_i[5]), .Z(n27574)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;
    defparam index_i_8__bdd_3_lut_23364_else_4_lut.init = 16'hf080;
    PFUMX i24401 (.BLUT(n26128), .ALUT(n26127), .C0(index_q[4]), .Z(n26129));
    LUT4 mux_229_Mux_5_i781_3_lut_4_lut_4_lut_else_4_lut (.A(index_i[3]), 
         .B(index_i[0]), .C(index_i[4]), .Z(n27474)) /* synthesis lut_function=(!(A (C)+!A (B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_5_i781_3_lut_4_lut_4_lut_else_4_lut.init = 16'h1f1f;
    LUT4 i19732_3_lut (.A(n29938), .B(n29955), .C(index_q[3]), .Z(n22087)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19732_3_lut.init = 16'hcaca;
    LUT4 i19911_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n22266)) /* synthesis lut_function=(!(A (B (D)+!B !(D))+!A (B ((D)+!C)+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19911_3_lut_4_lut_4_lut_4_lut.init = 16'h33c8;
    LUT4 mux_229_Mux_3_i262_rep_765 (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .Z(n27430)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_3_i262_rep_765.init = 16'h7c7c;
    LUT4 i19596_3_lut_else_4_lut (.A(index_q[4]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n29961)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C+!(D)))+!A !(B ((D)+!C)+!B (C (D)+!C !(D))))) */ ;
    defparam i19596_3_lut_else_4_lut.init = 16'h5685;
    LUT4 i11844_2_lut_3_lut_4_lut (.A(index_q[2]), .B(index_q[3]), .C(index_q[1]), 
         .D(index_q[0]), .Z(n844)) /* synthesis lut_function=(A ((C (D)+!C !(D))+!B)+!A (B+(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i11844_2_lut_3_lut_4_lut.init = 16'hf66f;
    LUT4 mux_230_Mux_2_i731_3_lut_3_lut_4_lut (.A(index_q[2]), .B(index_q[3]), 
         .C(index_q[1]), .D(index_q[0]), .Z(n731_adj_2670)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(B (C)+!B !(C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_2_i731_3_lut_3_lut_4_lut.init = 16'h69f0;
    LUT4 i19683_3_lut (.A(n29919), .B(n27277), .C(index_q[3]), .Z(n22038)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19683_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_0_i747_3_lut_4_lut_3_lut_4_lut (.A(index_q[2]), .B(index_q[3]), 
         .C(index_q[1]), .D(index_q[0]), .Z(n747_adj_2417)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (D))+!A (B (D)+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_0_i747_3_lut_4_lut_3_lut_4_lut.init = 16'h09f6;
    LUT4 i19731_3_lut (.A(n27277), .B(n29949), .C(index_q[3]), .Z(n22086)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19731_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_6_i924_3_lut_4_lut (.A(index_q[2]), .B(index_q[3]), 
         .C(index_q[4]), .D(n762_adj_2326), .Z(n924_adj_2715)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_6_i924_3_lut_4_lut.init = 16'h6f60;
    L6MUX21 i24393 (.D0(n26120), .D1(n26117), .SD(index_q[5]), .Z(n26121));
    LUT4 mux_229_Mux_0_i262_3_lut_3_lut_3_lut_rep_767 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27432)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_0_i262_3_lut_3_lut_3_lut_rep_767.init = 16'hc7c7;
    LUT4 i9480_2_lut_rep_651 (.A(index_i[2]), .B(index_i[3]), .Z(n27316)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9480_2_lut_rep_651.init = 16'h8888;
    LUT4 mux_229_Mux_5_i30_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n30)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A (B+!(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_5_i30_3_lut_4_lut.init = 16'hcc67;
    PFUMX i24391 (.BLUT(n26119), .ALUT(n26118), .C0(index_q[4]), .Z(n26120));
    PFUMX i26897 (.BLUT(n29961), .ALUT(n29962), .C0(index_q[0]), .Z(n29963));
    LUT4 mux_229_Mux_7_i924_3_lut_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[4]), .D(n27434), .Z(n924_adj_2716)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_7_i924_3_lut_3_lut_4_lut.init = 16'h878f;
    LUT4 i11906_2_lut_rep_446_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[4]), .D(n27434), .Z(n27111)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11906_2_lut_rep_446_3_lut_4_lut.init = 16'hf8f0;
    LUT4 index_i_6__bdd_3_lut_24155_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(n27429), .D(index_i[6]), .Z(n25796)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(D))+!A !(D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam index_i_6__bdd_3_lut_24155_4_lut.init = 16'h887f;
    LUT4 i12570_2_lut_rep_491_3_lut (.A(index_i[2]), .B(index_i[3]), .C(index_i[1]), 
         .Z(n27156)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12570_2_lut_rep_491_3_lut.init = 16'h8080;
    PFUMX i24388 (.BLUT(n27081), .ALUT(n26116), .C0(index_q[4]), .Z(n26117));
    LUT4 i19965_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n22320)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+(D)))+!A !(B (D)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19965_3_lut_4_lut_4_lut.init = 16'h99c7;
    LUT4 i6952_3_lut_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), .C(index_i[1]), 
         .D(index_i[0]), .Z(n157_adj_2527)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(D))+!A !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i6952_3_lut_3_lut_4_lut.init = 16'h7780;
    LUT4 i22381_3_lut (.A(n22086), .B(n22087), .C(index_q[4]), .Z(n22088)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22381_3_lut.init = 16'hcaca;
    LUT4 i20369_1_lut_2_lut (.A(index_i[2]), .B(index_i[3]), .Z(n22743)) /* synthesis lut_function=(!(A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20369_1_lut_2_lut.init = 16'h7777;
    LUT4 mux_229_Mux_0_i142_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n142_adj_2711)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C))+!A !(B (C (D)+!C !(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_0_i142_3_lut_4_lut_4_lut.init = 16'ha569;
    LUT4 i12556_2_lut_rep_452_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[4]), .D(n27429), .Z(n27117)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12556_2_lut_rep_452_3_lut_4_lut.init = 16'hf8f0;
    LUT4 n389_bdd_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n26727)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C))+!A (B (C (D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n389_bdd_3_lut_3_lut_4_lut.init = 16'h0fc7;
    LUT4 mux_230_Mux_3_i94_3_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[4]), .D(n93_adj_2687), .Z(n94_adj_2622)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_3_i94_3_lut_4_lut.init = 16'hf606;
    LUT4 index_q_6__bdd_4_lut_25288 (.A(index_q[6]), .B(index_q[5]), .C(index_q[1]), 
         .D(index_q[0]), .Z(n27669)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C))+!A (B (C)+!B !(C)))) */ ;
    defparam index_q_6__bdd_4_lut_25288.init = 16'h3cbc;
    L6MUX21 i24364 (.D0(n26095), .D1(n26092), .SD(index_q[5]), .Z(n26096));
    PFUMX i24362 (.BLUT(n26094), .ALUT(n26093), .C0(index_q[4]), .Z(n26095));
    LUT4 mux_229_Mux_0_i762_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n762_adj_2740)) /* synthesis lut_function=(A (B+!((D)+!C))+!A !(B (D)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_0_i762_3_lut_4_lut_4_lut.init = 16'h98fc;
    LUT4 mux_230_Mux_3_i62_3_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[4]), .D(n812_adj_2628), .Z(n62_adj_2784)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_3_i62_3_lut_4_lut.init = 16'h6f60;
    LUT4 index_q_6__bdd_1_lut_26535 (.A(index_q[5]), .Z(n27668)) /* synthesis lut_function=(!(A)) */ ;
    defparam index_q_6__bdd_1_lut_26535.init = 16'h5555;
    LUT4 mux_230_Mux_4_i828_3_lut_4_lut (.A(index_q[4]), .B(index_q[3]), 
         .C(n812_adj_2768), .D(n29950), .Z(n828_adj_2610)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_4_i828_3_lut_4_lut.init = 16'hf1e0;
    L6MUX21 i23497 (.D0(n25151), .D1(n25149), .SD(index_q[6]), .Z(n25152));
    LUT4 mux_230_Mux_5_i797_3_lut_4_lut (.A(index_q[4]), .B(index_q[3]), 
         .C(n27460), .D(n27274), .Z(n797_adj_2592)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_5_i797_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_230_Mux_11_i766_3_lut (.A(n638_adj_2427), .B(n765), .C(index_q[7]), 
         .Z(n766)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_11_i766_3_lut.init = 16'h3a3a;
    LUT4 i19353_3_lut (.A(n27256), .B(n29923), .C(index_i[3]), .Z(n21708)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19353_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_1_i763_3_lut_4_lut (.A(index_q[4]), .B(index_q[3]), 
         .C(n27551), .D(n27274), .Z(n763_adj_2403)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_1_i763_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_rep_652 (.A(index_q[3]), .B(index_q[2]), .Z(n27317)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i1_2_lut_rep_652.init = 16'h8888;
    LUT4 index_q_1__bdd_3_lut_4_lut (.A(index_q[3]), .B(index_q[2]), .C(index_q[4]), 
         .D(index_q[1]), .Z(n23305)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam index_q_1__bdd_3_lut_4_lut.init = 16'h878f;
    LUT4 i11480_2_lut_rep_769 (.A(index_i[0]), .B(index_i[1]), .Z(n27434)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11480_2_lut_rep_769.init = 16'heeee;
    LUT4 i12568_2_lut_rep_509_3_lut (.A(index_q[3]), .B(index_q[2]), .C(index_q[1]), 
         .Z(n27174)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i12568_2_lut_rep_509_3_lut.init = 16'h8080;
    LUT4 i19729_3_lut (.A(n29958), .B(n29929), .C(index_q[3]), .Z(n22084)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19729_3_lut.init = 16'hcaca;
    LUT4 i19728_3_lut (.A(n27297), .B(n619), .C(index_q[3]), .Z(n22083)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19728_3_lut.init = 16'hcaca;
    PFUMX i23495 (.BLUT(n924_adj_2790), .ALUT(n25150), .C0(index_q[5]), 
          .Z(n25151));
    PFUMX i24359 (.BLUT(n78_adj_2625), .ALUT(n26091), .C0(index_q[4]), 
          .Z(n26092));
    LUT4 i7918_3_lut_3_lut_4_lut (.A(index_q[3]), .B(index_q[2]), .C(index_q[1]), 
         .D(index_q[0]), .Z(n157_adj_2374)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(D))+!A !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i7918_3_lut_3_lut_4_lut.init = 16'h7780;
    LUT4 i22383_3_lut (.A(n22083), .B(n22084), .C(index_q[4]), .Z(n22085)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22383_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_8_i397_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n397_adj_2410)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_8_i397_3_lut_3_lut_4_lut.init = 16'hf10f;
    LUT4 n24852_bdd_3_lut_3_lut (.A(n1021_adj_2722), .B(index_q[8]), .C(n24852), 
         .Z(n24853)) /* synthesis lut_function=(A (B+(C))+!A !(B+!(C))) */ ;
    defparam n24852_bdd_3_lut_3_lut.init = 16'hb8b8;
    LUT4 i20582_3_lut (.A(n22953), .B(n22954), .C(index_i[8]), .Z(n22956)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20582_3_lut.init = 16'hcaca;
    LUT4 n27674_bdd_3_lut (.A(n27674), .B(n27671), .C(index_q[4]), .Z(n27675)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n27674_bdd_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_0_i985_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n985)) /* synthesis lut_function=(!(A (B+!(C))+!A (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_0_i985_3_lut_3_lut.init = 16'h2525;
    LUT4 index_q_2__bdd_4_lut (.A(index_q[2]), .B(index_q[1]), .C(index_q[3]), 
         .D(index_q[0]), .Z(n29960)) /* synthesis lut_function=(A (B ((D)+!C))+!A !(B+!(C+!(D)))) */ ;
    defparam index_q_2__bdd_4_lut.init = 16'h9819;
    LUT4 i9607_3_lut_3_lut_4_lut_3_lut_4_lut (.A(index_q[3]), .B(index_q[2]), 
         .C(index_q[1]), .D(index_q[0]), .Z(n762)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C (D)+!C !(D)))+!A !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i9607_3_lut_3_lut_4_lut_3_lut_4_lut.init = 16'h700f;
    LUT4 i12043_2_lut_rep_501_3_lut_4_lut (.A(index_q[3]), .B(index_q[2]), 
         .C(index_q[1]), .D(index_q[0]), .Z(n27166)) /* synthesis lut_function=(A (B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i12043_2_lut_rep_501_3_lut_4_lut.init = 16'h8880;
    LUT4 mux_229_Mux_3_i30_3_lut_3_lut_4_lut_3_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n30_adj_2460)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_3_i30_3_lut_3_lut_4_lut_3_lut_4_lut.init = 16'hfe11;
    LUT4 i12127_2_lut_2_lut_3_lut (.A(index_q[3]), .B(index_q[2]), .C(index_q[0]), 
         .Z(n14725)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i12127_2_lut_2_lut_3_lut.init = 16'h0808;
    LUT4 i9614_3_lut_4_lut_3_lut_4_lut (.A(index_q[3]), .B(index_q[2]), 
         .C(index_q[1]), .D(index_q[0]), .Z(n875_adj_2282)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(D))+!A !(D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i9614_3_lut_4_lut_3_lut_4_lut.init = 16'h887f;
    LUT4 i15938_3_lut_3_lut_4_lut (.A(index_q[3]), .B(index_q[2]), .C(index_q[1]), 
         .D(index_q[0]), .Z(n18124)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i15938_3_lut_3_lut_4_lut.init = 16'hf078;
    LUT4 i20355_1_lut_2_lut (.A(index_q[3]), .B(index_q[2]), .Z(n22729)) /* synthesis lut_function=(!(A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i20355_1_lut_2_lut.init = 16'h7777;
    LUT4 i1_2_lut_rep_530_3_lut_4_lut (.A(index_q[3]), .B(index_q[2]), .C(index_q[1]), 
         .D(index_q[0]), .Z(n27195)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i1_2_lut_rep_530_3_lut_4_lut.init = 16'h8000;
    LUT4 i21371_3_lut (.A(n23738), .B(n23739), .C(index_q[7]), .Z(n23745)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21371_3_lut.init = 16'hcaca;
    PFUMX i23493 (.BLUT(n25148), .ALUT(n27178), .C0(index_q[5]), .Z(n25149));
    LUT4 i11488_2_lut_rep_466_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n27131)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11488_2_lut_rep_466_3_lut_4_lut.init = 16'hfef0;
    LUT4 i19351_3_lut (.A(n27438), .B(n29956), .C(index_i[3]), .Z(n21706)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19351_3_lut.init = 16'hcaca;
    PFUMX i21185 (.BLUT(n23555), .ALUT(n23556), .C0(index_i[4]), .Z(n23559));
    LUT4 i21370_3_lut (.A(n23736), .B(n23737), .C(index_q[7]), .Z(n23744)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21370_3_lut.init = 16'hcaca;
    LUT4 i21996_3_lut (.A(n21705), .B(n21706), .C(index_i[4]), .Z(n21707)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21996_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_6_i908_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n908_adj_2549)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A (B (C (D)+!C !(D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_6_i908_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h1cf0;
    LUT4 i21375_3_lut (.A(n23746), .B(n23747), .C(index_q[8]), .Z(n23749)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21375_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_4_i541_3_lut_4_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n541_adj_2420)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_4_i541_3_lut_4_lut_3_lut_4_lut.init = 16'h0ef0;
    LUT4 i11837_2_lut_rep_669 (.A(index_q[1]), .B(index_q[2]), .Z(n27334)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i11837_2_lut_rep_669.init = 16'heeee;
    LUT4 mux_229_Mux_7_i506_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n506_adj_2777)) /* synthesis lut_function=(!(A (B (D)+!B ((D)+!C))+!A (B (D)+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_7_i506_3_lut_4_lut_4_lut_4_lut.init = 16'h01ec;
    PFUMX i21186 (.BLUT(n23557), .ALUT(n23558), .C0(index_i[4]), .Z(n23560));
    LUT4 mux_229_Mux_3_i252_3_lut_4_lut (.A(n27214), .B(index_i[3]), .C(index_i[4]), 
         .D(n15004), .Z(n252_adj_2779)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_3_i252_3_lut_4_lut.init = 16'h08f8;
    LUT4 i21327_3_lut (.A(n23696), .B(n23697), .C(index_q[7]), .Z(n23701)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21327_3_lut.init = 16'hcaca;
    LUT4 i20581_3_lut (.A(n22951), .B(n22952), .C(index_i[8]), .Z(n22955)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20581_3_lut.init = 16'hcaca;
    LUT4 i19720_3_lut (.A(n27280), .B(n356), .C(index_q[3]), .Z(n22075)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19720_3_lut.init = 16'hcaca;
    LUT4 mux_230_Mux_4_i236_3_lut_4_lut_3_lut_rep_645_4_lut (.A(index_q[1]), 
         .B(index_q[2]), .C(index_q[3]), .D(index_q[0]), .Z(n27310)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_4_i236_3_lut_4_lut_3_lut_rep_645_4_lut.init = 16'hf01f;
    LUT4 i21319_3_lut (.A(n23680), .B(n25526), .C(index_q[6]), .Z(n23693)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21319_3_lut.init = 16'hcaca;
    LUT4 i21318_3_lut (.A(n25520), .B(n23679), .C(index_q[6]), .Z(n23692)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21318_3_lut.init = 16'hcaca;
    LUT4 i22395_3_lut (.A(n22074), .B(n22075), .C(index_q[4]), .Z(n22076)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22395_3_lut.init = 16'hcaca;
    PFUMX i20695 (.BLUT(n221), .ALUT(n252_adj_2359), .C0(index_q[5]), 
          .Z(n23069));
    PFUMX i9445 (.BLUT(n12151), .ALUT(n12152), .C0(n22743), .Z(n11931));
    PFUMX i9657 (.BLUT(n12172), .ALUT(n12173), .C0(n22740), .Z(n12145));
    LUT4 i9491_3_lut_4_lut_4_lut (.A(index_i[0]), .B(n588), .C(index_i[4]), 
         .D(n27322), .Z(n11977)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B ((D)+!C)+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9491_3_lut_4_lut_4_lut.init = 16'h5c0c;
    LUT4 i1_2_lut_rep_655 (.A(index_i[5]), .B(index_i[6]), .Z(n27320)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_2_lut_rep_655.init = 16'heeee;
    LUT4 mux_230_Mux_9_i93_3_lut_3_lut_3_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .Z(n93)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_230_Mux_9_i93_3_lut_3_lut_3_lut.init = 16'hc1c1;
    LUT4 i1_3_lut_4_lut_adj_87 (.A(index_i[5]), .B(index_i[6]), .C(index_i[7]), 
         .D(n27321), .Z(n20713)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_3_lut_4_lut_adj_87.init = 16'hfffe;
    LUT4 i21316_3_lut (.A(n25712), .B(n23675), .C(index_q[6]), .Z(n23690)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21316_3_lut.init = 16'hcaca;
    LUT4 i8260_2_lut_rep_656 (.A(index_i[3]), .B(index_i[4]), .Z(n27321)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i8260_2_lut_rep_656.init = 16'h8888;
    LUT4 i12539_2_lut_3_lut (.A(index_i[3]), .B(index_i[4]), .C(index_i[5]), 
         .Z(n15146)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12539_2_lut_3_lut.init = 16'hf8f8;
    LUT4 i1_2_lut_3_lut (.A(index_i[3]), .B(index_i[4]), .C(index_i[5]), 
         .Z(n20888)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_2_lut_3_lut.init = 16'h8080;
    LUT4 i21205_3_lut_3_lut_4_lut (.A(index_i[3]), .B(index_i[4]), .C(n413_adj_2337), 
         .D(index_i[5]), .Z(n23579)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21205_3_lut_3_lut_4_lut.init = 16'h77f0;
    LUT4 i20845_3_lut (.A(n23216), .B(n23217), .C(index_q[8]), .Z(n23219)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20845_3_lut.init = 16'hcaca;
    LUT4 i12585_2_lut_3_lut_4_lut (.A(index_i[3]), .B(index_i[4]), .C(index_i[2]), 
         .D(n27429), .Z(n15194)) /* synthesis lut_function=(A (B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12585_2_lut_3_lut_4_lut.init = 16'h8880;
    LUT4 mux_229_Mux_6_i955_3_lut_4_lut (.A(n27214), .B(index_i[3]), .C(index_i[4]), 
         .D(n27072), .Z(n955_adj_2732)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_6_i955_3_lut_4_lut.init = 16'h8f80;
    LUT4 i20894_3_lut (.A(n23261), .B(n23262), .C(index_i[7]), .Z(n23268)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20894_3_lut.init = 16'hcaca;
    LUT4 i11996_2_lut_rep_493_3_lut (.A(index_q[1]), .B(index_q[2]), .C(index_q[0]), 
         .Z(n27158)) /* synthesis lut_function=(A (C)+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i11996_2_lut_rep_493_3_lut.init = 16'hf1f1;
    LUT4 i22135_3_lut (.A(n21702), .B(n21703), .C(index_i[4]), .Z(n21704)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22135_3_lut.init = 16'hcaca;
    PFUMX i9569 (.BLUT(n12165), .ALUT(n12166), .C0(n22729), .Z(n12055));
    PFUMX i25251 (.BLUT(n27623), .ALUT(n27622), .C0(index_i[2]), .Z(n27624));
    LUT4 i20893_3_lut (.A(n23259), .B(n23260), .C(index_i[7]), .Z(n23267)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20893_3_lut.init = 16'hcaca;
    LUT4 i19716_3_lut (.A(n14), .B(n27278), .C(index_q[3]), .Z(n22071)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19716_3_lut.init = 16'hcaca;
    LUT4 i11402_2_lut_rep_657 (.A(index_i[1]), .B(index_i[2]), .Z(n27322)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11402_2_lut_rep_657.init = 16'heeee;
    PFUMX i20725 (.BLUT(n158_adj_2375), .ALUT(n189_adj_2462), .C0(index_q[5]), 
          .Z(n23099));
    LUT4 i11639_2_lut_rep_518_3_lut (.A(index_q[1]), .B(index_q[2]), .C(index_q[3]), 
         .Z(n27183)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i11639_2_lut_rep_518_3_lut.init = 16'he0e0;
    LUT4 i20945_3_lut_4_lut (.A(n27214), .B(index_i[3]), .C(index_i[4]), 
         .D(n364_adj_2618), .Z(n23319)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20945_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_229_Mux_10_i62_3_lut_3_lut_4_lut (.A(n27214), .B(index_i[3]), 
         .C(n27159), .D(index_i[4]), .Z(n62_adj_2475)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_10_i62_3_lut_3_lut_4_lut.init = 16'hf077;
    LUT4 i11868_2_lut_rep_405_3_lut_4_lut (.A(n27214), .B(index_i[3]), .C(index_i[5]), 
         .D(index_i[4]), .Z(n27070)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11868_2_lut_rep_405_3_lut_4_lut.init = 16'hf080;
    LUT4 n954_bdd_3_lut_23936_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[4]), .D(index_i[3]), .Z(n25644)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C+(D)))+!A (B (C (D)+!C !(D))+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n954_bdd_3_lut_23936_4_lut_4_lut_4_lut.init = 16'hc10f;
    LUT4 i20750_3_lut (.A(n23119), .B(n23120), .C(index_q[7]), .Z(n23124)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20750_3_lut.init = 16'hcaca;
    LUT4 i19710_3_lut (.A(n29958), .B(n27425), .C(index_q[3]), .Z(n22065)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19710_3_lut.init = 16'hcaca;
    LUT4 i19342_3_lut (.A(n498), .B(n27257), .C(index_i[3]), .Z(n21697)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19342_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_11_i766_3_lut (.A(n638_adj_2419), .B(n765_adj_2772), 
         .C(index_i[7]), .Z(n766_adj_2791)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_11_i766_3_lut.init = 16'h3a3a;
    PFUMX i15904 (.BLUT(n18088), .ALUT(n18089), .C0(index_i[4]), .Z(n18090));
    LUT4 i22915_3_lut (.A(n766_adj_2791), .B(n20713), .C(index_i[8]), 
         .Z(n21757)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22915_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_3_i189_3_lut_3_lut_4_lut (.A(n27214), .B(index_i[3]), 
         .C(index_i[4]), .D(n27156), .Z(n189_adj_2778)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_3_i189_3_lut_3_lut_4_lut.init = 16'h08f8;
    PFUMX i21221 (.BLUT(n23591), .ALUT(n23592), .C0(index_i[4]), .Z(n23595));
    PFUMX i21222 (.BLUT(n23593), .ALUT(n23594), .C0(index_i[4]), .Z(n23596));
    PFUMX i21228 (.BLUT(n23598), .ALUT(n23599), .C0(index_i[4]), .Z(n23602));
    LUT4 i20020_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n22375)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)+!C !(D)))+!A (B (C+!(D))+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20020_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h0e30;
    PFUMX i23299 (.BLUT(n24882), .ALUT(n1022_adj_2774), .C0(index_q[9]), 
          .Z(quarter_wave_sample_register_q_15__N_2160[12]));
    LUT4 i19388_then_4_lut (.A(index_i[2]), .B(index_i[1]), .C(index_i[4]), 
         .D(index_i[3]), .Z(n27478)) /* synthesis lut_function=(A (B (C+(D))+!B !(C))+!A !(B (C+(D))+!B !(C+!(D)))) */ ;
    defparam i19388_then_4_lut.init = 16'h9a97;
    LUT4 mux_229_Mux_9_i93_3_lut_3_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .Z(n93_adj_2792)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_9_i93_3_lut_3_lut_3_lut.init = 16'hc1c1;
    LUT4 i12106_2_lut_rep_433_2_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .Z(n27098)) /* synthesis lut_function=(A (C)+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12106_2_lut_rep_433_2_lut_3_lut.init = 16'hf1f1;
    LUT4 i20686_3_lut (.A(n23053), .B(n23054), .C(index_q[7]), .Z(n23060)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20686_3_lut.init = 16'hcaca;
    LUT4 i20685_3_lut (.A(n23051), .B(n23052), .C(index_q[7]), .Z(n23059)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20685_3_lut.init = 16'hcaca;
    LUT4 i11896_2_lut_rep_535_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[3]), 
         .Z(n27200)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11896_2_lut_rep_535_3_lut.init = 16'he0e0;
    PFUMX i24259 (.BLUT(n25983), .ALUT(n25979), .C0(index_i[6]), .Z(n25984));
    LUT4 i19681_3_lut (.A(n27289), .B(n27277), .C(index_q[3]), .Z(n22036)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19681_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_3_i109_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n109_adj_2496)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (D)+!B !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_3_i109_3_lut_4_lut_4_lut.init = 16'hcf10;
    LUT4 i11897_2_lut_rep_455_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[4]), .D(index_i[3]), .Z(n27120)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11897_2_lut_rep_455_3_lut_4_lut.init = 16'hfef0;
    LUT4 i7267_2_lut_rep_658 (.A(index_q[3]), .B(index_q[4]), .Z(n27323)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i7267_2_lut_rep_658.init = 16'h8888;
    LUT4 i19596_3_lut_then_4_lut (.A(index_q[4]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n29962)) /* synthesis lut_function=(A (B (C)+!B !(C (D)+!C !(D)))+!A !(B (C)+!B !(C (D)+!C !(D)))) */ ;
    defparam i19596_3_lut_then_4_lut.init = 16'h96a5;
    LUT4 i20404_3_lut_3_lut_4_lut (.A(index_q[3]), .B(index_q[4]), .C(n413), 
         .D(index_q[5]), .Z(n22778)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i20404_3_lut_3_lut_4_lut.init = 16'h77f0;
    LUT4 i1_2_lut_rep_517_3_lut (.A(index_q[3]), .B(index_q[4]), .C(index_q[5]), 
         .Z(n27182)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i1_2_lut_rep_517_3_lut.init = 16'hf8f8;
    LUT4 i1_2_lut_3_lut_adj_88 (.A(index_q[3]), .B(index_q[4]), .C(index_q[5]), 
         .Z(n20896)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i1_2_lut_3_lut_adj_88.init = 16'h8080;
    LUT4 i19341_3_lut (.A(n27346), .B(n356_adj_2398), .C(index_i[3]), 
         .Z(n21696)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19341_3_lut.init = 16'hcaca;
    LUT4 i19798_3_lut_3_lut_4_lut (.A(n27213), .B(index_i[3]), .C(n93_adj_2792), 
         .D(index_i[4]), .Z(n22153)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19798_3_lut_3_lut_4_lut.init = 16'h11f0;
    LUT4 i19339_3_lut (.A(n27346), .B(n27257), .C(index_i[3]), .Z(n21694)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19339_3_lut.init = 16'hcaca;
    LUT4 i11640_2_lut_rep_451_3_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[4]), .D(index_q[3]), .Z(n27116)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i11640_2_lut_rep_451_3_lut_4_lut.init = 16'hfef0;
    LUT4 i19698_3_lut_3_lut_4_lut (.A(index_q[1]), .B(index_q[2]), .C(index_q[3]), 
         .D(index_q[0]), .Z(n22053)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i19698_3_lut_3_lut_4_lut.init = 16'h0fe0;
    LUT4 i19338_3_lut (.A(n356_adj_2398), .B(n204), .C(index_i[3]), .Z(n21693)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19338_3_lut.init = 16'hcaca;
    LUT4 n557_bdd_3_lut_23886_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[4]), .D(index_q[3]), .Z(n25596)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C+(D)))+!A (B (C (D)+!C !(D))+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam n557_bdd_3_lut_23886_4_lut_4_lut_4_lut.init = 16'hc10f;
    LUT4 i19774_3_lut_3_lut (.A(n27096), .B(index_i[4]), .C(n109_adj_2496), 
         .Z(n22129)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam i19774_3_lut_3_lut.init = 16'h7474;
    LUT4 i11887_3_lut_4_lut (.A(n27213), .B(index_i[3]), .C(n10667), .D(index_i[6]), 
         .Z(n765_adj_2772)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11887_3_lut_4_lut.init = 16'hffe0;
    LUT4 i8266_2_lut_rep_670 (.A(index_i[3]), .B(index_i[4]), .Z(n27335)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i8266_2_lut_rep_670.init = 16'heeee;
    LUT4 n124_bdd_3_lut_4_lut_adj_89 (.A(n27213), .B(index_i[3]), .C(index_i[4]), 
         .D(n93_adj_2792), .Z(n25782)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n124_bdd_3_lut_4_lut_adj_89.init = 16'hfe0e;
    LUT4 i19705_3_lut (.A(n29953), .B(n27274), .C(index_q[3]), .Z(n22060)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19705_3_lut.init = 16'hcaca;
    LUT4 i19704_3_lut (.A(n29948), .B(n356), .C(index_q[3]), .Z(n22059)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19704_3_lut.init = 16'hcaca;
    PFUMX i21229 (.BLUT(n23600), .ALUT(n23601), .C0(index_i[4]), .Z(n23603));
    PFUMX i24208 (.BLUT(n25921), .ALUT(n25918), .C0(index_i[6]), .Z(n22915));
    PFUMX i21235 (.BLUT(n23605), .ALUT(n23606), .C0(index_i[4]), .Z(n23609));
    PFUMX i23295 (.BLUT(n254_adj_2727), .ALUT(n24876), .C0(index_q[8]), 
          .Z(n24877));
    PFUMX i21236 (.BLUT(n23607), .ALUT(n23608), .C0(index_i[4]), .Z(n23610));
    LUT4 i22406_3_lut (.A(n22059), .B(n22060), .C(index_q[4]), .Z(n22061)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22406_3_lut.init = 16'hcaca;
    PFUMX i23278 (.BLUT(n24855), .ALUT(n24853), .C0(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_2160[10]));
    PFUMX i23276 (.BLUT(n21786), .ALUT(n24851), .C0(index_q[7]), .Z(n24852));
    PFUMX i23274 (.BLUT(n24849), .ALUT(n1022), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2145[12]));
    LUT4 i20844_3_lut (.A(n23214), .B(n23215), .C(index_q[8]), .Z(n23218)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20844_3_lut.init = 16'hcaca;
    LUT4 mux_229_Mux_10_i317_3_lut_3_lut_4_lut (.A(n27213), .B(index_i[3]), 
         .C(n27156), .D(index_i[4]), .Z(n317_adj_2752)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_229_Mux_10_i317_3_lut_3_lut_4_lut.init = 16'hf011;
    CCU2D add_417_5 (.A0(quarter_wave_sample_register_i[4]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[5]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17895), .COUT(n17896));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam add_417_5.INIT0 = 16'hf555;
    defparam add_417_5.INIT1 = 16'hf555;
    defparam add_417_5.INJECT1_0 = "NO";
    defparam add_417_5.INJECT1_1 = "NO";
    CCU2D add_417_3 (.A0(quarter_wave_sample_register_i[2]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[3]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17894), .COUT(n17895));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam add_417_3.INIT0 = 16'hf555;
    defparam add_417_3.INIT1 = 16'hf555;
    defparam add_417_3.INJECT1_0 = "NO";
    defparam add_417_3.INJECT1_1 = "NO";
    CCU2D add_417_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(quarter_wave_sample_register_i[0]), .B1(quarter_wave_sample_register_i[1]), 
          .C1(GND_net), .D1(GND_net), .COUT(n17894));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam add_417_1.INIT0 = 16'hF000;
    defparam add_417_1.INIT1 = 16'ha666;
    defparam add_417_1.INJECT1_0 = "NO";
    defparam add_417_1.INJECT1_1 = "NO";
    PFUMX i20645 (.BLUT(n23017), .ALUT(n23018), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2145[1]));
    LUT4 i9451_3_lut_4_lut (.A(index_i[3]), .B(index_i[4]), .C(n29915), 
         .D(n29956), .Z(n605_adj_2764)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9451_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i21179_3_lut (.A(n23550), .B(n23551), .C(index_i[7]), .Z(n23553)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21179_3_lut.init = 16'hcaca;
    LUT4 i21178_3_lut (.A(n23548), .B(n23549), .C(index_i[7]), .Z(n23552)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21178_3_lut.init = 16'hcaca;
    PFUMX i24129 (.BLUT(n25839), .ALUT(n27339), .C0(index_i[5]), .Z(n25840));
    PFUMX i24127 (.BLUT(n27247), .ALUT(n25837), .C0(index_i[2]), .Z(n25838));
    FD1P3AX phase_i_i0_i11 (.D(o_phase[11]), .SP(dac_clk_p_c_enable_488), 
            .CK(dac_clk_p_c), .Q(phase_i[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam phase_i_i0_i11.GSR = "DISABLED";
    L6MUX21 i24125 (.D0(n25835), .D1(n25832), .SD(index_i[5]), .Z(n25836));
    PFUMX i24123 (.BLUT(n25834), .ALUT(n25833), .C0(index_i[4]), .Z(n25835));
    FD1P3AX phase_i_i0_i10 (.D(o_phase[10]), .SP(dac_clk_p_c_enable_488), 
            .CK(dac_clk_p_c), .Q(phase_i[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam phase_i_i0_i10.GSR = "DISABLED";
    PFUMX i24120 (.BLUT(n25831), .ALUT(n25830), .C0(index_i[4]), .Z(n25832));
    PFUMX i20722 (.BLUT(n23094), .ALUT(n23095), .C0(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_2160[5]));
    L6MUX21 i24117 (.D0(n25828), .D1(n25826), .SD(index_i[5]), .Z(n25829));
    PFUMX i24115 (.BLUT(n25827), .ALUT(n285_adj_2489), .C0(index_i[4]), 
          .Z(n25828));
    PFUMX i24113 (.BLUT(n25825), .ALUT(n25824), .C0(index_i[4]), .Z(n25826));
    PFUMX i23270 (.BLUT(n254_adj_2728), .ALUT(n24843), .C0(index_i[8]), 
          .Z(n24844));
    PFUMX i20784 (.BLUT(n23156), .ALUT(n23157), .C0(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_2160[3]));
    L6MUX21 i24107 (.D0(n25818), .D1(n25815), .SD(index_i[5]), .Z(n25819));
    PFUMX i24105 (.BLUT(n15_adj_2503), .ALUT(n25816), .C0(index_i[4]), 
          .Z(n25818));
    PFUMX i24102 (.BLUT(n25814), .ALUT(n25813), .C0(index_i[4]), .Z(n25815));
    
endmodule
//
// Verilog Description of module \nco(OW=12)_U1 
//

module \nco(OW=12)_U1  (increment, o_phase, GND_net, dac_clk_p_c, i_sw0_c) /* synthesis syn_module_defined=1 */ ;
    input [30:0]increment;
    output [11:0]o_phase;
    input GND_net;
    input dac_clk_p_c;
    input i_sw0_c;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[49:58])
    
    wire n18029;
    wire [31:0]n133;
    
    wire n18028, n18027, n18026, n18025, n18024, n18023;
    wire [31:0]n233;
    
    wire n18022, n18021, n18020, n18019, n18018, n18017, n18016, 
        n18015;
    
    CCU2D phase_register_597_add_4_32 (.A0(increment[30]), .B0(o_phase[10]), 
          .C0(GND_net), .D0(GND_net), .A1(o_phase[11]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n18029), .S0(n133[30]), .S1(n133[31]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_597_add_4_32.INIT0 = 16'h5666;
    defparam phase_register_597_add_4_32.INIT1 = 16'hfaaa;
    defparam phase_register_597_add_4_32.INJECT1_0 = "NO";
    defparam phase_register_597_add_4_32.INJECT1_1 = "NO";
    CCU2D phase_register_597_add_4_30 (.A0(increment[28]), .B0(o_phase[8]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[29]), .B1(o_phase[9]), 
          .C1(GND_net), .D1(GND_net), .CIN(n18028), .COUT(n18029), .S0(n133[28]), 
          .S1(n133[29]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_597_add_4_30.INIT0 = 16'h5666;
    defparam phase_register_597_add_4_30.INIT1 = 16'h5666;
    defparam phase_register_597_add_4_30.INJECT1_0 = "NO";
    defparam phase_register_597_add_4_30.INJECT1_1 = "NO";
    CCU2D phase_register_597_add_4_28 (.A0(increment[26]), .B0(o_phase[6]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[27]), .B1(o_phase[7]), 
          .C1(GND_net), .D1(GND_net), .CIN(n18027), .COUT(n18028), .S0(n133[26]), 
          .S1(n133[27]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_597_add_4_28.INIT0 = 16'h5666;
    defparam phase_register_597_add_4_28.INIT1 = 16'h5666;
    defparam phase_register_597_add_4_28.INJECT1_0 = "NO";
    defparam phase_register_597_add_4_28.INJECT1_1 = "NO";
    CCU2D phase_register_597_add_4_26 (.A0(increment[24]), .B0(o_phase[4]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[25]), .B1(o_phase[5]), 
          .C1(GND_net), .D1(GND_net), .CIN(n18026), .COUT(n18027), .S0(n133[24]), 
          .S1(n133[25]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_597_add_4_26.INIT0 = 16'h5666;
    defparam phase_register_597_add_4_26.INIT1 = 16'h5666;
    defparam phase_register_597_add_4_26.INJECT1_0 = "NO";
    defparam phase_register_597_add_4_26.INJECT1_1 = "NO";
    CCU2D phase_register_597_add_4_24 (.A0(increment[22]), .B0(o_phase[2]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[23]), .B1(o_phase[3]), 
          .C1(GND_net), .D1(GND_net), .CIN(n18025), .COUT(n18026), .S0(n133[22]), 
          .S1(n133[23]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_597_add_4_24.INIT0 = 16'h5666;
    defparam phase_register_597_add_4_24.INIT1 = 16'h5666;
    defparam phase_register_597_add_4_24.INJECT1_0 = "NO";
    defparam phase_register_597_add_4_24.INJECT1_1 = "NO";
    CCU2D phase_register_597_add_4_22 (.A0(increment[20]), .B0(o_phase[0]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[21]), .B1(o_phase[1]), 
          .C1(GND_net), .D1(GND_net), .CIN(n18024), .COUT(n18025), .S0(n133[20]), 
          .S1(n133[21]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_597_add_4_22.INIT0 = 16'h5666;
    defparam phase_register_597_add_4_22.INIT1 = 16'h5666;
    defparam phase_register_597_add_4_22.INJECT1_0 = "NO";
    defparam phase_register_597_add_4_22.INJECT1_1 = "NO";
    CCU2D phase_register_597_add_4_20 (.A0(increment[18]), .B0(n233[18]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[19]), .B1(n233[19]), 
          .C1(GND_net), .D1(GND_net), .CIN(n18023), .COUT(n18024), .S0(n133[18]), 
          .S1(n133[19]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_597_add_4_20.INIT0 = 16'h5666;
    defparam phase_register_597_add_4_20.INIT1 = 16'h5666;
    defparam phase_register_597_add_4_20.INJECT1_0 = "NO";
    defparam phase_register_597_add_4_20.INJECT1_1 = "NO";
    CCU2D phase_register_597_add_4_18 (.A0(increment[16]), .B0(n233[16]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[17]), .B1(n233[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n18022), .COUT(n18023), .S0(n133[16]), 
          .S1(n133[17]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_597_add_4_18.INIT0 = 16'h5666;
    defparam phase_register_597_add_4_18.INIT1 = 16'h5666;
    defparam phase_register_597_add_4_18.INJECT1_0 = "NO";
    defparam phase_register_597_add_4_18.INJECT1_1 = "NO";
    CCU2D phase_register_597_add_4_16 (.A0(increment[14]), .B0(n233[14]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[15]), .B1(n233[15]), 
          .C1(GND_net), .D1(GND_net), .CIN(n18021), .COUT(n18022), .S0(n133[14]), 
          .S1(n133[15]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_597_add_4_16.INIT0 = 16'h5666;
    defparam phase_register_597_add_4_16.INIT1 = 16'h5666;
    defparam phase_register_597_add_4_16.INJECT1_0 = "NO";
    defparam phase_register_597_add_4_16.INJECT1_1 = "NO";
    CCU2D phase_register_597_add_4_14 (.A0(increment[12]), .B0(n233[12]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[13]), .B1(n233[13]), 
          .C1(GND_net), .D1(GND_net), .CIN(n18020), .COUT(n18021), .S0(n133[12]), 
          .S1(n133[13]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_597_add_4_14.INIT0 = 16'h5666;
    defparam phase_register_597_add_4_14.INIT1 = 16'h5666;
    defparam phase_register_597_add_4_14.INJECT1_0 = "NO";
    defparam phase_register_597_add_4_14.INJECT1_1 = "NO";
    CCU2D phase_register_597_add_4_12 (.A0(increment[10]), .B0(n233[10]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[11]), .B1(n233[11]), 
          .C1(GND_net), .D1(GND_net), .CIN(n18019), .COUT(n18020), .S0(n133[10]), 
          .S1(n133[11]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_597_add_4_12.INIT0 = 16'h5666;
    defparam phase_register_597_add_4_12.INIT1 = 16'h5666;
    defparam phase_register_597_add_4_12.INJECT1_0 = "NO";
    defparam phase_register_597_add_4_12.INJECT1_1 = "NO";
    CCU2D phase_register_597_add_4_10 (.A0(increment[8]), .B0(n233[8]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[9]), .B1(n233[9]), 
          .C1(GND_net), .D1(GND_net), .CIN(n18018), .COUT(n18019), .S0(n133[8]), 
          .S1(n133[9]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_597_add_4_10.INIT0 = 16'h5666;
    defparam phase_register_597_add_4_10.INIT1 = 16'h5666;
    defparam phase_register_597_add_4_10.INJECT1_0 = "NO";
    defparam phase_register_597_add_4_10.INJECT1_1 = "NO";
    CCU2D phase_register_597_add_4_8 (.A0(increment[6]), .B0(n233[6]), .C0(GND_net), 
          .D0(GND_net), .A1(increment[7]), .B1(n233[7]), .C1(GND_net), 
          .D1(GND_net), .CIN(n18017), .COUT(n18018), .S0(n133[6]), .S1(n133[7]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_597_add_4_8.INIT0 = 16'h5666;
    defparam phase_register_597_add_4_8.INIT1 = 16'h5666;
    defparam phase_register_597_add_4_8.INJECT1_0 = "NO";
    defparam phase_register_597_add_4_8.INJECT1_1 = "NO";
    CCU2D phase_register_597_add_4_6 (.A0(increment[4]), .B0(n233[4]), .C0(GND_net), 
          .D0(GND_net), .A1(increment[5]), .B1(n233[5]), .C1(GND_net), 
          .D1(GND_net), .CIN(n18016), .COUT(n18017), .S0(n133[4]), .S1(n133[5]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_597_add_4_6.INIT0 = 16'h5666;
    defparam phase_register_597_add_4_6.INIT1 = 16'h5666;
    defparam phase_register_597_add_4_6.INJECT1_0 = "NO";
    defparam phase_register_597_add_4_6.INJECT1_1 = "NO";
    CCU2D phase_register_597_add_4_4 (.A0(increment[2]), .B0(n233[2]), .C0(GND_net), 
          .D0(GND_net), .A1(increment[3]), .B1(n233[3]), .C1(GND_net), 
          .D1(GND_net), .CIN(n18015), .COUT(n18016), .S0(n133[2]), .S1(n133[3]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_597_add_4_4.INIT0 = 16'h5666;
    defparam phase_register_597_add_4_4.INIT1 = 16'h5666;
    defparam phase_register_597_add_4_4.INJECT1_0 = "NO";
    defparam phase_register_597_add_4_4.INJECT1_1 = "NO";
    CCU2D phase_register_597_add_4_2 (.A0(increment[0]), .B0(n233[0]), .C0(GND_net), 
          .D0(GND_net), .A1(increment[1]), .B1(n233[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n18015), .S1(n133[1]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_597_add_4_2.INIT0 = 16'h7000;
    defparam phase_register_597_add_4_2.INIT1 = 16'h5666;
    defparam phase_register_597_add_4_2.INJECT1_0 = "NO";
    defparam phase_register_597_add_4_2.INJECT1_1 = "NO";
    LUT4 i15863_2_lut (.A(increment[0]), .B(n233[0]), .Z(n133[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i15863_2_lut.init = 16'h6666;
    FD1S3DX phase_register_597__i0 (.D(n133[0]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[0])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_597__i0.GSR = "DISABLED";
    FD1S3DX phase_register_597__i31 (.D(n133[31]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_phase[11])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_597__i31.GSR = "DISABLED";
    FD1S3DX phase_register_597__i30 (.D(n133[30]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_phase[10])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_597__i30.GSR = "DISABLED";
    FD1S3DX phase_register_597__i29 (.D(n133[29]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_phase[9])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_597__i29.GSR = "DISABLED";
    FD1S3DX phase_register_597__i28 (.D(n133[28]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_phase[8])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_597__i28.GSR = "DISABLED";
    FD1S3DX phase_register_597__i27 (.D(n133[27]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_phase[7])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_597__i27.GSR = "DISABLED";
    FD1S3DX phase_register_597__i26 (.D(n133[26]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_phase[6])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_597__i26.GSR = "DISABLED";
    FD1S3DX phase_register_597__i25 (.D(n133[25]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_phase[5])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_597__i25.GSR = "DISABLED";
    FD1S3DX phase_register_597__i24 (.D(n133[24]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_phase[4])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_597__i24.GSR = "DISABLED";
    FD1S3DX phase_register_597__i23 (.D(n133[23]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_phase[3])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_597__i23.GSR = "DISABLED";
    FD1S3DX phase_register_597__i22 (.D(n133[22]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_phase[2])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_597__i22.GSR = "DISABLED";
    FD1S3DX phase_register_597__i21 (.D(n133[21]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_phase[1])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_597__i21.GSR = "DISABLED";
    FD1S3DX phase_register_597__i20 (.D(n133[20]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_phase[0])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_597__i20.GSR = "DISABLED";
    FD1S3DX phase_register_597__i19 (.D(n133[19]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[19])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_597__i19.GSR = "DISABLED";
    FD1S3DX phase_register_597__i18 (.D(n133[18]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[18])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_597__i18.GSR = "DISABLED";
    FD1S3DX phase_register_597__i17 (.D(n133[17]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[17])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_597__i17.GSR = "DISABLED";
    FD1S3DX phase_register_597__i16 (.D(n133[16]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[16])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_597__i16.GSR = "DISABLED";
    FD1S3DX phase_register_597__i15 (.D(n133[15]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[15])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_597__i15.GSR = "DISABLED";
    FD1S3DX phase_register_597__i14 (.D(n133[14]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[14])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_597__i14.GSR = "DISABLED";
    FD1S3DX phase_register_597__i13 (.D(n133[13]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[13])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_597__i13.GSR = "DISABLED";
    FD1S3DX phase_register_597__i12 (.D(n133[12]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[12])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_597__i12.GSR = "DISABLED";
    FD1S3DX phase_register_597__i11 (.D(n133[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[11])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_597__i11.GSR = "DISABLED";
    FD1S3DX phase_register_597__i10 (.D(n133[10]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[10])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_597__i10.GSR = "DISABLED";
    FD1S3DX phase_register_597__i9 (.D(n133[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[9])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_597__i9.GSR = "DISABLED";
    FD1S3DX phase_register_597__i8 (.D(n133[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[8])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_597__i8.GSR = "DISABLED";
    FD1S3DX phase_register_597__i7 (.D(n133[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[7])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_597__i7.GSR = "DISABLED";
    FD1S3DX phase_register_597__i6 (.D(n133[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[6])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_597__i6.GSR = "DISABLED";
    FD1S3DX phase_register_597__i5 (.D(n133[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[5])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_597__i5.GSR = "DISABLED";
    FD1S3DX phase_register_597__i4 (.D(n133[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[4])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_597__i4.GSR = "DISABLED";
    FD1S3DX phase_register_597__i3 (.D(n133[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[3])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_597__i3.GSR = "DISABLED";
    FD1S3DX phase_register_597__i2 (.D(n133[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[2])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_597__i2.GSR = "DISABLED";
    FD1S3DX phase_register_597__i1 (.D(n133[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[1])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_597__i1.GSR = "DISABLED";
    
endmodule
