// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.12.0.240.2
// Netlist written on Sun Apr 11 02:50:10 2021
//
// Verilog Description of module top
//

module top (i_ref_clk, i_wbu_uart_rx, o_wbu_uart_tx, i_sw0, i_sw1, 
            o_dac_a, o_dac_b, dac_clk_p, dac_clk_n, o_dac_cw_b, o_lo_i, 
            o_lo_q) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(4[8:11])
    input i_ref_clk;   // d:/documents/git_local/fm_modulator/rtl/top.v(26[12:21])
    input i_wbu_uart_rx;   // d:/documents/git_local/fm_modulator/rtl/top.v(28[12:25])
    output o_wbu_uart_tx;   // d:/documents/git_local/fm_modulator/rtl/top.v(29[13:26])
    input i_sw0;   // d:/documents/git_local/fm_modulator/rtl/top.v(31[12:17])
    input i_sw1;   // d:/documents/git_local/fm_modulator/rtl/top.v(31[19:24])
    output [9:0]o_dac_a;   // d:/documents/git_local/fm_modulator/rtl/top.v(33[38:45])
    output [9:0]o_dac_b;   // d:/documents/git_local/fm_modulator/rtl/top.v(33[47:54])
    output dac_clk_p;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[29:38])
    output dac_clk_n;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[40:49])
    output o_dac_cw_b;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[51:61])
    output o_lo_i;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[13:19])
    output o_lo_q;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[21:27])
    
    wire i_ref_clk_c /* synthesis is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(26[12:21])
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[29:38])
    wire lo_q /* synthesis is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(159[24:28])
    
    wire GND_net, VCC_net, i_wbu_uart_rx_c, o_wbu_uart_tx_c, i_sw0_c, 
        o_dac_a_c_9, o_dac_a_c_8, o_dac_a_c_7, o_dac_a_c_6, o_dac_a_c_5, 
        o_dac_a_c_4, o_dac_a_c_3, o_dac_a_c_2, o_dac_a_c_1, o_dac_a_c_0, 
        o_dac_b_c_9, o_dac_b_c_8, o_dac_b_c_7, o_dac_b_c_6, o_dac_b_c_5, 
        o_dac_b_c_4, o_dac_b_c_3, o_dac_b_c_2, o_dac_b_c_1, o_dac_b_c_0, 
        o_lo_i_c, o_lo_q_c, dac_clk_n_c, o_dac_cw_b_c, rx_stb;
    wire [7:0]rx_data;   // d:/documents/git_local/fm_modulator/rtl/top.v(58[12:19])
    
    wire tx_stb, tx_busy;
    wire [7:0]tx_data;   // d:/documents/git_local/fm_modulator/rtl/top.v(66[12:19])
    
    wire wb_cyc, wb_stb, wb_we;
    wire [29:0]wb_addr;   // d:/documents/git_local/fm_modulator/rtl/top.v(75[13:20])
    wire [31:0]wb_odata;   // d:/documents/git_local/fm_modulator/rtl/top.v(76[13:21])
    
    wire wb_ack, wb_err;
    wire [31:0]wb_idata;   // d:/documents/git_local/fm_modulator/rtl/top.v(81[12:20])
    
    wire wb_fm_ack;
    wire [31:0]wb_fm_data;   // d:/documents/git_local/fm_modulator/rtl/top.v(114[13:23])
    wire [7:0]wb_lo_data;   // d:/documents/git_local/fm_modulator/rtl/top.v(137[12:22])
    
    wire wb_lo_ack, pll_clk, pll_rst, pll_stb, pll_we, pll_ack;
    wire [7:0]pll_data_i;   // d:/documents/git_local/fm_modulator/rtl/top.v(143[12:22])
    wire [7:0]pll_data_o;   // d:/documents/git_local/fm_modulator/rtl/top.v(143[24:34])
    wire [4:0]pll_addr;   // d:/documents/git_local/fm_modulator/rtl/top.v(144[12:20])
    
    wire lo_i_en, lo_q_en, wb_control_ack;
    wire [31:0]wb_control_data;   // d:/documents/git_local/fm_modulator/rtl/top.v(203[13:28])
    
    wire none_sel, o_dac_a_9__N_1, wb_lo_data_7__N_34, wb_control_data_31__N_35, 
        wb_control_sel_N_78, wb_lo_sel_N_80;
    wire [31:0]wb_idata_31__N_36;
    wire [31:0]wb_idata_31__N_2;
    wire [23:0]chg_counter;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(97[17:28])
    
    wire chg_counter_23__N_173, n22828, n22822, n22816, n2;
    wire [31:0]\addr_space[1]_adj_3700 ;   // d:/documents/git_local/fm_modulator/rtl/control.v(22[12:22])
    wire [31:0]\addr_space[2]_adj_3701 ;   // d:/documents/git_local/fm_modulator/rtl/control.v(22[12:22])
    wire [31:0]\addr_space[3]_adj_3702 ;   // d:/documents/git_local/fm_modulator/rtl/control.v(22[12:22])
    wire [31:0]\addr_space[4]_adj_3703 ;   // d:/documents/git_local/fm_modulator/rtl/control.v(22[12:22])
    
    wire n22808;
    wire [31:0]o_wb_data_31__N_2456;
    
    wire n26570, n26569, n26568, n22782, n22780, n22774, n22470, 
        n26546, n26545, n21641, n26544, dac_clk_p_c_enable_277, n29065, 
        n22458, n22972, n22448, n22664, n22662, n22660, n22974, 
        n22650, n22976, n29302, n29300, n21662, dac_clk_p_c_enable_502, 
        n14148, n22526, n38, dac_clk_p_c_enable_439, n22966, n34, 
        dac_clk_p_c_enable_407, n29199, n29197, dac_clk_p_c_enable_375, 
        dac_clk_p_c_enable_241, dac_clk_p_c_enable_106, dac_clk_p_c_enable_471, 
        dac_clk_p_c_enable_243, n29155, n4, n22968, n32067, n26, 
        dac_clk_p_c_enable_227, n22940, n32066, n29081;
    
    VHI i2 (.Z(VCC_net));
    GSR GSR_INST (.GSR(i_sw0_c)) /* synthesis syn_instantiated=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(41[6:29])
    FD1S3JX wb_ack_36 (.D(n4), .CK(dac_clk_p_c), .PD(wb_control_ack), 
            .Q(wb_ack)) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(243[8] 244[59])
    defparam wb_ack_36.GSR = "DISABLED";
    \rxuartlite(CLOCKS_PER_BAUD=10000)  rxtransport (.\rx_data[0] (rx_data[0]), 
            .dac_clk_p_c(dac_clk_p_c), .rx_stb(rx_stb), .i_wbu_uart_rx_c(i_wbu_uart_rx_c), 
            .chg_counter({chg_counter}), .dac_clk_p_c_enable_277(dac_clk_p_c_enable_277), 
            .chg_counter_23__N_173(chg_counter_23__N_173), .GND_net(GND_net), 
            .\rx_data[6] (rx_data[6]), .\rx_data[5] (rx_data[5]), .\rx_data[4] (rx_data[4]), 
            .\rx_data[3] (rx_data[3]), .\rx_data[2] (rx_data[2]), .\rx_data[1] (rx_data[1])) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(60[57:105])
    PUR PUR_INST (.PUR(i_sw0_c)) /* synthesis syn_instantiated=1 */ ;
    defparam PUR_INST.RST_PULSE = 1;
    control control_inst (.dac_clk_p_c(dac_clk_p_c), .dac_clk_p_c_enable_227(dac_clk_p_c_enable_227), 
            .wb_odata({wb_odata}), .dac_clk_p_c_enable_243(dac_clk_p_c_enable_243), 
            .i_sw0_c(i_sw0_c), .lo_i_en(lo_i_en), .\addr_space[4][1] (\addr_space[4]_adj_3703 [1]), 
            .\addr_space[4][0] (\addr_space[4]_adj_3703 [0]), .dac_clk_p_c_enable_106(dac_clk_p_c_enable_106), 
            .dac_clk_p_c_enable_241(dac_clk_p_c_enable_241), .wb_control_data({wb_control_data}), 
            .o_wb_data_31__N_2456({Open_0, Open_1, Open_2, Open_3, Open_4, 
            Open_5, Open_6, Open_7, Open_8, Open_9, Open_10, Open_11, 
            Open_12, Open_13, Open_14, Open_15, Open_16, Open_17, 
            Open_18, Open_19, Open_20, Open_21, Open_22, Open_23, 
            Open_24, Open_25, Open_26, Open_27, Open_28, Open_29, 
            Open_30, o_wb_data_31__N_2456[0]}), .lo_q_en(lo_q_en), .\addr_space[1][1] (\addr_space[1]_adj_3700 [1]), 
            .\addr_space[1][0] (\addr_space[1]_adj_3700 [0]), .\addr_space[2][1] (\addr_space[2]_adj_3701 [1]), 
            .\addr_space[2][0] (\addr_space[2]_adj_3701 [0]), .\addr_space[3][1] (\addr_space[3]_adj_3702 [1]), 
            .n29300(n29300), .\wb_addr[2] (wb_addr[2]), .\addr_space[3][0] (\addr_space[3]_adj_3702 [0]), 
            .wb_control_ack(wb_control_ack), .wb_control_data_31__N_35(wb_control_data_31__N_35), 
            .n21662(n21662), .n29302(n29302), .n29065(n29065), .n22526(n22526), 
            .\o_wb_data_31__N_2456[1] (o_wb_data_31__N_2456[1]), .\wb_addr[1] (wb_addr[1]), 
            .\wb_addr[0] (wb_addr[0]), .lo_q(lo_q), .o_lo_q_c(o_lo_q_c)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(204[9] 216[2])
    PFUMX i24949 (.BLUT(n26569), .ALUT(n26568), .C0(wb_addr[1]), .Z(n26570));
    FD1S3IX wb_err_34 (.D(none_sel), .CK(dac_clk_p_c), .CD(n2), .Q(wb_err));   // d:/documents/git_local/fm_modulator/rtl/top.v(232[8] 233[33])
    defparam wb_err_34.GSR = "DISABLED";
    OB o_dac_a_pad_7 (.I(o_dac_a_c_7), .O(o_dac_a[7]));   // d:/documents/git_local/fm_modulator/rtl/top.v(33[38:45])
    OB o_dac_a_pad_8 (.I(o_dac_a_c_8), .O(o_dac_a[8]));   // d:/documents/git_local/fm_modulator/rtl/top.v(33[38:45])
    OB o_dac_a_pad_9 (.I(o_dac_a_c_9), .O(o_dac_a[9]));   // d:/documents/git_local/fm_modulator/rtl/top.v(33[38:45])
    OB o_wbu_uart_tx_pad (.I(o_wbu_uart_tx_c), .O(o_wbu_uart_tx));   // d:/documents/git_local/fm_modulator/rtl/top.v(29[13:26])
    LUT4 n26570_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4]_adj_3703 [0]), 
         .C(wb_addr[2]), .D(n26570), .Z(o_wb_data_31__N_2456[0])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n26570_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 i1_4_lut (.A(n26), .B(wb_addr[15]), .C(wb_addr[12]), .D(wb_addr[9]), 
         .Z(n22526)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(223[20:46])
    defparam i1_4_lut.init = 16'hfffb;
    LUT4 wb_cyc_I_0_2_lut (.A(wb_cyc), .B(wb_lo_sel_N_80), .Z(wb_lo_data_7__N_34)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(187[13:36])
    defparam wb_cyc_I_0_2_lut.init = 16'h2222;
    LUT4 i1_4_lut_adj_228 (.A(n22808), .B(n38), .C(n26), .D(wb_addr[12]), 
         .Z(wb_lo_sel_N_80)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(223[20:46])
    defparam i1_4_lut_adj_228.init = 16'hfffe;
    LUT4 i1_4_lut_adj_229 (.A(n22972), .B(n22974), .C(n22976), .D(chg_counter_23__N_173), 
         .Z(dac_clk_p_c_enable_277)) /* synthesis lut_function=((((D)+!C)+!B)+!A) */ ;
    defparam i1_4_lut_adj_229.init = 16'hff7f;
    LUT4 i20565_4_lut (.A(chg_counter[1]), .B(chg_counter[6]), .C(chg_counter[10]), 
         .D(chg_counter[4]), .Z(n22972)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i20565_4_lut.init = 16'h8000;
    LUT4 i20567_4_lut (.A(n22774), .B(n22966), .C(n22782), .D(n22780), 
         .Z(n22974)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i20567_4_lut.init = 16'h8000;
    LUT4 i20569_4_lut (.A(chg_counter[21]), .B(n22968), .C(n22940), .D(chg_counter[0]), 
         .Z(n22976)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i20569_4_lut.init = 16'h8000;
    LUT4 i1_2_lut (.A(chg_counter[16]), .B(chg_counter[3]), .Z(n22774)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i20559_4_lut (.A(chg_counter[12]), .B(chg_counter[20]), .C(chg_counter[5]), 
         .D(chg_counter[15]), .Z(n22966)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i20559_4_lut.init = 16'h8000;
    LUT4 i1_4_lut_adj_230 (.A(chg_counter[19]), .B(chg_counter[13]), .C(chg_counter[18]), 
         .D(chg_counter[2]), .Z(n22782)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_230.init = 16'h8000;
    LUT4 i1_2_lut_adj_231 (.A(chg_counter[14]), .B(chg_counter[23]), .Z(n22780)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_231.init = 16'h8888;
    LUT4 i20561_4_lut (.A(chg_counter[22]), .B(chg_counter[9]), .C(chg_counter[8]), 
         .D(chg_counter[7]), .Z(n22968)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i20561_4_lut.init = 16'h8000;
    LUT4 i20534_2_lut (.A(chg_counter[11]), .B(chg_counter[17]), .Z(n22940)) /* synthesis lut_function=(A (B)) */ ;
    defparam i20534_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_adj_232 (.A(wb_fm_ack), .B(wb_lo_ack), .Z(n4)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[12:58])
    defparam i1_2_lut_adj_232.init = 16'heeee;
    LUT4 i1_4_lut_adj_233 (.A(n29081), .B(wb_lo_sel_N_80), .C(wb_control_sel_N_78), 
         .D(n22470), .Z(none_sel)) /* synthesis lut_function=(A (B (C))+!A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(228[19:70])
    defparam i1_4_lut_adj_233.init = 16'hc080;
    LUT4 i1_4_lut_adj_234 (.A(n26), .B(wb_addr[15]), .C(wb_addr[12]), 
         .D(wb_addr[8]), .Z(n22470)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(223[20:46])
    defparam i1_4_lut_adj_234.init = 16'hfffb;
    LUT4 i1_4_lut_adj_235 (.A(n26), .B(n38), .C(n34), .D(n22816), .Z(wb_control_data_31__N_35)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut_adj_235.init = 16'h0100;
    LUT4 i1_4_lut_adj_236 (.A(wb_addr[12]), .B(wb_addr[9]), .C(n22822), 
         .D(wb_addr[8]), .Z(n22816)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_4_lut_adj_236.init = 16'h1000;
    LUT4 i1_2_lut_adj_237 (.A(wb_stb), .B(wb_addr[15]), .Z(n22822)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_237.init = 16'h8888;
    LUT4 i1_4_lut_adj_238 (.A(n29302), .B(n26), .C(wb_addr[15]), .D(n22448), 
         .Z(n22458)) /* synthesis lut_function=((B+((D)+!C))+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(223[20:46])
    defparam i1_4_lut_adj_238.init = 16'hffdf;
    LUT4 i24657_2_lut_3_lut (.A(n22458), .B(n29065), .C(n21641), .Z(dac_clk_p_c_enable_243)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(223[20:46])
    defparam i24657_2_lut_3_lut.init = 16'h0101;
    PFUMX i24923 (.BLUT(n26545), .ALUT(n26544), .C0(wb_addr[1]), .Z(n26546));
    LUT4 i1_4_lut_adj_239 (.A(n26), .B(n38), .C(n34), .D(n22828), .Z(o_dac_a_9__N_1)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut_adj_239.init = 16'h0100;
    LUT4 i1_4_lut_adj_240 (.A(wb_addr[12]), .B(wb_addr[8]), .C(n22822), 
         .D(wb_addr[9]), .Z(n22828)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_4_lut_adj_240.init = 16'h1000;
    LUT4 i1_3_lut (.A(wb_addr[9]), .B(wb_addr[12]), .C(i_sw0_c), .Z(n22448)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(223[20:46])
    defparam i1_3_lut.init = 16'hfefe;
    LUT4 i1_3_lut_4_lut (.A(wb_addr[9]), .B(n34), .C(wb_addr[8]), .D(wb_addr[15]), 
         .Z(n22808)) /* synthesis lut_function=((B+!(C (D)))+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(223[20:46])
    defparam i1_3_lut_4_lut.init = 16'hdfff;
    LUT4 i1_2_lut_rep_421_3_lut (.A(wb_addr[9]), .B(n34), .C(n38), .Z(n29081)) /* synthesis lut_function=((B+(C))+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(223[20:46])
    defparam i1_2_lut_rep_421_3_lut.init = 16'hfdfd;
    LUT4 i1_4_lut_adj_241 (.A(n22660), .B(n22662), .C(n22664), .D(n22650), 
         .Z(n38)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(223[20:46])
    defparam i1_4_lut_adj_241.init = 16'hfffe;
    LUT4 i1_2_lut_adj_242 (.A(wb_addr[27]), .B(wb_addr[14]), .Z(n22660)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(223[20:46])
    defparam i1_2_lut_adj_242.init = 16'heeee;
    LUT4 i1_4_lut_adj_243 (.A(wb_addr[17]), .B(wb_addr[11]), .C(wb_addr[23]), 
         .D(wb_addr[16]), .Z(n22662)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(223[20:46])
    defparam i1_4_lut_adj_243.init = 16'hfffe;
    LUT4 i1_4_lut_adj_244 (.A(wb_addr[25]), .B(wb_addr[24]), .C(wb_addr[26]), 
         .D(wb_addr[20]), .Z(n22664)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(223[20:46])
    defparam i1_4_lut_adj_244.init = 16'hfffe;
    LUT4 i1_2_lut_adj_245 (.A(wb_addr[19]), .B(wb_addr[18]), .Z(n22650)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(223[20:46])
    defparam i1_2_lut_adj_245.init = 16'heeee;
    LUT4 i1_4_lut_adj_246 (.A(wb_addr[28]), .B(wb_addr[13]), .C(wb_addr[10]), 
         .D(wb_addr[29]), .Z(n34)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(223[20:46])
    defparam i1_4_lut_adj_246.init = 16'hfffe;
    LUT4 lo_q_en_bdd_3_lut_24922 (.A(\addr_space[2]_adj_3701 [1]), .B(\addr_space[3]_adj_3702 [1]), 
         .C(wb_addr[0]), .Z(n26544)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam lo_q_en_bdd_3_lut_24922.init = 16'hcaca;
    LUT4 i6_2_lut (.A(wb_addr[22]), .B(wb_addr[21]), .Z(n26)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(223[20:46])
    defparam i6_2_lut.init = 16'heeee;
    LUT4 i1_2_lut_rep_642 (.A(wb_stb), .B(wb_we), .Z(n29302)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(207[17:41])
    defparam i1_2_lut_rep_642.init = 16'h8888;
    LUT4 lo_q_en_bdd_3_lut_25687 (.A(lo_q_en), .B(\addr_space[1]_adj_3700 [1]), 
         .C(wb_addr[0]), .Z(n26545)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam lo_q_en_bdd_3_lut_25687.init = 16'hcaca;
    LUT4 i1_3_lut_rep_405 (.A(wb_addr[8]), .B(n38), .C(n34), .Z(n29065)) /* synthesis lut_function=((B+(C))+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(223[20:46])
    defparam i1_3_lut_rep_405.init = 16'hfdfd;
    LUT4 i1_2_lut_4_lut (.A(wb_addr[8]), .B(n38), .C(n34), .D(n22526), 
         .Z(wb_control_sel_N_78)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(223[20:46])
    defparam i1_2_lut_4_lut.init = 16'hfffd;
    LUT4 lo_i_en_bdd_3_lut_24948 (.A(\addr_space[2]_adj_3701 [0]), .B(\addr_space[3]_adj_3702 [0]), 
         .C(wb_addr[0]), .Z(n26568)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam lo_i_en_bdd_3_lut_24948.init = 16'hcaca;
    LUT4 lo_i_en_bdd_3_lut (.A(lo_i_en), .B(\addr_space[1]_adj_3700 [0]), 
         .C(wb_addr[0]), .Z(n26569)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam lo_i_en_bdd_3_lut.init = 16'hcaca;
    LUT4 i11772_1_lut (.A(wb_idata[1]), .Z(n14148)) /* synthesis lut_function=(!(A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(246[8] 254[52])
    defparam i11772_1_lut.init = 16'h5555;
    LUT4 i24689_3_lut_4_lut (.A(n29302), .B(n22470), .C(n29081), .D(n29155), 
         .Z(dac_clk_p_c_enable_502)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(223[20:46])
    defparam i24689_3_lut_4_lut.init = 16'h0002;
    LUT4 i24680_2_lut_3_lut_4_lut (.A(n29302), .B(n22470), .C(n29199), 
         .D(n29081), .Z(dac_clk_p_c_enable_407)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(223[20:46])
    defparam i24680_2_lut_3_lut_4_lut.init = 16'h0002;
    LUT4 i24677_2_lut_3_lut_4_lut (.A(n29302), .B(n22470), .C(n21641), 
         .D(n29081), .Z(dac_clk_p_c_enable_439)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(223[20:46])
    defparam i24677_2_lut_3_lut_4_lut.init = 16'h0002;
    LUT4 i24674_2_lut_3_lut_4_lut (.A(n29302), .B(n22470), .C(n29197), 
         .D(n29081), .Z(dac_clk_p_c_enable_471)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(223[20:46])
    defparam i24674_2_lut_3_lut_4_lut.init = 16'h0002;
    LUT4 i24683_3_lut_4_lut (.A(n29302), .B(n22470), .C(n29081), .D(n21662), 
         .Z(dac_clk_p_c_enable_375)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(223[20:46])
    defparam i24683_3_lut_4_lut.init = 16'h0002;
    LUT4 wb_idata_31__I_0_i32_4_lut (.A(wb_control_data[31]), .B(wb_fm_data[31]), 
         .C(wb_fm_ack), .D(wb_control_ack), .Z(wb_idata_31__N_2[31])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(249[7] 254[52])
    defparam wb_idata_31__I_0_i32_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i31_4_lut (.A(wb_control_data[30]), .B(wb_fm_data[30]), 
         .C(wb_fm_ack), .D(wb_control_ack), .Z(wb_idata_31__N_2[30])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(249[7] 254[52])
    defparam wb_idata_31__I_0_i31_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i1_3_lut (.A(wb_idata_31__N_36[0]), .B(wb_fm_data[0]), 
         .C(wb_fm_ack), .Z(wb_idata_31__N_2[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(249[7] 254[52])
    defparam wb_idata_31__I_0_i1_3_lut.init = 16'hcaca;
    LUT4 mux_30_i1_4_lut (.A(wb_lo_data[0]), .B(wb_control_data[0]), .C(wb_control_ack), 
         .D(wb_lo_ack), .Z(wb_idata_31__N_36[0])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(251[7] 254[52])
    defparam mux_30_i1_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i30_4_lut (.A(wb_control_data[29]), .B(wb_fm_data[29]), 
         .C(wb_fm_ack), .D(wb_control_ack), .Z(wb_idata_31__N_2[29])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(249[7] 254[52])
    defparam wb_idata_31__I_0_i30_4_lut.init = 16'hcac0;
    LUT4 dac_clk_p_I_0_1_lut (.A(dac_clk_p_c), .Z(dac_clk_n_c)) /* synthesis lut_function=(!(A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(54[20:30])
    defparam dac_clk_p_I_0_1_lut.init = 16'h5555;
    hbbus genbus (.dac_clk_p_c(dac_clk_p_c), .wb_cyc(wb_cyc), .wb_we(wb_we), 
          .wb_odata({wb_odata}), .wb_stb(wb_stb), .wb_addr({wb_addr}), 
          .GND_net(GND_net), .wb_ack(wb_ack), .\wb_idata[0] (wb_idata[0]), 
          .\wb_idata[2] (wb_idata[2]), .\wb_idata[3] (wb_idata[3]), .\wb_idata[4] (wb_idata[4]), 
          .\wb_idata[5] (wb_idata[5]), .\wb_idata[6] (wb_idata[6]), .\wb_idata[7] (wb_idata[7]), 
          .\wb_idata[8] (wb_idata[8]), .\wb_idata[9] (wb_idata[9]), .\wb_idata[10] (wb_idata[10]), 
          .\wb_idata[11] (wb_idata[11]), .\wb_idata[12] (wb_idata[12]), 
          .\wb_idata[13] (wb_idata[13]), .\wb_idata[14] (wb_idata[14]), 
          .\wb_idata[15] (wb_idata[15]), .\wb_idata[16] (wb_idata[16]), 
          .\wb_idata[17] (wb_idata[17]), .\wb_idata[18] (wb_idata[18]), 
          .\wb_idata[19] (wb_idata[19]), .\wb_idata[20] (wb_idata[20]), 
          .\wb_idata[21] (wb_idata[21]), .\wb_idata[22] (wb_idata[22]), 
          .\wb_idata[23] (wb_idata[23]), .\wb_idata[24] (wb_idata[24]), 
          .\wb_idata[25] (wb_idata[25]), .\wb_idata[26] (wb_idata[26]), 
          .\wb_idata[27] (wb_idata[27]), .\wb_idata[28] (wb_idata[28]), 
          .wb_err(wb_err), .\wb_idata[29] (wb_idata[29]), .\wb_idata[30] (wb_idata[30]), 
          .\wb_idata[31] (wb_idata[31]), .n2(n2), .n14148(n14148), .n32067(n32067), 
          .VCC_net(VCC_net), .\rx_data[1] (rx_data[1]), .\rx_data[2] (rx_data[2]), 
          .\rx_data[0] (rx_data[0]), .\rx_data[3] (rx_data[3]), .\rx_data[5] (rx_data[5]), 
          .\rx_data[6] (rx_data[6]), .\rx_data[4] (rx_data[4]), .rx_stb(rx_stb), 
          .\tx_data[1] (tx_data[1]), .\tx_data[2] (tx_data[2]), .\tx_data[3] (tx_data[3]), 
          .\tx_data[4] (tx_data[4]), .\tx_data[5] (tx_data[5]), .\tx_data[6] (tx_data[6]), 
          .tx_stb(tx_stb), .\tx_data[0] (tx_data[0]), .tx_busy(tx_busy)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(84[7] 100[22])
    LUT4 wb_idata_31__I_0_i11_4_lut (.A(wb_control_data[10]), .B(wb_fm_data[10]), 
         .C(wb_fm_ack), .D(wb_control_ack), .Z(wb_idata_31__N_2[10])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(249[7] 254[52])
    defparam wb_idata_31__I_0_i11_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i29_4_lut (.A(wb_control_data[28]), .B(wb_fm_data[28]), 
         .C(wb_fm_ack), .D(wb_control_ack), .Z(wb_idata_31__N_2[28])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(249[7] 254[52])
    defparam wb_idata_31__I_0_i29_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i10_4_lut (.A(wb_control_data[9]), .B(wb_fm_data[9]), 
         .C(wb_fm_ack), .D(wb_control_ack), .Z(wb_idata_31__N_2[9])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(249[7] 254[52])
    defparam wb_idata_31__I_0_i10_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i28_4_lut (.A(wb_control_data[27]), .B(wb_fm_data[27]), 
         .C(wb_fm_ack), .D(wb_control_ack), .Z(wb_idata_31__N_2[27])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(249[7] 254[52])
    defparam wb_idata_31__I_0_i28_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i9_4_lut (.A(wb_control_data[8]), .B(wb_fm_data[8]), 
         .C(wb_fm_ack), .D(wb_control_ack), .Z(wb_idata_31__N_2[8])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(249[7] 254[52])
    defparam wb_idata_31__I_0_i9_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i27_4_lut (.A(wb_control_data[26]), .B(wb_fm_data[26]), 
         .C(wb_fm_ack), .D(wb_control_ack), .Z(wb_idata_31__N_2[26])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(249[7] 254[52])
    defparam wb_idata_31__I_0_i27_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i8_3_lut (.A(wb_idata_31__N_36[7]), .B(wb_fm_data[7]), 
         .C(wb_fm_ack), .Z(wb_idata_31__N_2[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(249[7] 254[52])
    defparam wb_idata_31__I_0_i8_3_lut.init = 16'hcaca;
    LUT4 mux_30_i8_4_lut (.A(wb_lo_data[7]), .B(wb_control_data[7]), .C(wb_control_ack), 
         .D(wb_lo_ack), .Z(wb_idata_31__N_36[7])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(251[7] 254[52])
    defparam mux_30_i8_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i26_4_lut (.A(wb_control_data[25]), .B(wb_fm_data[25]), 
         .C(wb_fm_ack), .D(wb_control_ack), .Z(wb_idata_31__N_2[25])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(249[7] 254[52])
    defparam wb_idata_31__I_0_i26_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i7_3_lut (.A(wb_idata_31__N_36[6]), .B(wb_fm_data[6]), 
         .C(wb_fm_ack), .Z(wb_idata_31__N_2[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(249[7] 254[52])
    defparam wb_idata_31__I_0_i7_3_lut.init = 16'hcaca;
    LUT4 mux_30_i7_4_lut (.A(wb_lo_data[6]), .B(wb_control_data[6]), .C(wb_control_ack), 
         .D(wb_lo_ack), .Z(wb_idata_31__N_36[6])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(251[7] 254[52])
    defparam mux_30_i7_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i25_4_lut (.A(wb_control_data[24]), .B(wb_fm_data[24]), 
         .C(wb_fm_ack), .D(wb_control_ack), .Z(wb_idata_31__N_2[24])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(249[7] 254[52])
    defparam wb_idata_31__I_0_i25_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i6_3_lut (.A(wb_idata_31__N_36[5]), .B(wb_fm_data[5]), 
         .C(wb_fm_ack), .Z(wb_idata_31__N_2[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(249[7] 254[52])
    defparam wb_idata_31__I_0_i6_3_lut.init = 16'hcaca;
    LUT4 mux_30_i6_4_lut (.A(wb_lo_data[5]), .B(wb_control_data[5]), .C(wb_control_ack), 
         .D(wb_lo_ack), .Z(wb_idata_31__N_36[5])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(251[7] 254[52])
    defparam mux_30_i6_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i24_4_lut (.A(wb_control_data[23]), .B(wb_fm_data[23]), 
         .C(wb_fm_ack), .D(wb_control_ack), .Z(wb_idata_31__N_2[23])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(249[7] 254[52])
    defparam wb_idata_31__I_0_i24_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i5_3_lut (.A(wb_idata_31__N_36[4]), .B(wb_fm_data[4]), 
         .C(wb_fm_ack), .Z(wb_idata_31__N_2[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(249[7] 254[52])
    defparam wb_idata_31__I_0_i5_3_lut.init = 16'hcaca;
    LUT4 mux_30_i5_4_lut (.A(wb_lo_data[4]), .B(wb_control_data[4]), .C(wb_control_ack), 
         .D(wb_lo_ack), .Z(wb_idata_31__N_36[4])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(251[7] 254[52])
    defparam mux_30_i5_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i23_4_lut (.A(wb_control_data[22]), .B(wb_fm_data[22]), 
         .C(wb_fm_ack), .D(wb_control_ack), .Z(wb_idata_31__N_2[22])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(249[7] 254[52])
    defparam wb_idata_31__I_0_i23_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i4_3_lut (.A(wb_idata_31__N_36[3]), .B(wb_fm_data[3]), 
         .C(wb_fm_ack), .Z(wb_idata_31__N_2[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(249[7] 254[52])
    defparam wb_idata_31__I_0_i4_3_lut.init = 16'hcaca;
    LUT4 mux_30_i4_4_lut (.A(wb_lo_data[3]), .B(wb_control_data[3]), .C(wb_control_ack), 
         .D(wb_lo_ack), .Z(wb_idata_31__N_36[3])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(251[7] 254[52])
    defparam mux_30_i4_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i22_4_lut (.A(wb_control_data[21]), .B(wb_fm_data[21]), 
         .C(wb_fm_ack), .D(wb_control_ack), .Z(wb_idata_31__N_2[21])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(249[7] 254[52])
    defparam wb_idata_31__I_0_i22_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i3_3_lut (.A(wb_idata_31__N_36[2]), .B(wb_fm_data[2]), 
         .C(wb_fm_ack), .Z(wb_idata_31__N_2[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(249[7] 254[52])
    defparam wb_idata_31__I_0_i3_3_lut.init = 16'hcaca;
    LUT4 mux_30_i3_4_lut (.A(wb_lo_data[2]), .B(wb_control_data[2]), .C(wb_control_ack), 
         .D(wb_lo_ack), .Z(wb_idata_31__N_36[2])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(251[7] 254[52])
    defparam mux_30_i3_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i21_4_lut (.A(wb_control_data[20]), .B(wb_fm_data[20]), 
         .C(wb_fm_ack), .D(wb_control_ack), .Z(wb_idata_31__N_2[20])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(249[7] 254[52])
    defparam wb_idata_31__I_0_i21_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i2_3_lut (.A(wb_idata_31__N_36[1]), .B(wb_fm_data[1]), 
         .C(wb_fm_ack), .Z(wb_idata_31__N_2[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(249[7] 254[52])
    defparam wb_idata_31__I_0_i2_3_lut.init = 16'hcaca;
    LUT4 mux_30_i2_4_lut (.A(wb_lo_data[1]), .B(wb_control_data[1]), .C(wb_control_ack), 
         .D(wb_lo_ack), .Z(wb_idata_31__N_36[1])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(251[7] 254[52])
    defparam mux_30_i2_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i20_4_lut (.A(wb_control_data[19]), .B(wb_fm_data[19]), 
         .C(wb_fm_ack), .D(wb_control_ack), .Z(wb_idata_31__N_2[19])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(249[7] 254[52])
    defparam wb_idata_31__I_0_i20_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i19_4_lut (.A(wb_control_data[18]), .B(wb_fm_data[18]), 
         .C(wb_fm_ack), .D(wb_control_ack), .Z(wb_idata_31__N_2[18])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(249[7] 254[52])
    defparam wb_idata_31__I_0_i19_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i18_4_lut (.A(wb_control_data[17]), .B(wb_fm_data[17]), 
         .C(wb_fm_ack), .D(wb_control_ack), .Z(wb_idata_31__N_2[17])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(249[7] 254[52])
    defparam wb_idata_31__I_0_i18_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i17_4_lut (.A(wb_control_data[16]), .B(wb_fm_data[16]), 
         .C(wb_fm_ack), .D(wb_control_ack), .Z(wb_idata_31__N_2[16])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(249[7] 254[52])
    defparam wb_idata_31__I_0_i17_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i16_4_lut (.A(wb_control_data[15]), .B(wb_fm_data[15]), 
         .C(wb_fm_ack), .D(wb_control_ack), .Z(wb_idata_31__N_2[15])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(249[7] 254[52])
    defparam wb_idata_31__I_0_i16_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i15_4_lut (.A(wb_control_data[14]), .B(wb_fm_data[14]), 
         .C(wb_fm_ack), .D(wb_control_ack), .Z(wb_idata_31__N_2[14])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(249[7] 254[52])
    defparam wb_idata_31__I_0_i15_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i14_4_lut (.A(wb_control_data[13]), .B(wb_fm_data[13]), 
         .C(wb_fm_ack), .D(wb_control_ack), .Z(wb_idata_31__N_2[13])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(249[7] 254[52])
    defparam wb_idata_31__I_0_i14_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i13_4_lut (.A(wb_control_data[12]), .B(wb_fm_data[12]), 
         .C(wb_fm_ack), .D(wb_control_ack), .Z(wb_idata_31__N_2[12])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(249[7] 254[52])
    defparam wb_idata_31__I_0_i13_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i12_4_lut (.A(wb_control_data[11]), .B(wb_fm_data[11]), 
         .C(wb_fm_ack), .D(wb_control_ack), .Z(wb_idata_31__N_2[11])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(249[7] 254[52])
    defparam wb_idata_31__I_0_i12_4_lut.init = 16'hcac0;
    LUT4 n26546_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4]_adj_3703 [1]), 
         .C(wb_addr[2]), .D(n26546), .Z(o_wb_data_31__N_2456[1])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n26546_bdd_3_lut_4_lut.init = 16'h8f80;
    VLO i1 (.Z(GND_net));
    TSALL TSALL_INST (.TSALL(GND_net));
    efb_inst efb_inst_0 (.dac_clk_p_c(dac_clk_p_c), .i_sw0_c(i_sw0_c), .wb_cyc(wb_cyc), 
            .wb_lo_data_7__N_34(wb_lo_data_7__N_34), .wb_we(wb_we), .\wb_addr[7] (wb_addr[7]), 
            .\wb_addr[6] (wb_addr[6]), .\wb_addr[5] (wb_addr[5]), .\wb_addr[4] (wb_addr[4]), 
            .\wb_addr[3] (wb_addr[3]), .\wb_addr[2] (wb_addr[2]), .\wb_addr[1] (wb_addr[1]), 
            .\wb_addr[0] (wb_addr[0]), .\wb_odata[7] (wb_odata[7]), .\wb_odata[6] (wb_odata[6]), 
            .\wb_odata[5] (wb_odata[5]), .\wb_odata[4] (wb_odata[4]), .\wb_odata[3] (wb_odata[3]), 
            .\wb_odata[2] (wb_odata[2]), .\wb_odata[1] (wb_odata[1]), .\wb_odata[0] (wb_odata[0]), 
            .pll_data_o({pll_data_o}), .pll_ack(pll_ack), .wb_lo_data({wb_lo_data}), 
            .wb_lo_ack(wb_lo_ack), .pll_clk(pll_clk), .pll_rst(pll_rst), 
            .pll_stb(pll_stb), .pll_we(pll_we), .pll_addr({pll_addr}), 
            .pll_data_i({pll_data_i}), .GND_net(GND_net), .VCC_net(VCC_net)) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(183[11] 195[4])
    sys_clk sys_clk_inst (.i_ref_clk_c(i_ref_clk_c), .dac_clk_p_c(dac_clk_p_c), 
            .GND_net(GND_net)) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(47[10:54])
    OB o_dac_a_pad_6 (.I(o_dac_a_c_6), .O(o_dac_a[6]));   // d:/documents/git_local/fm_modulator/rtl/top.v(33[38:45])
    dynamic_pll lo_gen (.i_ref_clk_c(i_ref_clk_c), .pll_clk(pll_clk), .pll_rst(pll_rst), 
            .pll_stb(pll_stb), .pll_we(pll_we), .pll_data_i({pll_data_i}), 
            .pll_addr({pll_addr}), .lo_q(lo_q), .pll_data_o({pll_data_o}), 
            .pll_ack(pll_ack), .GND_net(GND_net), .lo_i_en(lo_i_en), .o_lo_i_c(o_lo_i_c)) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(169[14] 181[5])
    LUT4 m1_lut (.Z(n32067)) /* synthesis lut_function=1, syn_instantiated=1 */ ;
    defparam m1_lut.init = 16'hffff;
    FD1S3AX wb_idata_i31 (.D(wb_idata_31__N_2[31]), .CK(dac_clk_p_c), .Q(wb_idata[31]));   // d:/documents/git_local/fm_modulator/rtl/top.v(246[8] 254[52])
    defparam wb_idata_i31.GSR = "DISABLED";
    FD1S3AX wb_idata_i30 (.D(wb_idata_31__N_2[30]), .CK(dac_clk_p_c), .Q(wb_idata[30]));   // d:/documents/git_local/fm_modulator/rtl/top.v(246[8] 254[52])
    defparam wb_idata_i30.GSR = "DISABLED";
    fm_generator_wb_slave fm_generator_wb_instance (.o_dac_b_c_0(o_dac_b_c_0), 
            .dac_clk_p_c(dac_clk_p_c), .wb_fm_data({wb_fm_data}), .i_sw0_c(i_sw0_c), 
            .o_dac_a_c_0(o_dac_a_c_0), .GND_net(GND_net), .\wb_addr[0] (wb_addr[0]), 
            .n29300(n29300), .\wb_addr[2] (wb_addr[2]), .\wb_addr[1] (wb_addr[1]), 
            .wb_fm_ack(wb_fm_ack), .o_dac_a_9__N_1(o_dac_a_9__N_1), .dac_clk_p_c_enable_502(dac_clk_p_c_enable_502), 
            .wb_odata({wb_odata}), .n21641(n21641), .n29065(n29065), .n22458(n22458), 
            .dac_clk_p_c_enable_227(dac_clk_p_c_enable_227), .o_dac_a_c_9(o_dac_a_c_9), 
            .dac_clk_p_c_enable_241(dac_clk_p_c_enable_241), .dac_clk_p_c_enable_106(dac_clk_p_c_enable_106), 
            .o_dac_a_c_8(o_dac_a_c_8), .o_dac_a_c_7(o_dac_a_c_7), .o_dac_a_c_6(o_dac_a_c_6), 
            .o_dac_a_c_5(o_dac_a_c_5), .o_dac_a_c_4(o_dac_a_c_4), .o_dac_a_c_3(o_dac_a_c_3), 
            .o_dac_a_c_2(o_dac_a_c_2), .o_dac_a_c_1(o_dac_a_c_1), .o_dac_b_c_9(o_dac_b_c_9), 
            .o_dac_b_c_8(o_dac_b_c_8), .o_dac_b_c_7(o_dac_b_c_7), .o_dac_b_c_6(o_dac_b_c_6), 
            .o_dac_b_c_5(o_dac_b_c_5), .o_dac_b_c_4(o_dac_b_c_4), .o_dac_b_c_3(o_dac_b_c_3), 
            .o_dac_b_c_2(o_dac_b_c_2), .o_dac_b_c_1(o_dac_b_c_1), .dac_clk_p_c_enable_375(dac_clk_p_c_enable_375), 
            .dac_clk_p_c_enable_407(dac_clk_p_c_enable_407), .dac_clk_p_c_enable_439(dac_clk_p_c_enable_439), 
            .dac_clk_p_c_enable_471(dac_clk_p_c_enable_471), .n21662(n21662), 
            .n29155(n29155), .n29197(n29197), .n29199(n29199), .o_dac_cw_b_c(o_dac_cw_b_c), 
            .n32067(n32067), .n32066(n32066)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(122[2] 134[2])
    LUT4 m0_lut (.Z(n32066)) /* synthesis lut_function=0, syn_instantiated=1 */ ;
    defparam m0_lut.init = 16'h0000;
    \txuartlite(TIMING_BITS=24,CLOCKS_PER_BAUD=10000)  txtransport (.dac_clk_p_c(dac_clk_p_c), 
            .o_wbu_uart_tx_c(o_wbu_uart_tx_c), .GND_net(GND_net), .tx_stb(tx_stb), 
            .tx_busy(tx_busy), .\tx_data[0] (tx_data[0]), .\tx_data[6] (tx_data[6]), 
            .\tx_data[5] (tx_data[5]), .\tx_data[4] (tx_data[4]), .\tx_data[3] (tx_data[3]), 
            .\tx_data[2] (tx_data[2]), .\tx_data[1] (tx_data[1]), .n32067(n32067)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(69[58:115])
    FD1S3AX wb_idata_i0 (.D(wb_idata_31__N_2[0]), .CK(dac_clk_p_c), .Q(wb_idata[0]));   // d:/documents/git_local/fm_modulator/rtl/top.v(246[8] 254[52])
    defparam wb_idata_i0.GSR = "DISABLED";
    FD1S3AX wb_idata_i29 (.D(wb_idata_31__N_2[29]), .CK(dac_clk_p_c), .Q(wb_idata[29]));   // d:/documents/git_local/fm_modulator/rtl/top.v(246[8] 254[52])
    defparam wb_idata_i29.GSR = "DISABLED";
    OB o_dac_a_pad_5 (.I(o_dac_a_c_5), .O(o_dac_a[5]));   // d:/documents/git_local/fm_modulator/rtl/top.v(33[38:45])
    OB o_dac_a_pad_4 (.I(o_dac_a_c_4), .O(o_dac_a[4]));   // d:/documents/git_local/fm_modulator/rtl/top.v(33[38:45])
    OB o_dac_a_pad_3 (.I(o_dac_a_c_3), .O(o_dac_a[3]));   // d:/documents/git_local/fm_modulator/rtl/top.v(33[38:45])
    OB o_dac_a_pad_2 (.I(o_dac_a_c_2), .O(o_dac_a[2]));   // d:/documents/git_local/fm_modulator/rtl/top.v(33[38:45])
    OB o_dac_a_pad_1 (.I(o_dac_a_c_1), .O(o_dac_a[1]));   // d:/documents/git_local/fm_modulator/rtl/top.v(33[38:45])
    OB o_dac_a_pad_0 (.I(o_dac_a_c_0), .O(o_dac_a[0]));   // d:/documents/git_local/fm_modulator/rtl/top.v(33[38:45])
    OB o_dac_b_pad_9 (.I(o_dac_b_c_9), .O(o_dac_b[9]));   // d:/documents/git_local/fm_modulator/rtl/top.v(33[47:54])
    OB o_dac_b_pad_8 (.I(o_dac_b_c_8), .O(o_dac_b[8]));   // d:/documents/git_local/fm_modulator/rtl/top.v(33[47:54])
    OB o_dac_b_pad_7 (.I(o_dac_b_c_7), .O(o_dac_b[7]));   // d:/documents/git_local/fm_modulator/rtl/top.v(33[47:54])
    OB o_dac_b_pad_6 (.I(o_dac_b_c_6), .O(o_dac_b[6]));   // d:/documents/git_local/fm_modulator/rtl/top.v(33[47:54])
    OB o_dac_b_pad_5 (.I(o_dac_b_c_5), .O(o_dac_b[5]));   // d:/documents/git_local/fm_modulator/rtl/top.v(33[47:54])
    OB o_dac_b_pad_4 (.I(o_dac_b_c_4), .O(o_dac_b[4]));   // d:/documents/git_local/fm_modulator/rtl/top.v(33[47:54])
    OB o_dac_b_pad_3 (.I(o_dac_b_c_3), .O(o_dac_b[3]));   // d:/documents/git_local/fm_modulator/rtl/top.v(33[47:54])
    OB o_dac_b_pad_2 (.I(o_dac_b_c_2), .O(o_dac_b[2]));   // d:/documents/git_local/fm_modulator/rtl/top.v(33[47:54])
    OB o_dac_b_pad_1 (.I(o_dac_b_c_1), .O(o_dac_b[1]));   // d:/documents/git_local/fm_modulator/rtl/top.v(33[47:54])
    OB o_dac_b_pad_0 (.I(o_dac_b_c_0), .O(o_dac_b[0]));   // d:/documents/git_local/fm_modulator/rtl/top.v(33[47:54])
    OB dac_clk_p_pad (.I(dac_clk_p_c), .O(dac_clk_p));   // d:/documents/git_local/fm_modulator/rtl/top.v(34[29:38])
    OB dac_clk_n_pad (.I(dac_clk_n_c), .O(dac_clk_n));   // d:/documents/git_local/fm_modulator/rtl/top.v(34[40:49])
    OB o_dac_cw_b_pad (.I(o_dac_cw_b_c), .O(o_dac_cw_b));   // d:/documents/git_local/fm_modulator/rtl/top.v(34[51:61])
    OB o_lo_i_pad (.I(o_lo_i_c), .O(o_lo_i));   // d:/documents/git_local/fm_modulator/rtl/top.v(34[13:19])
    OB o_lo_q_pad (.I(o_lo_q_c), .O(o_lo_q));   // d:/documents/git_local/fm_modulator/rtl/top.v(34[21:27])
    IB i_ref_clk_pad (.I(i_ref_clk), .O(i_ref_clk_c));   // d:/documents/git_local/fm_modulator/rtl/top.v(26[12:21])
    IB i_wbu_uart_rx_pad (.I(i_wbu_uart_rx), .O(i_wbu_uart_rx_c));   // d:/documents/git_local/fm_modulator/rtl/top.v(28[12:25])
    IB i_sw0_pad (.I(i_sw0), .O(i_sw0_c));   // d:/documents/git_local/fm_modulator/rtl/top.v(31[12:17])
    FD1S3AX wb_idata_i10 (.D(wb_idata_31__N_2[10]), .CK(dac_clk_p_c), .Q(wb_idata[10]));   // d:/documents/git_local/fm_modulator/rtl/top.v(246[8] 254[52])
    defparam wb_idata_i10.GSR = "DISABLED";
    FD1S3AX wb_idata_i28 (.D(wb_idata_31__N_2[28]), .CK(dac_clk_p_c), .Q(wb_idata[28]));   // d:/documents/git_local/fm_modulator/rtl/top.v(246[8] 254[52])
    defparam wb_idata_i28.GSR = "DISABLED";
    FD1S3AX wb_idata_i9 (.D(wb_idata_31__N_2[9]), .CK(dac_clk_p_c), .Q(wb_idata[9]));   // d:/documents/git_local/fm_modulator/rtl/top.v(246[8] 254[52])
    defparam wb_idata_i9.GSR = "DISABLED";
    FD1S3AX wb_idata_i27 (.D(wb_idata_31__N_2[27]), .CK(dac_clk_p_c), .Q(wb_idata[27]));   // d:/documents/git_local/fm_modulator/rtl/top.v(246[8] 254[52])
    defparam wb_idata_i27.GSR = "DISABLED";
    FD1S3AX wb_idata_i8 (.D(wb_idata_31__N_2[8]), .CK(dac_clk_p_c), .Q(wb_idata[8]));   // d:/documents/git_local/fm_modulator/rtl/top.v(246[8] 254[52])
    defparam wb_idata_i8.GSR = "DISABLED";
    FD1S3AX wb_idata_i26 (.D(wb_idata_31__N_2[26]), .CK(dac_clk_p_c), .Q(wb_idata[26]));   // d:/documents/git_local/fm_modulator/rtl/top.v(246[8] 254[52])
    defparam wb_idata_i26.GSR = "DISABLED";
    FD1S3AX wb_idata_i7 (.D(wb_idata_31__N_2[7]), .CK(dac_clk_p_c), .Q(wb_idata[7]));   // d:/documents/git_local/fm_modulator/rtl/top.v(246[8] 254[52])
    defparam wb_idata_i7.GSR = "DISABLED";
    FD1S3AX wb_idata_i25 (.D(wb_idata_31__N_2[25]), .CK(dac_clk_p_c), .Q(wb_idata[25]));   // d:/documents/git_local/fm_modulator/rtl/top.v(246[8] 254[52])
    defparam wb_idata_i25.GSR = "DISABLED";
    FD1S3AX wb_idata_i6 (.D(wb_idata_31__N_2[6]), .CK(dac_clk_p_c), .Q(wb_idata[6]));   // d:/documents/git_local/fm_modulator/rtl/top.v(246[8] 254[52])
    defparam wb_idata_i6.GSR = "DISABLED";
    FD1S3AX wb_idata_i24 (.D(wb_idata_31__N_2[24]), .CK(dac_clk_p_c), .Q(wb_idata[24]));   // d:/documents/git_local/fm_modulator/rtl/top.v(246[8] 254[52])
    defparam wb_idata_i24.GSR = "DISABLED";
    FD1S3AX wb_idata_i5 (.D(wb_idata_31__N_2[5]), .CK(dac_clk_p_c), .Q(wb_idata[5]));   // d:/documents/git_local/fm_modulator/rtl/top.v(246[8] 254[52])
    defparam wb_idata_i5.GSR = "DISABLED";
    FD1S3AX wb_idata_i23 (.D(wb_idata_31__N_2[23]), .CK(dac_clk_p_c), .Q(wb_idata[23]));   // d:/documents/git_local/fm_modulator/rtl/top.v(246[8] 254[52])
    defparam wb_idata_i23.GSR = "DISABLED";
    FD1S3AX wb_idata_i4 (.D(wb_idata_31__N_2[4]), .CK(dac_clk_p_c), .Q(wb_idata[4]));   // d:/documents/git_local/fm_modulator/rtl/top.v(246[8] 254[52])
    defparam wb_idata_i4.GSR = "DISABLED";
    FD1S3AX wb_idata_i22 (.D(wb_idata_31__N_2[22]), .CK(dac_clk_p_c), .Q(wb_idata[22]));   // d:/documents/git_local/fm_modulator/rtl/top.v(246[8] 254[52])
    defparam wb_idata_i22.GSR = "DISABLED";
    FD1S3AX wb_idata_i3 (.D(wb_idata_31__N_2[3]), .CK(dac_clk_p_c), .Q(wb_idata[3]));   // d:/documents/git_local/fm_modulator/rtl/top.v(246[8] 254[52])
    defparam wb_idata_i3.GSR = "DISABLED";
    FD1S3AX wb_idata_i21 (.D(wb_idata_31__N_2[21]), .CK(dac_clk_p_c), .Q(wb_idata[21]));   // d:/documents/git_local/fm_modulator/rtl/top.v(246[8] 254[52])
    defparam wb_idata_i21.GSR = "DISABLED";
    FD1S3AX wb_idata_i2 (.D(wb_idata_31__N_2[2]), .CK(dac_clk_p_c), .Q(wb_idata[2]));   // d:/documents/git_local/fm_modulator/rtl/top.v(246[8] 254[52])
    defparam wb_idata_i2.GSR = "DISABLED";
    FD1S3AX wb_idata_i20 (.D(wb_idata_31__N_2[20]), .CK(dac_clk_p_c), .Q(wb_idata[20]));   // d:/documents/git_local/fm_modulator/rtl/top.v(246[8] 254[52])
    defparam wb_idata_i20.GSR = "DISABLED";
    FD1S3AX wb_idata_i1 (.D(wb_idata_31__N_2[1]), .CK(dac_clk_p_c), .Q(wb_idata[1]));   // d:/documents/git_local/fm_modulator/rtl/top.v(246[8] 254[52])
    defparam wb_idata_i1.GSR = "DISABLED";
    FD1S3AX wb_idata_i19 (.D(wb_idata_31__N_2[19]), .CK(dac_clk_p_c), .Q(wb_idata[19]));   // d:/documents/git_local/fm_modulator/rtl/top.v(246[8] 254[52])
    defparam wb_idata_i19.GSR = "DISABLED";
    FD1S3AX wb_idata_i18 (.D(wb_idata_31__N_2[18]), .CK(dac_clk_p_c), .Q(wb_idata[18]));   // d:/documents/git_local/fm_modulator/rtl/top.v(246[8] 254[52])
    defparam wb_idata_i18.GSR = "DISABLED";
    FD1S3AX wb_idata_i17 (.D(wb_idata_31__N_2[17]), .CK(dac_clk_p_c), .Q(wb_idata[17]));   // d:/documents/git_local/fm_modulator/rtl/top.v(246[8] 254[52])
    defparam wb_idata_i17.GSR = "DISABLED";
    FD1S3AX wb_idata_i16 (.D(wb_idata_31__N_2[16]), .CK(dac_clk_p_c), .Q(wb_idata[16]));   // d:/documents/git_local/fm_modulator/rtl/top.v(246[8] 254[52])
    defparam wb_idata_i16.GSR = "DISABLED";
    FD1S3AX wb_idata_i15 (.D(wb_idata_31__N_2[15]), .CK(dac_clk_p_c), .Q(wb_idata[15]));   // d:/documents/git_local/fm_modulator/rtl/top.v(246[8] 254[52])
    defparam wb_idata_i15.GSR = "DISABLED";
    FD1S3AX wb_idata_i14 (.D(wb_idata_31__N_2[14]), .CK(dac_clk_p_c), .Q(wb_idata[14]));   // d:/documents/git_local/fm_modulator/rtl/top.v(246[8] 254[52])
    defparam wb_idata_i14.GSR = "DISABLED";
    FD1S3AX wb_idata_i13 (.D(wb_idata_31__N_2[13]), .CK(dac_clk_p_c), .Q(wb_idata[13]));   // d:/documents/git_local/fm_modulator/rtl/top.v(246[8] 254[52])
    defparam wb_idata_i13.GSR = "DISABLED";
    FD1S3AX wb_idata_i12 (.D(wb_idata_31__N_2[12]), .CK(dac_clk_p_c), .Q(wb_idata[12]));   // d:/documents/git_local/fm_modulator/rtl/top.v(246[8] 254[52])
    defparam wb_idata_i12.GSR = "DISABLED";
    FD1S3AX wb_idata_i11 (.D(wb_idata_31__N_2[11]), .CK(dac_clk_p_c), .Q(wb_idata[11]));   // d:/documents/git_local/fm_modulator/rtl/top.v(246[8] 254[52])
    defparam wb_idata_i11.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module \rxuartlite(CLOCKS_PER_BAUD=10000) 
//

module \rxuartlite(CLOCKS_PER_BAUD=10000)  (\rx_data[0] , dac_clk_p_c, rx_stb, 
            i_wbu_uart_rx_c, chg_counter, dac_clk_p_c_enable_277, chg_counter_23__N_173, 
            GND_net, \rx_data[6] , \rx_data[5] , \rx_data[4] , \rx_data[3] , 
            \rx_data[2] , \rx_data[1] ) /* synthesis syn_module_defined=1 */ ;
    output \rx_data[0] ;
    input dac_clk_p_c;
    output rx_stb;
    input i_wbu_uart_rx_c;
    output [23:0]chg_counter;
    input dac_clk_p_c_enable_277;
    output chg_counter_23__N_173;
    input GND_net;
    output \rx_data[6] ;
    output \rx_data[5] ;
    output \rx_data[4] ;
    output \rx_data[3] ;
    output \rx_data[2] ;
    output \rx_data[1] ;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[29:38])
    
    wire o_data_7__N_185;
    wire [7:0]data_reg;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(142[12:20])
    
    wire qq_uart, q_uart, ck_uart, half_baud_time, half_baud_time_N_224;
    wire [3:0]state;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(75[13:18])
    
    wire dac_clk_p_c_enable_637;
    wire [3:0]state_3__N_89;
    
    wire data_reg_7__N_183;
    wire [23:0]n8;
    wire [23:0]baud_counter;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(78[17:29])
    
    wire dac_clk_p_c_enable_629, baud_counter_23__N_212;
    wire [23:0]baud_counter_23__N_188;
    
    wire zero_baud_counter, dac_clk_p_c_enable_221, n16540, n19359;
    wire [23:0]n254;
    
    wire n19360, n19341, n19342, n29275, n29274, n171;
    wire [3:0]n174;
    
    wire n27375, n19358, n19357, n29158, zero_baud_counter_N_221, 
        n12839, n27550, n29358, n27551, n29077, n22728, n22162, 
        n22712, n22720, n22718, n22710, n22696, n22706, n22708, 
        n22698, n19364, n19363, n19775, half_baud_time_N_225, n19774, 
        n19773, n19772, n19771, n19770, n19769, n19768, n19767, 
        n19766, n19765, n19764, n19362, n164, n19356, n19355, 
        n19354, n19353, n19352, n19351, n19350, n19349, n19348, 
        n19347, n19346, n19345, n19344, n19343, n19361, dac_clk_p_c_enable_570, 
        n29113;
    
    FD1P3AX o_data__i1 (.D(data_reg[0]), .SP(o_data_7__N_185), .CK(dac_clk_p_c), 
            .Q(\rx_data[0] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(155[9] 161[18])
    defparam o_data__i1.GSR = "DISABLED";
    FD1S3AY qq_uart_70 (.D(q_uart), .CK(dac_clk_p_c), .Q(qq_uart)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(90[9] 91[66])
    defparam qq_uart_70.GSR = "DISABLED";
    FD1S3AY ck_uart_71 (.D(qq_uart), .CK(dac_clk_p_c), .Q(ck_uart)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(90[9] 91[66])
    defparam ck_uart_71.GSR = "DISABLED";
    FD1S3AX half_baud_time_73 (.D(half_baud_time_N_224), .CK(dac_clk_p_c), 
            .Q(half_baud_time)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(111[9] 112[70])
    defparam half_baud_time_73.GSR = "DISABLED";
    FD1P3AY state_i0 (.D(state_3__N_89[0]), .SP(dac_clk_p_c_enable_637), 
            .CK(dac_clk_p_c), .Q(state[0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(116[9] 134[5])
    defparam state_i0.GSR = "DISABLED";
    FD1S3AX o_wr_76 (.D(o_data_7__N_185), .CK(dac_clk_p_c), .Q(rx_stb)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(155[9] 161[18])
    defparam o_wr_76.GSR = "DISABLED";
    FD1S3AY q_uart_69 (.D(i_wbu_uart_rx_c), .CK(dac_clk_p_c), .Q(q_uart)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(90[9] 91[66])
    defparam q_uart_69.GSR = "DISABLED";
    FD1P3AX data_reg_i0_i0 (.D(data_reg[1]), .SP(data_reg_7__N_183), .CK(dac_clk_p_c), 
            .Q(data_reg[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(143[9] 145[42])
    defparam data_reg_i0_i0.GSR = "DISABLED";
    FD1P3IX chg_counter__i0 (.D(n8[0]), .SP(dac_clk_p_c_enable_277), .CD(chg_counter_23__N_173), 
            .CK(dac_clk_p_c), .Q(chg_counter[0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i0.GSR = "DISABLED";
    FD1P3JX baud_counter_i1 (.D(baud_counter_23__N_188[1]), .SP(dac_clk_p_c_enable_629), 
            .PD(baud_counter_23__N_212), .CK(dac_clk_p_c), .Q(baud_counter[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i1.GSR = "DISABLED";
    FD1P3JX baud_counter_i2 (.D(baud_counter_23__N_188[2]), .SP(dac_clk_p_c_enable_629), 
            .PD(baud_counter_23__N_212), .CK(dac_clk_p_c), .Q(baud_counter[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i2.GSR = "DISABLED";
    FD1P3JX baud_counter_i3 (.D(baud_counter_23__N_188[3]), .SP(dac_clk_p_c_enable_629), 
            .PD(baud_counter_23__N_212), .CK(dac_clk_p_c), .Q(baud_counter[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i3.GSR = "DISABLED";
    FD1P3JX baud_counter_i8 (.D(baud_counter_23__N_188[8]), .SP(dac_clk_p_c_enable_629), 
            .PD(baud_counter_23__N_212), .CK(dac_clk_p_c), .Q(baud_counter[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i8.GSR = "DISABLED";
    FD1P3JX baud_counter_i9 (.D(baud_counter_23__N_188[9]), .SP(dac_clk_p_c_enable_629), 
            .PD(baud_counter_23__N_212), .CK(dac_clk_p_c), .Q(baud_counter[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i9.GSR = "DISABLED";
    FD1P3JX baud_counter_i10 (.D(baud_counter_23__N_188[10]), .SP(dac_clk_p_c_enable_629), 
            .PD(baud_counter_23__N_212), .CK(dac_clk_p_c), .Q(baud_counter[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i10.GSR = "DISABLED";
    FD1P3JX baud_counter_i13 (.D(baud_counter_23__N_188[13]), .SP(dac_clk_p_c_enable_629), 
            .PD(baud_counter_23__N_212), .CK(dac_clk_p_c), .Q(baud_counter[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i13.GSR = "DISABLED";
    FD1P3AY zero_baud_counter_79 (.D(n16540), .SP(dac_clk_p_c_enable_221), 
            .CK(dac_clk_p_c), .Q(zero_baud_counter)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(187[9] 195[29])
    defparam zero_baud_counter_79.GSR = "DISABLED";
    CCU2D sub_49_add_2_15 (.A0(baud_counter[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n19359), .COUT(n19360), .S0(n254[13]), 
          .S1(n254[14]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_15.INIT0 = 16'h5555;
    defparam sub_49_add_2_15.INIT1 = 16'h5555;
    defparam sub_49_add_2_15.INJECT1_0 = "NO";
    defparam sub_49_add_2_15.INJECT1_1 = "NO";
    CCU2D add_8_3 (.A0(chg_counter[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(chg_counter[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n19341), .COUT(n19342), .S0(n8[1]), .S1(n8[2]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:36])
    defparam add_8_3.INIT0 = 16'h5aaa;
    defparam add_8_3.INIT1 = 16'h5aaa;
    defparam add_8_3.INJECT1_0 = "NO";
    defparam add_8_3.INJECT1_1 = "NO";
    LUT4 i1_3_lut_4_lut (.A(n29275), .B(n29274), .C(zero_baud_counter), 
         .D(n171), .Z(dac_clk_p_c_enable_637)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(125[11] 134[5])
    defparam i1_3_lut_4_lut.init = 16'hfff8;
    LUT4 i1275_3_lut_4_lut_4_lut (.A(state[1]), .B(state[2]), .C(state[0]), 
         .D(state[3]), .Z(n174[2])) /* synthesis lut_function=(A (B ((D)+!C)+!B !((D)+!C))+!A (B)) */ ;
    defparam i1275_3_lut_4_lut_4_lut.init = 16'hcc6c;
    CCU2D add_8_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(chg_counter[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n19341), .S1(n8[0]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:36])
    defparam add_8_1.INIT0 = 16'hF000;
    defparam add_8_1.INIT1 = 16'h5555;
    defparam add_8_1.INJECT1_0 = "NO";
    defparam add_8_1.INJECT1_1 = "NO";
    LUT4 state_3__bdd_4_lut (.A(state[3]), .B(ck_uart), .C(half_baud_time), 
         .D(state[2]), .Z(n27375)) /* synthesis lut_function=(A (B+!(C (D)))+!A (D)) */ ;
    defparam state_3__bdd_4_lut.init = 16'hdfaa;
    CCU2D sub_49_add_2_13 (.A0(baud_counter[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n19358), .COUT(n19359), .S0(n254[11]), 
          .S1(n254[12]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_13.INIT0 = 16'h5555;
    defparam sub_49_add_2_13.INIT1 = 16'h5555;
    defparam sub_49_add_2_13.INJECT1_0 = "NO";
    defparam sub_49_add_2_13.INJECT1_1 = "NO";
    LUT4 qq_uart_I_0_2_lut (.A(qq_uart), .B(ck_uart), .Z(chg_counter_23__N_173)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(100[6:24])
    defparam qq_uart_I_0_2_lut.init = 16'h6666;
    CCU2D sub_49_add_2_11 (.A0(baud_counter[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n19357), .COUT(n19358), .S0(n254[9]), .S1(n254[10]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_11.INIT0 = 16'h5555;
    defparam sub_49_add_2_11.INIT1 = 16'h5555;
    defparam sub_49_add_2_11.INJECT1_0 = "NO";
    defparam sub_49_add_2_11.INJECT1_1 = "NO";
    LUT4 i13253_3_lut_4_lut (.A(state[0]), .B(n29158), .C(zero_baud_counter_N_221), 
         .D(n254[1]), .Z(baud_counter_23__N_188[1])) /* synthesis lut_function=(A (B (C+(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(117[6:25])
    defparam i13253_3_lut_4_lut.init = 16'hddd0;
    LUT4 i1_2_lut_3_lut_4_lut (.A(state[0]), .B(n29158), .C(zero_baud_counter_N_221), 
         .D(baud_counter_23__N_212), .Z(n12839)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(117[6:25])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfff2;
    LUT4 i13249_3_lut_4_lut (.A(state[0]), .B(n29158), .C(zero_baud_counter_N_221), 
         .D(n254[2]), .Z(baud_counter_23__N_188[2])) /* synthesis lut_function=(A (B (C+(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(117[6:25])
    defparam i13249_3_lut_4_lut.init = 16'hddd0;
    LUT4 i13246_3_lut_4_lut (.A(state[0]), .B(n29158), .C(zero_baud_counter_N_221), 
         .D(n254[3]), .Z(baud_counter_23__N_188[3])) /* synthesis lut_function=(A (B (C+(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(117[6:25])
    defparam i13246_3_lut_4_lut.init = 16'hddd0;
    LUT4 i13241_3_lut_4_lut (.A(state[0]), .B(n29158), .C(zero_baud_counter_N_221), 
         .D(n254[8]), .Z(baud_counter_23__N_188[8])) /* synthesis lut_function=(A (B (C+(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(117[6:25])
    defparam i13241_3_lut_4_lut.init = 16'hddd0;
    LUT4 i13240_3_lut_4_lut (.A(state[0]), .B(n29158), .C(zero_baud_counter_N_221), 
         .D(n254[9]), .Z(baud_counter_23__N_188[9])) /* synthesis lut_function=(A (B (C+(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(117[6:25])
    defparam i13240_3_lut_4_lut.init = 16'hddd0;
    LUT4 i13239_3_lut_4_lut (.A(state[0]), .B(n29158), .C(zero_baud_counter_N_221), 
         .D(n254[10]), .Z(baud_counter_23__N_188[10])) /* synthesis lut_function=(A (B (C+(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(117[6:25])
    defparam i13239_3_lut_4_lut.init = 16'hddd0;
    LUT4 i13224_3_lut_4_lut (.A(state[0]), .B(n29158), .C(zero_baud_counter_N_221), 
         .D(n254[13]), .Z(baud_counter_23__N_188[13])) /* synthesis lut_function=(A (B (C+(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(117[6:25])
    defparam i13224_3_lut_4_lut.init = 16'hddd0;
    LUT4 i24605_3_lut_4_lut (.A(state[0]), .B(n29158), .C(zero_baud_counter_N_221), 
         .D(baud_counter_23__N_212), .Z(n16540)) /* synthesis lut_function=(!(A (B (C+(D))+!B (D))+!A (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(117[6:25])
    defparam i24605_3_lut_4_lut.init = 16'h002f;
    LUT4 i12417_3_lut_4_lut (.A(state[0]), .B(n29158), .C(zero_baud_counter_N_221), 
         .D(n254[0]), .Z(baud_counter_23__N_188[0])) /* synthesis lut_function=(A (B (C+(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(117[6:25])
    defparam i12417_3_lut_4_lut.init = 16'hddd0;
    LUT4 i1_3_lut_4_lut_adj_213 (.A(state[0]), .B(n29158), .C(ck_uart), 
         .D(zero_baud_counter), .Z(o_data_7__N_185)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(117[6:25])
    defparam i1_3_lut_4_lut_adj_213.init = 16'h1000;
    FD1P3IX chg_counter__i23 (.D(n8[23]), .SP(dac_clk_p_c_enable_277), .CD(chg_counter_23__N_173), 
            .CK(dac_clk_p_c), .Q(chg_counter[23])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i23.GSR = "DISABLED";
    FD1P3IX chg_counter__i22 (.D(n8[22]), .SP(dac_clk_p_c_enable_277), .CD(chg_counter_23__N_173), 
            .CK(dac_clk_p_c), .Q(chg_counter[22])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i22.GSR = "DISABLED";
    FD1P3IX chg_counter__i21 (.D(n8[21]), .SP(dac_clk_p_c_enable_277), .CD(chg_counter_23__N_173), 
            .CK(dac_clk_p_c), .Q(chg_counter[21])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i21.GSR = "DISABLED";
    FD1P3IX chg_counter__i20 (.D(n8[20]), .SP(dac_clk_p_c_enable_277), .CD(chg_counter_23__N_173), 
            .CK(dac_clk_p_c), .Q(chg_counter[20])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i20.GSR = "DISABLED";
    FD1P3IX chg_counter__i19 (.D(n8[19]), .SP(dac_clk_p_c_enable_277), .CD(chg_counter_23__N_173), 
            .CK(dac_clk_p_c), .Q(chg_counter[19])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i19.GSR = "DISABLED";
    FD1P3IX chg_counter__i18 (.D(n8[18]), .SP(dac_clk_p_c_enable_277), .CD(chg_counter_23__N_173), 
            .CK(dac_clk_p_c), .Q(chg_counter[18])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i18.GSR = "DISABLED";
    FD1P3IX chg_counter__i17 (.D(n8[17]), .SP(dac_clk_p_c_enable_277), .CD(chg_counter_23__N_173), 
            .CK(dac_clk_p_c), .Q(chg_counter[17])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i17.GSR = "DISABLED";
    FD1P3IX chg_counter__i16 (.D(n8[16]), .SP(dac_clk_p_c_enable_277), .CD(chg_counter_23__N_173), 
            .CK(dac_clk_p_c), .Q(chg_counter[16])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i16.GSR = "DISABLED";
    FD1P3IX chg_counter__i15 (.D(n8[15]), .SP(dac_clk_p_c_enable_277), .CD(chg_counter_23__N_173), 
            .CK(dac_clk_p_c), .Q(chg_counter[15])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i15.GSR = "DISABLED";
    FD1P3IX chg_counter__i14 (.D(n8[14]), .SP(dac_clk_p_c_enable_277), .CD(chg_counter_23__N_173), 
            .CK(dac_clk_p_c), .Q(chg_counter[14])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i14.GSR = "DISABLED";
    FD1P3IX chg_counter__i13 (.D(n8[13]), .SP(dac_clk_p_c_enable_277), .CD(chg_counter_23__N_173), 
            .CK(dac_clk_p_c), .Q(chg_counter[13])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i13.GSR = "DISABLED";
    LUT4 ck_uart_bdd_2_lut (.A(ck_uart), .B(half_baud_time), .Z(n27550)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam ck_uart_bdd_2_lut.init = 16'hbbbb;
    LUT4 ck_uart_bdd_4_lut_28815 (.A(ck_uart), .B(state[0]), .C(state[3]), 
         .D(n29358), .Z(n27551)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C)+!B !(C (D)))) */ ;
    defparam ck_uart_bdd_4_lut_28815.init = 16'he3f3;
    FD1P3IX chg_counter__i12 (.D(n8[12]), .SP(dac_clk_p_c_enable_277), .CD(chg_counter_23__N_173), 
            .CK(dac_clk_p_c), .Q(chg_counter[12])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i12.GSR = "DISABLED";
    FD1P3IX chg_counter__i11 (.D(n8[11]), .SP(dac_clk_p_c_enable_277), .CD(chg_counter_23__N_173), 
            .CK(dac_clk_p_c), .Q(chg_counter[11])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i11.GSR = "DISABLED";
    FD1P3IX chg_counter__i10 (.D(n8[10]), .SP(dac_clk_p_c_enable_277), .CD(chg_counter_23__N_173), 
            .CK(dac_clk_p_c), .Q(chg_counter[10])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i10.GSR = "DISABLED";
    FD1P3IX chg_counter__i9 (.D(n8[9]), .SP(dac_clk_p_c_enable_277), .CD(chg_counter_23__N_173), 
            .CK(dac_clk_p_c), .Q(chg_counter[9])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i9.GSR = "DISABLED";
    FD1P3IX chg_counter__i8 (.D(n8[8]), .SP(dac_clk_p_c_enable_277), .CD(chg_counter_23__N_173), 
            .CK(dac_clk_p_c), .Q(chg_counter[8])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i8.GSR = "DISABLED";
    FD1P3IX chg_counter__i7 (.D(n8[7]), .SP(dac_clk_p_c_enable_277), .CD(chg_counter_23__N_173), 
            .CK(dac_clk_p_c), .Q(chg_counter[7])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i7.GSR = "DISABLED";
    FD1P3IX chg_counter__i6 (.D(n8[6]), .SP(dac_clk_p_c_enable_277), .CD(chg_counter_23__N_173), 
            .CK(dac_clk_p_c), .Q(chg_counter[6])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i6.GSR = "DISABLED";
    FD1P3IX chg_counter__i5 (.D(n8[5]), .SP(dac_clk_p_c_enable_277), .CD(chg_counter_23__N_173), 
            .CK(dac_clk_p_c), .Q(chg_counter[5])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i5.GSR = "DISABLED";
    FD1P3IX chg_counter__i4 (.D(n8[4]), .SP(dac_clk_p_c_enable_277), .CD(chg_counter_23__N_173), 
            .CK(dac_clk_p_c), .Q(chg_counter[4])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i4.GSR = "DISABLED";
    FD1P3IX chg_counter__i3 (.D(n8[3]), .SP(dac_clk_p_c_enable_277), .CD(chg_counter_23__N_173), 
            .CK(dac_clk_p_c), .Q(chg_counter[3])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i3.GSR = "DISABLED";
    FD1P3IX chg_counter__i2 (.D(n8[2]), .SP(dac_clk_p_c_enable_277), .CD(chg_counter_23__N_173), 
            .CK(dac_clk_p_c), .Q(chg_counter[2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i2.GSR = "DISABLED";
    FD1P3IX chg_counter__i1 (.D(n8[1]), .SP(dac_clk_p_c_enable_277), .CD(chg_counter_23__N_173), 
            .CK(dac_clk_p_c), .Q(chg_counter[1])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i1.GSR = "DISABLED";
    FD1P3AX data_reg_i0_i7 (.D(qq_uart), .SP(data_reg_7__N_183), .CK(dac_clk_p_c), 
            .Q(data_reg[7])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(143[9] 145[42])
    defparam data_reg_i0_i7.GSR = "DISABLED";
    LUT4 i1_3_lut_4_lut_adj_214 (.A(baud_counter_23__N_212), .B(n29077), 
         .C(state[3]), .D(zero_baud_counter), .Z(dac_clk_p_c_enable_629)) /* synthesis lut_function=(A+!(B (C (D)))) */ ;
    defparam i1_3_lut_4_lut_adj_214.init = 16'hbfff;
    LUT4 zero_baud_counter_I_0_82_2_lut_3_lut_4_lut (.A(state[3]), .B(n29358), 
         .C(zero_baud_counter), .D(state[0]), .Z(data_reg_7__N_183)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(117[6:25])
    defparam zero_baud_counter_I_0_82_2_lut_3_lut_4_lut.init = 16'hf0d0;
    LUT4 i1_4_lut (.A(n29274), .B(ck_uart), .C(n22728), .D(state[1]), 
         .Z(baud_counter_23__N_212)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(125[11] 134[5])
    defparam i1_4_lut.init = 16'h2000;
    LUT4 zero_baud_counter_I_0_2_lut (.A(zero_baud_counter), .B(state[3]), 
         .Z(zero_baud_counter_N_221)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(175[11:52])
    defparam zero_baud_counter_I_0_2_lut.init = 16'h2222;
    LUT4 i1_2_lut (.A(state[2]), .B(half_baud_time), .Z(n22728)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(125[11] 134[5])
    defparam i1_2_lut.init = 16'h8888;
    FD1P3AX data_reg_i0_i6 (.D(data_reg[7]), .SP(data_reg_7__N_183), .CK(dac_clk_p_c), 
            .Q(data_reg[6])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(143[9] 145[42])
    defparam data_reg_i0_i6.GSR = "DISABLED";
    FD1P3AX data_reg_i0_i5 (.D(data_reg[6]), .SP(data_reg_7__N_183), .CK(dac_clk_p_c), 
            .Q(data_reg[5])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(143[9] 145[42])
    defparam data_reg_i0_i5.GSR = "DISABLED";
    FD1P3AX data_reg_i0_i4 (.D(data_reg[5]), .SP(data_reg_7__N_183), .CK(dac_clk_p_c), 
            .Q(data_reg[4])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(143[9] 145[42])
    defparam data_reg_i0_i4.GSR = "DISABLED";
    FD1P3AX data_reg_i0_i3 (.D(data_reg[4]), .SP(data_reg_7__N_183), .CK(dac_clk_p_c), 
            .Q(data_reg[3])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(143[9] 145[42])
    defparam data_reg_i0_i3.GSR = "DISABLED";
    FD1P3AX data_reg_i0_i2 (.D(data_reg[3]), .SP(data_reg_7__N_183), .CK(dac_clk_p_c), 
            .Q(data_reg[2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(143[9] 145[42])
    defparam data_reg_i0_i2.GSR = "DISABLED";
    FD1P3AX data_reg_i0_i1 (.D(data_reg[2]), .SP(data_reg_7__N_183), .CK(dac_clk_p_c), 
            .Q(data_reg[1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(143[9] 145[42])
    defparam data_reg_i0_i1.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_215 (.A(n22162), .B(n29077), .C(baud_counter_23__N_212), 
         .D(zero_baud_counter_N_221), .Z(dac_clk_p_c_enable_221)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;
    defparam i1_4_lut_adj_215.init = 16'hfff7;
    LUT4 i1_4_lut_adj_216 (.A(n22712), .B(n22720), .C(n22718), .D(n22710), 
         .Z(n22162)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(194[11:28])
    defparam i1_4_lut_adj_216.init = 16'hfffe;
    LUT4 i1_4_lut_adj_217 (.A(baud_counter[14]), .B(baud_counter[21]), .C(baud_counter[20]), 
         .D(baud_counter[3]), .Z(n22712)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(194[11:28])
    defparam i1_4_lut_adj_217.init = 16'hfffe;
    LUT4 i1_4_lut_adj_218 (.A(n22696), .B(baud_counter[0]), .C(n22706), 
         .D(baud_counter[8]), .Z(n22720)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(194[11:28])
    defparam i1_4_lut_adj_218.init = 16'hfffb;
    LUT4 i1_4_lut_adj_219 (.A(baud_counter[7]), .B(n22708), .C(n22698), 
         .D(baud_counter[22]), .Z(n22718)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(194[11:28])
    defparam i1_4_lut_adj_219.init = 16'hfffe;
    LUT4 i1_4_lut_adj_220 (.A(baud_counter[6]), .B(baud_counter[12]), .C(baud_counter[13]), 
         .D(baud_counter[5]), .Z(n22710)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(194[11:28])
    defparam i1_4_lut_adj_220.init = 16'hfffe;
    LUT4 i1_2_lut_adj_221 (.A(baud_counter[19]), .B(baud_counter[1]), .Z(n22696)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(194[11:28])
    defparam i1_2_lut_adj_221.init = 16'heeee;
    LUT4 i1_4_lut_adj_222 (.A(baud_counter[15]), .B(baud_counter[9]), .C(baud_counter[17]), 
         .D(baud_counter[23]), .Z(n22706)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(194[11:28])
    defparam i1_4_lut_adj_222.init = 16'hfffe;
    LUT4 i1_4_lut_adj_223 (.A(baud_counter[4]), .B(baud_counter[16]), .C(baud_counter[18]), 
         .D(baud_counter[2]), .Z(n22708)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(194[11:28])
    defparam i1_4_lut_adj_223.init = 16'hfffe;
    LUT4 i1_2_lut_adj_224 (.A(baud_counter[11]), .B(baud_counter[10]), .Z(n22698)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(194[11:28])
    defparam i1_2_lut_adj_224.init = 16'heeee;
    LUT4 state_3__bdd_3_lut_4_lut (.A(state[3]), .B(n27375), .C(state[1]), 
         .D(state[0]), .Z(state_3__N_89[3])) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C (D)))) */ ;
    defparam state_3__bdd_3_lut_4_lut.init = 16'hcaaa;
    CCU2D sub_49_add_2_25 (.A0(baud_counter[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n19364), .S0(n254[23]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_25.INIT0 = 16'h5555;
    defparam sub_49_add_2_25.INIT1 = 16'h0000;
    defparam sub_49_add_2_25.INJECT1_0 = "NO";
    defparam sub_49_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_49_add_2_23 (.A0(baud_counter[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n19363), .COUT(n19364), .S0(n254[21]), 
          .S1(n254[22]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_23.INIT0 = 16'h5555;
    defparam sub_49_add_2_23.INIT1 = 16'h5555;
    defparam sub_49_add_2_23.INJECT1_0 = "NO";
    defparam sub_49_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_542_add_2_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n19775), .S0(half_baud_time_N_225));
    defparam sub_542_add_2_cout.INIT0 = 16'h0000;
    defparam sub_542_add_2_cout.INIT1 = 16'h0000;
    defparam sub_542_add_2_cout.INJECT1_0 = "NO";
    defparam sub_542_add_2_cout.INJECT1_1 = "NO";
    CCU2D sub_542_add_2_24 (.A0(chg_counter[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n19774), .COUT(n19775));
    defparam sub_542_add_2_24.INIT0 = 16'h5555;
    defparam sub_542_add_2_24.INIT1 = 16'h5555;
    defparam sub_542_add_2_24.INJECT1_0 = "NO";
    defparam sub_542_add_2_24.INJECT1_1 = "NO";
    CCU2D sub_542_add_2_22 (.A0(chg_counter[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n19773), .COUT(n19774));
    defparam sub_542_add_2_22.INIT0 = 16'h5555;
    defparam sub_542_add_2_22.INIT1 = 16'h5555;
    defparam sub_542_add_2_22.INJECT1_0 = "NO";
    defparam sub_542_add_2_22.INJECT1_1 = "NO";
    CCU2D sub_542_add_2_20 (.A0(chg_counter[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n19772), .COUT(n19773));
    defparam sub_542_add_2_20.INIT0 = 16'h5555;
    defparam sub_542_add_2_20.INIT1 = 16'h5555;
    defparam sub_542_add_2_20.INJECT1_0 = "NO";
    defparam sub_542_add_2_20.INJECT1_1 = "NO";
    CCU2D sub_542_add_2_18 (.A0(chg_counter[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n19771), .COUT(n19772));
    defparam sub_542_add_2_18.INIT0 = 16'h5555;
    defparam sub_542_add_2_18.INIT1 = 16'h5555;
    defparam sub_542_add_2_18.INJECT1_0 = "NO";
    defparam sub_542_add_2_18.INJECT1_1 = "NO";
    CCU2D sub_542_add_2_16 (.A0(chg_counter[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n19770), .COUT(n19771));
    defparam sub_542_add_2_16.INIT0 = 16'h5555;
    defparam sub_542_add_2_16.INIT1 = 16'h5555;
    defparam sub_542_add_2_16.INJECT1_0 = "NO";
    defparam sub_542_add_2_16.INJECT1_1 = "NO";
    CCU2D sub_542_add_2_14 (.A0(chg_counter[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n19769), .COUT(n19770));
    defparam sub_542_add_2_14.INIT0 = 16'h5aaa;
    defparam sub_542_add_2_14.INIT1 = 16'h5555;
    defparam sub_542_add_2_14.INJECT1_0 = "NO";
    defparam sub_542_add_2_14.INJECT1_1 = "NO";
    CCU2D sub_542_add_2_12 (.A0(chg_counter[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n19768), .COUT(n19769));
    defparam sub_542_add_2_12.INIT0 = 16'h5555;
    defparam sub_542_add_2_12.INIT1 = 16'h5555;
    defparam sub_542_add_2_12.INJECT1_0 = "NO";
    defparam sub_542_add_2_12.INJECT1_1 = "NO";
    LUT4 i1_2_lut_adj_225 (.A(ck_uart), .B(half_baud_time_N_225), .Z(half_baud_time_N_224)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(112[21:31])
    defparam i1_2_lut_adj_225.init = 16'h4444;
    CCU2D sub_542_add_2_10 (.A0(chg_counter[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n19767), .COUT(n19768));
    defparam sub_542_add_2_10.INIT0 = 16'h5aaa;
    defparam sub_542_add_2_10.INIT1 = 16'h5aaa;
    defparam sub_542_add_2_10.INJECT1_0 = "NO";
    defparam sub_542_add_2_10.INJECT1_1 = "NO";
    CCU2D sub_542_add_2_8 (.A0(chg_counter[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n19766), .COUT(n19767));
    defparam sub_542_add_2_8.INIT0 = 16'h5555;
    defparam sub_542_add_2_8.INIT1 = 16'h5aaa;
    defparam sub_542_add_2_8.INJECT1_0 = "NO";
    defparam sub_542_add_2_8.INJECT1_1 = "NO";
    CCU2D sub_542_add_2_6 (.A0(chg_counter[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n19765), .COUT(n19766));
    defparam sub_542_add_2_6.INIT0 = 16'h5555;
    defparam sub_542_add_2_6.INIT1 = 16'h5555;
    defparam sub_542_add_2_6.INJECT1_0 = "NO";
    defparam sub_542_add_2_6.INJECT1_1 = "NO";
    CCU2D sub_542_add_2_4 (.A0(chg_counter[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n19764), .COUT(n19765));
    defparam sub_542_add_2_4.INIT0 = 16'h5aaa;
    defparam sub_542_add_2_4.INIT1 = 16'h5555;
    defparam sub_542_add_2_4.INJECT1_0 = "NO";
    defparam sub_542_add_2_4.INJECT1_1 = "NO";
    CCU2D sub_542_add_2_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(chg_counter[1]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n19764));
    defparam sub_542_add_2_2.INIT0 = 16'h0000;
    defparam sub_542_add_2_2.INIT1 = 16'h5aaa;
    defparam sub_542_add_2_2.INJECT1_0 = "NO";
    defparam sub_542_add_2_2.INJECT1_1 = "NO";
    CCU2D sub_49_add_2_21 (.A0(baud_counter[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n19362), .COUT(n19363), .S0(n254[19]), 
          .S1(n254[20]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_21.INIT0 = 16'h5555;
    defparam sub_49_add_2_21.INIT1 = 16'h5555;
    defparam sub_49_add_2_21.INJECT1_0 = "NO";
    defparam sub_49_add_2_21.INJECT1_1 = "NO";
    LUT4 i1_2_lut_adj_226 (.A(ck_uart), .B(half_baud_time), .Z(n164)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(112[21:31])
    defparam i1_2_lut_adj_226.init = 16'h4444;
    CCU2D sub_49_add_2_9 (.A0(baud_counter[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n19356), .COUT(n19357), .S0(n254[7]), .S1(n254[8]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_9.INIT0 = 16'h5555;
    defparam sub_49_add_2_9.INIT1 = 16'h5555;
    defparam sub_49_add_2_9.INJECT1_0 = "NO";
    defparam sub_49_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_49_add_2_7 (.A0(baud_counter[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n19355), .COUT(n19356), .S0(n254[5]), .S1(n254[6]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_7.INIT0 = 16'h5555;
    defparam sub_49_add_2_7.INIT1 = 16'h5555;
    defparam sub_49_add_2_7.INJECT1_0 = "NO";
    defparam sub_49_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_49_add_2_5 (.A0(baud_counter[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n19354), .COUT(n19355), .S0(n254[3]), .S1(n254[4]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_5.INIT0 = 16'h5555;
    defparam sub_49_add_2_5.INIT1 = 16'h5555;
    defparam sub_49_add_2_5.INJECT1_0 = "NO";
    defparam sub_49_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_49_add_2_3 (.A0(baud_counter[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n19353), .COUT(n19354), .S0(n254[1]), .S1(n254[2]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_3.INIT0 = 16'h5555;
    defparam sub_49_add_2_3.INIT1 = 16'h5555;
    defparam sub_49_add_2_3.INJECT1_0 = "NO";
    defparam sub_49_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_49_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(baud_counter[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n19353), .S1(n254[0]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_1.INIT0 = 16'hF000;
    defparam sub_49_add_2_1.INIT1 = 16'h5555;
    defparam sub_49_add_2_1.INJECT1_0 = "NO";
    defparam sub_49_add_2_1.INJECT1_1 = "NO";
    CCU2D add_8_25 (.A0(chg_counter[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n19352), .S0(n8[23]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:36])
    defparam add_8_25.INIT0 = 16'h5aaa;
    defparam add_8_25.INIT1 = 16'h0000;
    defparam add_8_25.INJECT1_0 = "NO";
    defparam add_8_25.INJECT1_1 = "NO";
    CCU2D add_8_23 (.A0(chg_counter[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n19351), .COUT(n19352), .S0(n8[21]), .S1(n8[22]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:36])
    defparam add_8_23.INIT0 = 16'h5aaa;
    defparam add_8_23.INIT1 = 16'h5aaa;
    defparam add_8_23.INJECT1_0 = "NO";
    defparam add_8_23.INJECT1_1 = "NO";
    CCU2D add_8_21 (.A0(chg_counter[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n19350), .COUT(n19351), .S0(n8[19]), .S1(n8[20]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:36])
    defparam add_8_21.INIT0 = 16'h5aaa;
    defparam add_8_21.INIT1 = 16'h5aaa;
    defparam add_8_21.INJECT1_0 = "NO";
    defparam add_8_21.INJECT1_1 = "NO";
    CCU2D add_8_19 (.A0(chg_counter[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n19349), .COUT(n19350), .S0(n8[17]), .S1(n8[18]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:36])
    defparam add_8_19.INIT0 = 16'h5aaa;
    defparam add_8_19.INIT1 = 16'h5aaa;
    defparam add_8_19.INJECT1_0 = "NO";
    defparam add_8_19.INJECT1_1 = "NO";
    CCU2D add_8_17 (.A0(chg_counter[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n19348), .COUT(n19349), .S0(n8[15]), .S1(n8[16]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:36])
    defparam add_8_17.INIT0 = 16'h5aaa;
    defparam add_8_17.INIT1 = 16'h5aaa;
    defparam add_8_17.INJECT1_0 = "NO";
    defparam add_8_17.INJECT1_1 = "NO";
    CCU2D add_8_15 (.A0(chg_counter[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n19347), .COUT(n19348), .S0(n8[13]), .S1(n8[14]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:36])
    defparam add_8_15.INIT0 = 16'h5aaa;
    defparam add_8_15.INIT1 = 16'h5aaa;
    defparam add_8_15.INJECT1_0 = "NO";
    defparam add_8_15.INJECT1_1 = "NO";
    CCU2D add_8_13 (.A0(chg_counter[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n19346), .COUT(n19347), .S0(n8[11]), .S1(n8[12]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:36])
    defparam add_8_13.INIT0 = 16'h5aaa;
    defparam add_8_13.INIT1 = 16'h5aaa;
    defparam add_8_13.INJECT1_0 = "NO";
    defparam add_8_13.INJECT1_1 = "NO";
    CCU2D add_8_11 (.A0(chg_counter[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(chg_counter[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n19345), .COUT(n19346), .S0(n8[9]), .S1(n8[10]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:36])
    defparam add_8_11.INIT0 = 16'h5aaa;
    defparam add_8_11.INIT1 = 16'h5aaa;
    defparam add_8_11.INJECT1_0 = "NO";
    defparam add_8_11.INJECT1_1 = "NO";
    CCU2D add_8_9 (.A0(chg_counter[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(chg_counter[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n19344), .COUT(n19345), .S0(n8[7]), .S1(n8[8]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:36])
    defparam add_8_9.INIT0 = 16'h5aaa;
    defparam add_8_9.INIT1 = 16'h5aaa;
    defparam add_8_9.INJECT1_0 = "NO";
    defparam add_8_9.INJECT1_1 = "NO";
    CCU2D add_8_7 (.A0(chg_counter[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(chg_counter[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n19343), .COUT(n19344), .S0(n8[5]), .S1(n8[6]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:36])
    defparam add_8_7.INIT0 = 16'h5aaa;
    defparam add_8_7.INIT1 = 16'h5aaa;
    defparam add_8_7.INJECT1_0 = "NO";
    defparam add_8_7.INJECT1_1 = "NO";
    CCU2D sub_49_add_2_19 (.A0(baud_counter[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n19361), .COUT(n19362), .S0(n254[17]), 
          .S1(n254[18]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_19.INIT0 = 16'h5555;
    defparam sub_49_add_2_19.INIT1 = 16'h5555;
    defparam sub_49_add_2_19.INJECT1_0 = "NO";
    defparam sub_49_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_49_add_2_17 (.A0(baud_counter[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n19360), .COUT(n19361), .S0(n254[15]), 
          .S1(n254[16]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_17.INIT0 = 16'h5555;
    defparam sub_49_add_2_17.INIT1 = 16'h5555;
    defparam sub_49_add_2_17.INJECT1_0 = "NO";
    defparam sub_49_add_2_17.INJECT1_1 = "NO";
    FD1P3IX baud_counter_i23 (.D(n254[23]), .SP(dac_clk_p_c_enable_570), 
            .CD(n12839), .CK(dac_clk_p_c), .Q(baud_counter[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i23.GSR = "DISABLED";
    FD1P3IX baud_counter_i22 (.D(n254[22]), .SP(dac_clk_p_c_enable_570), 
            .CD(n12839), .CK(dac_clk_p_c), .Q(baud_counter[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i22.GSR = "DISABLED";
    FD1P3IX baud_counter_i21 (.D(n254[21]), .SP(dac_clk_p_c_enable_570), 
            .CD(n12839), .CK(dac_clk_p_c), .Q(baud_counter[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i21.GSR = "DISABLED";
    FD1P3IX baud_counter_i20 (.D(n254[20]), .SP(dac_clk_p_c_enable_570), 
            .CD(n12839), .CK(dac_clk_p_c), .Q(baud_counter[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i20.GSR = "DISABLED";
    FD1P3IX baud_counter_i19 (.D(n254[19]), .SP(dac_clk_p_c_enable_570), 
            .CD(n12839), .CK(dac_clk_p_c), .Q(baud_counter[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i19.GSR = "DISABLED";
    FD1P3IX baud_counter_i18 (.D(n254[18]), .SP(dac_clk_p_c_enable_570), 
            .CD(n12839), .CK(dac_clk_p_c), .Q(baud_counter[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i18.GSR = "DISABLED";
    FD1P3IX baud_counter_i17 (.D(n254[17]), .SP(dac_clk_p_c_enable_570), 
            .CD(n12839), .CK(dac_clk_p_c), .Q(baud_counter[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i17.GSR = "DISABLED";
    FD1P3IX baud_counter_i16 (.D(n254[16]), .SP(dac_clk_p_c_enable_570), 
            .CD(n12839), .CK(dac_clk_p_c), .Q(baud_counter[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i16.GSR = "DISABLED";
    FD1P3IX baud_counter_i15 (.D(n254[15]), .SP(dac_clk_p_c_enable_570), 
            .CD(n12839), .CK(dac_clk_p_c), .Q(baud_counter[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i15.GSR = "DISABLED";
    FD1P3IX baud_counter_i14 (.D(n254[14]), .SP(dac_clk_p_c_enable_570), 
            .CD(n12839), .CK(dac_clk_p_c), .Q(baud_counter[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i14.GSR = "DISABLED";
    FD1P3IX baud_counter_i12 (.D(n254[12]), .SP(dac_clk_p_c_enable_570), 
            .CD(n12839), .CK(dac_clk_p_c), .Q(baud_counter[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i12.GSR = "DISABLED";
    FD1P3IX baud_counter_i11 (.D(n254[11]), .SP(dac_clk_p_c_enable_570), 
            .CD(n12839), .CK(dac_clk_p_c), .Q(baud_counter[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i11.GSR = "DISABLED";
    FD1P3IX baud_counter_i7 (.D(n254[7]), .SP(dac_clk_p_c_enable_570), .CD(n12839), 
            .CK(dac_clk_p_c), .Q(baud_counter[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i7.GSR = "DISABLED";
    FD1P3IX baud_counter_i6 (.D(n254[6]), .SP(dac_clk_p_c_enable_570), .CD(n12839), 
            .CK(dac_clk_p_c), .Q(baud_counter[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i6.GSR = "DISABLED";
    FD1P3IX baud_counter_i5 (.D(n254[5]), .SP(dac_clk_p_c_enable_570), .CD(n12839), 
            .CK(dac_clk_p_c), .Q(baud_counter[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i5.GSR = "DISABLED";
    FD1P3IX baud_counter_i4 (.D(n254[4]), .SP(dac_clk_p_c_enable_570), .CD(n12839), 
            .CK(dac_clk_p_c), .Q(baud_counter[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i4.GSR = "DISABLED";
    LUT4 i11320_1_lut (.A(zero_baud_counter), .Z(dac_clk_p_c_enable_570)) /* synthesis lut_function=(!(A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(187[9] 195[29])
    defparam i11320_1_lut.init = 16'h5555;
    CCU2D add_8_5 (.A0(chg_counter[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(chg_counter[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n19342), .COUT(n19343), .S0(n8[3]), .S1(n8[4]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:36])
    defparam add_8_5.INIT0 = 16'h5aaa;
    defparam add_8_5.INIT1 = 16'h5aaa;
    defparam add_8_5.INJECT1_0 = "NO";
    defparam add_8_5.INJECT1_1 = "NO";
    LUT4 i1_3_lut_4_lut_adj_227 (.A(state[0]), .B(n29358), .C(ck_uart), 
         .D(state[3]), .Z(n171)) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;
    defparam i1_3_lut_4_lut_adj_227.init = 16'he000;
    LUT4 i1_2_lut_rep_698 (.A(state[1]), .B(state[2]), .Z(n29358)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(117[6:25])
    defparam i1_2_lut_rep_698.init = 16'heeee;
    LUT4 i1268_3_lut_4_lut_3_lut_3_lut (.A(state[1]), .B(state[3]), .C(state[0]), 
         .Z(n174[1])) /* synthesis lut_function=(A (B+!(C))+!A !(B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(117[6:25])
    defparam i1268_3_lut_4_lut_3_lut_3_lut.init = 16'h9a9a;
    LUT4 i1_2_lut_rep_498_3_lut (.A(state[1]), .B(state[2]), .C(state[3]), 
         .Z(n29158)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(117[6:25])
    defparam i1_2_lut_rep_498_3_lut.init = 16'hefef;
    LUT4 i1_rep_417_3_lut_4_lut (.A(state[1]), .B(state[2]), .C(state[0]), 
         .D(state[3]), .Z(n29077)) /* synthesis lut_function=(A+(B+!(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(117[6:25])
    defparam i1_rep_417_3_lut_4_lut.init = 16'hefff;
    LUT4 state_3__I_0_80_i3_4_lut (.A(n164), .B(n174[2]), .C(n29113), 
         .D(n171), .Z(state_3__N_89[2])) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A !(B+(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(125[11] 134[5])
    defparam state_3__I_0_80_i3_4_lut.init = 16'h5f5c;
    LUT4 state_3__I_0_80_i2_4_lut (.A(n164), .B(n174[1]), .C(n29113), 
         .D(n171), .Z(state_3__N_89[1])) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A !(B+(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(125[11] 134[5])
    defparam state_3__I_0_80_i2_4_lut.init = 16'h5f5c;
    LUT4 i1_2_lut_rep_614 (.A(state[0]), .B(state[3]), .Z(n29274)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_614.init = 16'h8888;
    LUT4 i1_2_lut_rep_615 (.A(state[1]), .B(state[2]), .Z(n29275)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(125[11] 134[5])
    defparam i1_2_lut_rep_615.init = 16'h8888;
    PFUMX i25798 (.BLUT(n27551), .ALUT(n27550), .C0(n29113), .Z(state_3__N_89[0]));
    LUT4 i1_2_lut_rep_453_3_lut_4_lut (.A(state[1]), .B(state[2]), .C(state[3]), 
         .D(state[0]), .Z(n29113)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(125[11] 134[5])
    defparam i1_2_lut_rep_453_3_lut_4_lut.init = 16'h8000;
    FD1P3JX baud_counter_i0 (.D(baud_counter_23__N_188[0]), .SP(dac_clk_p_c_enable_629), 
            .PD(baud_counter_23__N_212), .CK(dac_clk_p_c), .Q(baud_counter[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i0.GSR = "DISABLED";
    FD1P3AY state_i3 (.D(state_3__N_89[3]), .SP(dac_clk_p_c_enable_637), 
            .CK(dac_clk_p_c), .Q(state[3])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(116[9] 134[5])
    defparam state_i3.GSR = "DISABLED";
    FD1P3AY state_i2 (.D(state_3__N_89[2]), .SP(dac_clk_p_c_enable_637), 
            .CK(dac_clk_p_c), .Q(state[2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(116[9] 134[5])
    defparam state_i2.GSR = "DISABLED";
    FD1P3AY state_i1 (.D(state_3__N_89[1]), .SP(dac_clk_p_c_enable_637), 
            .CK(dac_clk_p_c), .Q(state[1])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(116[9] 134[5])
    defparam state_i1.GSR = "DISABLED";
    FD1P3AX o_data__i7 (.D(data_reg[6]), .SP(o_data_7__N_185), .CK(dac_clk_p_c), 
            .Q(\rx_data[6] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(155[9] 161[18])
    defparam o_data__i7.GSR = "DISABLED";
    FD1P3AX o_data__i6 (.D(data_reg[5]), .SP(o_data_7__N_185), .CK(dac_clk_p_c), 
            .Q(\rx_data[5] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(155[9] 161[18])
    defparam o_data__i6.GSR = "DISABLED";
    FD1P3AX o_data__i5 (.D(data_reg[4]), .SP(o_data_7__N_185), .CK(dac_clk_p_c), 
            .Q(\rx_data[4] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(155[9] 161[18])
    defparam o_data__i5.GSR = "DISABLED";
    FD1P3AX o_data__i4 (.D(data_reg[3]), .SP(o_data_7__N_185), .CK(dac_clk_p_c), 
            .Q(\rx_data[3] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(155[9] 161[18])
    defparam o_data__i4.GSR = "DISABLED";
    FD1P3AX o_data__i3 (.D(data_reg[2]), .SP(o_data_7__N_185), .CK(dac_clk_p_c), 
            .Q(\rx_data[2] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(155[9] 161[18])
    defparam o_data__i3.GSR = "DISABLED";
    FD1P3AX o_data__i2 (.D(data_reg[1]), .SP(o_data_7__N_185), .CK(dac_clk_p_c), 
            .Q(\rx_data[1] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=7, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=60, LSE_RLINE=60 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(155[9] 161[18])
    defparam o_data__i2.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module control
//

module control (dac_clk_p_c, dac_clk_p_c_enable_227, wb_odata, dac_clk_p_c_enable_243, 
            i_sw0_c, lo_i_en, \addr_space[4][1] , \addr_space[4][0] , 
            dac_clk_p_c_enable_106, dac_clk_p_c_enable_241, wb_control_data, 
            o_wb_data_31__N_2456, lo_q_en, \addr_space[1][1] , \addr_space[1][0] , 
            \addr_space[2][1] , \addr_space[2][0] , \addr_space[3][1] , 
            n29300, \wb_addr[2] , \addr_space[3][0] , wb_control_ack, 
            wb_control_data_31__N_35, n21662, n29302, n29065, n22526, 
            \o_wb_data_31__N_2456[1] , \wb_addr[1] , \wb_addr[0] , lo_q, 
            o_lo_q_c) /* synthesis syn_module_defined=1 */ ;
    input dac_clk_p_c;
    input dac_clk_p_c_enable_227;
    input [31:0]wb_odata;
    input dac_clk_p_c_enable_243;
    input i_sw0_c;
    output lo_i_en;
    output \addr_space[4][1] ;
    output \addr_space[4][0] ;
    input dac_clk_p_c_enable_106;
    input dac_clk_p_c_enable_241;
    output [31:0]wb_control_data;
    input [31:0]o_wb_data_31__N_2456;
    output lo_q_en;
    output \addr_space[1][1] ;
    output \addr_space[1][0] ;
    output \addr_space[2][1] ;
    output \addr_space[2][0] ;
    output \addr_space[3][1] ;
    input n29300;
    input \wb_addr[2] ;
    output \addr_space[3][0] ;
    output wb_control_ack;
    input wb_control_data_31__N_35;
    input n21662;
    input n29302;
    input n29065;
    input n22526;
    input \o_wb_data_31__N_2456[1] ;
    input \wb_addr[1] ;
    input \wb_addr[0] ;
    input lo_q;
    output o_lo_q_c;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[29:38])
    wire lo_q /* synthesis is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(159[24:28])
    wire [31:0]\addr_space[4] ;   // d:/documents/git_local/fm_modulator/rtl/control.v(22[12:22])
    wire [31:0]\addr_space[2] ;   // d:/documents/git_local/fm_modulator/rtl/control.v(22[12:22])
    wire [31:0]\addr_space[0] ;   // d:/documents/git_local/fm_modulator/rtl/control.v(22[12:22])
    
    wire dac_clk_p_c_enable_79;
    wire [31:0]\addr_space[1] ;   // d:/documents/git_local/fm_modulator/rtl/control.v(22[12:22])
    wire [31:0]\addr_space[3] ;   // d:/documents/git_local/fm_modulator/rtl/control.v(22[12:22])
    
    wire n26891;
    wire [31:0]o_wb_data_31__N_2456_c;
    
    wire n26886, n26875, n26863, n26858, n26842, n26831, n26826, 
        n26817, n26812, n26807, n26802, n26789, n26777, n26759, 
        n26699, n26700, n26750, n26704, n26705, n26709, n26710, 
        n26714, n26715, n26739, n26732, n26733, n26737, n26738, 
        n26734, n26939, n26938, n26940, n26748, n26934, n26933, 
        n26935, n26929, n26928, n26930, n26749, n26924, n26923, 
        n26925, n26716, n26711, n26706, n26701, n26919, n26918, 
        n26920, n26757, n26758, n26914, n26913, n26915, n26909, 
        n26908, n26910, n26775, n26776, n26895, n26894, n26896, 
        n26890, n26889, n26787, n26788, n26885, n26884, n26801, 
        n26800, n26805, n26806, n26810, n26811, n26874, n26873, 
        n26815, n26816, n26825, n26824, n26829, n26862, n26861, 
        n26830, n26857, n26856, n26841, n26840;
    
    FD1P3AX \addr_space_4[[22__424  (.D(wb_odata[22]), .SP(dac_clk_p_c_enable_227), 
            .CK(dac_clk_p_c), .Q(\addr_space[4] [22])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_4[[22__424 .GSR = "DISABLED";
    FD1P3AX \addr_space_4[[21__426  (.D(wb_odata[21]), .SP(dac_clk_p_c_enable_227), 
            .CK(dac_clk_p_c), .Q(\addr_space[4] [21])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_4[[21__426 .GSR = "DISABLED";
    FD1P3AX \addr_space_4[[20__428  (.D(wb_odata[20]), .SP(dac_clk_p_c_enable_227), 
            .CK(dac_clk_p_c), .Q(\addr_space[4] [20])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_4[[20__428 .GSR = "DISABLED";
    FD1P3AX \addr_space_4[[19__430  (.D(wb_odata[19]), .SP(dac_clk_p_c_enable_227), 
            .CK(dac_clk_p_c), .Q(\addr_space[4] [19])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_4[[19__430 .GSR = "DISABLED";
    FD1P3AX \addr_space_4[[18__432  (.D(wb_odata[18]), .SP(dac_clk_p_c_enable_227), 
            .CK(dac_clk_p_c), .Q(\addr_space[4] [18])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_4[[18__432 .GSR = "DISABLED";
    FD1P3AX \addr_space_4[[17__434  (.D(wb_odata[17]), .SP(dac_clk_p_c_enable_227), 
            .CK(dac_clk_p_c), .Q(\addr_space[4] [17])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_4[[17__434 .GSR = "DISABLED";
    FD1P3AX \addr_space_4[[16__436  (.D(wb_odata[16]), .SP(dac_clk_p_c_enable_227), 
            .CK(dac_clk_p_c), .Q(\addr_space[4] [16])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_4[[16__436 .GSR = "DISABLED";
    FD1P3AX \addr_space_4[[15__438  (.D(wb_odata[15]), .SP(dac_clk_p_c_enable_227), 
            .CK(dac_clk_p_c), .Q(\addr_space[4] [15])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_4[[15__438 .GSR = "DISABLED";
    FD1P3AX \addr_space_2[[8__324  (.D(wb_odata[8]), .SP(dac_clk_p_c_enable_243), 
            .CK(dac_clk_p_c), .Q(\addr_space[2] [8])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_2[[8__324 .GSR = "DISABLED";
    FD1P3AX \addr_space_4[[14__440  (.D(wb_odata[14]), .SP(dac_clk_p_c_enable_227), 
            .CK(dac_clk_p_c), .Q(\addr_space[4] [14])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_4[[14__440 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[30__181  (.D(wb_odata[30]), .SP(dac_clk_p_c_enable_79), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [30])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_0[[30__181 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[29__182  (.D(wb_odata[29]), .SP(dac_clk_p_c_enable_79), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [29])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_0[[29__182 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[28__183  (.D(wb_odata[28]), .SP(dac_clk_p_c_enable_79), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [28])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_0[[28__183 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[27__184  (.D(wb_odata[27]), .SP(dac_clk_p_c_enable_79), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [27])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_0[[27__184 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[26__185  (.D(wb_odata[26]), .SP(dac_clk_p_c_enable_79), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [26])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_0[[26__185 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[25__186  (.D(wb_odata[25]), .SP(dac_clk_p_c_enable_79), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [25])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_0[[25__186 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[24__187  (.D(wb_odata[24]), .SP(dac_clk_p_c_enable_79), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [24])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_0[[24__187 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[23__188  (.D(wb_odata[23]), .SP(dac_clk_p_c_enable_79), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [23])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_0[[23__188 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[22__189  (.D(wb_odata[22]), .SP(dac_clk_p_c_enable_79), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [22])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_0[[22__189 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[21__190  (.D(wb_odata[21]), .SP(dac_clk_p_c_enable_79), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [21])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_0[[21__190 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[20__191  (.D(wb_odata[20]), .SP(dac_clk_p_c_enable_79), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [20])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_0[[20__191 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[19__192  (.D(wb_odata[19]), .SP(dac_clk_p_c_enable_79), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [19])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_0[[19__192 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[18__193  (.D(wb_odata[18]), .SP(dac_clk_p_c_enable_79), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [18])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_0[[18__193 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[17__194  (.D(wb_odata[17]), .SP(dac_clk_p_c_enable_79), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [17])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_0[[17__194 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[16__195  (.D(wb_odata[16]), .SP(dac_clk_p_c_enable_79), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [16])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_0[[16__195 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[15__196  (.D(wb_odata[15]), .SP(dac_clk_p_c_enable_79), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [15])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_0[[15__196 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[14__197  (.D(wb_odata[14]), .SP(dac_clk_p_c_enable_79), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [14])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_0[[14__197 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[13__198  (.D(wb_odata[13]), .SP(dac_clk_p_c_enable_79), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [13])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_0[[13__198 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[12__199  (.D(wb_odata[12]), .SP(dac_clk_p_c_enable_79), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [12])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_0[[12__199 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[11__200  (.D(wb_odata[11]), .SP(dac_clk_p_c_enable_79), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [11])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_0[[11__200 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[10__201  (.D(wb_odata[10]), .SP(dac_clk_p_c_enable_79), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [10])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_0[[10__201 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[9__202  (.D(wb_odata[9]), .SP(dac_clk_p_c_enable_79), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [9])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_0[[9__202 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[8__203  (.D(wb_odata[8]), .SP(dac_clk_p_c_enable_79), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [8])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_0[[8__203 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[7__204  (.D(wb_odata[7]), .SP(dac_clk_p_c_enable_79), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [7])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_0[[7__204 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[6__205  (.D(wb_odata[6]), .SP(dac_clk_p_c_enable_79), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [6])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_0[[6__205 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[5__206  (.D(wb_odata[5]), .SP(dac_clk_p_c_enable_79), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [5])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_0[[5__206 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[4__207  (.D(wb_odata[4]), .SP(dac_clk_p_c_enable_79), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [4])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_0[[4__207 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[3__208  (.D(wb_odata[3]), .SP(dac_clk_p_c_enable_79), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [3])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_0[[3__208 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[2__209  (.D(wb_odata[2]), .SP(dac_clk_p_c_enable_79), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_0[[2__209 .GSR = "DISABLED";
    FD1P3BX \addr_space_0[[0__212  (.D(wb_odata[0]), .SP(dac_clk_p_c_enable_79), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(lo_i_en)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_0[[0__212 .GSR = "DISABLED";
    FD1P3AX \addr_space_4[[13__442  (.D(wb_odata[13]), .SP(dac_clk_p_c_enable_227), 
            .CK(dac_clk_p_c), .Q(\addr_space[4] [13])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_4[[13__442 .GSR = "DISABLED";
    FD1P3AX \addr_space_4[[12__444  (.D(wb_odata[12]), .SP(dac_clk_p_c_enable_227), 
            .CK(dac_clk_p_c), .Q(\addr_space[4] [12])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_4[[12__444 .GSR = "DISABLED";
    FD1P3AX \addr_space_4[[11__446  (.D(wb_odata[11]), .SP(dac_clk_p_c_enable_227), 
            .CK(dac_clk_p_c), .Q(\addr_space[4] [11])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_4[[11__446 .GSR = "DISABLED";
    FD1P3AX \addr_space_4[[10__448  (.D(wb_odata[10]), .SP(dac_clk_p_c_enable_227), 
            .CK(dac_clk_p_c), .Q(\addr_space[4] [10])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_4[[10__448 .GSR = "DISABLED";
    FD1P3AX \addr_space_4[[9__450  (.D(wb_odata[9]), .SP(dac_clk_p_c_enable_227), 
            .CK(dac_clk_p_c), .Q(\addr_space[4] [9])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_4[[9__450 .GSR = "DISABLED";
    FD1P3AX \addr_space_4[[8__452  (.D(wb_odata[8]), .SP(dac_clk_p_c_enable_227), 
            .CK(dac_clk_p_c), .Q(\addr_space[4] [8])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_4[[8__452 .GSR = "DISABLED";
    FD1P3AX \addr_space_4[[7__454  (.D(wb_odata[7]), .SP(dac_clk_p_c_enable_227), 
            .CK(dac_clk_p_c), .Q(\addr_space[4] [7])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_4[[7__454 .GSR = "DISABLED";
    FD1P3AX \addr_space_4[[6__456  (.D(wb_odata[6]), .SP(dac_clk_p_c_enable_227), 
            .CK(dac_clk_p_c), .Q(\addr_space[4] [6])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_4[[6__456 .GSR = "DISABLED";
    FD1P3AX \addr_space_4[[5__458  (.D(wb_odata[5]), .SP(dac_clk_p_c_enable_227), 
            .CK(dac_clk_p_c), .Q(\addr_space[4] [5])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_4[[5__458 .GSR = "DISABLED";
    FD1P3AX \addr_space_4[[4__460  (.D(wb_odata[4]), .SP(dac_clk_p_c_enable_227), 
            .CK(dac_clk_p_c), .Q(\addr_space[4] [4])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_4[[4__460 .GSR = "DISABLED";
    FD1P3AX \addr_space_4[[3__462  (.D(wb_odata[3]), .SP(dac_clk_p_c_enable_227), 
            .CK(dac_clk_p_c), .Q(\addr_space[4] [3])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_4[[3__462 .GSR = "DISABLED";
    FD1P3AX \addr_space_4[[2__464  (.D(wb_odata[2]), .SP(dac_clk_p_c_enable_227), 
            .CK(dac_clk_p_c), .Q(\addr_space[4] [2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_4[[2__464 .GSR = "DISABLED";
    FD1P3AX \addr_space_4[[1__466  (.D(wb_odata[1]), .SP(dac_clk_p_c_enable_227), 
            .CK(dac_clk_p_c), .Q(\addr_space[4][1] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_4[[1__466 .GSR = "DISABLED";
    FD1P3AX \addr_space_4[[0__468  (.D(wb_odata[0]), .SP(dac_clk_p_c_enable_227), 
            .CK(dac_clk_p_c), .Q(\addr_space[4][0] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_4[[0__468 .GSR = "DISABLED";
    FD1P3AX \addr_space_1[[31__214  (.D(wb_odata[31]), .SP(dac_clk_p_c_enable_106), 
            .CK(dac_clk_p_c), .Q(\addr_space[1] [31])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_1[[31__214 .GSR = "DISABLED";
    FD1P3AX \addr_space_1[[30__216  (.D(wb_odata[30]), .SP(dac_clk_p_c_enable_106), 
            .CK(dac_clk_p_c), .Q(\addr_space[1] [30])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_1[[30__216 .GSR = "DISABLED";
    FD1P3AX \addr_space_2[[7__326  (.D(wb_odata[7]), .SP(dac_clk_p_c_enable_243), 
            .CK(dac_clk_p_c), .Q(\addr_space[2] [7])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_2[[7__326 .GSR = "DISABLED";
    FD1P3AX \addr_space_1[[29__218  (.D(wb_odata[29]), .SP(dac_clk_p_c_enable_106), 
            .CK(dac_clk_p_c), .Q(\addr_space[1] [29])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_1[[29__218 .GSR = "DISABLED";
    FD1P3AX \addr_space_2[[6__328  (.D(wb_odata[6]), .SP(dac_clk_p_c_enable_243), 
            .CK(dac_clk_p_c), .Q(\addr_space[2] [6])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_2[[6__328 .GSR = "DISABLED";
    FD1P3AX \addr_space_1[[28__220  (.D(wb_odata[28]), .SP(dac_clk_p_c_enable_106), 
            .CK(dac_clk_p_c), .Q(\addr_space[1] [28])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_1[[28__220 .GSR = "DISABLED";
    FD1P3AX \addr_space_1[[27__222  (.D(wb_odata[27]), .SP(dac_clk_p_c_enable_106), 
            .CK(dac_clk_p_c), .Q(\addr_space[1] [27])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_1[[27__222 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[10__384  (.D(wb_odata[10]), .SP(dac_clk_p_c_enable_241), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [10])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_3[[10__384 .GSR = "DISABLED";
    FD1P3AX \addr_space_2[[5__330  (.D(wb_odata[5]), .SP(dac_clk_p_c_enable_243), 
            .CK(dac_clk_p_c), .Q(\addr_space[2] [5])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_2[[5__330 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[9__386  (.D(wb_odata[9]), .SP(dac_clk_p_c_enable_241), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [9])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_3[[9__386 .GSR = "DISABLED";
    FD1S3AX o_wb_data_i0 (.D(o_wb_data_31__N_2456[0]), .CK(dac_clk_p_c), 
            .Q(wb_control_data[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(34[8] 36[4])
    defparam o_wb_data_i0.GSR = "DISABLED";
    FD1P3AX \addr_space_2[[4__332  (.D(wb_odata[4]), .SP(dac_clk_p_c_enable_243), 
            .CK(dac_clk_p_c), .Q(\addr_space[2] [4])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_2[[4__332 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[31__180  (.D(wb_odata[31]), .SP(dac_clk_p_c_enable_79), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [31])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_0[[31__180 .GSR = "DISABLED";
    FD1P3BX \addr_space_0[[1__211  (.D(wb_odata[1]), .SP(dac_clk_p_c_enable_79), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(lo_q_en)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_0[[1__211 .GSR = "DISABLED";
    FD1P3AX \addr_space_1[[26__224  (.D(wb_odata[26]), .SP(dac_clk_p_c_enable_106), 
            .CK(dac_clk_p_c), .Q(\addr_space[1] [26])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_1[[26__224 .GSR = "DISABLED";
    FD1P3AX \addr_space_1[[25__226  (.D(wb_odata[25]), .SP(dac_clk_p_c_enable_106), 
            .CK(dac_clk_p_c), .Q(\addr_space[1] [25])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_1[[25__226 .GSR = "DISABLED";
    FD1P3AX \addr_space_1[[24__228  (.D(wb_odata[24]), .SP(dac_clk_p_c_enable_106), 
            .CK(dac_clk_p_c), .Q(\addr_space[1] [24])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_1[[24__228 .GSR = "DISABLED";
    FD1P3AX \addr_space_1[[23__230  (.D(wb_odata[23]), .SP(dac_clk_p_c_enable_106), 
            .CK(dac_clk_p_c), .Q(\addr_space[1] [23])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_1[[23__230 .GSR = "DISABLED";
    FD1P3AX \addr_space_1[[22__232  (.D(wb_odata[22]), .SP(dac_clk_p_c_enable_106), 
            .CK(dac_clk_p_c), .Q(\addr_space[1] [22])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_1[[22__232 .GSR = "DISABLED";
    FD1P3AX \addr_space_1[[21__234  (.D(wb_odata[21]), .SP(dac_clk_p_c_enable_106), 
            .CK(dac_clk_p_c), .Q(\addr_space[1] [21])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_1[[21__234 .GSR = "DISABLED";
    FD1P3AX \addr_space_1[[20__236  (.D(wb_odata[20]), .SP(dac_clk_p_c_enable_106), 
            .CK(dac_clk_p_c), .Q(\addr_space[1] [20])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_1[[20__236 .GSR = "DISABLED";
    FD1P3AX \addr_space_1[[19__238  (.D(wb_odata[19]), .SP(dac_clk_p_c_enable_106), 
            .CK(dac_clk_p_c), .Q(\addr_space[1] [19])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_1[[19__238 .GSR = "DISABLED";
    FD1P3AX \addr_space_1[[18__240  (.D(wb_odata[18]), .SP(dac_clk_p_c_enable_106), 
            .CK(dac_clk_p_c), .Q(\addr_space[1] [18])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_1[[18__240 .GSR = "DISABLED";
    FD1P3AX \addr_space_1[[17__242  (.D(wb_odata[17]), .SP(dac_clk_p_c_enable_106), 
            .CK(dac_clk_p_c), .Q(\addr_space[1] [17])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_1[[17__242 .GSR = "DISABLED";
    FD1P3AX \addr_space_1[[16__244  (.D(wb_odata[16]), .SP(dac_clk_p_c_enable_106), 
            .CK(dac_clk_p_c), .Q(\addr_space[1] [16])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_1[[16__244 .GSR = "DISABLED";
    FD1P3AX \addr_space_1[[15__246  (.D(wb_odata[15]), .SP(dac_clk_p_c_enable_106), 
            .CK(dac_clk_p_c), .Q(\addr_space[1] [15])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_1[[15__246 .GSR = "DISABLED";
    FD1P3AX \addr_space_1[[14__248  (.D(wb_odata[14]), .SP(dac_clk_p_c_enable_106), 
            .CK(dac_clk_p_c), .Q(\addr_space[1] [14])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_1[[14__248 .GSR = "DISABLED";
    FD1P3AX \addr_space_1[[13__250  (.D(wb_odata[13]), .SP(dac_clk_p_c_enable_106), 
            .CK(dac_clk_p_c), .Q(\addr_space[1] [13])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_1[[13__250 .GSR = "DISABLED";
    FD1P3AX \addr_space_1[[12__252  (.D(wb_odata[12]), .SP(dac_clk_p_c_enable_106), 
            .CK(dac_clk_p_c), .Q(\addr_space[1] [12])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_1[[12__252 .GSR = "DISABLED";
    FD1P3AX \addr_space_1[[11__254  (.D(wb_odata[11]), .SP(dac_clk_p_c_enable_106), 
            .CK(dac_clk_p_c), .Q(\addr_space[1] [11])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_1[[11__254 .GSR = "DISABLED";
    FD1P3AX \addr_space_1[[10__256  (.D(wb_odata[10]), .SP(dac_clk_p_c_enable_106), 
            .CK(dac_clk_p_c), .Q(\addr_space[1] [10])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_1[[10__256 .GSR = "DISABLED";
    FD1P3AX \addr_space_1[[9__258  (.D(wb_odata[9]), .SP(dac_clk_p_c_enable_106), 
            .CK(dac_clk_p_c), .Q(\addr_space[1] [9])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_1[[9__258 .GSR = "DISABLED";
    FD1P3AX \addr_space_1[[8__260  (.D(wb_odata[8]), .SP(dac_clk_p_c_enable_106), 
            .CK(dac_clk_p_c), .Q(\addr_space[1] [8])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_1[[8__260 .GSR = "DISABLED";
    FD1P3AX \addr_space_1[[7__262  (.D(wb_odata[7]), .SP(dac_clk_p_c_enable_106), 
            .CK(dac_clk_p_c), .Q(\addr_space[1] [7])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_1[[7__262 .GSR = "DISABLED";
    FD1P3AX \addr_space_1[[6__264  (.D(wb_odata[6]), .SP(dac_clk_p_c_enable_106), 
            .CK(dac_clk_p_c), .Q(\addr_space[1] [6])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_1[[6__264 .GSR = "DISABLED";
    FD1P3AX \addr_space_1[[5__266  (.D(wb_odata[5]), .SP(dac_clk_p_c_enable_106), 
            .CK(dac_clk_p_c), .Q(\addr_space[1] [5])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_1[[5__266 .GSR = "DISABLED";
    FD1P3AX \addr_space_1[[4__268  (.D(wb_odata[4]), .SP(dac_clk_p_c_enable_106), 
            .CK(dac_clk_p_c), .Q(\addr_space[1] [4])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_1[[4__268 .GSR = "DISABLED";
    FD1P3AX \addr_space_1[[3__270  (.D(wb_odata[3]), .SP(dac_clk_p_c_enable_106), 
            .CK(dac_clk_p_c), .Q(\addr_space[1] [3])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_1[[3__270 .GSR = "DISABLED";
    FD1P3AX \addr_space_1[[2__272  (.D(wb_odata[2]), .SP(dac_clk_p_c_enable_106), 
            .CK(dac_clk_p_c), .Q(\addr_space[1] [2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_1[[2__272 .GSR = "DISABLED";
    FD1P3AX \addr_space_1[[1__274  (.D(wb_odata[1]), .SP(dac_clk_p_c_enable_106), 
            .CK(dac_clk_p_c), .Q(\addr_space[1][1] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_1[[1__274 .GSR = "DISABLED";
    FD1P3AX \addr_space_1[[0__276  (.D(wb_odata[0]), .SP(dac_clk_p_c_enable_106), 
            .CK(dac_clk_p_c), .Q(\addr_space[1][0] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_1[[0__276 .GSR = "DISABLED";
    FD1P3AX \addr_space_2[[31__278  (.D(wb_odata[31]), .SP(dac_clk_p_c_enable_243), 
            .CK(dac_clk_p_c), .Q(\addr_space[2] [31])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_2[[31__278 .GSR = "DISABLED";
    FD1P3AX \addr_space_2[[30__280  (.D(wb_odata[30]), .SP(dac_clk_p_c_enable_243), 
            .CK(dac_clk_p_c), .Q(\addr_space[2] [30])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_2[[30__280 .GSR = "DISABLED";
    FD1P3AX \addr_space_2[[29__282  (.D(wb_odata[29]), .SP(dac_clk_p_c_enable_243), 
            .CK(dac_clk_p_c), .Q(\addr_space[2] [29])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_2[[29__282 .GSR = "DISABLED";
    FD1P3AX \addr_space_2[[28__284  (.D(wb_odata[28]), .SP(dac_clk_p_c_enable_243), 
            .CK(dac_clk_p_c), .Q(\addr_space[2] [28])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_2[[28__284 .GSR = "DISABLED";
    FD1P3AX \addr_space_2[[27__286  (.D(wb_odata[27]), .SP(dac_clk_p_c_enable_243), 
            .CK(dac_clk_p_c), .Q(\addr_space[2] [27])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_2[[27__286 .GSR = "DISABLED";
    FD1P3AX \addr_space_2[[26__288  (.D(wb_odata[26]), .SP(dac_clk_p_c_enable_243), 
            .CK(dac_clk_p_c), .Q(\addr_space[2] [26])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_2[[26__288 .GSR = "DISABLED";
    FD1P3AX \addr_space_2[[25__290  (.D(wb_odata[25]), .SP(dac_clk_p_c_enable_243), 
            .CK(dac_clk_p_c), .Q(\addr_space[2] [25])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_2[[25__290 .GSR = "DISABLED";
    FD1P3AX \addr_space_2[[24__292  (.D(wb_odata[24]), .SP(dac_clk_p_c_enable_243), 
            .CK(dac_clk_p_c), .Q(\addr_space[2] [24])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_2[[24__292 .GSR = "DISABLED";
    FD1P3AX \addr_space_2[[23__294  (.D(wb_odata[23]), .SP(dac_clk_p_c_enable_243), 
            .CK(dac_clk_p_c), .Q(\addr_space[2] [23])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_2[[23__294 .GSR = "DISABLED";
    FD1P3AX \addr_space_2[[22__296  (.D(wb_odata[22]), .SP(dac_clk_p_c_enable_243), 
            .CK(dac_clk_p_c), .Q(\addr_space[2] [22])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_2[[22__296 .GSR = "DISABLED";
    FD1P3AX \addr_space_2[[21__298  (.D(wb_odata[21]), .SP(dac_clk_p_c_enable_243), 
            .CK(dac_clk_p_c), .Q(\addr_space[2] [21])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_2[[21__298 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[8__388  (.D(wb_odata[8]), .SP(dac_clk_p_c_enable_241), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [8])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_3[[8__388 .GSR = "DISABLED";
    FD1P3AX \addr_space_2[[3__334  (.D(wb_odata[3]), .SP(dac_clk_p_c_enable_243), 
            .CK(dac_clk_p_c), .Q(\addr_space[2] [3])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_2[[3__334 .GSR = "DISABLED";
    FD1P3AX \addr_space_2[[9__322  (.D(wb_odata[9]), .SP(dac_clk_p_c_enable_243), 
            .CK(dac_clk_p_c), .Q(\addr_space[2] [9])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_2[[9__322 .GSR = "DISABLED";
    FD1P3AX \addr_space_2[[20__300  (.D(wb_odata[20]), .SP(dac_clk_p_c_enable_243), 
            .CK(dac_clk_p_c), .Q(\addr_space[2] [20])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_2[[20__300 .GSR = "DISABLED";
    FD1P3AX \addr_space_2[[2__336  (.D(wb_odata[2]), .SP(dac_clk_p_c_enable_243), 
            .CK(dac_clk_p_c), .Q(\addr_space[2] [2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_2[[2__336 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[7__390  (.D(wb_odata[7]), .SP(dac_clk_p_c_enable_241), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [7])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_3[[7__390 .GSR = "DISABLED";
    FD1P3AX \addr_space_2[[1__338  (.D(wb_odata[1]), .SP(dac_clk_p_c_enable_243), 
            .CK(dac_clk_p_c), .Q(\addr_space[2][1] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_2[[1__338 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[6__392  (.D(wb_odata[6]), .SP(dac_clk_p_c_enable_241), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [6])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_3[[6__392 .GSR = "DISABLED";
    FD1P3AX \addr_space_2[[0__340  (.D(wb_odata[0]), .SP(dac_clk_p_c_enable_243), 
            .CK(dac_clk_p_c), .Q(\addr_space[2][0] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_2[[0__340 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[5__394  (.D(wb_odata[5]), .SP(dac_clk_p_c_enable_241), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [5])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_3[[5__394 .GSR = "DISABLED";
    FD1P3AX \addr_space_2[[19__302  (.D(wb_odata[19]), .SP(dac_clk_p_c_enable_243), 
            .CK(dac_clk_p_c), .Q(\addr_space[2] [19])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_2[[19__302 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[31__342  (.D(wb_odata[31]), .SP(dac_clk_p_c_enable_241), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [31])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_3[[31__342 .GSR = "DISABLED";
    FD1P3AX \addr_space_2[[18__304  (.D(wb_odata[18]), .SP(dac_clk_p_c_enable_243), 
            .CK(dac_clk_p_c), .Q(\addr_space[2] [18])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_2[[18__304 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[4__396  (.D(wb_odata[4]), .SP(dac_clk_p_c_enable_241), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [4])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_3[[4__396 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[30__344  (.D(wb_odata[30]), .SP(dac_clk_p_c_enable_241), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [30])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_3[[30__344 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[29__346  (.D(wb_odata[29]), .SP(dac_clk_p_c_enable_241), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [29])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_3[[29__346 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[3__398  (.D(wb_odata[3]), .SP(dac_clk_p_c_enable_241), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [3])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_3[[3__398 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[28__348  (.D(wb_odata[28]), .SP(dac_clk_p_c_enable_241), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [28])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_3[[28__348 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[2__400  (.D(wb_odata[2]), .SP(dac_clk_p_c_enable_241), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_3[[2__400 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[27__350  (.D(wb_odata[27]), .SP(dac_clk_p_c_enable_241), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [27])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_3[[27__350 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[1__402  (.D(wb_odata[1]), .SP(dac_clk_p_c_enable_241), 
            .CK(dac_clk_p_c), .Q(\addr_space[3][1] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_3[[1__402 .GSR = "DISABLED";
    LUT4 n26891_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4] [10]), .C(\wb_addr[2] ), 
         .D(n26891), .Z(o_wb_data_31__N_2456_c[10])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n26891_bdd_3_lut_4_lut.init = 16'h8f80;
    FD1P3AX \addr_space_2[[17__306  (.D(wb_odata[17]), .SP(dac_clk_p_c_enable_243), 
            .CK(dac_clk_p_c), .Q(\addr_space[2] [17])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_2[[17__306 .GSR = "DISABLED";
    FD1P3AX \addr_space_2[[16__308  (.D(wb_odata[16]), .SP(dac_clk_p_c_enable_243), 
            .CK(dac_clk_p_c), .Q(\addr_space[2] [16])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_2[[16__308 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[26__352  (.D(wb_odata[26]), .SP(dac_clk_p_c_enable_241), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [26])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_3[[26__352 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[0__404  (.D(wb_odata[0]), .SP(dac_clk_p_c_enable_241), 
            .CK(dac_clk_p_c), .Q(\addr_space[3][0] )) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_3[[0__404 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[25__354  (.D(wb_odata[25]), .SP(dac_clk_p_c_enable_241), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [25])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_3[[25__354 .GSR = "DISABLED";
    FD1P3AX \addr_space_4[[31__406  (.D(wb_odata[31]), .SP(dac_clk_p_c_enable_227), 
            .CK(dac_clk_p_c), .Q(\addr_space[4] [31])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_4[[31__406 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[24__356  (.D(wb_odata[24]), .SP(dac_clk_p_c_enable_241), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [24])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_3[[24__356 .GSR = "DISABLED";
    FD1P3AX \addr_space_4[[30__408  (.D(wb_odata[30]), .SP(dac_clk_p_c_enable_227), 
            .CK(dac_clk_p_c), .Q(\addr_space[4] [30])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_4[[30__408 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[23__358  (.D(wb_odata[23]), .SP(dac_clk_p_c_enable_241), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [23])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_3[[23__358 .GSR = "DISABLED";
    FD1S3IX o_wb_ack_470 (.D(wb_control_data_31__N_35), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(wb_control_ack)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(38[8] 43[4])
    defparam o_wb_ack_470.GSR = "DISABLED";
    FD1P3AX \addr_space_4[[29__410  (.D(wb_odata[29]), .SP(dac_clk_p_c_enable_227), 
            .CK(dac_clk_p_c), .Q(\addr_space[4] [29])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_4[[29__410 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[22__360  (.D(wb_odata[22]), .SP(dac_clk_p_c_enable_241), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [22])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_3[[22__360 .GSR = "DISABLED";
    FD1P3AX \addr_space_4[[28__412  (.D(wb_odata[28]), .SP(dac_clk_p_c_enable_227), 
            .CK(dac_clk_p_c), .Q(\addr_space[4] [28])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_4[[28__412 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[21__362  (.D(wb_odata[21]), .SP(dac_clk_p_c_enable_241), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [21])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_3[[21__362 .GSR = "DISABLED";
    FD1P3AX \addr_space_4[[27__414  (.D(wb_odata[27]), .SP(dac_clk_p_c_enable_227), 
            .CK(dac_clk_p_c), .Q(\addr_space[4] [27])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_4[[27__414 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[20__364  (.D(wb_odata[20]), .SP(dac_clk_p_c_enable_241), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [20])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_3[[20__364 .GSR = "DISABLED";
    FD1P3AX \addr_space_4[[26__416  (.D(wb_odata[26]), .SP(dac_clk_p_c_enable_227), 
            .CK(dac_clk_p_c), .Q(\addr_space[4] [26])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_4[[26__416 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[19__366  (.D(wb_odata[19]), .SP(dac_clk_p_c_enable_241), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [19])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_3[[19__366 .GSR = "DISABLED";
    FD1P3AX \addr_space_4[[25__418  (.D(wb_odata[25]), .SP(dac_clk_p_c_enable_227), 
            .CK(dac_clk_p_c), .Q(\addr_space[4] [25])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_4[[25__418 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[18__368  (.D(wb_odata[18]), .SP(dac_clk_p_c_enable_241), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [18])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_3[[18__368 .GSR = "DISABLED";
    FD1P3AX \addr_space_4[[24__420  (.D(wb_odata[24]), .SP(dac_clk_p_c_enable_227), 
            .CK(dac_clk_p_c), .Q(\addr_space[4] [24])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_4[[24__420 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[17__370  (.D(wb_odata[17]), .SP(dac_clk_p_c_enable_241), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [17])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_3[[17__370 .GSR = "DISABLED";
    FD1P3AX \addr_space_4[[23__422  (.D(wb_odata[23]), .SP(dac_clk_p_c_enable_227), 
            .CK(dac_clk_p_c), .Q(\addr_space[4] [23])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_4[[23__422 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[16__372  (.D(wb_odata[16]), .SP(dac_clk_p_c_enable_241), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [16])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_3[[16__372 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[15__374  (.D(wb_odata[15]), .SP(dac_clk_p_c_enable_241), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [15])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_3[[15__374 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[14__376  (.D(wb_odata[14]), .SP(dac_clk_p_c_enable_241), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [14])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_3[[14__376 .GSR = "DISABLED";
    FD1P3AX \addr_space_2[[15__310  (.D(wb_odata[15]), .SP(dac_clk_p_c_enable_243), 
            .CK(dac_clk_p_c), .Q(\addr_space[2] [15])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_2[[15__310 .GSR = "DISABLED";
    FD1P3AX \addr_space_2[[14__312  (.D(wb_odata[14]), .SP(dac_clk_p_c_enable_243), 
            .CK(dac_clk_p_c), .Q(\addr_space[2] [14])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_2[[14__312 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[13__378  (.D(wb_odata[13]), .SP(dac_clk_p_c_enable_241), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [13])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_3[[13__378 .GSR = "DISABLED";
    FD1P3AX \addr_space_2[[13__314  (.D(wb_odata[13]), .SP(dac_clk_p_c_enable_243), 
            .CK(dac_clk_p_c), .Q(\addr_space[2] [13])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_2[[13__314 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[12__380  (.D(wb_odata[12]), .SP(dac_clk_p_c_enable_241), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [12])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_3[[12__380 .GSR = "DISABLED";
    FD1P3AX \addr_space_2[[12__316  (.D(wb_odata[12]), .SP(dac_clk_p_c_enable_243), 
            .CK(dac_clk_p_c), .Q(\addr_space[2] [12])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_2[[12__316 .GSR = "DISABLED";
    LUT4 n26886_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4] [11]), .C(\wb_addr[2] ), 
         .D(n26886), .Z(o_wb_data_31__N_2456_c[11])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n26886_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 n26875_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4] [12]), .C(\wb_addr[2] ), 
         .D(n26875), .Z(o_wb_data_31__N_2456_c[12])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n26875_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 n26863_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4] [13]), .C(\wb_addr[2] ), 
         .D(n26863), .Z(o_wb_data_31__N_2456_c[13])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n26863_bdd_3_lut_4_lut.init = 16'h8f80;
    FD1P3AX \addr_space_3[[11__382  (.D(wb_odata[11]), .SP(dac_clk_p_c_enable_241), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [11])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_3[[11__382 .GSR = "DISABLED";
    FD1P3AX \addr_space_2[[11__318  (.D(wb_odata[11]), .SP(dac_clk_p_c_enable_243), 
            .CK(dac_clk_p_c), .Q(\addr_space[2] [11])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_2[[11__318 .GSR = "DISABLED";
    LUT4 n26858_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4] [14]), .C(\wb_addr[2] ), 
         .D(n26858), .Z(o_wb_data_31__N_2456_c[14])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n26858_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 i24654_4_lut (.A(n21662), .B(n29302), .C(n29065), .D(n22526), 
         .Z(dac_clk_p_c_enable_79)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(28[3] 30[6])
    defparam i24654_4_lut.init = 16'h0004;
    FD1P3AX \addr_space_2[[10__320  (.D(wb_odata[10]), .SP(dac_clk_p_c_enable_243), 
            .CK(dac_clk_p_c), .Q(\addr_space[2] [10])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam \addr_space_2[[10__320 .GSR = "DISABLED";
    LUT4 n26842_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4] [15]), .C(\wb_addr[2] ), 
         .D(n26842), .Z(o_wb_data_31__N_2456_c[15])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n26842_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 n26831_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4] [16]), .C(\wb_addr[2] ), 
         .D(n26831), .Z(o_wb_data_31__N_2456_c[16])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n26831_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 n26826_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4] [17]), .C(\wb_addr[2] ), 
         .D(n26826), .Z(o_wb_data_31__N_2456_c[17])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n26826_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 n26817_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4] [18]), .C(\wb_addr[2] ), 
         .D(n26817), .Z(o_wb_data_31__N_2456_c[18])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n26817_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 n26812_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4] [19]), .C(\wb_addr[2] ), 
         .D(n26812), .Z(o_wb_data_31__N_2456_c[19])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n26812_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 n26807_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4] [20]), .C(\wb_addr[2] ), 
         .D(n26807), .Z(o_wb_data_31__N_2456_c[20])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n26807_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 n26802_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4] [21]), .C(\wb_addr[2] ), 
         .D(n26802), .Z(o_wb_data_31__N_2456_c[21])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n26802_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 n26789_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4] [22]), .C(\wb_addr[2] ), 
         .D(n26789), .Z(o_wb_data_31__N_2456_c[22])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n26789_bdd_3_lut_4_lut.init = 16'h8f80;
    FD1S3AX o_wb_data_i31 (.D(o_wb_data_31__N_2456_c[31]), .CK(dac_clk_p_c), 
            .Q(wb_control_data[31])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(34[8] 36[4])
    defparam o_wb_data_i31.GSR = "DISABLED";
    FD1S3AX o_wb_data_i30 (.D(o_wb_data_31__N_2456_c[30]), .CK(dac_clk_p_c), 
            .Q(wb_control_data[30])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(34[8] 36[4])
    defparam o_wb_data_i30.GSR = "DISABLED";
    FD1S3AX o_wb_data_i29 (.D(o_wb_data_31__N_2456_c[29]), .CK(dac_clk_p_c), 
            .Q(wb_control_data[29])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(34[8] 36[4])
    defparam o_wb_data_i29.GSR = "DISABLED";
    FD1S3AX o_wb_data_i28 (.D(o_wb_data_31__N_2456_c[28]), .CK(dac_clk_p_c), 
            .Q(wb_control_data[28])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(34[8] 36[4])
    defparam o_wb_data_i28.GSR = "DISABLED";
    FD1S3AX o_wb_data_i27 (.D(o_wb_data_31__N_2456_c[27]), .CK(dac_clk_p_c), 
            .Q(wb_control_data[27])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(34[8] 36[4])
    defparam o_wb_data_i27.GSR = "DISABLED";
    FD1S3AX o_wb_data_i26 (.D(o_wb_data_31__N_2456_c[26]), .CK(dac_clk_p_c), 
            .Q(wb_control_data[26])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(34[8] 36[4])
    defparam o_wb_data_i26.GSR = "DISABLED";
    FD1S3AX o_wb_data_i25 (.D(o_wb_data_31__N_2456_c[25]), .CK(dac_clk_p_c), 
            .Q(wb_control_data[25])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(34[8] 36[4])
    defparam o_wb_data_i25.GSR = "DISABLED";
    FD1S3AX o_wb_data_i24 (.D(o_wb_data_31__N_2456_c[24]), .CK(dac_clk_p_c), 
            .Q(wb_control_data[24])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(34[8] 36[4])
    defparam o_wb_data_i24.GSR = "DISABLED";
    FD1S3AX o_wb_data_i23 (.D(o_wb_data_31__N_2456_c[23]), .CK(dac_clk_p_c), 
            .Q(wb_control_data[23])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(34[8] 36[4])
    defparam o_wb_data_i23.GSR = "DISABLED";
    FD1S3AX o_wb_data_i22 (.D(o_wb_data_31__N_2456_c[22]), .CK(dac_clk_p_c), 
            .Q(wb_control_data[22])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(34[8] 36[4])
    defparam o_wb_data_i22.GSR = "DISABLED";
    FD1S3AX o_wb_data_i21 (.D(o_wb_data_31__N_2456_c[21]), .CK(dac_clk_p_c), 
            .Q(wb_control_data[21])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(34[8] 36[4])
    defparam o_wb_data_i21.GSR = "DISABLED";
    FD1S3AX o_wb_data_i20 (.D(o_wb_data_31__N_2456_c[20]), .CK(dac_clk_p_c), 
            .Q(wb_control_data[20])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(34[8] 36[4])
    defparam o_wb_data_i20.GSR = "DISABLED";
    FD1S3AX o_wb_data_i19 (.D(o_wb_data_31__N_2456_c[19]), .CK(dac_clk_p_c), 
            .Q(wb_control_data[19])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(34[8] 36[4])
    defparam o_wb_data_i19.GSR = "DISABLED";
    FD1S3AX o_wb_data_i18 (.D(o_wb_data_31__N_2456_c[18]), .CK(dac_clk_p_c), 
            .Q(wb_control_data[18])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(34[8] 36[4])
    defparam o_wb_data_i18.GSR = "DISABLED";
    FD1S3AX o_wb_data_i17 (.D(o_wb_data_31__N_2456_c[17]), .CK(dac_clk_p_c), 
            .Q(wb_control_data[17])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(34[8] 36[4])
    defparam o_wb_data_i17.GSR = "DISABLED";
    FD1S3AX o_wb_data_i16 (.D(o_wb_data_31__N_2456_c[16]), .CK(dac_clk_p_c), 
            .Q(wb_control_data[16])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(34[8] 36[4])
    defparam o_wb_data_i16.GSR = "DISABLED";
    FD1S3AX o_wb_data_i15 (.D(o_wb_data_31__N_2456_c[15]), .CK(dac_clk_p_c), 
            .Q(wb_control_data[15])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(34[8] 36[4])
    defparam o_wb_data_i15.GSR = "DISABLED";
    FD1S3AX o_wb_data_i14 (.D(o_wb_data_31__N_2456_c[14]), .CK(dac_clk_p_c), 
            .Q(wb_control_data[14])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(34[8] 36[4])
    defparam o_wb_data_i14.GSR = "DISABLED";
    FD1S3AX o_wb_data_i13 (.D(o_wb_data_31__N_2456_c[13]), .CK(dac_clk_p_c), 
            .Q(wb_control_data[13])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(34[8] 36[4])
    defparam o_wb_data_i13.GSR = "DISABLED";
    FD1S3AX o_wb_data_i12 (.D(o_wb_data_31__N_2456_c[12]), .CK(dac_clk_p_c), 
            .Q(wb_control_data[12])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(34[8] 36[4])
    defparam o_wb_data_i12.GSR = "DISABLED";
    LUT4 n26777_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4] [23]), .C(\wb_addr[2] ), 
         .D(n26777), .Z(o_wb_data_31__N_2456_c[23])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n26777_bdd_3_lut_4_lut.init = 16'h8f80;
    FD1S3AX o_wb_data_i11 (.D(o_wb_data_31__N_2456_c[11]), .CK(dac_clk_p_c), 
            .Q(wb_control_data[11])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(34[8] 36[4])
    defparam o_wb_data_i11.GSR = "DISABLED";
    FD1S3AX o_wb_data_i10 (.D(o_wb_data_31__N_2456_c[10]), .CK(dac_clk_p_c), 
            .Q(wb_control_data[10])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(34[8] 36[4])
    defparam o_wb_data_i10.GSR = "DISABLED";
    FD1S3AX o_wb_data_i9 (.D(o_wb_data_31__N_2456_c[9]), .CK(dac_clk_p_c), 
            .Q(wb_control_data[9])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(34[8] 36[4])
    defparam o_wb_data_i9.GSR = "DISABLED";
    FD1S3AX o_wb_data_i8 (.D(o_wb_data_31__N_2456_c[8]), .CK(dac_clk_p_c), 
            .Q(wb_control_data[8])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(34[8] 36[4])
    defparam o_wb_data_i8.GSR = "DISABLED";
    FD1S3AX o_wb_data_i7 (.D(o_wb_data_31__N_2456_c[7]), .CK(dac_clk_p_c), 
            .Q(wb_control_data[7])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(34[8] 36[4])
    defparam o_wb_data_i7.GSR = "DISABLED";
    FD1S3AX o_wb_data_i6 (.D(o_wb_data_31__N_2456_c[6]), .CK(dac_clk_p_c), 
            .Q(wb_control_data[6])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(34[8] 36[4])
    defparam o_wb_data_i6.GSR = "DISABLED";
    FD1S3AX o_wb_data_i5 (.D(o_wb_data_31__N_2456_c[5]), .CK(dac_clk_p_c), 
            .Q(wb_control_data[5])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(34[8] 36[4])
    defparam o_wb_data_i5.GSR = "DISABLED";
    FD1S3AX o_wb_data_i4 (.D(o_wb_data_31__N_2456_c[4]), .CK(dac_clk_p_c), 
            .Q(wb_control_data[4])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(34[8] 36[4])
    defparam o_wb_data_i4.GSR = "DISABLED";
    FD1S3AX o_wb_data_i3 (.D(o_wb_data_31__N_2456_c[3]), .CK(dac_clk_p_c), 
            .Q(wb_control_data[3])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(34[8] 36[4])
    defparam o_wb_data_i3.GSR = "DISABLED";
    FD1S3AX o_wb_data_i2 (.D(o_wb_data_31__N_2456_c[2]), .CK(dac_clk_p_c), 
            .Q(wb_control_data[2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(34[8] 36[4])
    defparam o_wb_data_i2.GSR = "DISABLED";
    FD1S3AX o_wb_data_i1 (.D(\o_wb_data_31__N_2456[1] ), .CK(dac_clk_p_c), 
            .Q(wb_control_data[1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=2, LSE_LLINE=204, LSE_RLINE=216 */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(34[8] 36[4])
    defparam o_wb_data_i1.GSR = "DISABLED";
    LUT4 n26759_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4] [24]), .C(\wb_addr[2] ), 
         .D(n26759), .Z(o_wb_data_31__N_2456_c[24])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n26759_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 \addr_space_0[[31__bdd_3_lut_25053  (.A(\addr_space[1] [31]), .B(\addr_space[3] [31]), 
         .C(\wb_addr[1] ), .Z(n26699)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[31__bdd_3_lut_25053 .init = 16'hcaca;
    LUT4 \addr_space_0[[31__bdd_3_lut_26939  (.A(\addr_space[0] [31]), .B(\addr_space[2] [31]), 
         .C(\wb_addr[1] ), .Z(n26700)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[31__bdd_3_lut_26939 .init = 16'hcaca;
    LUT4 n26750_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4] [25]), .C(\wb_addr[2] ), 
         .D(n26750), .Z(o_wb_data_31__N_2456_c[25])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n26750_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 \addr_space_0[[30__bdd_3_lut_25057  (.A(\addr_space[1] [30]), .B(\addr_space[3] [30]), 
         .C(\wb_addr[1] ), .Z(n26704)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[30__bdd_3_lut_25057 .init = 16'hcaca;
    LUT4 \addr_space_0[[30__bdd_3_lut_26935  (.A(\addr_space[0] [30]), .B(\addr_space[2] [30]), 
         .C(\wb_addr[1] ), .Z(n26705)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[30__bdd_3_lut_26935 .init = 16'hcaca;
    LUT4 \addr_space_0[[29__bdd_3_lut_25061  (.A(\addr_space[1] [29]), .B(\addr_space[3] [29]), 
         .C(\wb_addr[1] ), .Z(n26709)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[29__bdd_3_lut_25061 .init = 16'hcaca;
    LUT4 \addr_space_0[[29__bdd_3_lut_26931  (.A(\addr_space[0] [29]), .B(\addr_space[2] [29]), 
         .C(\wb_addr[1] ), .Z(n26710)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[29__bdd_3_lut_26931 .init = 16'hcaca;
    LUT4 \addr_space_0[[28__bdd_3_lut_25065  (.A(\addr_space[1] [28]), .B(\addr_space[3] [28]), 
         .C(\wb_addr[1] ), .Z(n26714)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[28__bdd_3_lut_25065 .init = 16'hcaca;
    LUT4 \addr_space_0[[28__bdd_3_lut_26908  (.A(\addr_space[0] [28]), .B(\addr_space[2] [28]), 
         .C(\wb_addr[1] ), .Z(n26715)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[28__bdd_3_lut_26908 .init = 16'hcaca;
    LUT4 n26739_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4] [26]), .C(\wb_addr[2] ), 
         .D(n26739), .Z(o_wb_data_31__N_2456_c[26])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n26739_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 \addr_space_0[[27__bdd_3_lut_25084  (.A(\addr_space[1] [27]), .B(\addr_space[3] [27]), 
         .C(\wb_addr[1] ), .Z(n26732)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[27__bdd_3_lut_25084 .init = 16'hcaca;
    LUT4 \addr_space_0[[27__bdd_3_lut_26817  (.A(\addr_space[0] [27]), .B(\addr_space[2] [27]), 
         .C(\wb_addr[1] ), .Z(n26733)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[27__bdd_3_lut_26817 .init = 16'hcaca;
    LUT4 \addr_space_0[[26__bdd_3_lut_25088  (.A(\addr_space[1] [26]), .B(\addr_space[3] [26]), 
         .C(\wb_addr[1] ), .Z(n26737)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[26__bdd_3_lut_25088 .init = 16'hcaca;
    LUT4 \addr_space_0[[26__bdd_3_lut_26798  (.A(\addr_space[0] [26]), .B(\addr_space[2] [26]), 
         .C(\wb_addr[1] ), .Z(n26738)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[26__bdd_3_lut_26798 .init = 16'hcaca;
    LUT4 n26734_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4] [27]), .C(\wb_addr[2] ), 
         .D(n26734), .Z(o_wb_data_31__N_2456_c[27])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n26734_bdd_3_lut_4_lut.init = 16'h8f80;
    PFUMX i25263 (.BLUT(n26939), .ALUT(n26938), .C0(\wb_addr[0] ), .Z(n26940));
    LUT4 \addr_space_0[[25__bdd_3_lut_25099  (.A(\addr_space[1] [25]), .B(\addr_space[3] [25]), 
         .C(\wb_addr[1] ), .Z(n26748)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[25__bdd_3_lut_25099 .init = 16'hcaca;
    PFUMX i25259 (.BLUT(n26934), .ALUT(n26933), .C0(\wb_addr[0] ), .Z(n26935));
    PFUMX i25255 (.BLUT(n26929), .ALUT(n26928), .C0(\wb_addr[0] ), .Z(n26930));
    LUT4 \addr_space_0[[25__bdd_3_lut_26246  (.A(\addr_space[0] [25]), .B(\addr_space[2] [25]), 
         .C(\wb_addr[1] ), .Z(n26749)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[25__bdd_3_lut_26246 .init = 16'hcaca;
    PFUMX i25251 (.BLUT(n26924), .ALUT(n26923), .C0(\wb_addr[0] ), .Z(n26925));
    LUT4 n26716_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4] [28]), .C(\wb_addr[2] ), 
         .D(n26716), .Z(o_wb_data_31__N_2456_c[28])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n26716_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 n26711_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4] [29]), .C(\wb_addr[2] ), 
         .D(n26711), .Z(o_wb_data_31__N_2456_c[29])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n26711_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 n26706_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4] [30]), .C(\wb_addr[2] ), 
         .D(n26706), .Z(o_wb_data_31__N_2456_c[30])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n26706_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 n26701_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4] [31]), .C(\wb_addr[2] ), 
         .D(n26701), .Z(o_wb_data_31__N_2456_c[31])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n26701_bdd_3_lut_4_lut.init = 16'h8f80;
    PFUMX i25247 (.BLUT(n26919), .ALUT(n26918), .C0(\wb_addr[0] ), .Z(n26920));
    LUT4 \addr_space_0[[24__bdd_3_lut_25107  (.A(\addr_space[1] [24]), .B(\addr_space[3] [24]), 
         .C(\wb_addr[1] ), .Z(n26757)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[24__bdd_3_lut_25107 .init = 16'hcaca;
    LUT4 \addr_space_0[[24__bdd_3_lut_25958  (.A(\addr_space[0] [24]), .B(\addr_space[2] [24]), 
         .C(\wb_addr[1] ), .Z(n26758)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[24__bdd_3_lut_25958 .init = 16'hcaca;
    PFUMX i25243 (.BLUT(n26914), .ALUT(n26913), .C0(\wb_addr[0] ), .Z(n26915));
    PFUMX i25239 (.BLUT(n26909), .ALUT(n26908), .C0(\wb_addr[0] ), .Z(n26910));
    LUT4 \addr_space_0[[23__bdd_3_lut_25123  (.A(\addr_space[1] [23]), .B(\addr_space[3] [23]), 
         .C(\wb_addr[1] ), .Z(n26775)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[23__bdd_3_lut_25123 .init = 16'hcaca;
    LUT4 \addr_space_0[[23__bdd_3_lut_25949  (.A(\addr_space[0] [23]), .B(\addr_space[2] [23]), 
         .C(\wb_addr[1] ), .Z(n26776)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[23__bdd_3_lut_25949 .init = 16'hcaca;
    PFUMX i25226 (.BLUT(n26895), .ALUT(n26894), .C0(\wb_addr[0] ), .Z(n26896));
    PFUMX i25222 (.BLUT(n26890), .ALUT(n26889), .C0(\wb_addr[0] ), .Z(n26891));
    LUT4 \addr_space_0[[22__bdd_3_lut_25132  (.A(\addr_space[1] [22]), .B(\addr_space[3] [22]), 
         .C(\wb_addr[1] ), .Z(n26787)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[22__bdd_3_lut_25132 .init = 16'hcaca;
    LUT4 \addr_space_0[[22__bdd_3_lut_25938  (.A(\addr_space[0] [22]), .B(\addr_space[2] [22]), 
         .C(\wb_addr[1] ), .Z(n26788)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[22__bdd_3_lut_25938 .init = 16'hcaca;
    PFUMX i25218 (.BLUT(n26885), .ALUT(n26884), .C0(\wb_addr[0] ), .Z(n26886));
    LUT4 \addr_space_0[[21__bdd_3_lut_25926  (.A(\addr_space[0] [21]), .B(\addr_space[2] [21]), 
         .C(\wb_addr[1] ), .Z(n26801)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[21__bdd_3_lut_25926 .init = 16'hcaca;
    LUT4 \addr_space_0[[21__bdd_3_lut_25142  (.A(\addr_space[1] [21]), .B(\addr_space[3] [21]), 
         .C(\wb_addr[1] ), .Z(n26800)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[21__bdd_3_lut_25142 .init = 16'hcaca;
    LUT4 \addr_space_0[[20__bdd_3_lut_25146  (.A(\addr_space[1] [20]), .B(\addr_space[3] [20]), 
         .C(\wb_addr[1] ), .Z(n26805)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[20__bdd_3_lut_25146 .init = 16'hcaca;
    LUT4 \addr_space_0[[20__bdd_3_lut_25913  (.A(\addr_space[0] [20]), .B(\addr_space[2] [20]), 
         .C(\wb_addr[1] ), .Z(n26806)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[20__bdd_3_lut_25913 .init = 16'hcaca;
    LUT4 \addr_space_0[[19__bdd_3_lut_25150  (.A(\addr_space[1] [19]), .B(\addr_space[3] [19]), 
         .C(\wb_addr[1] ), .Z(n26810)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[19__bdd_3_lut_25150 .init = 16'hcaca;
    LUT4 \addr_space_0[[19__bdd_3_lut_25909  (.A(\addr_space[0] [19]), .B(\addr_space[2] [19]), 
         .C(\wb_addr[1] ), .Z(n26811)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[19__bdd_3_lut_25909 .init = 16'hcaca;
    PFUMX i25209 (.BLUT(n26874), .ALUT(n26873), .C0(\wb_addr[0] ), .Z(n26875));
    LUT4 \addr_space_0[[18__bdd_3_lut_25154  (.A(\addr_space[1] [18]), .B(\addr_space[3] [18]), 
         .C(\wb_addr[1] ), .Z(n26815)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[18__bdd_3_lut_25154 .init = 16'hcaca;
    LUT4 \addr_space_0[[18__bdd_3_lut_25902  (.A(\addr_space[0] [18]), .B(\addr_space[2] [18]), 
         .C(\wb_addr[1] ), .Z(n26816)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[18__bdd_3_lut_25902 .init = 16'hcaca;
    LUT4 \addr_space_0[[17__bdd_3_lut_25876  (.A(\addr_space[0] [17]), .B(\addr_space[2] [17]), 
         .C(\wb_addr[1] ), .Z(n26825)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[17__bdd_3_lut_25876 .init = 16'hcaca;
    LUT4 \addr_space_0[[17__bdd_3_lut_25162  (.A(\addr_space[1] [17]), .B(\addr_space[3] [17]), 
         .C(\wb_addr[1] ), .Z(n26824)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[17__bdd_3_lut_25162 .init = 16'hcaca;
    LUT4 \addr_space_0[[16__bdd_3_lut_25166  (.A(\addr_space[1] [16]), .B(\addr_space[3] [16]), 
         .C(\wb_addr[1] ), .Z(n26829)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[16__bdd_3_lut_25166 .init = 16'hcaca;
    PFUMX i25198 (.BLUT(n26862), .ALUT(n26861), .C0(\wb_addr[0] ), .Z(n26863));
    LUT4 \addr_space_0[[16__bdd_3_lut_25869  (.A(\addr_space[0] [16]), .B(\addr_space[2] [16]), 
         .C(\wb_addr[1] ), .Z(n26830)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[16__bdd_3_lut_25869 .init = 16'hcaca;
    PFUMX i25194 (.BLUT(n26857), .ALUT(n26856), .C0(\wb_addr[0] ), .Z(n26858));
    LUT4 \addr_space_0[[15__bdd_3_lut_25863  (.A(\addr_space[0] [15]), .B(\addr_space[2] [15]), 
         .C(\wb_addr[1] ), .Z(n26841)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[15__bdd_3_lut_25863 .init = 16'hcaca;
    LUT4 \addr_space_0[[15__bdd_3_lut_25177  (.A(\addr_space[1] [15]), .B(\addr_space[3] [15]), 
         .C(\wb_addr[1] ), .Z(n26840)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[15__bdd_3_lut_25177 .init = 16'hcaca;
    PFUMX i25178 (.BLUT(n26841), .ALUT(n26840), .C0(\wb_addr[0] ), .Z(n26842));
    LUT4 \addr_space_0[[14__bdd_3_lut_25193  (.A(\addr_space[1] [14]), .B(\addr_space[3] [14]), 
         .C(\wb_addr[1] ), .Z(n26856)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[14__bdd_3_lut_25193 .init = 16'hcaca;
    LUT4 \addr_space_0[[14__bdd_3_lut_25800  (.A(\addr_space[0] [14]), .B(\addr_space[2] [14]), 
         .C(\wb_addr[1] ), .Z(n26857)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[14__bdd_3_lut_25800 .init = 16'hcaca;
    LUT4 \addr_space_0[[13__bdd_3_lut_25197  (.A(\addr_space[1] [13]), .B(\addr_space[3] [13]), 
         .C(\wb_addr[1] ), .Z(n26861)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[13__bdd_3_lut_25197 .init = 16'hcaca;
    LUT4 \addr_space_0[[13__bdd_3_lut_25794  (.A(\addr_space[0] [13]), .B(\addr_space[2] [13]), 
         .C(\wb_addr[1] ), .Z(n26862)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[13__bdd_3_lut_25794 .init = 16'hcaca;
    PFUMX i25167 (.BLUT(n26830), .ALUT(n26829), .C0(\wb_addr[0] ), .Z(n26831));
    LUT4 \addr_space_0[[12__bdd_3_lut_25208  (.A(\addr_space[1] [12]), .B(\addr_space[3] [12]), 
         .C(\wb_addr[1] ), .Z(n26873)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[12__bdd_3_lut_25208 .init = 16'hcaca;
    LUT4 \addr_space_0[[12__bdd_3_lut_25781  (.A(\addr_space[0] [12]), .B(\addr_space[2] [12]), 
         .C(\wb_addr[1] ), .Z(n26874)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[12__bdd_3_lut_25781 .init = 16'hcaca;
    LUT4 \addr_space_0[[11__bdd_3_lut_25752  (.A(\addr_space[0] [11]), .B(\addr_space[2] [11]), 
         .C(\wb_addr[1] ), .Z(n26885)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[11__bdd_3_lut_25752 .init = 16'hcaca;
    PFUMX i25163 (.BLUT(n26825), .ALUT(n26824), .C0(\wb_addr[0] ), .Z(n26826));
    LUT4 \addr_space_0[[11__bdd_3_lut_25217  (.A(\addr_space[1] [11]), .B(\addr_space[3] [11]), 
         .C(\wb_addr[1] ), .Z(n26884)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[11__bdd_3_lut_25217 .init = 16'hcaca;
    PFUMX i25155 (.BLUT(n26816), .ALUT(n26815), .C0(\wb_addr[0] ), .Z(n26817));
    PFUMX i25151 (.BLUT(n26811), .ALUT(n26810), .C0(\wb_addr[0] ), .Z(n26812));
    LUT4 \addr_space_0[[10__bdd_3_lut_25221  (.A(\addr_space[1] [10]), .B(\addr_space[3] [10]), 
         .C(\wb_addr[1] ), .Z(n26889)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[10__bdd_3_lut_25221 .init = 16'hcaca;
    LUT4 \addr_space_0[[10__bdd_3_lut_25739  (.A(\addr_space[0] [10]), .B(\addr_space[2] [10]), 
         .C(\wb_addr[1] ), .Z(n26890)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[10__bdd_3_lut_25739 .init = 16'hcaca;
    PFUMX i25147 (.BLUT(n26806), .ALUT(n26805), .C0(\wb_addr[0] ), .Z(n26807));
    LUT4 \addr_space_0[[9__bdd_3_lut_25225  (.A(\addr_space[1] [9]), .B(\addr_space[3] [9]), 
         .C(\wb_addr[1] ), .Z(n26894)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[9__bdd_3_lut_25225 .init = 16'hcaca;
    LUT4 \addr_space_0[[9__bdd_3_lut_25728  (.A(\addr_space[0] [9]), .B(\addr_space[2] [9]), 
         .C(\wb_addr[1] ), .Z(n26895)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[9__bdd_3_lut_25728 .init = 16'hcaca;
    LUT4 \addr_space_0[[8__bdd_3_lut_25719  (.A(\addr_space[0] [8]), .B(\addr_space[2] [8]), 
         .C(\wb_addr[1] ), .Z(n26909)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[8__bdd_3_lut_25719 .init = 16'hcaca;
    LUT4 \addr_space_0[[8__bdd_3_lut_25238  (.A(\addr_space[1] [8]), .B(\addr_space[3] [8]), 
         .C(\wb_addr[1] ), .Z(n26908)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[8__bdd_3_lut_25238 .init = 16'hcaca;
    LUT4 \addr_space_0[[7__bdd_3_lut_25242  (.A(\addr_space[1] [7]), .B(\addr_space[3] [7]), 
         .C(\wb_addr[1] ), .Z(n26913)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[7__bdd_3_lut_25242 .init = 16'hcaca;
    LUT4 \addr_space_0[[7__bdd_3_lut_25705  (.A(\addr_space[0] [7]), .B(\addr_space[2] [7]), 
         .C(\wb_addr[1] ), .Z(n26914)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[7__bdd_3_lut_25705 .init = 16'hcaca;
    PFUMX i25143 (.BLUT(n26801), .ALUT(n26800), .C0(\wb_addr[0] ), .Z(n26802));
    PFUMX i25133 (.BLUT(n26788), .ALUT(n26787), .C0(\wb_addr[0] ), .Z(n26789));
    LUT4 \addr_space_0[[6__bdd_3_lut_25246  (.A(\addr_space[1] [6]), .B(\addr_space[3] [6]), 
         .C(\wb_addr[1] ), .Z(n26918)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[6__bdd_3_lut_25246 .init = 16'hcaca;
    LUT4 \addr_space_0[[6__bdd_3_lut_25699  (.A(\addr_space[0] [6]), .B(\addr_space[2] [6]), 
         .C(\wb_addr[1] ), .Z(n26919)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[6__bdd_3_lut_25699 .init = 16'hcaca;
    LUT4 \addr_space_0[[5__bdd_3_lut_25250  (.A(\addr_space[1] [5]), .B(\addr_space[3] [5]), 
         .C(\wb_addr[1] ), .Z(n26923)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[5__bdd_3_lut_25250 .init = 16'hcaca;
    LUT4 \addr_space_0[[5__bdd_3_lut_25695  (.A(\addr_space[0] [5]), .B(\addr_space[2] [5]), 
         .C(\wb_addr[1] ), .Z(n26924)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[5__bdd_3_lut_25695 .init = 16'hcaca;
    LUT4 \addr_space_0[[4__bdd_3_lut_25254  (.A(\addr_space[1] [4]), .B(\addr_space[3] [4]), 
         .C(\wb_addr[1] ), .Z(n26928)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[4__bdd_3_lut_25254 .init = 16'hcaca;
    LUT4 \addr_space_0[[4__bdd_3_lut_25691  (.A(\addr_space[0] [4]), .B(\addr_space[2] [4]), 
         .C(\wb_addr[1] ), .Z(n26929)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[4__bdd_3_lut_25691 .init = 16'hcaca;
    LUT4 \addr_space_0[[3__bdd_3_lut_25258  (.A(\addr_space[1] [3]), .B(\addr_space[3] [3]), 
         .C(\wb_addr[1] ), .Z(n26933)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[3__bdd_3_lut_25258 .init = 16'hcaca;
    LUT4 \addr_space_0[[3__bdd_3_lut_25683  (.A(\addr_space[0] [3]), .B(\addr_space[2] [3]), 
         .C(\wb_addr[1] ), .Z(n26934)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[3__bdd_3_lut_25683 .init = 16'hcaca;
    PFUMX i25124 (.BLUT(n26776), .ALUT(n26775), .C0(\wb_addr[0] ), .Z(n26777));
    LUT4 \addr_space_0[[2__bdd_3_lut_25262  (.A(\addr_space[1] [2]), .B(\addr_space[3] [2]), 
         .C(\wb_addr[1] ), .Z(n26938)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[2__bdd_3_lut_25262 .init = 16'hcaca;
    LUT4 \addr_space_0[[2__bdd_3_lut_25671  (.A(\addr_space[0] [2]), .B(\addr_space[2] [2]), 
         .C(\wb_addr[1] ), .Z(n26939)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[2__bdd_3_lut_25671 .init = 16'hcaca;
    PFUMX i25108 (.BLUT(n26758), .ALUT(n26757), .C0(\wb_addr[0] ), .Z(n26759));
    PFUMX i25100 (.BLUT(n26749), .ALUT(n26748), .C0(\wb_addr[0] ), .Z(n26750));
    LUT4 n26915_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4] [7]), .C(\wb_addr[2] ), 
         .D(n26915), .Z(o_wb_data_31__N_2456_c[7])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n26915_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 n26910_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4] [8]), .C(\wb_addr[2] ), 
         .D(n26910), .Z(o_wb_data_31__N_2456_c[8])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n26910_bdd_3_lut_4_lut.init = 16'h8f80;
    PFUMX i25089 (.BLUT(n26738), .ALUT(n26737), .C0(\wb_addr[0] ), .Z(n26739));
    PFUMX i25085 (.BLUT(n26733), .ALUT(n26732), .C0(\wb_addr[0] ), .Z(n26734));
    PFUMX i25066 (.BLUT(n26715), .ALUT(n26714), .C0(\wb_addr[0] ), .Z(n26716));
    LUT4 i1_2_lut (.A(lo_q_en), .B(lo_q), .Z(o_lo_q_c)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/control.v(27[11] 31[5])
    defparam i1_2_lut.init = 16'h8888;
    PFUMX i25062 (.BLUT(n26710), .ALUT(n26709), .C0(\wb_addr[0] ), .Z(n26711));
    PFUMX i25058 (.BLUT(n26705), .ALUT(n26704), .C0(\wb_addr[0] ), .Z(n26706));
    PFUMX i25054 (.BLUT(n26700), .ALUT(n26699), .C0(\wb_addr[0] ), .Z(n26701));
    LUT4 n26940_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4] [2]), .C(\wb_addr[2] ), 
         .D(n26940), .Z(o_wb_data_31__N_2456_c[2])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n26940_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 n26935_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4] [3]), .C(\wb_addr[2] ), 
         .D(n26935), .Z(o_wb_data_31__N_2456_c[3])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n26935_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 n26930_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4] [4]), .C(\wb_addr[2] ), 
         .D(n26930), .Z(o_wb_data_31__N_2456_c[4])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n26930_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 n26925_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4] [5]), .C(\wb_addr[2] ), 
         .D(n26925), .Z(o_wb_data_31__N_2456_c[5])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n26925_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 n26896_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4] [9]), .C(\wb_addr[2] ), 
         .D(n26896), .Z(o_wb_data_31__N_2456_c[9])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n26896_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 n26920_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4] [6]), .C(\wb_addr[2] ), 
         .D(n26920), .Z(o_wb_data_31__N_2456_c[6])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n26920_bdd_3_lut_4_lut.init = 16'h8f80;
    
endmodule
//
// Verilog Description of module hbbus
//

module hbbus (dac_clk_p_c, wb_cyc, wb_we, wb_odata, wb_stb, wb_addr, 
            GND_net, wb_ack, \wb_idata[0] , \wb_idata[2] , \wb_idata[3] , 
            \wb_idata[4] , \wb_idata[5] , \wb_idata[6] , \wb_idata[7] , 
            \wb_idata[8] , \wb_idata[9] , \wb_idata[10] , \wb_idata[11] , 
            \wb_idata[12] , \wb_idata[13] , \wb_idata[14] , \wb_idata[15] , 
            \wb_idata[16] , \wb_idata[17] , \wb_idata[18] , \wb_idata[19] , 
            \wb_idata[20] , \wb_idata[21] , \wb_idata[22] , \wb_idata[23] , 
            \wb_idata[24] , \wb_idata[25] , \wb_idata[26] , \wb_idata[27] , 
            \wb_idata[28] , wb_err, \wb_idata[29] , \wb_idata[30] , 
            \wb_idata[31] , n2, n14148, n32067, VCC_net, \rx_data[1] , 
            \rx_data[2] , \rx_data[0] , \rx_data[3] , \rx_data[5] , 
            \rx_data[6] , \rx_data[4] , rx_stb, \tx_data[1] , \tx_data[2] , 
            \tx_data[3] , \tx_data[4] , \tx_data[5] , \tx_data[6] , 
            tx_stb, \tx_data[0] , tx_busy) /* synthesis syn_module_defined=1 */ ;
    input dac_clk_p_c;
    output wb_cyc;
    output wb_we;
    output [31:0]wb_odata;
    output wb_stb;
    output [29:0]wb_addr;
    input GND_net;
    input wb_ack;
    input \wb_idata[0] ;
    input \wb_idata[2] ;
    input \wb_idata[3] ;
    input \wb_idata[4] ;
    input \wb_idata[5] ;
    input \wb_idata[6] ;
    input \wb_idata[7] ;
    input \wb_idata[8] ;
    input \wb_idata[9] ;
    input \wb_idata[10] ;
    input \wb_idata[11] ;
    input \wb_idata[12] ;
    input \wb_idata[13] ;
    input \wb_idata[14] ;
    input \wb_idata[15] ;
    input \wb_idata[16] ;
    input \wb_idata[17] ;
    input \wb_idata[18] ;
    input \wb_idata[19] ;
    input \wb_idata[20] ;
    input \wb_idata[21] ;
    input \wb_idata[22] ;
    input \wb_idata[23] ;
    input \wb_idata[24] ;
    input \wb_idata[25] ;
    input \wb_idata[26] ;
    input \wb_idata[27] ;
    input \wb_idata[28] ;
    input wb_err;
    input \wb_idata[29] ;
    input \wb_idata[30] ;
    input \wb_idata[31] ;
    output n2;
    input n14148;
    input n32067;
    input VCC_net;
    input \rx_data[1] ;
    input \rx_data[2] ;
    input \rx_data[0] ;
    input \rx_data[3] ;
    input \rx_data[5] ;
    input \rx_data[6] ;
    input \rx_data[4] ;
    input rx_stb;
    output \tx_data[1] ;
    output \tx_data[2] ;
    output \tx_data[3] ;
    output \tx_data[4] ;
    output \tx_data[5] ;
    output \tx_data[6] ;
    output tx_stb;
    output \tx_data[0] ;
    input tx_busy;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[29:38])
    wire [33:0]iw_word;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(71[14:21])
    
    wire ow_stb;
    wire [33:0]ow_word;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(73[14:21])
    
    wire n32126, iw_stb, n32125;
    wire [4:0]hb_bits;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(79[13:20])
    
    wire dac_clk_p_c_enable_312, hb_busy, w_reset;
    wire [33:0]idl_word;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(77[14:22])
    
    wire nl_busy, hx_stb, idl_stb, dac_clk_p_c_enable_548, cmd_loaded, 
        dac_clk_p_c_enable_166, cmd_loaded_N_535, o_pck_stb_N_532;
    wire [4:0]dec_bits;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(69[13:21])
    
    wire dac_clk_p_c_enable_517;
    wire [33:0]n14;
    wire [7:0]w_gx_char;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbgenhex.v(80[12:21])
    
    wire int_stb, n29458;
    wire [33:0]int_word;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(75[14:22])
    
    hbexec wbexec (.dac_clk_p_c(dac_clk_p_c), .wb_cyc(wb_cyc), .wb_we(wb_we), 
           .wb_odata({wb_odata}), .iw_word({iw_word}), .ow_stb(ow_stb), 
           .ow_word({ow_word}), .n32126(n32126), .iw_stb(iw_stb), .wb_stb(wb_stb), 
           .wb_addr({wb_addr}), .GND_net(GND_net), .wb_ack(wb_ack), .\wb_idata[0] (\wb_idata[0] ), 
           .\wb_idata[2] (\wb_idata[2] ), .\wb_idata[3] (\wb_idata[3] ), 
           .\wb_idata[4] (\wb_idata[4] ), .\wb_idata[5] (\wb_idata[5] ), 
           .\wb_idata[6] (\wb_idata[6] ), .\wb_idata[7] (\wb_idata[7] ), 
           .\wb_idata[8] (\wb_idata[8] ), .\wb_idata[9] (\wb_idata[9] ), 
           .\wb_idata[10] (\wb_idata[10] ), .\wb_idata[11] (\wb_idata[11] ), 
           .\wb_idata[12] (\wb_idata[12] ), .\wb_idata[13] (\wb_idata[13] ), 
           .\wb_idata[14] (\wb_idata[14] ), .\wb_idata[15] (\wb_idata[15] ), 
           .\wb_idata[16] (\wb_idata[16] ), .\wb_idata[17] (\wb_idata[17] ), 
           .\wb_idata[18] (\wb_idata[18] ), .\wb_idata[19] (\wb_idata[19] ), 
           .\wb_idata[20] (\wb_idata[20] ), .\wb_idata[21] (\wb_idata[21] ), 
           .\wb_idata[22] (\wb_idata[22] ), .\wb_idata[23] (\wb_idata[23] ), 
           .\wb_idata[24] (\wb_idata[24] ), .\wb_idata[25] (\wb_idata[25] ), 
           .\wb_idata[26] (\wb_idata[26] ), .\wb_idata[27] (\wb_idata[27] ), 
           .\wb_idata[28] (\wb_idata[28] ), .wb_err(wb_err), .\wb_idata[29] (\wb_idata[29] ), 
           .\wb_idata[30] (\wb_idata[30] ), .\wb_idata[31] (\wb_idata[31] ), 
           .n2(n2), .n32125(n32125), .n14148(n14148)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(105[15] 109[15])
    hbdeword unpackx (.hb_bits({hb_bits}), .dac_clk_p_c(dac_clk_p_c), .dac_clk_p_c_enable_312(dac_clk_p_c_enable_312), 
            .n32067(n32067), .n32126(n32126), .hb_busy(hb_busy), .w_reset(w_reset), 
            .idl_word({idl_word}), .n32125(n32125), .nl_busy(nl_busy), 
            .hx_stb(hx_stb), .idl_stb(idl_stb)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(127[11] 129[29])
    hbpack packxi (.iw_word({iw_word}), .dac_clk_p_c(dac_clk_p_c), .dac_clk_p_c_enable_548(dac_clk_p_c_enable_548), 
           .n32126(n32126), .cmd_loaded(cmd_loaded), .dac_clk_p_c_enable_166(dac_clk_p_c_enable_166), 
           .w_reset(w_reset), .cmd_loaded_N_535(cmd_loaded_N_535), .iw_stb(iw_stb), 
           .o_pck_stb_N_532(o_pck_stb_N_532), .\dec_bits[0] (dec_bits[0]), 
           .\dec_bits[4] (dec_bits[4]), .dac_clk_p_c_enable_517(dac_clk_p_c_enable_517), 
           .\dec_bits[1] (dec_bits[1]), .n45(n14[3]), .n46(n14[2])) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(99[9] 100[38])
    hbgenhex genhex (.hx_stb(hx_stb), .dac_clk_p_c(dac_clk_p_c), .n32126(n32126), 
            .hb_busy(hb_busy), .hb_bits({hb_bits}), .\w_gx_char[0] (w_gx_char[0]), 
            .\w_gx_char[1] (w_gx_char[1]), .\w_gx_char[2] (w_gx_char[2]), 
            .\w_gx_char[3] (w_gx_char[3]), .\w_gx_char[4] (w_gx_char[4]), 
            .\w_gx_char[5] (w_gx_char[5]), .\w_gx_char[6] (w_gx_char[6]), 
            .dac_clk_p_c_enable_312(dac_clk_p_c_enable_312), .GND_net(GND_net), 
            .VCC_net(VCC_net), .nl_busy(nl_busy), .n32125(n32125)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(132[11] 133[29])
    hbdechex dechxi (.dec_bits({dec_bits[4], Open_31, Open_32, Open_33, 
            dec_bits[0]}), .dac_clk_p_c(dac_clk_p_c), .w_reset(w_reset), 
            .n32126(n32126), .\rx_data[1] (\rx_data[1] ), .\rx_data[2] (\rx_data[2] ), 
            .\rx_data[0] (\rx_data[0] ), .\rx_data[3] (\rx_data[3] ), .\rx_data[5] (\rx_data[5] ), 
            .\rx_data[6] (\rx_data[6] ), .\rx_data[4] (\rx_data[4] ), .rx_stb(rx_stb), 
            .\dec_bits[1] (dec_bits[1]), .n32125(n32125), .dac_clk_p_c_enable_548(dac_clk_p_c_enable_548), 
            .dac_clk_p_c_enable_517(dac_clk_p_c_enable_517), .n45(n14[3]), 
            .n46(n14[2]), .dac_clk_p_c_enable_166(dac_clk_p_c_enable_166), 
            .cmd_loaded_N_535(cmd_loaded_N_535), .cmd_loaded(cmd_loaded), 
            .o_pck_stb_N_532(o_pck_stb_N_532)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(93[11] 95[30])
    hbnewline addnl (.\tx_data[1] (\tx_data[1] ), .dac_clk_p_c(dac_clk_p_c), 
            .w_reset(w_reset), .\tx_data[2] (\tx_data[2] ), .\tx_data[3] (\tx_data[3] ), 
            .\tx_data[4] (\tx_data[4] ), .\tx_data[5] (\tx_data[5] ), .\tx_data[6] (\tx_data[6] ), 
            .n32126(n32126), .tx_stb(tx_stb), .\tx_data[0] (\tx_data[0] ), 
            .\w_gx_char[2] (w_gx_char[2]), .\w_gx_char[3] (w_gx_char[3]), 
            .\w_gx_char[0] (w_gx_char[0]), .\w_gx_char[4] (w_gx_char[4]), 
            .\w_gx_char[1] (w_gx_char[1]), .\w_gx_char[5] (w_gx_char[5]), 
            .\w_gx_char[6] (w_gx_char[6]), .tx_busy(tx_busy), .nl_busy(nl_busy), 
            .hx_stb(hx_stb), .n32125(n32125)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(138[12] 139[40])
    hbints addints (.int_stb(int_stb), .dac_clk_p_c(dac_clk_p_c), .n32126(n32126), 
           .n32125(n32125), .n29458(n29458), .int_word({int_word}), .ow_word({ow_word}), 
           .ow_stb(ow_stb)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(114[9] 116[32])
    hbidle addidles (.idl_word({idl_word}), .dac_clk_p_c(dac_clk_p_c), .int_word({int_word}), 
           .idl_stb(idl_stb), .hb_busy(hb_busy), .n29458(n29458), .int_stb(int_stb), 
           .n32126(n32126), .n32125(n32125)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(121[9] 123[31])
    
endmodule
//
// Verilog Description of module hbexec
//

module hbexec (dac_clk_p_c, wb_cyc, wb_we, wb_odata, iw_word, ow_stb, 
            ow_word, n32126, iw_stb, wb_stb, wb_addr, GND_net, wb_ack, 
            \wb_idata[0] , \wb_idata[2] , \wb_idata[3] , \wb_idata[4] , 
            \wb_idata[5] , \wb_idata[6] , \wb_idata[7] , \wb_idata[8] , 
            \wb_idata[9] , \wb_idata[10] , \wb_idata[11] , \wb_idata[12] , 
            \wb_idata[13] , \wb_idata[14] , \wb_idata[15] , \wb_idata[16] , 
            \wb_idata[17] , \wb_idata[18] , \wb_idata[19] , \wb_idata[20] , 
            \wb_idata[21] , \wb_idata[22] , \wb_idata[23] , \wb_idata[24] , 
            \wb_idata[25] , \wb_idata[26] , \wb_idata[27] , \wb_idata[28] , 
            wb_err, \wb_idata[29] , \wb_idata[30] , \wb_idata[31] , 
            n2, n32125, n14148) /* synthesis syn_module_defined=1 */ ;
    input dac_clk_p_c;
    output wb_cyc;
    output wb_we;
    output [31:0]wb_odata;
    input [33:0]iw_word;
    output ow_stb;
    output [33:0]ow_word;
    input n32126;
    input iw_stb;
    output wb_stb;
    output [29:0]wb_addr;
    input GND_net;
    input wb_ack;
    input \wb_idata[0] ;
    input \wb_idata[2] ;
    input \wb_idata[3] ;
    input \wb_idata[4] ;
    input \wb_idata[5] ;
    input \wb_idata[6] ;
    input \wb_idata[7] ;
    input \wb_idata[8] ;
    input \wb_idata[9] ;
    input \wb_idata[10] ;
    input \wb_idata[11] ;
    input \wb_idata[12] ;
    input \wb_idata[13] ;
    input \wb_idata[14] ;
    input \wb_idata[15] ;
    input \wb_idata[16] ;
    input \wb_idata[17] ;
    input \wb_idata[18] ;
    input \wb_idata[19] ;
    input \wb_idata[20] ;
    input \wb_idata[21] ;
    input \wb_idata[22] ;
    input \wb_idata[23] ;
    input \wb_idata[24] ;
    input \wb_idata[25] ;
    input \wb_idata[26] ;
    input \wb_idata[27] ;
    input \wb_idata[28] ;
    input wb_err;
    input \wb_idata[29] ;
    input \wb_idata[30] ;
    input \wb_idata[31] ;
    output n2;
    input n32125;
    input n14148;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[29:38])
    
    wire newaddr, newaddr_N_757, inc, dac_clk_p_c_enable_60, i_cmd_word_0__N_762, 
        o_cmd_busy_N_698, i_cmd_wr, n29398, o_rsp_stb_N_754;
    wire [33:0]n338;
    wire [33:0]o_rsp_word_33__N_718;
    
    wire n29457, n19882, n19187, n19185;
    wire [29:0]n125;
    
    wire n19881, n19191, n19189, n19880, n19195, n19193, n19879, 
        n19199, n19197, n19878, n19203, n19201, n19877, n19207, 
        n19205, n19876, n19211, n19209, n19875, n19215, n19213, 
        n19874, n19219, n19217, n19873, n19223, n19221, n21661, 
        n24010, n19872, n19227, n19225, n19871, n19231, n19229, 
        n19870, n19235, n19233, n19869, n19239, n19237, n19868, 
        n19242, n19241;
    wire [32:0]n1639;
    
    wire n3, dac_clk_p_c_enable_631, o_cmd_busy_N_708, n29456, o_cmd_busy_N_700, 
        dac_clk_p_c_enable_640, n22149;
    
    FD1S3IX newaddr_72 (.D(newaddr_N_757), .CK(dac_clk_p_c), .CD(wb_cyc), 
            .Q(newaddr)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(192[9] 236[5])
    defparam newaddr_72.GSR = "DISABLED";
    FD1P3AX inc_71 (.D(i_cmd_word_0__N_762), .SP(dac_clk_p_c_enable_60), 
            .CK(dac_clk_p_c), .Q(inc)) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(192[9] 236[5])
    defparam inc_71.GSR = "DISABLED";
    FD1P3AX o_wb_we_69 (.D(i_cmd_wr), .SP(o_cmd_busy_N_698), .CK(dac_clk_p_c), 
            .Q(wb_we)) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(184[9] 186[26])
    defparam o_wb_we_69.GSR = "DISABLED";
    FD1S3AX o_wb_data_i0 (.D(iw_word[0]), .CK(dac_clk_p_c), .Q(wb_odata[0])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i0.GSR = "DISABLED";
    FD1S3JX o_rsp_stb_74 (.D(o_rsp_stb_N_754), .CK(dac_clk_p_c), .PD(n29398), 
            .Q(ow_stb)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_stb_74.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i0 (.D(n338[0]), .CK(dac_clk_p_c), .CD(n29398), 
            .Q(ow_word[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i0.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i2 (.D(n338[2]), .CK(dac_clk_p_c), .CD(n29398), 
            .Q(ow_word[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i2.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i3 (.D(n338[3]), .CK(dac_clk_p_c), .CD(n29398), 
            .Q(ow_word[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i3.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i4 (.D(n338[4]), .CK(dac_clk_p_c), .CD(n29398), 
            .Q(ow_word[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i4.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i5 (.D(n338[5]), .CK(dac_clk_p_c), .CD(n29398), 
            .Q(ow_word[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i5.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i6 (.D(n338[6]), .CK(dac_clk_p_c), .CD(n29398), 
            .Q(ow_word[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i6.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i7 (.D(n338[7]), .CK(dac_clk_p_c), .CD(n29398), 
            .Q(ow_word[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i7.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i8 (.D(n338[8]), .CK(dac_clk_p_c), .CD(n29398), 
            .Q(ow_word[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i8.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i9 (.D(n338[9]), .CK(dac_clk_p_c), .CD(n29398), 
            .Q(ow_word[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i9.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i10 (.D(n338[10]), .CK(dac_clk_p_c), .CD(n29398), 
            .Q(ow_word[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i10.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i11 (.D(n338[11]), .CK(dac_clk_p_c), .CD(n29398), 
            .Q(ow_word[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i11.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i12 (.D(n338[12]), .CK(dac_clk_p_c), .CD(n29398), 
            .Q(ow_word[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i12.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i13 (.D(n338[13]), .CK(dac_clk_p_c), .CD(n29398), 
            .Q(ow_word[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i13.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i14 (.D(n338[14]), .CK(dac_clk_p_c), .CD(n29398), 
            .Q(ow_word[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i14.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i15 (.D(n338[15]), .CK(dac_clk_p_c), .CD(n29398), 
            .Q(ow_word[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i15.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i16 (.D(n338[16]), .CK(dac_clk_p_c), .CD(n29398), 
            .Q(ow_word[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i16.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i17 (.D(n338[17]), .CK(dac_clk_p_c), .CD(n29398), 
            .Q(ow_word[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i17.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i18 (.D(n338[18]), .CK(dac_clk_p_c), .CD(n29398), 
            .Q(ow_word[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i18.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i19 (.D(n338[19]), .CK(dac_clk_p_c), .CD(n29398), 
            .Q(ow_word[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i19.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i20 (.D(n338[20]), .CK(dac_clk_p_c), .CD(n29398), 
            .Q(ow_word[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i20.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i21 (.D(n338[21]), .CK(dac_clk_p_c), .CD(n29398), 
            .Q(ow_word[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i21.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i22 (.D(n338[22]), .CK(dac_clk_p_c), .CD(n29398), 
            .Q(ow_word[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i22.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i23 (.D(n338[23]), .CK(dac_clk_p_c), .CD(n29398), 
            .Q(ow_word[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i23.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i24 (.D(n338[24]), .CK(dac_clk_p_c), .CD(n29398), 
            .Q(ow_word[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i24.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i25 (.D(n338[25]), .CK(dac_clk_p_c), .CD(n29398), 
            .Q(ow_word[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i25.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i26 (.D(n338[26]), .CK(dac_clk_p_c), .CD(n29398), 
            .Q(ow_word[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i26.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i27 (.D(n338[27]), .CK(dac_clk_p_c), .CD(n29398), 
            .Q(ow_word[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i27.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i28 (.D(n338[28]), .CK(dac_clk_p_c), .CD(n29398), 
            .Q(ow_word[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i28.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i29 (.D(o_rsp_word_33__N_718[29]), .CK(dac_clk_p_c), 
            .CD(n32126), .Q(ow_word[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i29.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i30 (.D(n338[30]), .CK(dac_clk_p_c), .CD(n29398), 
            .Q(ow_word[30])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i30.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i31 (.D(n338[31]), .CK(dac_clk_p_c), .CD(n29398), 
            .Q(ow_word[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i31.GSR = "DISABLED";
    FD1S3JX o_rsp_word_i32 (.D(n338[32]), .CK(dac_clk_p_c), .PD(n29398), 
            .Q(ow_word[32])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i32.GSR = "DISABLED";
    FD1S3JX o_rsp_word_i33 (.D(o_cmd_busy_N_698), .CK(dac_clk_p_c), .PD(n29398), 
            .Q(ow_word[33])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i33.GSR = "DISABLED";
    LUT4 i20555_2_lut_rep_797 (.A(iw_word[33]), .B(iw_stb), .Z(n29457)) /* synthesis lut_function=(A (B)) */ ;
    defparam i20555_2_lut_rep_797.init = 16'h8888;
    LUT4 i1_3_lut_rep_540_4_lut (.A(iw_word[33]), .B(iw_stb), .C(wb_cyc), 
         .D(iw_word[32]), .Z(dac_clk_p_c_enable_60)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_3_lut_rep_540_4_lut.init = 16'h0008;
    CCU2D o_wb_addr_858_add_4_31 (.A0(n19187), .B0(iw_word[1]), .C0(dac_clk_p_c_enable_60), 
          .D0(iw_word[30]), .A1(n19185), .B1(iw_word[1]), .C1(dac_clk_p_c_enable_60), 
          .D1(iw_word[31]), .CIN(n19882), .S0(n125[28]), .S1(n125[29]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_858_add_4_31.INIT0 = 16'h5aaa;
    defparam o_wb_addr_858_add_4_31.INIT1 = 16'h5aaa;
    defparam o_wb_addr_858_add_4_31.INJECT1_0 = "NO";
    defparam o_wb_addr_858_add_4_31.INJECT1_1 = "NO";
    CCU2D o_wb_addr_858_add_4_29 (.A0(n19191), .B0(iw_word[1]), .C0(dac_clk_p_c_enable_60), 
          .D0(iw_word[28]), .A1(n19189), .B1(iw_word[1]), .C1(dac_clk_p_c_enable_60), 
          .D1(iw_word[29]), .CIN(n19881), .COUT(n19882), .S0(n125[26]), 
          .S1(n125[27]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_858_add_4_29.INIT0 = 16'h5aaa;
    defparam o_wb_addr_858_add_4_29.INIT1 = 16'h5aaa;
    defparam o_wb_addr_858_add_4_29.INJECT1_0 = "NO";
    defparam o_wb_addr_858_add_4_29.INJECT1_1 = "NO";
    CCU2D o_wb_addr_858_add_4_27 (.A0(n19195), .B0(iw_word[1]), .C0(dac_clk_p_c_enable_60), 
          .D0(iw_word[26]), .A1(n19193), .B1(iw_word[1]), .C1(dac_clk_p_c_enable_60), 
          .D1(iw_word[27]), .CIN(n19880), .COUT(n19881), .S0(n125[24]), 
          .S1(n125[25]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_858_add_4_27.INIT0 = 16'h5aaa;
    defparam o_wb_addr_858_add_4_27.INIT1 = 16'h5aaa;
    defparam o_wb_addr_858_add_4_27.INJECT1_0 = "NO";
    defparam o_wb_addr_858_add_4_27.INJECT1_1 = "NO";
    CCU2D o_wb_addr_858_add_4_25 (.A0(n19199), .B0(iw_word[1]), .C0(dac_clk_p_c_enable_60), 
          .D0(iw_word[24]), .A1(n19197), .B1(iw_word[1]), .C1(dac_clk_p_c_enable_60), 
          .D1(iw_word[25]), .CIN(n19879), .COUT(n19880), .S0(n125[22]), 
          .S1(n125[23]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_858_add_4_25.INIT0 = 16'h5aaa;
    defparam o_wb_addr_858_add_4_25.INIT1 = 16'h5aaa;
    defparam o_wb_addr_858_add_4_25.INJECT1_0 = "NO";
    defparam o_wb_addr_858_add_4_25.INJECT1_1 = "NO";
    CCU2D o_wb_addr_858_add_4_23 (.A0(n19203), .B0(iw_word[1]), .C0(dac_clk_p_c_enable_60), 
          .D0(iw_word[22]), .A1(n19201), .B1(iw_word[1]), .C1(dac_clk_p_c_enable_60), 
          .D1(iw_word[23]), .CIN(n19878), .COUT(n19879), .S0(n125[20]), 
          .S1(n125[21]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_858_add_4_23.INIT0 = 16'h5aaa;
    defparam o_wb_addr_858_add_4_23.INIT1 = 16'h5aaa;
    defparam o_wb_addr_858_add_4_23.INJECT1_0 = "NO";
    defparam o_wb_addr_858_add_4_23.INJECT1_1 = "NO";
    CCU2D o_wb_addr_858_add_4_21 (.A0(n19207), .B0(iw_word[1]), .C0(dac_clk_p_c_enable_60), 
          .D0(iw_word[20]), .A1(n19205), .B1(iw_word[1]), .C1(dac_clk_p_c_enable_60), 
          .D1(iw_word[21]), .CIN(n19877), .COUT(n19878), .S0(n125[18]), 
          .S1(n125[19]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_858_add_4_21.INIT0 = 16'h5aaa;
    defparam o_wb_addr_858_add_4_21.INIT1 = 16'h5aaa;
    defparam o_wb_addr_858_add_4_21.INJECT1_0 = "NO";
    defparam o_wb_addr_858_add_4_21.INJECT1_1 = "NO";
    CCU2D o_wb_addr_858_add_4_19 (.A0(n19211), .B0(iw_word[1]), .C0(dac_clk_p_c_enable_60), 
          .D0(iw_word[18]), .A1(n19209), .B1(iw_word[1]), .C1(dac_clk_p_c_enable_60), 
          .D1(iw_word[19]), .CIN(n19876), .COUT(n19877), .S0(n125[16]), 
          .S1(n125[17]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_858_add_4_19.INIT0 = 16'h5aaa;
    defparam o_wb_addr_858_add_4_19.INIT1 = 16'h5aaa;
    defparam o_wb_addr_858_add_4_19.INJECT1_0 = "NO";
    defparam o_wb_addr_858_add_4_19.INJECT1_1 = "NO";
    CCU2D o_wb_addr_858_add_4_17 (.A0(n19215), .B0(iw_word[1]), .C0(dac_clk_p_c_enable_60), 
          .D0(iw_word[16]), .A1(n19213), .B1(iw_word[1]), .C1(dac_clk_p_c_enable_60), 
          .D1(iw_word[17]), .CIN(n19875), .COUT(n19876), .S0(n125[14]), 
          .S1(n125[15]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_858_add_4_17.INIT0 = 16'h5aaa;
    defparam o_wb_addr_858_add_4_17.INIT1 = 16'h5aaa;
    defparam o_wb_addr_858_add_4_17.INJECT1_0 = "NO";
    defparam o_wb_addr_858_add_4_17.INJECT1_1 = "NO";
    CCU2D o_wb_addr_858_add_4_15 (.A0(n19219), .B0(iw_word[1]), .C0(dac_clk_p_c_enable_60), 
          .D0(iw_word[14]), .A1(n19217), .B1(iw_word[1]), .C1(dac_clk_p_c_enable_60), 
          .D1(iw_word[15]), .CIN(n19874), .COUT(n19875), .S0(n125[12]), 
          .S1(n125[13]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_858_add_4_15.INIT0 = 16'h5aaa;
    defparam o_wb_addr_858_add_4_15.INIT1 = 16'h5aaa;
    defparam o_wb_addr_858_add_4_15.INJECT1_0 = "NO";
    defparam o_wb_addr_858_add_4_15.INJECT1_1 = "NO";
    CCU2D o_wb_addr_858_add_4_13 (.A0(n19223), .B0(iw_word[1]), .C0(dac_clk_p_c_enable_60), 
          .D0(iw_word[12]), .A1(n19221), .B1(iw_word[1]), .C1(dac_clk_p_c_enable_60), 
          .D1(iw_word[13]), .CIN(n19873), .COUT(n19874), .S0(n125[10]), 
          .S1(n125[11]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_858_add_4_13.INIT0 = 16'h5aaa;
    defparam o_wb_addr_858_add_4_13.INIT1 = 16'h5aaa;
    defparam o_wb_addr_858_add_4_13.INJECT1_0 = "NO";
    defparam o_wb_addr_858_add_4_13.INJECT1_1 = "NO";
    FD1P3IX o_wb_stb_68 (.D(n24010), .SP(o_cmd_busy_N_698), .CD(n21661), 
            .CK(dac_clk_p_c), .Q(wb_stb)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(121[9] 168[5])
    defparam o_wb_stb_68.GSR = "DISABLED";
    FD1S3AX o_wb_data_i31 (.D(iw_word[31]), .CK(dac_clk_p_c), .Q(wb_odata[31])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i31.GSR = "DISABLED";
    CCU2D o_wb_addr_858_add_4_11 (.A0(n19227), .B0(iw_word[1]), .C0(dac_clk_p_c_enable_60), 
          .D0(iw_word[10]), .A1(n19225), .B1(iw_word[1]), .C1(dac_clk_p_c_enable_60), 
          .D1(iw_word[11]), .CIN(n19872), .COUT(n19873), .S0(n125[8]), 
          .S1(n125[9]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_858_add_4_11.INIT0 = 16'h5aaa;
    defparam o_wb_addr_858_add_4_11.INIT1 = 16'h5aaa;
    defparam o_wb_addr_858_add_4_11.INJECT1_0 = "NO";
    defparam o_wb_addr_858_add_4_11.INJECT1_1 = "NO";
    CCU2D o_wb_addr_858_add_4_9 (.A0(n19231), .B0(iw_word[1]), .C0(dac_clk_p_c_enable_60), 
          .D0(iw_word[8]), .A1(n19229), .B1(iw_word[1]), .C1(dac_clk_p_c_enable_60), 
          .D1(iw_word[9]), .CIN(n19871), .COUT(n19872), .S0(n125[6]), 
          .S1(n125[7]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_858_add_4_9.INIT0 = 16'h5aaa;
    defparam o_wb_addr_858_add_4_9.INIT1 = 16'h5aaa;
    defparam o_wb_addr_858_add_4_9.INJECT1_0 = "NO";
    defparam o_wb_addr_858_add_4_9.INJECT1_1 = "NO";
    CCU2D o_wb_addr_858_add_4_7 (.A0(n19235), .B0(iw_word[1]), .C0(dac_clk_p_c_enable_60), 
          .D0(iw_word[6]), .A1(n19233), .B1(iw_word[1]), .C1(dac_clk_p_c_enable_60), 
          .D1(iw_word[7]), .CIN(n19870), .COUT(n19871), .S0(n125[4]), 
          .S1(n125[5]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_858_add_4_7.INIT0 = 16'h5aaa;
    defparam o_wb_addr_858_add_4_7.INIT1 = 16'h5aaa;
    defparam o_wb_addr_858_add_4_7.INJECT1_0 = "NO";
    defparam o_wb_addr_858_add_4_7.INJECT1_1 = "NO";
    CCU2D o_wb_addr_858_add_4_5 (.A0(n19239), .B0(iw_word[1]), .C0(dac_clk_p_c_enable_60), 
          .D0(iw_word[4]), .A1(n19237), .B1(iw_word[1]), .C1(dac_clk_p_c_enable_60), 
          .D1(iw_word[5]), .CIN(n19869), .COUT(n19870), .S0(n125[2]), 
          .S1(n125[3]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_858_add_4_5.INIT0 = 16'h5aaa;
    defparam o_wb_addr_858_add_4_5.INIT1 = 16'h5aaa;
    defparam o_wb_addr_858_add_4_5.INJECT1_0 = "NO";
    defparam o_wb_addr_858_add_4_5.INJECT1_1 = "NO";
    CCU2D o_wb_addr_858_add_4_3 (.A0(n19242), .B0(dac_clk_p_c_enable_60), 
          .C0(iw_word[1]), .D0(wb_addr[0]), .A1(n19241), .B1(iw_word[1]), 
          .C1(dac_clk_p_c_enable_60), .D1(iw_word[3]), .CIN(n19868), .COUT(n19869), 
          .S0(n125[0]), .S1(n125[1]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_858_add_4_3.INIT0 = 16'h59aa;
    defparam o_wb_addr_858_add_4_3.INIT1 = 16'h5aaa;
    defparam o_wb_addr_858_add_4_3.INJECT1_0 = "NO";
    defparam o_wb_addr_858_add_4_3.INJECT1_1 = "NO";
    CCU2D o_wb_addr_858_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(iw_word[1]), .B1(dac_clk_p_c_enable_60), .C1(GND_net), 
          .D1(GND_net), .COUT(n19868));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_858_add_4_1.INIT0 = 16'hF000;
    defparam o_wb_addr_858_add_4_1.INIT1 = 16'hffff;
    defparam o_wb_addr_858_add_4_1.INJECT1_0 = "NO";
    defparam o_wb_addr_858_add_4_1.INJECT1_1 = "NO";
    LUT4 i_cmd_word_0__I_0_1_lut (.A(iw_word[0]), .Z(i_cmd_word_0__N_762)) /* synthesis lut_function=(!(A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(214[11:25])
    defparam i_cmd_word_0__I_0_1_lut.init = 16'h5555;
    LUT4 o_cmd_busy_I_0_1_lut (.A(wb_cyc), .Z(o_cmd_busy_N_698)) /* synthesis lut_function=(!(A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(194[21:34])
    defparam o_cmd_busy_I_0_1_lut.init = 16'h5555;
    FD1S3AX o_wb_data_i30 (.D(iw_word[30]), .CK(dac_clk_p_c), .Q(wb_odata[30])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i30.GSR = "DISABLED";
    FD1S3AX o_wb_data_i29 (.D(iw_word[29]), .CK(dac_clk_p_c), .Q(wb_odata[29])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i29.GSR = "DISABLED";
    FD1S3AX o_wb_data_i28 (.D(iw_word[28]), .CK(dac_clk_p_c), .Q(wb_odata[28])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i28.GSR = "DISABLED";
    FD1S3AX o_wb_data_i27 (.D(iw_word[27]), .CK(dac_clk_p_c), .Q(wb_odata[27])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i27.GSR = "DISABLED";
    FD1S3AX o_wb_data_i26 (.D(iw_word[26]), .CK(dac_clk_p_c), .Q(wb_odata[26])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i26.GSR = "DISABLED";
    FD1S3AX o_wb_data_i25 (.D(iw_word[25]), .CK(dac_clk_p_c), .Q(wb_odata[25])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i25.GSR = "DISABLED";
    FD1S3AX o_wb_data_i24 (.D(iw_word[24]), .CK(dac_clk_p_c), .Q(wb_odata[24])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i24.GSR = "DISABLED";
    FD1S3AX o_wb_data_i23 (.D(iw_word[23]), .CK(dac_clk_p_c), .Q(wb_odata[23])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i23.GSR = "DISABLED";
    FD1S3AX o_wb_data_i22 (.D(iw_word[22]), .CK(dac_clk_p_c), .Q(wb_odata[22])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i22.GSR = "DISABLED";
    FD1S3AX o_wb_data_i21 (.D(iw_word[21]), .CK(dac_clk_p_c), .Q(wb_odata[21])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i21.GSR = "DISABLED";
    FD1S3AX o_wb_data_i20 (.D(iw_word[20]), .CK(dac_clk_p_c), .Q(wb_odata[20])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i20.GSR = "DISABLED";
    FD1S3AX o_wb_data_i19 (.D(iw_word[19]), .CK(dac_clk_p_c), .Q(wb_odata[19])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i19.GSR = "DISABLED";
    FD1S3AX o_wb_data_i18 (.D(iw_word[18]), .CK(dac_clk_p_c), .Q(wb_odata[18])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i18.GSR = "DISABLED";
    FD1S3AX o_wb_data_i17 (.D(iw_word[17]), .CK(dac_clk_p_c), .Q(wb_odata[17])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i17.GSR = "DISABLED";
    FD1S3AX o_wb_data_i16 (.D(iw_word[16]), .CK(dac_clk_p_c), .Q(wb_odata[16])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i16.GSR = "DISABLED";
    FD1S3AX o_wb_data_i15 (.D(iw_word[15]), .CK(dac_clk_p_c), .Q(wb_odata[15])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i15.GSR = "DISABLED";
    FD1S3AX o_wb_data_i14 (.D(iw_word[14]), .CK(dac_clk_p_c), .Q(wb_odata[14])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i14.GSR = "DISABLED";
    FD1S3AX o_wb_data_i13 (.D(iw_word[13]), .CK(dac_clk_p_c), .Q(wb_odata[13])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i13.GSR = "DISABLED";
    FD1S3AX o_wb_data_i12 (.D(iw_word[12]), .CK(dac_clk_p_c), .Q(wb_odata[12])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i12.GSR = "DISABLED";
    FD1S3AX o_wb_data_i11 (.D(iw_word[11]), .CK(dac_clk_p_c), .Q(wb_odata[11])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i11.GSR = "DISABLED";
    FD1S3AX o_wb_data_i10 (.D(iw_word[10]), .CK(dac_clk_p_c), .Q(wb_odata[10])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i10.GSR = "DISABLED";
    FD1S3AX o_wb_data_i9 (.D(iw_word[9]), .CK(dac_clk_p_c), .Q(wb_odata[9])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i9.GSR = "DISABLED";
    FD1S3AX o_wb_data_i8 (.D(iw_word[8]), .CK(dac_clk_p_c), .Q(wb_odata[8])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i8.GSR = "DISABLED";
    FD1S3AX o_wb_data_i7 (.D(iw_word[7]), .CK(dac_clk_p_c), .Q(wb_odata[7])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i7.GSR = "DISABLED";
    FD1S3AX o_wb_data_i6 (.D(iw_word[6]), .CK(dac_clk_p_c), .Q(wb_odata[6])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i6.GSR = "DISABLED";
    FD1S3AX o_wb_data_i5 (.D(iw_word[5]), .CK(dac_clk_p_c), .Q(wb_odata[5])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i5.GSR = "DISABLED";
    FD1S3AX o_wb_data_i4 (.D(iw_word[4]), .CK(dac_clk_p_c), .Q(wb_odata[4])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i4.GSR = "DISABLED";
    FD1S3AX o_wb_data_i3 (.D(iw_word[3]), .CK(dac_clk_p_c), .Q(wb_odata[3])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i3.GSR = "DISABLED";
    FD1S3AX o_wb_data_i2 (.D(iw_word[2]), .CK(dac_clk_p_c), .Q(wb_odata[2])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i2.GSR = "DISABLED";
    FD1S3AX o_wb_data_i1 (.D(iw_word[1]), .CK(dac_clk_p_c), .Q(wb_odata[1])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i1.GSR = "DISABLED";
    LUT4 newaddr_I_0_3_lut (.A(newaddr), .B(wb_ack), .C(wb_cyc), .Z(o_rsp_stb_N_754)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam newaddr_I_0_3_lut.init = 16'hcaca;
    LUT4 mux_59_i1_4_lut (.A(inc), .B(\wb_idata[0] ), .C(wb_cyc), .D(wb_we), 
         .Z(n338[0])) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A (B (C (D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i1_4_lut.init = 16'h05c5;
    LUT4 mux_59_i3_4_lut (.A(wb_addr[0]), .B(\wb_idata[2] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[2])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i3_4_lut.init = 16'h0aca;
    LUT4 mux_59_i4_4_lut (.A(wb_addr[1]), .B(\wb_idata[3] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[3])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i4_4_lut.init = 16'h0aca;
    LUT4 mux_59_i5_4_lut (.A(wb_addr[2]), .B(\wb_idata[4] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[4])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i5_4_lut.init = 16'h0aca;
    LUT4 mux_59_i6_4_lut (.A(wb_addr[3]), .B(\wb_idata[5] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[5])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i6_4_lut.init = 16'h0aca;
    LUT4 mux_59_i7_4_lut (.A(wb_addr[4]), .B(\wb_idata[6] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[6])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i7_4_lut.init = 16'h0aca;
    LUT4 mux_59_i8_4_lut (.A(wb_addr[5]), .B(\wb_idata[7] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[7])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i8_4_lut.init = 16'h0aca;
    LUT4 mux_59_i9_4_lut (.A(wb_addr[6]), .B(\wb_idata[8] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[8])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i9_4_lut.init = 16'h0aca;
    LUT4 mux_59_i10_4_lut (.A(wb_addr[7]), .B(\wb_idata[9] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[9])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i10_4_lut.init = 16'h0aca;
    LUT4 mux_59_i11_4_lut (.A(wb_addr[8]), .B(\wb_idata[10] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[10])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i11_4_lut.init = 16'h0aca;
    LUT4 mux_59_i12_4_lut (.A(wb_addr[9]), .B(\wb_idata[11] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[11])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i12_4_lut.init = 16'h0aca;
    LUT4 mux_59_i13_4_lut (.A(wb_addr[10]), .B(\wb_idata[12] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[12])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i13_4_lut.init = 16'h0aca;
    LUT4 mux_59_i14_4_lut (.A(wb_addr[11]), .B(\wb_idata[13] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[13])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i14_4_lut.init = 16'h0aca;
    LUT4 mux_59_i15_4_lut (.A(wb_addr[12]), .B(\wb_idata[14] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[14])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i15_4_lut.init = 16'h0aca;
    LUT4 mux_59_i16_4_lut (.A(wb_addr[13]), .B(\wb_idata[15] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[15])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i16_4_lut.init = 16'h0aca;
    LUT4 mux_59_i17_4_lut (.A(wb_addr[14]), .B(\wb_idata[16] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[16])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i17_4_lut.init = 16'h0aca;
    LUT4 mux_59_i18_4_lut (.A(wb_addr[15]), .B(\wb_idata[17] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[17])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i18_4_lut.init = 16'h0aca;
    LUT4 mux_59_i19_4_lut (.A(wb_addr[16]), .B(\wb_idata[18] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[18])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i19_4_lut.init = 16'h0aca;
    LUT4 mux_59_i20_4_lut (.A(wb_addr[17]), .B(\wb_idata[19] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[19])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i20_4_lut.init = 16'h0aca;
    LUT4 mux_59_i21_4_lut (.A(wb_addr[18]), .B(\wb_idata[20] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[20])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i21_4_lut.init = 16'h0aca;
    LUT4 mux_59_i22_4_lut (.A(wb_addr[19]), .B(\wb_idata[21] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[21])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i22_4_lut.init = 16'h0aca;
    LUT4 mux_59_i23_4_lut (.A(wb_addr[20]), .B(\wb_idata[22] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[22])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i23_4_lut.init = 16'h0aca;
    LUT4 mux_59_i24_4_lut (.A(wb_addr[21]), .B(\wb_idata[23] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[23])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i24_4_lut.init = 16'h0aca;
    LUT4 mux_59_i25_4_lut (.A(wb_addr[22]), .B(\wb_idata[24] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[24])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i25_4_lut.init = 16'h0aca;
    LUT4 mux_59_i26_4_lut (.A(wb_addr[23]), .B(\wb_idata[25] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[25])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i26_4_lut.init = 16'h0aca;
    LUT4 mux_59_i27_4_lut (.A(wb_addr[24]), .B(\wb_idata[26] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[26])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i27_4_lut.init = 16'h0aca;
    LUT4 mux_59_i28_4_lut (.A(wb_addr[25]), .B(\wb_idata[27] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[27])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i28_4_lut.init = 16'h0aca;
    LUT4 mux_59_i29_4_lut (.A(wb_addr[26]), .B(\wb_idata[28] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[28])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i29_4_lut.init = 16'h0aca;
    LUT4 i12571_4_lut (.A(wb_addr[27]), .B(wb_err), .C(n1639[29]), .D(wb_cyc), 
         .Z(o_rsp_word_33__N_718[29])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(287[11] 309[5])
    defparam i12571_4_lut.init = 16'hfcee;
    LUT4 i12597_2_lut (.A(\wb_idata[29] ), .B(wb_we), .Z(n1639[29])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(299[4:47])
    defparam i12597_2_lut.init = 16'h2222;
    LUT4 mux_59_i31_4_lut (.A(wb_addr[28]), .B(\wb_idata[30] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[30])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i31_4_lut.init = 16'h0aca;
    LUT4 mux_59_i32_4_lut (.A(wb_addr[29]), .B(\wb_idata[31] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[31])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i32_4_lut.init = 16'h0aca;
    LUT4 i12572_2_lut (.A(wb_we), .B(wb_cyc), .Z(n338[32])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam i12572_2_lut.init = 16'h8888;
    LUT4 i2_1_lut (.A(wb_stb), .Z(n2)) /* synthesis lut_function=(!(A)) */ ;
    defparam i2_1_lut.init = 16'h5555;
    LUT4 i17724_2_lut (.A(wb_addr[28]), .B(n3), .Z(n19187)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i17724_2_lut.init = 16'h8888;
    LUT4 i17725_2_lut (.A(wb_addr[29]), .B(n3), .Z(n19185)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i17725_2_lut.init = 16'h8888;
    LUT4 i1_4_lut (.A(n29457), .B(iw_word[1]), .C(wb_cyc), .D(iw_word[32]), 
         .Z(n3)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(110[35:71])
    defparam i1_4_lut.init = 16'hfffd;
    LUT4 i17722_2_lut (.A(wb_addr[26]), .B(n3), .Z(n19191)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i17722_2_lut.init = 16'h8888;
    LUT4 i17723_2_lut (.A(wb_addr[27]), .B(n3), .Z(n19189)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i17723_2_lut.init = 16'h8888;
    LUT4 i17719_2_lut (.A(wb_addr[24]), .B(n3), .Z(n19195)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i17719_2_lut.init = 16'h8888;
    LUT4 i17720_2_lut (.A(wb_addr[25]), .B(n3), .Z(n19193)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i17720_2_lut.init = 16'h8888;
    LUT4 i17704_2_lut (.A(wb_addr[22]), .B(n3), .Z(n19199)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i17704_2_lut.init = 16'h8888;
    LUT4 i17718_2_lut (.A(wb_addr[23]), .B(n3), .Z(n19197)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i17718_2_lut.init = 16'h8888;
    LUT4 i17665_2_lut (.A(wb_addr[20]), .B(n3), .Z(n19203)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i17665_2_lut.init = 16'h8888;
    LUT4 i17708_2_lut (.A(wb_addr[21]), .B(n3), .Z(n19201)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i17708_2_lut.init = 16'h8888;
    LUT4 i17709_2_lut (.A(wb_addr[18]), .B(n3), .Z(n19207)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i17709_2_lut.init = 16'h8888;
    LUT4 i17664_2_lut (.A(wb_addr[19]), .B(n3), .Z(n19205)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i17664_2_lut.init = 16'h8888;
    LUT4 i17672_2_lut (.A(wb_addr[16]), .B(n3), .Z(n19211)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i17672_2_lut.init = 16'h8888;
    LUT4 i17706_2_lut (.A(wb_addr[17]), .B(n3), .Z(n19209)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i17706_2_lut.init = 16'h8888;
    LUT4 i17710_2_lut (.A(wb_addr[14]), .B(n3), .Z(n19215)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i17710_2_lut.init = 16'h8888;
    LUT4 i17670_2_lut (.A(wb_addr[15]), .B(n3), .Z(n19213)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i17670_2_lut.init = 16'h8888;
    LUT4 i17676_2_lut (.A(wb_addr[12]), .B(n3), .Z(n19219)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i17676_2_lut.init = 16'h8888;
    LUT4 i17705_2_lut (.A(wb_addr[13]), .B(n3), .Z(n19217)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i17705_2_lut.init = 16'h8888;
    LUT4 i17666_2_lut (.A(wb_addr[10]), .B(n3), .Z(n19223)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i17666_2_lut.init = 16'h8888;
    LUT4 i17671_2_lut (.A(wb_addr[11]), .B(n3), .Z(n19221)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i17671_2_lut.init = 16'h8888;
    LUT4 i12447_2_lut_4_lut (.A(iw_word[32]), .B(wb_cyc), .C(n29457), 
         .D(wb_stb), .Z(dac_clk_p_c_enable_631)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C+(D)))) */ ;
    defparam i12447_2_lut_4_lut.init = 16'hff10;
    LUT4 i17707_2_lut (.A(wb_addr[8]), .B(n3), .Z(n19227)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i17707_2_lut.init = 16'h8888;
    LUT4 i17711_2_lut (.A(wb_addr[9]), .B(n3), .Z(n19225)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i17711_2_lut.init = 16'h8888;
    LUT4 i17696_2_lut (.A(wb_addr[6]), .B(n3), .Z(n19231)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i17696_2_lut.init = 16'h8888;
    LUT4 i17697_2_lut (.A(wb_addr[7]), .B(n3), .Z(n19229)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i17697_2_lut.init = 16'h8888;
    LUT4 i17685_2_lut (.A(wb_addr[4]), .B(n3), .Z(n19235)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i17685_2_lut.init = 16'h8888;
    LUT4 i17686_2_lut (.A(wb_addr[5]), .B(n3), .Z(n19233)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i17686_2_lut.init = 16'h8888;
    LUT4 i17677_2_lut (.A(wb_addr[2]), .B(n3), .Z(n19239)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i17677_2_lut.init = 16'h8888;
    LUT4 i17684_2_lut (.A(wb_addr[3]), .B(n3), .Z(n19237)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i17684_2_lut.init = 16'h8888;
    LUT4 i17674_3_lut (.A(inc), .B(iw_word[2]), .C(dac_clk_p_c_enable_60), 
         .Z(n19242)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i17674_3_lut.init = 16'hcaca;
    LUT4 i17675_2_lut (.A(wb_addr[1]), .B(n3), .Z(n19241)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i17675_2_lut.init = 16'h8888;
    LUT4 i3_4_lut (.A(n32125), .B(iw_word[32]), .C(iw_stb), .D(iw_word[33]), 
         .Z(newaddr_N_757)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i3_4_lut.init = 16'h1000;
    FD1P3AX o_wb_addr_858__i29 (.D(n125[29]), .SP(dac_clk_p_c_enable_631), 
            .CK(dac_clk_p_c), .Q(wb_addr[29])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_858__i29.GSR = "DISABLED";
    FD1P3AX o_wb_addr_858__i28 (.D(n125[28]), .SP(dac_clk_p_c_enable_631), 
            .CK(dac_clk_p_c), .Q(wb_addr[28])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_858__i28.GSR = "DISABLED";
    FD1P3AX o_wb_addr_858__i27 (.D(n125[27]), .SP(dac_clk_p_c_enable_631), 
            .CK(dac_clk_p_c), .Q(wb_addr[27])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_858__i27.GSR = "DISABLED";
    FD1P3AX o_wb_addr_858__i26 (.D(n125[26]), .SP(dac_clk_p_c_enable_631), 
            .CK(dac_clk_p_c), .Q(wb_addr[26])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_858__i26.GSR = "DISABLED";
    FD1P3AX o_wb_addr_858__i25 (.D(n125[25]), .SP(dac_clk_p_c_enable_631), 
            .CK(dac_clk_p_c), .Q(wb_addr[25])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_858__i25.GSR = "DISABLED";
    FD1P3AX o_wb_addr_858__i24 (.D(n125[24]), .SP(dac_clk_p_c_enable_631), 
            .CK(dac_clk_p_c), .Q(wb_addr[24])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_858__i24.GSR = "DISABLED";
    FD1P3AX o_wb_addr_858__i23 (.D(n125[23]), .SP(dac_clk_p_c_enable_631), 
            .CK(dac_clk_p_c), .Q(wb_addr[23])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_858__i23.GSR = "DISABLED";
    FD1P3AX o_wb_addr_858__i22 (.D(n125[22]), .SP(dac_clk_p_c_enable_631), 
            .CK(dac_clk_p_c), .Q(wb_addr[22])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_858__i22.GSR = "DISABLED";
    FD1P3AX o_wb_addr_858__i21 (.D(n125[21]), .SP(dac_clk_p_c_enable_631), 
            .CK(dac_clk_p_c), .Q(wb_addr[21])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_858__i21.GSR = "DISABLED";
    FD1P3AX o_wb_addr_858__i20 (.D(n125[20]), .SP(dac_clk_p_c_enable_631), 
            .CK(dac_clk_p_c), .Q(wb_addr[20])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_858__i20.GSR = "DISABLED";
    FD1P3AX o_wb_addr_858__i19 (.D(n125[19]), .SP(dac_clk_p_c_enable_631), 
            .CK(dac_clk_p_c), .Q(wb_addr[19])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_858__i19.GSR = "DISABLED";
    FD1P3AX o_wb_addr_858__i18 (.D(n125[18]), .SP(dac_clk_p_c_enable_631), 
            .CK(dac_clk_p_c), .Q(wb_addr[18])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_858__i18.GSR = "DISABLED";
    FD1P3AX o_wb_addr_858__i17 (.D(n125[17]), .SP(dac_clk_p_c_enable_631), 
            .CK(dac_clk_p_c), .Q(wb_addr[17])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_858__i17.GSR = "DISABLED";
    FD1P3AX o_wb_addr_858__i16 (.D(n125[16]), .SP(dac_clk_p_c_enable_631), 
            .CK(dac_clk_p_c), .Q(wb_addr[16])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_858__i16.GSR = "DISABLED";
    FD1P3AX o_wb_addr_858__i15 (.D(n125[15]), .SP(dac_clk_p_c_enable_631), 
            .CK(dac_clk_p_c), .Q(wb_addr[15])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_858__i15.GSR = "DISABLED";
    FD1P3AX o_wb_addr_858__i14 (.D(n125[14]), .SP(dac_clk_p_c_enable_631), 
            .CK(dac_clk_p_c), .Q(wb_addr[14])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_858__i14.GSR = "DISABLED";
    FD1P3AX o_wb_addr_858__i13 (.D(n125[13]), .SP(dac_clk_p_c_enable_631), 
            .CK(dac_clk_p_c), .Q(wb_addr[13])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_858__i13.GSR = "DISABLED";
    FD1P3AX o_wb_addr_858__i12 (.D(n125[12]), .SP(dac_clk_p_c_enable_631), 
            .CK(dac_clk_p_c), .Q(wb_addr[12])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_858__i12.GSR = "DISABLED";
    FD1P3AX o_wb_addr_858__i11 (.D(n125[11]), .SP(dac_clk_p_c_enable_631), 
            .CK(dac_clk_p_c), .Q(wb_addr[11])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_858__i11.GSR = "DISABLED";
    FD1P3AX o_wb_addr_858__i10 (.D(n125[10]), .SP(dac_clk_p_c_enable_631), 
            .CK(dac_clk_p_c), .Q(wb_addr[10])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_858__i10.GSR = "DISABLED";
    FD1P3AX o_wb_addr_858__i9 (.D(n125[9]), .SP(dac_clk_p_c_enable_631), 
            .CK(dac_clk_p_c), .Q(wb_addr[9])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_858__i9.GSR = "DISABLED";
    FD1P3AX o_wb_addr_858__i8 (.D(n125[8]), .SP(dac_clk_p_c_enable_631), 
            .CK(dac_clk_p_c), .Q(wb_addr[8])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_858__i8.GSR = "DISABLED";
    FD1P3AX o_wb_addr_858__i7 (.D(n125[7]), .SP(dac_clk_p_c_enable_631), 
            .CK(dac_clk_p_c), .Q(wb_addr[7])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_858__i7.GSR = "DISABLED";
    FD1P3AX o_wb_addr_858__i6 (.D(n125[6]), .SP(dac_clk_p_c_enable_631), 
            .CK(dac_clk_p_c), .Q(wb_addr[6])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_858__i6.GSR = "DISABLED";
    FD1P3AX o_wb_addr_858__i5 (.D(n125[5]), .SP(dac_clk_p_c_enable_631), 
            .CK(dac_clk_p_c), .Q(wb_addr[5])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_858__i5.GSR = "DISABLED";
    FD1P3AX o_wb_addr_858__i4 (.D(n125[4]), .SP(dac_clk_p_c_enable_631), 
            .CK(dac_clk_p_c), .Q(wb_addr[4])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_858__i4.GSR = "DISABLED";
    FD1P3AX o_wb_addr_858__i3 (.D(n125[3]), .SP(dac_clk_p_c_enable_631), 
            .CK(dac_clk_p_c), .Q(wb_addr[3])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_858__i3.GSR = "DISABLED";
    FD1P3AX o_wb_addr_858__i2 (.D(n125[2]), .SP(dac_clk_p_c_enable_631), 
            .CK(dac_clk_p_c), .Q(wb_addr[2])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_858__i2.GSR = "DISABLED";
    FD1P3AX o_wb_addr_858__i1 (.D(n125[1]), .SP(dac_clk_p_c_enable_631), 
            .CK(dac_clk_p_c), .Q(wb_addr[1])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_858__i1.GSR = "DISABLED";
    LUT4 i1_2_lut_3_lut_4_lut (.A(wb_err), .B(wb_cyc), .C(wb_stb), .D(n32125), 
         .Z(n21661)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(122[17:41])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfff8;
    LUT4 i1_2_lut_rep_469_3_lut (.A(wb_err), .B(wb_cyc), .C(n32125), .Z(o_cmd_busy_N_708)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(122[17:41])
    defparam i1_2_lut_rep_469_3_lut.init = 16'hf8f8;
    LUT4 i1_2_lut_rep_796 (.A(iw_stb), .B(iw_word[33]), .Z(n29456)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i1_2_lut_rep_796.init = 16'h2222;
    LUT4 i1_2_lut_3_lut (.A(iw_stb), .B(iw_word[33]), .C(iw_word[32]), 
         .Z(i_cmd_wr)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_3_lut.init = 16'h2020;
    LUT4 i21528_3_lut_3_lut (.A(iw_stb), .B(iw_word[33]), .C(wb_stb), 
         .Z(n24010)) /* synthesis lut_function=(A ((C)+!B)+!A (C)) */ ;
    defparam i21528_3_lut_3_lut.init = 16'hf2f2;
    LUT4 i1_4_lut_adj_212 (.A(n29456), .B(o_cmd_busy_N_708), .C(wb_ack), 
         .D(o_cmd_busy_N_700), .Z(dac_clk_p_c_enable_640)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+!((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(122[6:41])
    defparam i1_4_lut_adj_212.init = 16'heefc;
    LUT4 i24666_2_lut (.A(wb_cyc), .B(wb_stb), .Z(o_cmd_busy_N_700)) /* synthesis lut_function=(!(A+(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(149[11] 168[5])
    defparam i24666_2_lut.init = 16'h1111;
    FD1S3IX o_rsp_word_i1 (.D(n22149), .CK(dac_clk_p_c), .CD(n14148), 
            .Q(ow_word[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i1.GSR = "DISABLED";
    LUT4 i7657_2_lut_rep_738 (.A(wb_err), .B(n32125), .Z(n29398)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(283[11] 309[5])
    defparam i7657_2_lut_rep_738.init = 16'heeee;
    LUT4 i24578_3_lut_4_lut (.A(wb_err), .B(n32125), .C(wb_we), .D(wb_cyc), 
         .Z(n22149)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(283[11] 309[5])
    defparam i24578_3_lut_4_lut.init = 16'h0100;
    FD1P3AX o_wb_addr_858__i0 (.D(n125[0]), .SP(dac_clk_p_c_enable_631), 
            .CK(dac_clk_p_c), .Q(wb_addr[0])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_858__i0.GSR = "DISABLED";
    FD1P3IX o_wb_cyc_67 (.D(o_cmd_busy_N_700), .SP(dac_clk_p_c_enable_640), 
            .CD(o_cmd_busy_N_708), .CK(dac_clk_p_c), .Q(wb_cyc)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(121[9] 168[5])
    defparam o_wb_cyc_67.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module hbdeword
//

module hbdeword (hb_bits, dac_clk_p_c, dac_clk_p_c_enable_312, n32067, 
            n32126, hb_busy, w_reset, idl_word, n32125, nl_busy, 
            hx_stb, idl_stb) /* synthesis syn_module_defined=1 */ ;
    output [4:0]hb_bits;
    input dac_clk_p_c;
    input dac_clk_p_c_enable_312;
    input n32067;
    input n32126;
    output hb_busy;
    input w_reset;
    input [33:0]idl_word;
    input n32125;
    input nl_busy;
    input hx_stb;
    input idl_stb;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[29:38])
    
    wire dac_clk_p_c_enable_647;
    wire [4:0]o_dw_bits_4__N_955;
    wire [3:0]r_len;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(58[12:17])
    
    wire n29196;
    wire [3:0]n13;
    
    wire n14220, dac_clk_p_c_enable_168;
    wire [3:0]r_len_3__N_996;
    
    wire o_dw_busy_N_1036;
    wire [31:0]r_word;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(59[13:19])
    wire [31:0]r_word_31__N_964;
    
    wire n12776, n26463, n12780, n29366, n29364, n22051, n28875, 
        n29452;
    
    FD1P3AX o_dw_bits_i2 (.D(o_dw_bits_4__N_955[2]), .SP(dac_clk_p_c_enable_647), 
            .CK(dac_clk_p_c), .Q(hb_bits[2])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(95[9] 103[41])
    defparam o_dw_bits_i2.GSR = "DISABLED";
    FD1P3AX o_dw_bits_i1 (.D(o_dw_bits_4__N_955[1]), .SP(dac_clk_p_c_enable_647), 
            .CK(dac_clk_p_c), .Q(hb_bits[1])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(95[9] 103[41])
    defparam o_dw_bits_i1.GSR = "DISABLED";
    FD1P3IX r_len__i0 (.D(n13[0]), .SP(dac_clk_p_c_enable_312), .CD(n29196), 
            .CK(dac_clk_p_c), .Q(r_len[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(64[9] 81[6])
    defparam r_len__i0.GSR = "DISABLED";
    FD1P3IX o_dw_bits_i4 (.D(n32067), .SP(dac_clk_p_c_enable_647), .CD(n14220), 
            .CK(dac_clk_p_c), .Q(hb_bits[4])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(95[9] 103[41])
    defparam o_dw_bits_i4.GSR = "DISABLED";
    FD1P3AX o_dw_bits_i0 (.D(o_dw_bits_4__N_955[0]), .SP(dac_clk_p_c_enable_647), 
            .CK(dac_clk_p_c), .Q(hb_bits[0])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(95[9] 103[41])
    defparam o_dw_bits_i0.GSR = "DISABLED";
    FD1P3IX r_len__i3 (.D(r_len_3__N_996[3]), .SP(dac_clk_p_c_enable_168), 
            .CD(n32126), .CK(dac_clk_p_c), .Q(r_len[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(64[9] 81[6])
    defparam r_len__i3.GSR = "DISABLED";
    FD1P3IX o_dw_stb_36 (.D(o_dw_busy_N_1036), .SP(dac_clk_p_c_enable_168), 
            .CD(w_reset), .CK(dac_clk_p_c), .Q(hb_busy)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(64[9] 81[6])
    defparam o_dw_stb_36.GSR = "DISABLED";
    FD1P3IX r_word_i1 (.D(idl_word[1]), .SP(dac_clk_p_c_enable_647), .CD(n14220), 
            .CK(dac_clk_p_c), .Q(r_word[1])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i1.GSR = "DISABLED";
    FD1P3IX r_word_i2 (.D(idl_word[2]), .SP(dac_clk_p_c_enable_647), .CD(n14220), 
            .CK(dac_clk_p_c), .Q(r_word[2])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i2.GSR = "DISABLED";
    FD1P3IX r_word_i3 (.D(idl_word[3]), .SP(dac_clk_p_c_enable_647), .CD(n14220), 
            .CK(dac_clk_p_c), .Q(r_word[3])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i3.GSR = "DISABLED";
    FD1P3AX r_word_i31 (.D(r_word_31__N_964[31]), .SP(dac_clk_p_c_enable_647), 
            .CK(dac_clk_p_c), .Q(r_word[31])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i31.GSR = "DISABLED";
    FD1P3IX r_word_i0 (.D(idl_word[0]), .SP(dac_clk_p_c_enable_647), .CD(n14220), 
            .CK(dac_clk_p_c), .Q(r_word[0])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i0.GSR = "DISABLED";
    FD1P3AX r_word_i30 (.D(r_word_31__N_964[30]), .SP(dac_clk_p_c_enable_647), 
            .CK(dac_clk_p_c), .Q(r_word[30])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i30.GSR = "DISABLED";
    FD1P3AX r_word_i29 (.D(r_word_31__N_964[29]), .SP(dac_clk_p_c_enable_647), 
            .CK(dac_clk_p_c), .Q(r_word[29])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i29.GSR = "DISABLED";
    FD1P3AX r_word_i28 (.D(r_word_31__N_964[28]), .SP(dac_clk_p_c_enable_647), 
            .CK(dac_clk_p_c), .Q(r_word[28])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i28.GSR = "DISABLED";
    FD1P3AX r_word_i27 (.D(r_word_31__N_964[27]), .SP(dac_clk_p_c_enable_647), 
            .CK(dac_clk_p_c), .Q(r_word[27])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i27.GSR = "DISABLED";
    FD1P3AX r_word_i26 (.D(r_word_31__N_964[26]), .SP(dac_clk_p_c_enable_647), 
            .CK(dac_clk_p_c), .Q(r_word[26])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i26.GSR = "DISABLED";
    FD1P3AX r_word_i25 (.D(r_word_31__N_964[25]), .SP(dac_clk_p_c_enable_647), 
            .CK(dac_clk_p_c), .Q(r_word[25])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i25.GSR = "DISABLED";
    FD1P3AX r_word_i24 (.D(r_word_31__N_964[24]), .SP(dac_clk_p_c_enable_647), 
            .CK(dac_clk_p_c), .Q(r_word[24])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i24.GSR = "DISABLED";
    FD1P3AX r_word_i23 (.D(r_word_31__N_964[23]), .SP(dac_clk_p_c_enable_647), 
            .CK(dac_clk_p_c), .Q(r_word[23])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i23.GSR = "DISABLED";
    FD1P3AX r_word_i22 (.D(r_word_31__N_964[22]), .SP(dac_clk_p_c_enable_647), 
            .CK(dac_clk_p_c), .Q(r_word[22])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i22.GSR = "DISABLED";
    FD1P3AX r_word_i21 (.D(r_word_31__N_964[21]), .SP(dac_clk_p_c_enable_647), 
            .CK(dac_clk_p_c), .Q(r_word[21])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i21.GSR = "DISABLED";
    FD1P3AX r_word_i20 (.D(r_word_31__N_964[20]), .SP(dac_clk_p_c_enable_647), 
            .CK(dac_clk_p_c), .Q(r_word[20])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i20.GSR = "DISABLED";
    FD1P3AX r_word_i19 (.D(r_word_31__N_964[19]), .SP(dac_clk_p_c_enable_647), 
            .CK(dac_clk_p_c), .Q(r_word[19])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i19.GSR = "DISABLED";
    FD1P3AX r_word_i18 (.D(r_word_31__N_964[18]), .SP(dac_clk_p_c_enable_647), 
            .CK(dac_clk_p_c), .Q(r_word[18])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i18.GSR = "DISABLED";
    FD1P3AX r_word_i17 (.D(r_word_31__N_964[17]), .SP(dac_clk_p_c_enable_647), 
            .CK(dac_clk_p_c), .Q(r_word[17])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i17.GSR = "DISABLED";
    FD1P3AX r_word_i16 (.D(r_word_31__N_964[16]), .SP(dac_clk_p_c_enable_647), 
            .CK(dac_clk_p_c), .Q(r_word[16])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i16.GSR = "DISABLED";
    FD1P3AX r_word_i15 (.D(r_word_31__N_964[15]), .SP(dac_clk_p_c_enable_647), 
            .CK(dac_clk_p_c), .Q(r_word[15])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i15.GSR = "DISABLED";
    FD1P3AX r_word_i14 (.D(r_word_31__N_964[14]), .SP(dac_clk_p_c_enable_647), 
            .CK(dac_clk_p_c), .Q(r_word[14])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i14.GSR = "DISABLED";
    FD1P3AX r_word_i13 (.D(r_word_31__N_964[13]), .SP(dac_clk_p_c_enable_647), 
            .CK(dac_clk_p_c), .Q(r_word[13])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i13.GSR = "DISABLED";
    FD1P3AX r_word_i12 (.D(r_word_31__N_964[12]), .SP(dac_clk_p_c_enable_647), 
            .CK(dac_clk_p_c), .Q(r_word[12])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i12.GSR = "DISABLED";
    FD1P3AX r_word_i11 (.D(r_word_31__N_964[11]), .SP(dac_clk_p_c_enable_647), 
            .CK(dac_clk_p_c), .Q(r_word[11])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i11.GSR = "DISABLED";
    FD1P3AX r_word_i10 (.D(r_word_31__N_964[10]), .SP(dac_clk_p_c_enable_647), 
            .CK(dac_clk_p_c), .Q(r_word[10])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i10.GSR = "DISABLED";
    FD1P3AX r_word_i9 (.D(r_word_31__N_964[9]), .SP(dac_clk_p_c_enable_647), 
            .CK(dac_clk_p_c), .Q(r_word[9])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i9.GSR = "DISABLED";
    FD1P3AX r_word_i8 (.D(r_word_31__N_964[8]), .SP(dac_clk_p_c_enable_647), 
            .CK(dac_clk_p_c), .Q(r_word[8])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i8.GSR = "DISABLED";
    FD1P3AX r_word_i7 (.D(r_word_31__N_964[7]), .SP(dac_clk_p_c_enable_647), 
            .CK(dac_clk_p_c), .Q(r_word[7])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i7.GSR = "DISABLED";
    FD1P3AX r_word_i6 (.D(r_word_31__N_964[6]), .SP(dac_clk_p_c_enable_647), 
            .CK(dac_clk_p_c), .Q(r_word[6])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i6.GSR = "DISABLED";
    FD1P3AX r_word_i5 (.D(r_word_31__N_964[5]), .SP(dac_clk_p_c_enable_647), 
            .CK(dac_clk_p_c), .Q(r_word[5])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i5.GSR = "DISABLED";
    FD1P3AX r_word_i4 (.D(r_word_31__N_964[4]), .SP(dac_clk_p_c_enable_647), 
            .CK(dac_clk_p_c), .Q(r_word[4])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i4.GSR = "DISABLED";
    LUT4 i1_3_lut_4_lut_3_lut_4_lut (.A(r_len[0]), .B(r_len[1]), .C(r_len[2]), 
         .D(r_len[3]), .Z(n12776)) /* synthesis lut_function=(A (B)+!A !(B+!(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(80[14:26])
    defparam i1_3_lut_4_lut_3_lut_4_lut.init = 16'h9998;
    LUT4 r_word_29__bdd_3_lut_24851 (.A(idl_word[30]), .B(idl_word[33]), 
         .C(idl_word[32]), .Z(n26463)) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam r_word_29__bdd_3_lut_24851.init = 16'h8c8c;
    FD1P3IX r_len__i2 (.D(n12780), .SP(dac_clk_p_c_enable_312), .CD(n29196), 
            .CK(dac_clk_p_c), .Q(r_len[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(64[9] 81[6])
    defparam r_len__i2.GSR = "DISABLED";
    FD1P3IX r_len__i1 (.D(n12776), .SP(dac_clk_p_c_enable_312), .CD(n29196), 
            .CK(dac_clk_p_c), .Q(r_len[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(64[9] 81[6])
    defparam r_len__i1.GSR = "DISABLED";
    LUT4 o_dw_bits_4__I_0_i3_4_lut (.A(r_word[30]), .B(idl_word[31]), .C(n29366), 
         .D(n29364), .Z(o_dw_bits_4__N_955[2])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(102[12] 103[41])
    defparam o_dw_bits_4__I_0_i3_4_lut.init = 16'hca0a;
    LUT4 mux_15_i4_4_lut (.A(r_len[3]), .B(n29364), .C(n29366), .D(n22051), 
         .Z(r_len_3__N_996[3])) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(76[12] 81[6])
    defparam mux_15_i4_4_lut.init = 16'h3a35;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n29366), .B(n32125), .C(nl_busy), .D(hx_stb), 
         .Z(dac_clk_p_c_enable_168)) /* synthesis lut_function=(A+(B+!(C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'hefff;
    LUT4 r_word_28__bdd_3_lut_26923 (.A(idl_word[29]), .B(idl_word[32]), 
         .C(idl_word[33]), .Z(n28875)) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam r_word_28__bdd_3_lut_26923.init = 16'h8c8c;
    LUT4 i3_4_lut_rep_792 (.A(r_len[0]), .B(r_len[1]), .C(r_len[2]), .D(r_len[3]), 
         .Z(n29452)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(78[16:31])
    defparam i3_4_lut_rep_792.init = 16'hfffe;
    LUT4 i1_2_lut_4_lut (.A(r_len[0]), .B(r_len[1]), .C(r_len[2]), .D(r_len[3]), 
         .Z(n13[0])) /* synthesis lut_function=(!(A+!(B+(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(78[16:31])
    defparam i1_2_lut_4_lut.init = 16'h5554;
    LUT4 i1_3_lut_3_lut_4_lut (.A(r_len[0]), .B(r_len[1]), .C(r_len[3]), 
         .D(r_len[2]), .Z(n12780)) /* synthesis lut_function=(A (D)+!A (B (D)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(80[14:26])
    defparam i1_3_lut_3_lut_4_lut.init = 16'hee10;
    LUT4 i1_4_lut_4_lut (.A(r_len[0]), .B(r_len[1]), .C(r_len[3]), .D(r_len[2]), 
         .Z(n22051)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(80[14:26])
    defparam i1_4_lut_4_lut.init = 16'hffef;
    LUT4 i12434_2_lut_rep_704 (.A(idl_word[32]), .B(idl_word[33]), .Z(n29364)) /* synthesis lut_function=(A (B)) */ ;
    defparam i12434_2_lut_rep_704.init = 16'h8888;
    LUT4 o_dw_bits_4__I_0_i4_3_lut_4_lut (.A(idl_word[32]), .B(idl_word[33]), 
         .C(n29366), .D(r_word[31]), .Z(o_dw_bits_4__N_955[3])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam o_dw_bits_4__I_0_i4_3_lut_4_lut.init = 16'h8f80;
    LUT4 i_stb_I_0_2_lut_rep_706 (.A(idl_stb), .B(hb_busy), .Z(n29366)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam i_stb_I_0_2_lut_rep_706.init = 16'h2222;
    LUT4 i24602_2_lut_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(nl_busy), 
         .D(hx_stb), .Z(n14220)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam i24602_2_lut_3_lut_4_lut.init = 16'h0ddd;
    LUT4 r_word_31__I_0_i32_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[31]), 
         .D(r_word[27]), .Z(r_word_31__N_964[31])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i32_3_lut_4_lut.init = 16'hfd20;
    LUT4 i1_2_lut_3_lut_4_lut_adj_211 (.A(idl_stb), .B(hb_busy), .C(nl_busy), 
         .D(hx_stb), .Z(dac_clk_p_c_enable_647)) /* synthesis lut_function=(!(A (B (C (D)))+!A (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam i1_2_lut_3_lut_4_lut_adj_211.init = 16'h2fff;
    LUT4 i12443_2_lut_3_lut (.A(idl_stb), .B(hb_busy), .C(n29452), .Z(o_dw_busy_N_1036)) /* synthesis lut_function=(A ((C)+!B)+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam i12443_2_lut_3_lut.init = 16'hf2f2;
    LUT4 i1_2_lut_rep_536_3_lut (.A(idl_stb), .B(hb_busy), .C(n32125), 
         .Z(n29196)) /* synthesis lut_function=(A ((C)+!B)+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam i1_2_lut_rep_536_3_lut.init = 16'hf2f2;
    LUT4 r_word_28__bdd_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(n28875), 
         .D(r_word[28]), .Z(o_dw_bits_4__N_955[0])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_28__bdd_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_29__bdd_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(n26463), 
         .D(r_word[29]), .Z(o_dw_bits_4__N_955[1])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_29__bdd_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i31_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[30]), 
         .D(r_word[26]), .Z(r_word_31__N_964[30])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i31_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i30_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[29]), 
         .D(r_word[25]), .Z(r_word_31__N_964[29])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i30_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i29_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[28]), 
         .D(r_word[24]), .Z(r_word_31__N_964[28])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i29_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i28_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[27]), 
         .D(r_word[23]), .Z(r_word_31__N_964[27])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i28_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i27_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[26]), 
         .D(r_word[22]), .Z(r_word_31__N_964[26])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i27_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i26_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[25]), 
         .D(r_word[21]), .Z(r_word_31__N_964[25])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i26_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i25_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[24]), 
         .D(r_word[20]), .Z(r_word_31__N_964[24])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i25_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i24_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[23]), 
         .D(r_word[19]), .Z(r_word_31__N_964[23])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i24_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i23_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[22]), 
         .D(r_word[18]), .Z(r_word_31__N_964[22])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i23_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i22_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[21]), 
         .D(r_word[17]), .Z(r_word_31__N_964[21])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i22_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i21_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[20]), 
         .D(r_word[16]), .Z(r_word_31__N_964[20])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i21_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i20_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[19]), 
         .D(r_word[15]), .Z(r_word_31__N_964[19])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i20_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i19_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[18]), 
         .D(r_word[14]), .Z(r_word_31__N_964[18])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i19_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i18_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[17]), 
         .D(r_word[13]), .Z(r_word_31__N_964[17])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i18_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i17_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[16]), 
         .D(r_word[12]), .Z(r_word_31__N_964[16])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i17_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i16_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[15]), 
         .D(r_word[11]), .Z(r_word_31__N_964[15])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i16_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i15_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[14]), 
         .D(r_word[10]), .Z(r_word_31__N_964[14])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i15_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i14_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[13]), 
         .D(r_word[9]), .Z(r_word_31__N_964[13])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i14_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i13_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[12]), 
         .D(r_word[8]), .Z(r_word_31__N_964[12])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i13_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i12_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[11]), 
         .D(r_word[7]), .Z(r_word_31__N_964[11])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i12_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i11_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[10]), 
         .D(r_word[6]), .Z(r_word_31__N_964[10])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i11_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i10_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[9]), 
         .D(r_word[5]), .Z(r_word_31__N_964[9])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i10_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i9_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[8]), 
         .D(r_word[4]), .Z(r_word_31__N_964[8])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i9_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i8_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[7]), 
         .D(r_word[3]), .Z(r_word_31__N_964[7])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i8_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i7_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[6]), 
         .D(r_word[2]), .Z(r_word_31__N_964[6])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i7_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i6_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[5]), 
         .D(r_word[1]), .Z(r_word_31__N_964[5])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i6_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i5_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[4]), 
         .D(r_word[0]), .Z(r_word_31__N_964[4])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i5_3_lut_4_lut.init = 16'hfd20;
    FD1P3AX o_dw_bits_i3 (.D(o_dw_bits_4__N_955[3]), .SP(dac_clk_p_c_enable_647), 
            .CK(dac_clk_p_c), .Q(hb_bits[3])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(95[9] 103[41])
    defparam o_dw_bits_i3.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module hbpack
//

module hbpack (iw_word, dac_clk_p_c, dac_clk_p_c_enable_548, n32126, 
            cmd_loaded, dac_clk_p_c_enable_166, w_reset, cmd_loaded_N_535, 
            iw_stb, o_pck_stb_N_532, \dec_bits[0] , \dec_bits[4] , dac_clk_p_c_enable_517, 
            \dec_bits[1] , n45, n46) /* synthesis syn_module_defined=1 */ ;
    output [33:0]iw_word;
    input dac_clk_p_c;
    input dac_clk_p_c_enable_548;
    input n32126;
    output cmd_loaded;
    input dac_clk_p_c_enable_166;
    input w_reset;
    input cmd_loaded_N_535;
    output iw_stb;
    input o_pck_stb_N_532;
    input \dec_bits[0] ;
    input \dec_bits[4] ;
    input dac_clk_p_c_enable_517;
    input \dec_bits[1] ;
    input n45;
    input n46;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[29:38])
    wire [33:0]r_word;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(71[13:19])
    wire [33:0]n14;
    
    FD1P3IX o_pck_word__i0 (.D(r_word[0]), .SP(dac_clk_p_c_enable_548), 
            .CD(n32126), .CK(dac_clk_p_c), .Q(iw_word[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i0.GSR = "DISABLED";
    FD1P3IX cmd_loaded_23 (.D(cmd_loaded_N_535), .SP(dac_clk_p_c_enable_166), 
            .CD(w_reset), .CK(dac_clk_p_c), .Q(cmd_loaded)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(74[9] 80[23])
    defparam cmd_loaded_23.GSR = "DISABLED";
    FD1S3IX o_pck_stb_24 (.D(o_pck_stb_N_532), .CK(dac_clk_p_c), .CD(n32126), 
            .Q(iw_stb)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(83[9] 84[65])
    defparam o_pck_stb_24.GSR = "DISABLED";
    FD1P3IX r_word__i0 (.D(n14[0]), .SP(dac_clk_p_c_enable_548), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i0.GSR = "DISABLED";
    FD1P3IX o_pck_word__i33 (.D(r_word[33]), .SP(dac_clk_p_c_enable_548), 
            .CD(w_reset), .CK(dac_clk_p_c), .Q(iw_word[33])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i33.GSR = "DISABLED";
    FD1P3IX o_pck_word__i32 (.D(r_word[32]), .SP(dac_clk_p_c_enable_548), 
            .CD(w_reset), .CK(dac_clk_p_c), .Q(iw_word[32])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i32.GSR = "DISABLED";
    FD1P3IX o_pck_word__i31 (.D(r_word[31]), .SP(dac_clk_p_c_enable_548), 
            .CD(w_reset), .CK(dac_clk_p_c), .Q(iw_word[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i31.GSR = "DISABLED";
    FD1P3IX o_pck_word__i30 (.D(r_word[30]), .SP(dac_clk_p_c_enable_548), 
            .CD(w_reset), .CK(dac_clk_p_c), .Q(iw_word[30])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i30.GSR = "DISABLED";
    FD1P3IX o_pck_word__i29 (.D(r_word[29]), .SP(dac_clk_p_c_enable_548), 
            .CD(w_reset), .CK(dac_clk_p_c), .Q(iw_word[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i29.GSR = "DISABLED";
    FD1P3IX o_pck_word__i28 (.D(r_word[28]), .SP(dac_clk_p_c_enable_548), 
            .CD(w_reset), .CK(dac_clk_p_c), .Q(iw_word[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i28.GSR = "DISABLED";
    FD1P3IX o_pck_word__i27 (.D(r_word[27]), .SP(dac_clk_p_c_enable_548), 
            .CD(w_reset), .CK(dac_clk_p_c), .Q(iw_word[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i27.GSR = "DISABLED";
    FD1P3IX o_pck_word__i26 (.D(r_word[26]), .SP(dac_clk_p_c_enable_548), 
            .CD(w_reset), .CK(dac_clk_p_c), .Q(iw_word[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i26.GSR = "DISABLED";
    FD1P3IX o_pck_word__i25 (.D(r_word[25]), .SP(dac_clk_p_c_enable_548), 
            .CD(w_reset), .CK(dac_clk_p_c), .Q(iw_word[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i25.GSR = "DISABLED";
    FD1P3IX o_pck_word__i24 (.D(r_word[24]), .SP(dac_clk_p_c_enable_548), 
            .CD(w_reset), .CK(dac_clk_p_c), .Q(iw_word[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i24.GSR = "DISABLED";
    FD1P3IX o_pck_word__i23 (.D(r_word[23]), .SP(dac_clk_p_c_enable_548), 
            .CD(w_reset), .CK(dac_clk_p_c), .Q(iw_word[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i23.GSR = "DISABLED";
    FD1P3IX o_pck_word__i22 (.D(r_word[22]), .SP(dac_clk_p_c_enable_548), 
            .CD(w_reset), .CK(dac_clk_p_c), .Q(iw_word[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i22.GSR = "DISABLED";
    FD1P3IX o_pck_word__i21 (.D(r_word[21]), .SP(dac_clk_p_c_enable_548), 
            .CD(w_reset), .CK(dac_clk_p_c), .Q(iw_word[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i21.GSR = "DISABLED";
    FD1P3IX o_pck_word__i20 (.D(r_word[20]), .SP(dac_clk_p_c_enable_548), 
            .CD(w_reset), .CK(dac_clk_p_c), .Q(iw_word[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i20.GSR = "DISABLED";
    FD1P3IX o_pck_word__i19 (.D(r_word[19]), .SP(dac_clk_p_c_enable_548), 
            .CD(w_reset), .CK(dac_clk_p_c), .Q(iw_word[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i19.GSR = "DISABLED";
    FD1P3IX o_pck_word__i18 (.D(r_word[18]), .SP(dac_clk_p_c_enable_548), 
            .CD(n32126), .CK(dac_clk_p_c), .Q(iw_word[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i18.GSR = "DISABLED";
    FD1P3IX o_pck_word__i17 (.D(r_word[17]), .SP(dac_clk_p_c_enable_548), 
            .CD(w_reset), .CK(dac_clk_p_c), .Q(iw_word[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i17.GSR = "DISABLED";
    FD1P3IX o_pck_word__i16 (.D(r_word[16]), .SP(dac_clk_p_c_enable_548), 
            .CD(n32126), .CK(dac_clk_p_c), .Q(iw_word[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i16.GSR = "DISABLED";
    FD1P3IX o_pck_word__i15 (.D(r_word[15]), .SP(dac_clk_p_c_enable_548), 
            .CD(n32126), .CK(dac_clk_p_c), .Q(iw_word[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i15.GSR = "DISABLED";
    FD1P3IX o_pck_word__i14 (.D(r_word[14]), .SP(dac_clk_p_c_enable_548), 
            .CD(n32126), .CK(dac_clk_p_c), .Q(iw_word[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i14.GSR = "DISABLED";
    FD1P3IX o_pck_word__i13 (.D(r_word[13]), .SP(dac_clk_p_c_enable_548), 
            .CD(n32126), .CK(dac_clk_p_c), .Q(iw_word[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i13.GSR = "DISABLED";
    FD1P3IX o_pck_word__i12 (.D(r_word[12]), .SP(dac_clk_p_c_enable_548), 
            .CD(n32126), .CK(dac_clk_p_c), .Q(iw_word[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i12.GSR = "DISABLED";
    FD1P3IX o_pck_word__i11 (.D(r_word[11]), .SP(dac_clk_p_c_enable_548), 
            .CD(n32126), .CK(dac_clk_p_c), .Q(iw_word[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i11.GSR = "DISABLED";
    FD1P3IX o_pck_word__i10 (.D(r_word[10]), .SP(dac_clk_p_c_enable_548), 
            .CD(n32126), .CK(dac_clk_p_c), .Q(iw_word[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i10.GSR = "DISABLED";
    FD1P3IX o_pck_word__i9 (.D(r_word[9]), .SP(dac_clk_p_c_enable_548), 
            .CD(n32126), .CK(dac_clk_p_c), .Q(iw_word[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i9.GSR = "DISABLED";
    FD1P3IX o_pck_word__i8 (.D(r_word[8]), .SP(dac_clk_p_c_enable_548), 
            .CD(n32126), .CK(dac_clk_p_c), .Q(iw_word[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i8.GSR = "DISABLED";
    FD1P3IX o_pck_word__i7 (.D(r_word[7]), .SP(dac_clk_p_c_enable_548), 
            .CD(n32126), .CK(dac_clk_p_c), .Q(iw_word[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i7.GSR = "DISABLED";
    FD1P3IX o_pck_word__i6 (.D(r_word[6]), .SP(dac_clk_p_c_enable_548), 
            .CD(n32126), .CK(dac_clk_p_c), .Q(iw_word[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i6.GSR = "DISABLED";
    FD1P3IX o_pck_word__i5 (.D(r_word[5]), .SP(dac_clk_p_c_enable_548), 
            .CD(n32126), .CK(dac_clk_p_c), .Q(iw_word[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i5.GSR = "DISABLED";
    FD1P3IX o_pck_word__i4 (.D(r_word[4]), .SP(dac_clk_p_c_enable_548), 
            .CD(n32126), .CK(dac_clk_p_c), .Q(iw_word[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i4.GSR = "DISABLED";
    FD1P3IX o_pck_word__i3 (.D(r_word[3]), .SP(dac_clk_p_c_enable_548), 
            .CD(n32126), .CK(dac_clk_p_c), .Q(iw_word[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i3.GSR = "DISABLED";
    FD1P3IX o_pck_word__i2 (.D(r_word[2]), .SP(dac_clk_p_c_enable_548), 
            .CD(n32126), .CK(dac_clk_p_c), .Q(iw_word[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i2.GSR = "DISABLED";
    FD1P3IX o_pck_word__i1 (.D(r_word[1]), .SP(dac_clk_p_c_enable_548), 
            .CD(n32126), .CK(dac_clk_p_c), .Q(iw_word[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i1.GSR = "DISABLED";
    LUT4 i12429_2_lut (.A(\dec_bits[0] ), .B(\dec_bits[4] ), .Z(n14[0])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i12429_2_lut.init = 16'h2222;
    FD1P3IX r_word__i33 (.D(\dec_bits[1] ), .SP(dac_clk_p_c_enable_517), 
            .CD(n32126), .CK(dac_clk_p_c), .Q(r_word[33])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i33.GSR = "DISABLED";
    FD1P3IX r_word__i32 (.D(\dec_bits[0] ), .SP(dac_clk_p_c_enable_517), 
            .CD(n32126), .CK(dac_clk_p_c), .Q(r_word[32])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i32.GSR = "DISABLED";
    FD1P3IX r_word__i31 (.D(n14[31]), .SP(dac_clk_p_c_enable_548), .CD(n32126), 
            .CK(dac_clk_p_c), .Q(r_word[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i31.GSR = "DISABLED";
    FD1P3IX r_word__i30 (.D(n14[30]), .SP(dac_clk_p_c_enable_548), .CD(n32126), 
            .CK(dac_clk_p_c), .Q(r_word[30])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i30.GSR = "DISABLED";
    FD1P3IX r_word__i29 (.D(n14[29]), .SP(dac_clk_p_c_enable_548), .CD(n32126), 
            .CK(dac_clk_p_c), .Q(r_word[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i29.GSR = "DISABLED";
    FD1P3IX r_word__i28 (.D(n14[28]), .SP(dac_clk_p_c_enable_548), .CD(n32126), 
            .CK(dac_clk_p_c), .Q(r_word[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i28.GSR = "DISABLED";
    FD1P3IX r_word__i27 (.D(n14[27]), .SP(dac_clk_p_c_enable_548), .CD(n32126), 
            .CK(dac_clk_p_c), .Q(r_word[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i27.GSR = "DISABLED";
    FD1P3IX r_word__i26 (.D(n14[26]), .SP(dac_clk_p_c_enable_548), .CD(n32126), 
            .CK(dac_clk_p_c), .Q(r_word[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i26.GSR = "DISABLED";
    FD1P3IX r_word__i25 (.D(n14[25]), .SP(dac_clk_p_c_enable_548), .CD(n32126), 
            .CK(dac_clk_p_c), .Q(r_word[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i25.GSR = "DISABLED";
    FD1P3IX r_word__i24 (.D(n14[24]), .SP(dac_clk_p_c_enable_548), .CD(n32126), 
            .CK(dac_clk_p_c), .Q(r_word[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i24.GSR = "DISABLED";
    FD1P3IX r_word__i23 (.D(n14[23]), .SP(dac_clk_p_c_enable_548), .CD(n32126), 
            .CK(dac_clk_p_c), .Q(r_word[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i23.GSR = "DISABLED";
    FD1P3IX r_word__i22 (.D(n14[22]), .SP(dac_clk_p_c_enable_548), .CD(n32126), 
            .CK(dac_clk_p_c), .Q(r_word[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i22.GSR = "DISABLED";
    FD1P3IX r_word__i21 (.D(n14[21]), .SP(dac_clk_p_c_enable_548), .CD(n32126), 
            .CK(dac_clk_p_c), .Q(r_word[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i21.GSR = "DISABLED";
    FD1P3IX r_word__i20 (.D(n14[20]), .SP(dac_clk_p_c_enable_548), .CD(n32126), 
            .CK(dac_clk_p_c), .Q(r_word[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i20.GSR = "DISABLED";
    FD1P3IX r_word__i19 (.D(n14[19]), .SP(dac_clk_p_c_enable_548), .CD(n32126), 
            .CK(dac_clk_p_c), .Q(r_word[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i19.GSR = "DISABLED";
    FD1P3IX r_word__i18 (.D(n14[18]), .SP(dac_clk_p_c_enable_548), .CD(n32126), 
            .CK(dac_clk_p_c), .Q(r_word[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i18.GSR = "DISABLED";
    FD1P3IX r_word__i17 (.D(n14[17]), .SP(dac_clk_p_c_enable_548), .CD(n32126), 
            .CK(dac_clk_p_c), .Q(r_word[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i17.GSR = "DISABLED";
    FD1P3IX r_word__i16 (.D(n14[16]), .SP(dac_clk_p_c_enable_548), .CD(n32126), 
            .CK(dac_clk_p_c), .Q(r_word[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i16.GSR = "DISABLED";
    FD1P3IX r_word__i15 (.D(n14[15]), .SP(dac_clk_p_c_enable_548), .CD(n32126), 
            .CK(dac_clk_p_c), .Q(r_word[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i15.GSR = "DISABLED";
    FD1P3IX r_word__i14 (.D(n14[14]), .SP(dac_clk_p_c_enable_548), .CD(n32126), 
            .CK(dac_clk_p_c), .Q(r_word[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i14.GSR = "DISABLED";
    FD1P3IX r_word__i13 (.D(n14[13]), .SP(dac_clk_p_c_enable_548), .CD(n32126), 
            .CK(dac_clk_p_c), .Q(r_word[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i13.GSR = "DISABLED";
    FD1P3IX r_word__i12 (.D(n14[12]), .SP(dac_clk_p_c_enable_548), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i12.GSR = "DISABLED";
    FD1P3IX r_word__i11 (.D(n14[11]), .SP(dac_clk_p_c_enable_548), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i11.GSR = "DISABLED";
    FD1P3IX r_word__i10 (.D(n14[10]), .SP(dac_clk_p_c_enable_548), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i10.GSR = "DISABLED";
    FD1P3IX r_word__i9 (.D(n14[9]), .SP(dac_clk_p_c_enable_548), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i9.GSR = "DISABLED";
    FD1P3IX r_word__i8 (.D(n14[8]), .SP(dac_clk_p_c_enable_548), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i8.GSR = "DISABLED";
    FD1P3IX r_word__i7 (.D(n14[7]), .SP(dac_clk_p_c_enable_548), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i7.GSR = "DISABLED";
    FD1P3IX r_word__i6 (.D(n14[6]), .SP(dac_clk_p_c_enable_548), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i6.GSR = "DISABLED";
    FD1P3IX r_word__i5 (.D(n14[5]), .SP(dac_clk_p_c_enable_548), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i5.GSR = "DISABLED";
    FD1P3IX r_word__i4 (.D(n14[4]), .SP(dac_clk_p_c_enable_548), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i4.GSR = "DISABLED";
    FD1P3IX r_word__i3 (.D(n45), .SP(dac_clk_p_c_enable_548), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i3.GSR = "DISABLED";
    FD1P3IX r_word__i2 (.D(n46), .SP(dac_clk_p_c_enable_548), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i2.GSR = "DISABLED";
    FD1P3IX r_word__i1 (.D(n14[1]), .SP(dac_clk_p_c_enable_548), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i1.GSR = "DISABLED";
    LUT4 i12625_2_lut (.A(r_word[27]), .B(\dec_bits[4] ), .Z(n14[31])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i12625_2_lut.init = 16'h2222;
    LUT4 i12626_2_lut (.A(r_word[26]), .B(\dec_bits[4] ), .Z(n14[30])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i12626_2_lut.init = 16'h2222;
    LUT4 i12627_2_lut (.A(r_word[25]), .B(\dec_bits[4] ), .Z(n14[29])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i12627_2_lut.init = 16'h2222;
    LUT4 i12628_2_lut (.A(r_word[24]), .B(\dec_bits[4] ), .Z(n14[28])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i12628_2_lut.init = 16'h2222;
    LUT4 i12629_2_lut (.A(r_word[23]), .B(\dec_bits[4] ), .Z(n14[27])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i12629_2_lut.init = 16'h2222;
    LUT4 i12630_2_lut (.A(r_word[22]), .B(\dec_bits[4] ), .Z(n14[26])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i12630_2_lut.init = 16'h2222;
    LUT4 i12631_2_lut (.A(r_word[21]), .B(\dec_bits[4] ), .Z(n14[25])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i12631_2_lut.init = 16'h2222;
    LUT4 i12632_2_lut (.A(r_word[20]), .B(\dec_bits[4] ), .Z(n14[24])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i12632_2_lut.init = 16'h2222;
    LUT4 i12633_2_lut (.A(r_word[19]), .B(\dec_bits[4] ), .Z(n14[23])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i12633_2_lut.init = 16'h2222;
    LUT4 i12634_2_lut (.A(r_word[18]), .B(\dec_bits[4] ), .Z(n14[22])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i12634_2_lut.init = 16'h2222;
    LUT4 i12635_2_lut (.A(r_word[17]), .B(\dec_bits[4] ), .Z(n14[21])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i12635_2_lut.init = 16'h2222;
    LUT4 i12636_2_lut (.A(r_word[16]), .B(\dec_bits[4] ), .Z(n14[20])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i12636_2_lut.init = 16'h2222;
    LUT4 i12637_2_lut (.A(r_word[15]), .B(\dec_bits[4] ), .Z(n14[19])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i12637_2_lut.init = 16'h2222;
    LUT4 i12638_2_lut (.A(r_word[14]), .B(\dec_bits[4] ), .Z(n14[18])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i12638_2_lut.init = 16'h2222;
    LUT4 i12639_2_lut (.A(r_word[13]), .B(\dec_bits[4] ), .Z(n14[17])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i12639_2_lut.init = 16'h2222;
    LUT4 i12640_2_lut (.A(r_word[12]), .B(\dec_bits[4] ), .Z(n14[16])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i12640_2_lut.init = 16'h2222;
    LUT4 i12641_2_lut (.A(r_word[11]), .B(\dec_bits[4] ), .Z(n14[15])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i12641_2_lut.init = 16'h2222;
    LUT4 i12642_2_lut (.A(r_word[10]), .B(\dec_bits[4] ), .Z(n14[14])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i12642_2_lut.init = 16'h2222;
    LUT4 i12643_2_lut (.A(r_word[9]), .B(\dec_bits[4] ), .Z(n14[13])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i12643_2_lut.init = 16'h2222;
    LUT4 i12644_2_lut (.A(r_word[8]), .B(\dec_bits[4] ), .Z(n14[12])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i12644_2_lut.init = 16'h2222;
    LUT4 i12645_2_lut (.A(r_word[7]), .B(\dec_bits[4] ), .Z(n14[11])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i12645_2_lut.init = 16'h2222;
    LUT4 i12646_2_lut (.A(r_word[6]), .B(\dec_bits[4] ), .Z(n14[10])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i12646_2_lut.init = 16'h2222;
    LUT4 i12647_2_lut (.A(r_word[5]), .B(\dec_bits[4] ), .Z(n14[9])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i12647_2_lut.init = 16'h2222;
    LUT4 i12648_2_lut (.A(r_word[4]), .B(\dec_bits[4] ), .Z(n14[8])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i12648_2_lut.init = 16'h2222;
    LUT4 i12649_2_lut (.A(r_word[3]), .B(\dec_bits[4] ), .Z(n14[7])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i12649_2_lut.init = 16'h2222;
    LUT4 i12671_2_lut (.A(r_word[2]), .B(\dec_bits[4] ), .Z(n14[6])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i12671_2_lut.init = 16'h2222;
    LUT4 i12672_2_lut (.A(r_word[1]), .B(\dec_bits[4] ), .Z(n14[5])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i12672_2_lut.init = 16'h2222;
    LUT4 i12673_2_lut (.A(r_word[0]), .B(\dec_bits[4] ), .Z(n14[4])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i12673_2_lut.init = 16'h2222;
    LUT4 i12674_2_lut (.A(\dec_bits[1] ), .B(\dec_bits[4] ), .Z(n14[1])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i12674_2_lut.init = 16'h2222;
    
endmodule
//
// Verilog Description of module hbgenhex
//

module hbgenhex (hx_stb, dac_clk_p_c, n32126, hb_busy, hb_bits, \w_gx_char[0] , 
            \w_gx_char[1] , \w_gx_char[2] , \w_gx_char[3] , \w_gx_char[4] , 
            \w_gx_char[5] , \w_gx_char[6] , dac_clk_p_c_enable_312, GND_net, 
            VCC_net, nl_busy, n32125) /* synthesis syn_module_defined=1 */ ;
    output hx_stb;
    input dac_clk_p_c;
    input n32126;
    input hb_busy;
    input [4:0]hb_bits;
    output \w_gx_char[0] ;
    output \w_gx_char[1] ;
    output \w_gx_char[2] ;
    output \w_gx_char[3] ;
    output \w_gx_char[4] ;
    output \w_gx_char[5] ;
    output \w_gx_char[6] ;
    output dac_clk_p_c_enable_312;
    input GND_net;
    input VCC_net;
    input nl_busy;
    input n32125;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[29:38])
    
    wire dac_clk_p_c_enable_66;
    
    FD1P3IX o_gx_stb_13 (.D(hb_busy), .SP(dac_clk_p_c_enable_66), .CD(n32126), 
            .CK(dac_clk_p_c), .Q(hx_stb)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=132, LSE_RLINE=133 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbgenhex.v(74[9] 78[21])
    defparam o_gx_stb_13.GSR = "DISABLED";
    SP8KC mux_60 (.DI0(GND_net), .DI1(GND_net), .DI2(GND_net), .DI3(GND_net), 
          .DI4(GND_net), .DI5(GND_net), .DI6(GND_net), .DI7(GND_net), 
          .DI8(GND_net), .AD0(GND_net), .AD1(GND_net), .AD2(GND_net), 
          .AD3(hb_bits[0]), .AD4(hb_bits[1]), .AD5(hb_bits[2]), .AD6(hb_bits[3]), 
          .AD7(hb_bits[4]), .AD8(GND_net), .AD9(GND_net), .AD10(GND_net), 
          .AD11(GND_net), .AD12(GND_net), .CE(dac_clk_p_c_enable_312), 
          .OCE(VCC_net), .CLK(dac_clk_p_c), .WE(GND_net), .CS0(GND_net), 
          .CS1(GND_net), .CS2(GND_net), .RST(GND_net), .DO0(\w_gx_char[0] ), 
          .DO1(\w_gx_char[1] ), .DO2(\w_gx_char[2] ), .DO3(\w_gx_char[3] ), 
          .DO4(\w_gx_char[4] ), .DO5(\w_gx_char[5] ), .DO6(\w_gx_char[6] ));
    defparam mux_60.DATA_WIDTH = 9;
    defparam mux_60.REGMODE = "NOREG";
    defparam mux_60.CSDECODE = "0b000";
    defparam mux_60.WRITEMODE = "NORMAL";
    defparam mux_60.GSR = "DISABLED";
    defparam mux_60.RESETMODE = "ASYNC";
    defparam mux_60.ASYNC_RESET_RELEASE = "SYNC";
    defparam mux_60.INIT_DATA = "STATIC";
    defparam mux_60.INITVAL_00 = "0x01A0D01A0D0B44908A5401A0D01A0D0A641096520CC650C8630C4610723806E3606A340663206230";
    defparam mux_60.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_60.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_60.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_60.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_60.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_60.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_60.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_60.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_60.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_60.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_60.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_60.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_60.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_60.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_60.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_60.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_60.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_60.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_60.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_60.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_60.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_60.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_60.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_60.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_60.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_60.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_60.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_60.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_60.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_60.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_60.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    LUT4 i24589_2_lut_rep_511 (.A(hx_stb), .B(nl_busy), .Z(dac_clk_p_c_enable_312)) /* synthesis lut_function=(!(A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(76[16:26])
    defparam i24589_2_lut_rep_511.init = 16'h7777;
    LUT4 i1134_2_lut_3_lut (.A(hx_stb), .B(nl_busy), .C(n32125), .Z(dac_clk_p_c_enable_66)) /* synthesis lut_function=(((C)+!B)+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(76[16:26])
    defparam i1134_2_lut_3_lut.init = 16'hf7f7;
    
endmodule
//
// Verilog Description of module hbdechex
//

module hbdechex (dec_bits, dac_clk_p_c, w_reset, n32126, \rx_data[1] , 
            \rx_data[2] , \rx_data[0] , \rx_data[3] , \rx_data[5] , 
            \rx_data[6] , \rx_data[4] , rx_stb, \dec_bits[1] , n32125, 
            dac_clk_p_c_enable_548, dac_clk_p_c_enable_517, n45, n46, 
            dac_clk_p_c_enable_166, cmd_loaded_N_535, cmd_loaded, o_pck_stb_N_532) /* synthesis syn_module_defined=1 */ ;
    output [4:0]dec_bits;
    input dac_clk_p_c;
    output w_reset;
    output n32126;
    input \rx_data[1] ;
    input \rx_data[2] ;
    input \rx_data[0] ;
    input \rx_data[3] ;
    input \rx_data[5] ;
    input \rx_data[6] ;
    input \rx_data[4] ;
    input rx_stb;
    output \dec_bits[1] ;
    output n32125;
    output dac_clk_p_c_enable_548;
    output dac_clk_p_c_enable_517;
    output n45;
    output n46;
    output dac_clk_p_c_enable_166;
    output cmd_loaded_N_535;
    input cmd_loaded;
    output o_pck_stb_N_532;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[29:38])
    wire [4:0]o_dh_bits_4__N_363;
    
    wire dec_stb, o_dh_stb_N_390, o_reset_N_392, n4, n29449, n31063, 
        n31065, n32017, n21770, n22272, n55, n50, n29094, n22129, 
        n47, n22790, n29411, n22312, n9;
    wire [4:0]dec_bits_c;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(69[13:21])
    
    wire n27668, n27667, n27670, n27669, n27671, n19, n27699, 
        n22344, n41, n31062, n31061, n32057, n29093, n29410, n29543, 
        n29542, n29450, n29187, n29544, n49, n22280, n29191, n22278, 
        n42, n62, n34, n29303, n53, n21615;
    
    FD1S3AX o_dh_bits_i0 (.D(o_dh_bits_4__N_363[0]), .CK(dac_clk_p_c), .Q(dec_bits[0])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=11, LSE_RCOL=30, LSE_LLINE=93, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(60[9] 100[5])
    defparam o_dh_bits_i0.GSR = "DISABLED";
    FD1S3AX o_dh_stb_35 (.D(o_dh_stb_N_390), .CK(dac_clk_p_c), .Q(dec_stb)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=11, LSE_RCOL=30, LSE_LLINE=93, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(57[9] 58[47])
    defparam o_dh_stb_35.GSR = "DISABLED";
    FD1S3AY o_reset_34 (.D(o_reset_N_392), .CK(dac_clk_p_c), .Q(w_reset)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=9, LSE_LCOL=11, LSE_RCOL=30, LSE_LLINE=93, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(53[9] 54[46])
    defparam o_reset_34.GSR = "DISABLED";
    FD1S3AY o_reset_34_rep_858 (.D(o_reset_N_392), .CK(dac_clk_p_c), .Q(n32126)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=9, LSE_LCOL=11, LSE_RCOL=30, LSE_LLINE=93, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(53[9] 54[46])
    defparam o_reset_34_rep_858.GSR = "DISABLED";
    LUT4 i1_3_lut_4_lut_3_lut (.A(\rx_data[1] ), .B(\rx_data[2] ), .C(\rx_data[0] ), 
         .Z(n4)) /* synthesis lut_function=(!(A ((C)+!B))) */ ;
    defparam i1_3_lut_4_lut_3_lut.init = 16'h5d5d;
    LUT4 i1_3_lut_rep_789 (.A(\rx_data[1] ), .B(\rx_data[2] ), .C(\rx_data[0] ), 
         .Z(n29449)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_3_lut_rep_789.init = 16'h1010;
    LUT4 n31063_bdd_4_lut (.A(n31063), .B(\rx_data[3] ), .C(n31065), .D(\rx_data[5] ), 
         .Z(n32017)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A ((D)+!C))) */ ;
    defparam n31063_bdd_4_lut.init = 16'h22f0;
    LUT4 i1_4_lut (.A(n21770), .B(\rx_data[6] ), .C(n22272), .D(n55), 
         .Z(o_dh_bits_4__N_363[0])) /* synthesis lut_function=((B (C+(D))+!B (C))+!A) */ ;
    defparam i1_4_lut.init = 16'hfdf5;
    LUT4 i1_4_lut_adj_197 (.A(n32017), .B(\rx_data[6] ), .C(n50), .D(n29094), 
         .Z(n22272)) /* synthesis lut_function=(A+(B (C)+!B (C+!(D)))) */ ;
    defparam i1_4_lut_adj_197.init = 16'hfafb;
    LUT4 i1_4_lut_adj_198 (.A(\rx_data[5] ), .B(\rx_data[4] ), .C(\rx_data[3] ), 
         .D(\rx_data[6] ), .Z(n22129)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(71[3:8])
    defparam i1_4_lut_adj_198.init = 16'hfff7;
    LUT4 i1_3_lut (.A(\rx_data[4] ), .B(\rx_data[3] ), .C(n47), .Z(n55)) /* synthesis lut_function=(A (B+!(C))+!A (B)) */ ;
    defparam i1_3_lut.init = 16'hcece;
    LUT4 i1_4_lut_adj_199 (.A(\rx_data[5] ), .B(\rx_data[2] ), .C(\rx_data[1] ), 
         .D(\rx_data[0] ), .Z(n47)) /* synthesis lut_function=(!(A+!(B (C (D)+!C !(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(65[3] 99[10])
    defparam i1_4_lut_adj_199.init = 16'h5014;
    LUT4 i_stb_I_0_58_4_lut (.A(rx_stb), .B(n22790), .C(n29411), .D(n22312), 
         .Z(o_dh_stb_N_390)) /* synthesis lut_function=(!((B (C (D)))+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(58[15:46])
    defparam i_stb_I_0_58_4_lut.init = 16'h2aaa;
    LUT4 i1_3_lut_adj_200 (.A(\rx_data[2] ), .B(\rx_data[3] ), .C(\rx_data[6] ), 
         .Z(n22790)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut_adj_200.init = 16'h8080;
    FD1S3AX o_dh_bits_i4 (.D(o_dh_bits_4__N_363[4]), .CK(dac_clk_p_c), .Q(dec_bits[4])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=11, LSE_RCOL=30, LSE_LLINE=93, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(60[9] 100[5])
    defparam o_dh_bits_i4.GSR = "DISABLED";
    LUT4 i1_2_lut (.A(\rx_data[0] ), .B(\rx_data[1] ), .Z(n22312)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i1_3_lut_adj_201 (.A(\rx_data[0] ), .B(\rx_data[2] ), .C(\rx_data[1] ), 
         .Z(n9)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(54[23:45])
    defparam i1_3_lut_adj_201.init = 16'hfbfb;
    FD1S3AX o_dh_bits_i3 (.D(o_dh_bits_4__N_363[3]), .CK(dac_clk_p_c), .Q(dec_bits_c[3])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=11, LSE_RCOL=30, LSE_LLINE=93, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(60[9] 100[5])
    defparam o_dh_bits_i3.GSR = "DISABLED";
    FD1S3AX o_dh_bits_i2 (.D(o_dh_bits_4__N_363[2]), .CK(dac_clk_p_c), .Q(dec_bits_c[2])) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=11, LSE_RCOL=30, LSE_LLINE=93, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(60[9] 100[5])
    defparam o_dh_bits_i2.GSR = "DISABLED";
    FD1S3AX o_dh_bits_i1 (.D(o_dh_bits_4__N_363[1]), .CK(dac_clk_p_c), .Q(\dec_bits[1] )) /* synthesis LSE_LINE_FILE_ID=9, LSE_LCOL=11, LSE_RCOL=30, LSE_LLINE=93, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(60[9] 100[5])
    defparam o_dh_bits_i1.GSR = "DISABLED";
    LUT4 rx_data_0__bdd_4_lut_26297 (.A(\rx_data[0] ), .B(\rx_data[2] ), 
         .C(\rx_data[1] ), .D(\rx_data[4] ), .Z(n27668)) /* synthesis lut_function=(!(A (B+!(C (D)+!C !(D)))+!A ((C+!(D))+!B))) */ ;
    defparam rx_data_0__bdd_4_lut_26297.init = 16'h2402;
    LUT4 rx_data_0__bdd_3_lut_25908 (.A(\rx_data[0] ), .B(\rx_data[1] ), 
         .C(\rx_data[4] ), .Z(n27667)) /* synthesis lut_function=(!(A (B+(C))+!A ((C)+!B))) */ ;
    defparam rx_data_0__bdd_3_lut_25908.init = 16'h0606;
    LUT4 rx_data_0__bdd_3_lut_26296 (.A(\rx_data[1] ), .B(\rx_data[5] ), 
         .C(\rx_data[4] ), .Z(n27670)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam rx_data_0__bdd_3_lut_26296.init = 16'h8080;
    LUT4 n27670_bdd_3_lut (.A(n27670), .B(n27669), .C(\rx_data[6] ), .Z(n27671)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n27670_bdd_3_lut.init = 16'hcaca;
    LUT4 n19_bdd_4_lut (.A(n19), .B(\rx_data[2] ), .C(\rx_data[1] ), .D(\rx_data[0] ), 
         .Z(n27699)) /* synthesis lut_function=(!((B (C (D))+!B !(C+(D)))+!A)) */ ;
    defparam n19_bdd_4_lut.init = 16'h2aa8;
    LUT4 i1_2_lut_4_lut (.A(\rx_data[1] ), .B(\rx_data[2] ), .C(\rx_data[0] ), 
         .D(\rx_data[4] ), .Z(n22344)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C+(D)))) */ ;
    defparam i1_2_lut_4_lut.init = 16'hff10;
    LUT4 n506_bdd_2_lut_25921_3_lut (.A(n27671), .B(\rx_data[3] ), .C(n41), 
         .Z(o_dh_bits_4__N_363[1])) /* synthesis lut_function=(!(A (B (C))+!A (C))) */ ;
    defparam n506_bdd_2_lut_25921_3_lut.init = 16'h2f2f;
    LUT4 rx_data_0__bdd_4_lut_28621 (.A(\rx_data[0] ), .B(\rx_data[1] ), 
         .C(\rx_data[4] ), .D(\rx_data[6] ), .Z(n31062)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A ((C+!(D))+!B))) */ ;
    defparam rx_data_0__bdd_4_lut_28621.init = 16'h0480;
    LUT4 rx_data_0__bdd_3_lut_28215 (.A(\rx_data[0] ), .B(\rx_data[4] ), 
         .C(\rx_data[6] ), .Z(n31061)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B+!(C)))) */ ;
    defparam rx_data_0__bdd_3_lut_28215.init = 16'h1818;
    LUT4 rx_data_0__bdd_3_lut_28620 (.A(\rx_data[0] ), .B(\rx_data[1] ), 
         .C(\rx_data[4] ), .Z(n31065)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam rx_data_0__bdd_3_lut_28620.init = 16'h8080;
    FD1S3AY o_reset_34_rep_857 (.D(o_reset_N_392), .CK(dac_clk_p_c), .Q(n32125)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=9, LSE_LCOL=11, LSE_RCOL=30, LSE_LLINE=93, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(53[9] 54[46])
    defparam o_reset_34_rep_857.GSR = "DISABLED";
    LUT4 i1_4_lut_4_lut_rep_856 (.A(\rx_data[5] ), .B(\rx_data[2] ), .C(\rx_data[1] ), 
         .D(\rx_data[0] ), .Z(n32057)) /* synthesis lut_function=(!((B (C (D))+!B !(C+(D)))+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(65[3] 99[10])
    defparam i1_4_lut_4_lut_rep_856.init = 16'h2aa8;
    LUT4 i1_2_lut_rep_433_4_lut_4_lut (.A(\rx_data[5] ), .B(\rx_data[2] ), 
         .C(\rx_data[1] ), .D(\rx_data[0] ), .Z(n29093)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C+(D)))+!A (B+(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(65[3] 99[10])
    defparam i1_2_lut_rep_433_4_lut_4_lut.init = 16'h2ba8;
    LUT4 i1_4_lut_4_lut_then_4_lut (.A(n29410), .B(\rx_data[0] ), .C(\rx_data[1] ), 
         .D(\rx_data[2] ), .Z(n29543)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(71[3:8])
    defparam i1_4_lut_4_lut_then_4_lut.init = 16'hfeff;
    LUT4 i1_4_lut_4_lut_else_4_lut (.A(n29410), .B(\rx_data[0] ), .C(\rx_data[1] ), 
         .D(\rx_data[2] ), .Z(n29542)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(71[3:8])
    defparam i1_4_lut_4_lut_else_4_lut.init = 16'hfffb;
    LUT4 i_stb_I_0_2_lut_3_lut_4_lut (.A(n29410), .B(\rx_data[4] ), .C(rx_stb), 
         .D(n9), .Z(o_reset_N_392)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(71[3:8])
    defparam i_stb_I_0_2_lut_3_lut_4_lut.init = 16'h0040;
    LUT4 i1_3_lut_4_lut (.A(\rx_data[0] ), .B(n29450), .C(\rx_data[3] ), 
         .D(n22129), .Z(n50)) /* synthesis lut_function=(!((B+!(C+!(D)))+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(69[3:8])
    defparam i1_3_lut_4_lut.init = 16'h2022;
    LUT4 i24717_4_lut (.A(n29187), .B(n41), .C(n29544), .D(n4), .Z(o_dh_bits_4__N_363[4])) /* synthesis lut_function=(!(A (B (C))+!A (B (C (D))))) */ ;
    defparam i24717_4_lut.init = 16'h3f7f;
    LUT4 i1_4_lut_adj_202 (.A(n22344), .B(n49), .C(n22280), .D(n32057), 
         .Z(o_dh_bits_4__N_363[3])) /* synthesis lut_function=(A (B+(C))+!A (B+(C+!(D)))) */ ;
    defparam i1_4_lut_adj_202.init = 16'hfcfd;
    LUT4 i53_4_lut (.A(n29411), .B(n55), .C(\rx_data[6] ), .D(n29191), 
         .Z(n49)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B+!(C))) */ ;
    defparam i53_4_lut.init = 16'hc5cf;
    LUT4 i1_4_lut_adj_203 (.A(n27699), .B(\rx_data[1] ), .C(\rx_data[2] ), 
         .D(\rx_data[3] ), .Z(n22280)) /* synthesis lut_function=(A+!(B+(C+!(D)))) */ ;
    defparam i1_4_lut_adj_203.init = 16'habaa;
    LUT4 i1_4_lut_adj_204 (.A(n22278), .B(n21770), .C(n19), .D(n42), 
         .Z(o_dh_bits_4__N_363[2])) /* synthesis lut_function=(A+((C (D))+!B)) */ ;
    defparam i1_4_lut_adj_204.init = 16'hfbbb;
    LUT4 i1_4_lut_adj_205 (.A(n62), .B(\rx_data[2] ), .C(n22129), .D(n34), 
         .Z(n22278)) /* synthesis lut_function=(A+(B ((D)+!C))) */ ;
    defparam i1_4_lut_adj_205.init = 16'heeae;
    LUT4 i1_4_lut_adj_206 (.A(\rx_data[1] ), .B(n29303), .C(n19), .D(\rx_data[0] ), 
         .Z(n34)) /* synthesis lut_function=(!(A+!(B (C+!(D))+!B (C)))) */ ;
    defparam i1_4_lut_adj_206.init = 16'h5054;
    LUT4 i1_2_lut_rep_790 (.A(\rx_data[2] ), .B(\rx_data[1] ), .Z(n29450)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(65[3] 99[10])
    defparam i1_2_lut_rep_790.init = 16'heeee;
    LUT4 i19378_2_lut_rep_434_3_lut_4_lut (.A(\rx_data[2] ), .B(\rx_data[1] ), 
         .C(\rx_data[5] ), .D(\rx_data[3] ), .Z(n29094)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(65[3] 99[10])
    defparam i19378_2_lut_rep_434_3_lut_4_lut.init = 16'h10f0;
    LUT4 i19425_3_lut_4_lut (.A(n29449), .B(n32057), .C(\rx_data[6] ), 
         .D(\rx_data[4] ), .Z(n21770)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(65[3] 99[10])
    defparam i19425_3_lut_4_lut.init = 16'hffe0;
    LUT4 i64_3_lut_4_lut (.A(\rx_data[5] ), .B(n29191), .C(\rx_data[6] ), 
         .D(n55), .Z(n62)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C)) */ ;
    defparam i64_3_lut_4_lut.init = 16'hf707;
    LUT4 i66_3_lut_3_lut (.A(\rx_data[2] ), .B(\rx_data[1] ), .C(\rx_data[0] ), 
         .Z(n42)) /* synthesis lut_function=(!(A (C)+!A !(B (C)))) */ ;
    defparam i66_3_lut_3_lut.init = 16'h4a4a;
    LUT4 i1_2_lut_rep_643 (.A(\rx_data[4] ), .B(\rx_data[5] ), .Z(n29303)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i1_2_lut_rep_643.init = 16'h2222;
    LUT4 i1_3_lut_4_lut_adj_207 (.A(\rx_data[4] ), .B(\rx_data[5] ), .C(\rx_data[6] ), 
         .D(\rx_data[3] ), .Z(n19)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(71[3:8])
    defparam i1_3_lut_4_lut_adj_207.init = 16'h0040;
    LUT4 i24595_2_lut_rep_531_3_lut (.A(\rx_data[2] ), .B(\rx_data[1] ), 
         .C(\rx_data[3] ), .Z(n29191)) /* synthesis lut_function=(!(A (C)+!A (B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(65[3] 99[10])
    defparam i24595_2_lut_rep_531_3_lut.init = 16'h1f1f;
    LUT4 i1_2_lut_rep_791 (.A(n32125), .B(dec_stb), .Z(dac_clk_p_c_enable_548)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(53[9] 54[46])
    defparam i1_2_lut_rep_791.init = 16'heeee;
    LUT4 i8004_2_lut_3_lut (.A(n32125), .B(dec_stb), .C(dec_bits[4]), 
         .Z(dac_clk_p_c_enable_517)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(53[9] 54[46])
    defparam i8004_2_lut_3_lut.init = 16'he0e0;
    LUT4 i1_2_lut_adj_208 (.A(dec_bits[4]), .B(dec_bits_c[3]), .Z(n45)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(60[9] 100[5])
    defparam i1_2_lut_adj_208.init = 16'h4444;
    LUT4 i1_2_lut_adj_209 (.A(dec_bits[4]), .B(dec_bits_c[2]), .Z(n46)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(60[9] 100[5])
    defparam i1_2_lut_adj_209.init = 16'h4444;
    LUT4 i1_4_lut_4_lut (.A(\rx_data[3] ), .B(\rx_data[4] ), .C(n47), 
         .D(n29093), .Z(n53)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(65[3] 99[10])
    defparam i1_4_lut_4_lut.init = 16'h5140;
    PFUMX i27113 (.BLUT(n29542), .ALUT(n29543), .C0(\rx_data[4] ), .Z(n29544));
    LUT4 i1_2_lut_3_lut (.A(dec_stb), .B(dec_bits[4]), .C(n32125), .Z(dac_clk_p_c_enable_166)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(60[9] 100[5])
    defparam i1_2_lut_3_lut.init = 16'hf8f8;
    PFUMX i83 (.BLUT(n21615), .ALUT(n53), .C0(\rx_data[6] ), .Z(n41));
    LUT4 i2_3_lut_4_lut (.A(dec_stb), .B(dec_bits[4]), .C(dec_bits_c[2]), 
         .D(dec_bits_c[3]), .Z(cmd_loaded_N_535)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(60[9] 100[5])
    defparam i2_3_lut_4_lut.init = 16'h0008;
    LUT4 i1_2_lut_3_lut_adj_210 (.A(dec_stb), .B(dec_bits[4]), .C(cmd_loaded), 
         .Z(o_pck_stb_N_532)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(60[9] 100[5])
    defparam i1_2_lut_3_lut_adj_210.init = 16'h8080;
    PFUMX i28213 (.BLUT(n31062), .ALUT(n31061), .C0(\rx_data[2] ), .Z(n31063));
    PFUMX i25906 (.BLUT(n27668), .ALUT(n27667), .C0(\rx_data[5] ), .Z(n27669));
    LUT4 i1_3_lut_rep_750 (.A(\rx_data[6] ), .B(\rx_data[3] ), .C(\rx_data[5] ), 
         .Z(n29410)) /* synthesis lut_function=((B+(C))+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(71[3:8])
    defparam i1_3_lut_rep_750.init = 16'hfdfd;
    LUT4 i1_2_lut_rep_527_4_lut (.A(\rx_data[6] ), .B(\rx_data[3] ), .C(\rx_data[5] ), 
         .D(\rx_data[4] ), .Z(n29187)) /* synthesis lut_function=((B+(C+!(D)))+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(71[3:8])
    defparam i1_2_lut_rep_527_4_lut.init = 16'hfdff;
    LUT4 i1_2_lut_rep_751 (.A(\rx_data[4] ), .B(\rx_data[5] ), .Z(n29411)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(65[3] 99[10])
    defparam i1_2_lut_rep_751.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_4_lut (.A(\rx_data[4] ), .B(\rx_data[5] ), .C(n29450), 
         .D(\rx_data[3] ), .Z(n21615)) /* synthesis lut_function=(!(((C (D))+!B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(65[3] 99[10])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0888;
    
endmodule
//
// Verilog Description of module hbnewline
//

module hbnewline (\tx_data[1] , dac_clk_p_c, w_reset, \tx_data[2] , 
            \tx_data[3] , \tx_data[4] , \tx_data[5] , \tx_data[6] , 
            n32126, tx_stb, \tx_data[0] , \w_gx_char[2] , \w_gx_char[3] , 
            \w_gx_char[0] , \w_gx_char[4] , \w_gx_char[1] , \w_gx_char[5] , 
            \w_gx_char[6] , tx_busy, nl_busy, hx_stb, n32125) /* synthesis syn_module_defined=1 */ ;
    output \tx_data[1] ;
    input dac_clk_p_c;
    input w_reset;
    output \tx_data[2] ;
    output \tx_data[3] ;
    output \tx_data[4] ;
    output \tx_data[5] ;
    output \tx_data[6] ;
    input n32126;
    output tx_stb;
    output \tx_data[0] ;
    input \w_gx_char[2] ;
    input \w_gx_char[3] ;
    input \w_gx_char[0] ;
    input \w_gx_char[4] ;
    input \w_gx_char[1] ;
    input \w_gx_char[5] ;
    input \w_gx_char[6] ;
    input tx_busy;
    output nl_busy;
    input hx_stb;
    input n32125;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[29:38])
    
    wire dac_clk_p_c_enable_600;
    wire [6:0]o_nl_byte_6__N_1069;
    wire [6:0]o_nl_byte_6__N_1062;
    
    wire last_cr, last_cr_N_1090, loaded, loaded_N_1101, o_nl_stb_N_1082, 
        cr_state;
    wire [6:0]n32;
    
    wire n22338, n13159, n29399, cr_state_N_1098, n29564, n29563, 
        n28950, n28949;
    
    FD1P3JX o_nl_byte_i2 (.D(o_nl_byte_6__N_1069[1]), .SP(dac_clk_p_c_enable_600), 
            .PD(w_reset), .CK(dac_clk_p_c), .Q(\tx_data[1] )) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=9, LSE_LCOL=12, LSE_RCOL=40, LSE_LLINE=138, LSE_RLINE=139 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam o_nl_byte_i2.GSR = "DISABLED";
    FD1P3JX o_nl_byte_i3 (.D(o_nl_byte_6__N_1069[2]), .SP(dac_clk_p_c_enable_600), 
            .PD(w_reset), .CK(dac_clk_p_c), .Q(\tx_data[2] )) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=9, LSE_LCOL=12, LSE_RCOL=40, LSE_LLINE=138, LSE_RLINE=139 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam o_nl_byte_i3.GSR = "DISABLED";
    FD1P3AY o_nl_byte_i4 (.D(o_nl_byte_6__N_1062[3]), .SP(dac_clk_p_c_enable_600), 
            .CK(dac_clk_p_c), .Q(\tx_data[3] )) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=9, LSE_LCOL=12, LSE_RCOL=40, LSE_LLINE=138, LSE_RLINE=139 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam o_nl_byte_i4.GSR = "DISABLED";
    FD1P3JX o_nl_byte_i5 (.D(o_nl_byte_6__N_1069[4]), .SP(dac_clk_p_c_enable_600), 
            .PD(w_reset), .CK(dac_clk_p_c), .Q(\tx_data[4] )) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=9, LSE_LCOL=12, LSE_RCOL=40, LSE_LLINE=138, LSE_RLINE=139 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam o_nl_byte_i5.GSR = "DISABLED";
    FD1P3JX o_nl_byte_i6 (.D(o_nl_byte_6__N_1069[5]), .SP(dac_clk_p_c_enable_600), 
            .PD(w_reset), .CK(dac_clk_p_c), .Q(\tx_data[5] )) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=9, LSE_LCOL=12, LSE_RCOL=40, LSE_LLINE=138, LSE_RLINE=139 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam o_nl_byte_i6.GSR = "DISABLED";
    FD1P3JX o_nl_byte_i7 (.D(o_nl_byte_6__N_1069[6]), .SP(dac_clk_p_c_enable_600), 
            .PD(w_reset), .CK(dac_clk_p_c), .Q(\tx_data[6] )) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=9, LSE_LCOL=12, LSE_RCOL=40, LSE_LLINE=138, LSE_RLINE=139 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam o_nl_byte_i7.GSR = "DISABLED";
    FD1S3JX last_cr_45 (.D(last_cr_N_1090), .CK(dac_clk_p_c), .PD(n32126), 
            .Q(last_cr)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=9, LSE_LCOL=12, LSE_RCOL=40, LSE_LLINE=138, LSE_RLINE=139 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam last_cr_45.GSR = "DISABLED";
    FD1P3IX loaded_47 (.D(loaded_N_1101), .SP(dac_clk_p_c_enable_600), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(loaded)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=12, LSE_RCOL=40, LSE_LLINE=138, LSE_RLINE=139 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam loaded_47.GSR = "DISABLED";
    FD1S3IX o_nl_stb_46 (.D(o_nl_stb_N_1082), .CK(dac_clk_p_c), .CD(n32126), 
            .Q(tx_stb)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=12, LSE_RCOL=40, LSE_LLINE=138, LSE_RLINE=139 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam o_nl_stb_46.GSR = "DISABLED";
    FD1P3JX o_nl_byte_i1 (.D(o_nl_byte_6__N_1069[0]), .SP(dac_clk_p_c_enable_600), 
            .PD(n32126), .CK(dac_clk_p_c), .Q(\tx_data[0] )) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=9, LSE_LCOL=12, LSE_RCOL=40, LSE_LLINE=138, LSE_RLINE=139 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam o_nl_byte_i1.GSR = "DISABLED";
    LUT4 i12488_2_lut (.A(cr_state), .B(last_cr), .Z(n32[5])) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(108[13] 119[7])
    defparam i12488_2_lut.init = 16'h4444;
    LUT4 i1_4_lut (.A(\w_gx_char[2] ), .B(\w_gx_char[3] ), .C(\w_gx_char[0] ), 
         .D(n22338), .Z(n13159)) /* synthesis lut_function=((((D)+!C)+!B)+!A) */ ;
    defparam i1_4_lut.init = 16'hff7f;
    LUT4 i1_4_lut_adj_195 (.A(\w_gx_char[4] ), .B(\w_gx_char[1] ), .C(\w_gx_char[5] ), 
         .D(\w_gx_char[6] ), .Z(n22338)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_195.init = 16'hfffe;
    LUT4 i22_4_lut (.A(cr_state), .B(tx_stb), .C(tx_busy), .D(loaded), 
         .Z(nl_busy)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(90[16:37])
    defparam i22_4_lut.init = 16'hca0a;
    LUT4 mux_24_i2_3_lut_4_lut (.A(hx_stb), .B(nl_busy), .C(\w_gx_char[1] ), 
         .D(last_cr), .Z(o_nl_byte_6__N_1069[1])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(90[16:37])
    defparam mux_24_i2_3_lut_4_lut.init = 16'hfd20;
    LUT4 i1_3_lut_4_lut (.A(hx_stb), .B(nl_busy), .C(n32125), .D(tx_busy), 
         .Z(dac_clk_p_c_enable_600)) /* synthesis lut_function=(A ((C+!(D))+!B)+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(90[16:37])
    defparam i1_3_lut_4_lut.init = 16'hf2ff;
    LUT4 mux_24_i3_3_lut_4_lut (.A(hx_stb), .B(nl_busy), .C(\w_gx_char[2] ), 
         .D(n29399), .Z(o_nl_byte_6__N_1069[2])) /* synthesis lut_function=(!(A (B (D)+!B !(C))+!A (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(90[16:37])
    defparam mux_24_i3_3_lut_4_lut.init = 16'h20fd;
    LUT4 i1_3_lut_4_lut_adj_196 (.A(hx_stb), .B(nl_busy), .C(n32125), 
         .D(\w_gx_char[3] ), .Z(o_nl_byte_6__N_1062[3])) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(90[16:37])
    defparam i1_3_lut_4_lut_adj_196.init = 16'hfffd;
    LUT4 mux_24_i5_3_lut_4_lut (.A(hx_stb), .B(nl_busy), .C(\w_gx_char[4] ), 
         .D(n32[5]), .Z(o_nl_byte_6__N_1069[4])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(90[16:37])
    defparam mux_24_i5_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_24_i6_3_lut_4_lut (.A(hx_stb), .B(nl_busy), .C(\w_gx_char[5] ), 
         .D(n32[5]), .Z(o_nl_byte_6__N_1069[5])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(90[16:37])
    defparam mux_24_i6_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_24_i7_3_lut_4_lut (.A(hx_stb), .B(nl_busy), .C(\w_gx_char[6] ), 
         .D(n32[5]), .Z(o_nl_byte_6__N_1069[6])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(90[16:37])
    defparam mux_24_i7_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_24_i1_3_lut_4_lut (.A(hx_stb), .B(nl_busy), .C(\w_gx_char[0] ), 
         .D(n29399), .Z(o_nl_byte_6__N_1069[0])) /* synthesis lut_function=(!(A (B (D)+!B !(C))+!A (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(90[16:37])
    defparam mux_24_i1_3_lut_4_lut.init = 16'h20fd;
    LUT4 cr_state_I_40_3_lut_4_lut (.A(hx_stb), .B(nl_busy), .C(n13159), 
         .D(last_cr), .Z(cr_state_N_1098)) /* synthesis lut_function=(!(A (B (D)+!B (C))+!A (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(90[16:37])
    defparam cr_state_I_40_3_lut_4_lut.init = 16'h02df;
    LUT4 last_cr_I_38_4_lut_then_4_lut (.A(n13159), .B(nl_busy), .C(last_cr), 
         .D(hx_stb), .Z(n29564)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (B (C)+!B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(97[12] 120[6])
    defparam last_cr_I_38_4_lut_then_4_lut.init = 16'hd1f0;
    LUT4 last_cr_I_38_4_lut_else_4_lut (.A(n13159), .B(nl_busy), .C(last_cr), 
         .D(hx_stb), .Z(n29563)) /* synthesis lut_function=(A (B (C+!(D))+!B !(D))+!A ((C+!(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(97[12] 120[6])
    defparam last_cr_I_38_4_lut_else_4_lut.init = 16'hd1ff;
    PFUMX i27004 (.BLUT(n28950), .ALUT(n28949), .C0(tx_busy), .Z(o_nl_stb_N_1082));
    LUT4 last_cr_bdd_3_lut (.A(last_cr), .B(hx_stb), .C(cr_state), .Z(n28950)) /* synthesis lut_function=(A (B+(C))+!A !(B (C))) */ ;
    defparam last_cr_bdd_3_lut.init = 16'hbdbd;
    LUT4 last_cr_bdd_2_lut (.A(hx_stb), .B(tx_stb), .Z(n28949)) /* synthesis lut_function=(A+(B)) */ ;
    defparam last_cr_bdd_2_lut.init = 16'heeee;
    PFUMX i27127 (.BLUT(n29563), .ALUT(n29564), .C0(tx_busy), .Z(last_cr_N_1090));
    FD1P3IX cr_state_44 (.D(cr_state_N_1098), .SP(dac_clk_p_c_enable_600), 
            .CD(n32126), .CK(dac_clk_p_c), .Q(cr_state)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=12, LSE_RCOL=40, LSE_LLINE=138, LSE_RLINE=139 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam cr_state_44.GSR = "DISABLED";
    LUT4 i12445_2_lut_rep_739 (.A(cr_state), .B(last_cr), .Z(n29399)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(108[13] 119[7])
    defparam i12445_2_lut_rep_739.init = 16'h8888;
    LUT4 i12446_2_lut_3_lut_4_lut (.A(cr_state), .B(last_cr), .C(nl_busy), 
         .D(hx_stb), .Z(loaded_N_1101)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A !(C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(108[13] 119[7])
    defparam i12446_2_lut_3_lut_4_lut.init = 16'h8f88;
    
endmodule
//
// Verilog Description of module hbints
//

module hbints (int_stb, dac_clk_p_c, n32126, n32125, n29458, int_word, 
            ow_word, ow_stb) /* synthesis syn_module_defined=1 */ ;
    output int_stb;
    input dac_clk_p_c;
    input n32126;
    input n32125;
    input n29458;
    output [33:0]int_word;
    input [33:0]ow_word;
    input ow_stb;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[29:38])
    
    wire dac_clk_p_c_enable_174, n29327, loaded, dac_clk_p_c_enable_179, 
        dac_clk_p_c_enable_644, n14152;
    
    FD1P3IX o_int_stb_58 (.D(n29327), .SP(dac_clk_p_c_enable_174), .CD(n32126), 
            .CK(dac_clk_p_c), .Q(int_stb)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(90[9] 98[22])
    defparam o_int_stb_58.GSR = "DISABLED";
    FD1P3IX loaded_57 (.D(n29327), .SP(dac_clk_p_c_enable_179), .CD(n32126), 
            .CK(dac_clk_p_c), .Q(loaded)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(81[9] 87[19])
    defparam loaded_57.GSR = "DISABLED";
    LUT4 i1_3_lut_4_lut (.A(n32125), .B(n29327), .C(loaded), .D(n29458), 
         .Z(dac_clk_p_c_enable_174)) /* synthesis lut_function=(A+(B+!(C (D)))) */ ;
    defparam i1_3_lut_4_lut.init = 16'hefff;
    FD1P3JX o_int_word_i33 (.D(ow_word[33]), .SP(dac_clk_p_c_enable_644), 
            .PD(n14152), .CK(dac_clk_p_c), .Q(int_word[33])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i33.GSR = "DISABLED";
    LUT4 i1_2_lut_3_lut_4_lut (.A(int_stb), .B(n29458), .C(n29327), .D(n32125), 
         .Z(dac_clk_p_c_enable_179)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(77[12:34])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfff2;
    FD1P3JX o_int_word_i32 (.D(ow_word[32]), .SP(dac_clk_p_c_enable_644), 
            .PD(n14152), .CK(dac_clk_p_c), .Q(int_word[32])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i32.GSR = "DISABLED";
    LUT4 i_stb_I_0_3_lut_rep_667 (.A(ow_stb), .B(int_stb), .C(loaded), 
         .Z(n29327)) /* synthesis lut_function=(!((B (C))+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(93[12:34])
    defparam i_stb_I_0_3_lut_rep_667.init = 16'h2a2a;
    LUT4 i1_2_lut_3_lut_4_lut_adj_194 (.A(ow_stb), .B(int_stb), .C(loaded), 
         .D(n29458), .Z(dac_clk_p_c_enable_644)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(93[12:34])
    defparam i1_2_lut_3_lut_4_lut_adj_194.init = 16'h3bff;
    LUT4 i24583_2_lut_3_lut_4_lut (.A(ow_stb), .B(int_stb), .C(loaded), 
         .D(n29458), .Z(n14152)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A (B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(93[12:34])
    defparam i24583_2_lut_3_lut_4_lut.init = 16'h11d5;
    FD1P3IX o_int_word_i8 (.D(ow_word[8]), .SP(dac_clk_p_c_enable_644), 
            .CD(n14152), .CK(dac_clk_p_c), .Q(int_word[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i8.GSR = "DISABLED";
    FD1P3IX o_int_word_i31 (.D(ow_word[31]), .SP(dac_clk_p_c_enable_644), 
            .CD(n14152), .CK(dac_clk_p_c), .Q(int_word[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i31.GSR = "DISABLED";
    FD1P3JX o_int_word_i30 (.D(ow_word[30]), .SP(dac_clk_p_c_enable_644), 
            .PD(n14152), .CK(dac_clk_p_c), .Q(int_word[30])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i30.GSR = "DISABLED";
    FD1P3IX o_int_word_i29 (.D(ow_word[29]), .SP(dac_clk_p_c_enable_644), 
            .CD(n14152), .CK(dac_clk_p_c), .Q(int_word[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i29.GSR = "DISABLED";
    FD1P3IX o_int_word_i7 (.D(ow_word[7]), .SP(dac_clk_p_c_enable_644), 
            .CD(n14152), .CK(dac_clk_p_c), .Q(int_word[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i7.GSR = "DISABLED";
    FD1P3IX o_int_word_i28 (.D(ow_word[28]), .SP(dac_clk_p_c_enable_644), 
            .CD(n14152), .CK(dac_clk_p_c), .Q(int_word[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i28.GSR = "DISABLED";
    FD1P3IX o_int_word_i6 (.D(ow_word[6]), .SP(dac_clk_p_c_enable_644), 
            .CD(n14152), .CK(dac_clk_p_c), .Q(int_word[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i6.GSR = "DISABLED";
    FD1P3IX o_int_word_i27 (.D(ow_word[27]), .SP(dac_clk_p_c_enable_644), 
            .CD(n14152), .CK(dac_clk_p_c), .Q(int_word[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i27.GSR = "DISABLED";
    FD1P3IX o_int_word_i5 (.D(ow_word[5]), .SP(dac_clk_p_c_enable_644), 
            .CD(n14152), .CK(dac_clk_p_c), .Q(int_word[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i5.GSR = "DISABLED";
    FD1P3IX o_int_word_i26 (.D(ow_word[26]), .SP(dac_clk_p_c_enable_644), 
            .CD(n14152), .CK(dac_clk_p_c), .Q(int_word[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i26.GSR = "DISABLED";
    FD1P3IX o_int_word_i4 (.D(ow_word[4]), .SP(dac_clk_p_c_enable_644), 
            .CD(n14152), .CK(dac_clk_p_c), .Q(int_word[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i4.GSR = "DISABLED";
    FD1P3IX o_int_word_i3 (.D(ow_word[3]), .SP(dac_clk_p_c_enable_644), 
            .CD(n14152), .CK(dac_clk_p_c), .Q(int_word[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i3.GSR = "DISABLED";
    FD1P3IX o_int_word_i25 (.D(ow_word[25]), .SP(dac_clk_p_c_enable_644), 
            .CD(n14152), .CK(dac_clk_p_c), .Q(int_word[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i25.GSR = "DISABLED";
    FD1P3IX o_int_word_i24 (.D(ow_word[24]), .SP(dac_clk_p_c_enable_644), 
            .CD(n14152), .CK(dac_clk_p_c), .Q(int_word[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i24.GSR = "DISABLED";
    FD1P3IX o_int_word_i2 (.D(ow_word[2]), .SP(dac_clk_p_c_enable_644), 
            .CD(n14152), .CK(dac_clk_p_c), .Q(int_word[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i2.GSR = "DISABLED";
    FD1P3IX o_int_word_i23 (.D(ow_word[23]), .SP(dac_clk_p_c_enable_644), 
            .CD(n14152), .CK(dac_clk_p_c), .Q(int_word[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i23.GSR = "DISABLED";
    FD1P3IX o_int_word_i1 (.D(ow_word[1]), .SP(dac_clk_p_c_enable_644), 
            .CD(n14152), .CK(dac_clk_p_c), .Q(int_word[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i1.GSR = "DISABLED";
    FD1P3IX o_int_word_i0 (.D(ow_word[0]), .SP(dac_clk_p_c_enable_644), 
            .CD(n14152), .CK(dac_clk_p_c), .Q(int_word[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i0.GSR = "DISABLED";
    FD1P3IX o_int_word_i22 (.D(ow_word[22]), .SP(dac_clk_p_c_enable_644), 
            .CD(n14152), .CK(dac_clk_p_c), .Q(int_word[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i22.GSR = "DISABLED";
    FD1P3IX o_int_word_i21 (.D(ow_word[21]), .SP(dac_clk_p_c_enable_644), 
            .CD(n14152), .CK(dac_clk_p_c), .Q(int_word[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i21.GSR = "DISABLED";
    FD1P3IX o_int_word_i20 (.D(ow_word[20]), .SP(dac_clk_p_c_enable_644), 
            .CD(n14152), .CK(dac_clk_p_c), .Q(int_word[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i20.GSR = "DISABLED";
    FD1P3IX o_int_word_i19 (.D(ow_word[19]), .SP(dac_clk_p_c_enable_644), 
            .CD(n14152), .CK(dac_clk_p_c), .Q(int_word[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i19.GSR = "DISABLED";
    FD1P3IX o_int_word_i18 (.D(ow_word[18]), .SP(dac_clk_p_c_enable_644), 
            .CD(n14152), .CK(dac_clk_p_c), .Q(int_word[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i18.GSR = "DISABLED";
    FD1P3IX o_int_word_i17 (.D(ow_word[17]), .SP(dac_clk_p_c_enable_644), 
            .CD(n14152), .CK(dac_clk_p_c), .Q(int_word[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i17.GSR = "DISABLED";
    FD1P3IX o_int_word_i16 (.D(ow_word[16]), .SP(dac_clk_p_c_enable_644), 
            .CD(n14152), .CK(dac_clk_p_c), .Q(int_word[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i16.GSR = "DISABLED";
    FD1P3IX o_int_word_i15 (.D(ow_word[15]), .SP(dac_clk_p_c_enable_644), 
            .CD(n14152), .CK(dac_clk_p_c), .Q(int_word[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i15.GSR = "DISABLED";
    FD1P3IX o_int_word_i14 (.D(ow_word[14]), .SP(dac_clk_p_c_enable_644), 
            .CD(n14152), .CK(dac_clk_p_c), .Q(int_word[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i14.GSR = "DISABLED";
    FD1P3IX o_int_word_i13 (.D(ow_word[13]), .SP(dac_clk_p_c_enable_644), 
            .CD(n14152), .CK(dac_clk_p_c), .Q(int_word[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i13.GSR = "DISABLED";
    FD1P3IX o_int_word_i12 (.D(ow_word[12]), .SP(dac_clk_p_c_enable_644), 
            .CD(n14152), .CK(dac_clk_p_c), .Q(int_word[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i12.GSR = "DISABLED";
    FD1P3IX o_int_word_i9 (.D(ow_word[9]), .SP(dac_clk_p_c_enable_644), 
            .CD(n14152), .CK(dac_clk_p_c), .Q(int_word[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i9.GSR = "DISABLED";
    FD1P3IX o_int_word_i11 (.D(ow_word[11]), .SP(dac_clk_p_c_enable_644), 
            .CD(n14152), .CK(dac_clk_p_c), .Q(int_word[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i11.GSR = "DISABLED";
    FD1P3IX o_int_word_i10 (.D(ow_word[10]), .SP(dac_clk_p_c_enable_644), 
            .CD(n14152), .CK(dac_clk_p_c), .Q(int_word[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i10.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module hbidle
//

module hbidle (idl_word, dac_clk_p_c, int_word, idl_stb, hb_busy, 
            n29458, int_stb, n32126, n32125) /* synthesis syn_module_defined=1 */ ;
    output [33:0]idl_word;
    input dac_clk_p_c;
    input [33:0]int_word;
    output idl_stb;
    input hb_busy;
    output n29458;
    input int_stb;
    input n32126;
    input n32125;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[29:38])
    
    wire dac_clk_p_c_enable_646, n14199, n29203, dac_clk_p_c_enable_173;
    
    FD1P3IX o_idl_word_i10 (.D(int_word[10]), .SP(dac_clk_p_c_enable_646), 
            .CD(n14199), .CK(dac_clk_p_c), .Q(idl_word[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i10.GSR = "DISABLED";
    FD1P3IX o_idl_word_i9 (.D(int_word[9]), .SP(dac_clk_p_c_enable_646), 
            .CD(n14199), .CK(dac_clk_p_c), .Q(idl_word[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i9.GSR = "DISABLED";
    FD1P3IX o_idl_word_i8 (.D(int_word[8]), .SP(dac_clk_p_c_enable_646), 
            .CD(n14199), .CK(dac_clk_p_c), .Q(idl_word[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i8.GSR = "DISABLED";
    LUT4 o_idl_stb_I_0_30_2_lut_rep_798 (.A(idl_stb), .B(hb_busy), .Z(n29458)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(97[22:43])
    defparam o_idl_stb_I_0_30_2_lut_rep_798.init = 16'h8888;
    LUT4 o_int_stb_I_0_66_2_lut_rep_543_3_lut (.A(idl_stb), .B(hb_busy), 
         .C(int_stb), .Z(n29203)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(97[22:43])
    defparam o_int_stb_I_0_66_2_lut_rep_543_3_lut.init = 16'h7070;
    LUT4 i1_2_lut_3_lut_3_lut (.A(idl_stb), .B(hb_busy), .C(int_stb), 
         .Z(dac_clk_p_c_enable_646)) /* synthesis lut_function=(!(A (B)+!A !((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(97[22:43])
    defparam i1_2_lut_3_lut_3_lut.init = 16'h7373;
    FD1P3IX o_idl_stb_28 (.D(n29203), .SP(dac_clk_p_c_enable_173), .CD(n32126), 
            .CK(dac_clk_p_c), .Q(idl_stb)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(80[9] 88[22])
    defparam o_idl_stb_28.GSR = "DISABLED";
    LUT4 i1_3_lut_4_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(n32125), .D(int_stb), 
         .Z(dac_clk_p_c_enable_173)) /* synthesis lut_function=(A ((C)+!B)+!A ((C+(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(97[22:43])
    defparam i1_3_lut_4_lut_4_lut.init = 16'hf7f3;
    FD1P3JX o_idl_word_i33 (.D(int_word[33]), .SP(dac_clk_p_c_enable_646), 
            .PD(n14199), .CK(dac_clk_p_c), .Q(idl_word[33])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i33.GSR = "DISABLED";
    FD1P3JX o_idl_word_i32 (.D(int_word[32]), .SP(dac_clk_p_c_enable_646), 
            .PD(n14199), .CK(dac_clk_p_c), .Q(idl_word[32])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i32.GSR = "DISABLED";
    FD1P3IX o_idl_word_i7 (.D(int_word[7]), .SP(dac_clk_p_c_enable_646), 
            .CD(n14199), .CK(dac_clk_p_c), .Q(idl_word[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i7.GSR = "DISABLED";
    FD1P3IX o_idl_word_i6 (.D(int_word[6]), .SP(dac_clk_p_c_enable_646), 
            .CD(n14199), .CK(dac_clk_p_c), .Q(idl_word[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i6.GSR = "DISABLED";
    FD1P3IX o_idl_word_i5 (.D(int_word[5]), .SP(dac_clk_p_c_enable_646), 
            .CD(n14199), .CK(dac_clk_p_c), .Q(idl_word[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i5.GSR = "DISABLED";
    FD1P3IX o_idl_word_i4 (.D(int_word[4]), .SP(dac_clk_p_c_enable_646), 
            .CD(n14199), .CK(dac_clk_p_c), .Q(idl_word[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i4.GSR = "DISABLED";
    FD1P3IX o_idl_word_i3 (.D(int_word[3]), .SP(dac_clk_p_c_enable_646), 
            .CD(n14199), .CK(dac_clk_p_c), .Q(idl_word[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i3.GSR = "DISABLED";
    FD1P3IX o_idl_word_i2 (.D(int_word[2]), .SP(dac_clk_p_c_enable_646), 
            .CD(n14199), .CK(dac_clk_p_c), .Q(idl_word[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i2.GSR = "DISABLED";
    FD1P3IX o_idl_word_i1 (.D(int_word[1]), .SP(dac_clk_p_c_enable_646), 
            .CD(n14199), .CK(dac_clk_p_c), .Q(idl_word[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i1.GSR = "DISABLED";
    FD1P3IX o_idl_word_i0 (.D(int_word[0]), .SP(dac_clk_p_c_enable_646), 
            .CD(n14199), .CK(dac_clk_p_c), .Q(idl_word[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i0.GSR = "DISABLED";
    LUT4 i24671_2_lut (.A(hb_busy), .B(int_stb), .Z(n14199)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i24671_2_lut.init = 16'h1111;
    FD1P3IX o_idl_word_i31 (.D(int_word[31]), .SP(dac_clk_p_c_enable_646), 
            .CD(n14199), .CK(dac_clk_p_c), .Q(idl_word[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i31.GSR = "DISABLED";
    FD1P3JX o_idl_word_i30 (.D(int_word[30]), .SP(dac_clk_p_c_enable_646), 
            .PD(n14199), .CK(dac_clk_p_c), .Q(idl_word[30])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i30.GSR = "DISABLED";
    FD1P3JX o_idl_word_i29 (.D(int_word[29]), .SP(dac_clk_p_c_enable_646), 
            .PD(n14199), .CK(dac_clk_p_c), .Q(idl_word[29])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i29.GSR = "DISABLED";
    FD1P3IX o_idl_word_i28 (.D(int_word[28]), .SP(dac_clk_p_c_enable_646), 
            .CD(n14199), .CK(dac_clk_p_c), .Q(idl_word[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i28.GSR = "DISABLED";
    FD1P3IX o_idl_word_i27 (.D(int_word[27]), .SP(dac_clk_p_c_enable_646), 
            .CD(n14199), .CK(dac_clk_p_c), .Q(idl_word[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i27.GSR = "DISABLED";
    FD1P3IX o_idl_word_i26 (.D(int_word[26]), .SP(dac_clk_p_c_enable_646), 
            .CD(n14199), .CK(dac_clk_p_c), .Q(idl_word[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i26.GSR = "DISABLED";
    FD1P3IX o_idl_word_i25 (.D(int_word[25]), .SP(dac_clk_p_c_enable_646), 
            .CD(n14199), .CK(dac_clk_p_c), .Q(idl_word[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i25.GSR = "DISABLED";
    FD1P3IX o_idl_word_i24 (.D(int_word[24]), .SP(dac_clk_p_c_enable_646), 
            .CD(n14199), .CK(dac_clk_p_c), .Q(idl_word[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i24.GSR = "DISABLED";
    FD1P3IX o_idl_word_i23 (.D(int_word[23]), .SP(dac_clk_p_c_enable_646), 
            .CD(n14199), .CK(dac_clk_p_c), .Q(idl_word[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i23.GSR = "DISABLED";
    FD1P3IX o_idl_word_i22 (.D(int_word[22]), .SP(dac_clk_p_c_enable_646), 
            .CD(n14199), .CK(dac_clk_p_c), .Q(idl_word[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i22.GSR = "DISABLED";
    FD1P3IX o_idl_word_i21 (.D(int_word[21]), .SP(dac_clk_p_c_enable_646), 
            .CD(n14199), .CK(dac_clk_p_c), .Q(idl_word[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i21.GSR = "DISABLED";
    FD1P3IX o_idl_word_i20 (.D(int_word[20]), .SP(dac_clk_p_c_enable_646), 
            .CD(n14199), .CK(dac_clk_p_c), .Q(idl_word[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i20.GSR = "DISABLED";
    FD1P3IX o_idl_word_i19 (.D(int_word[19]), .SP(dac_clk_p_c_enable_646), 
            .CD(n14199), .CK(dac_clk_p_c), .Q(idl_word[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i19.GSR = "DISABLED";
    FD1P3IX o_idl_word_i18 (.D(int_word[18]), .SP(dac_clk_p_c_enable_646), 
            .CD(n14199), .CK(dac_clk_p_c), .Q(idl_word[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i18.GSR = "DISABLED";
    FD1P3IX o_idl_word_i17 (.D(int_word[17]), .SP(dac_clk_p_c_enable_646), 
            .CD(n14199), .CK(dac_clk_p_c), .Q(idl_word[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i17.GSR = "DISABLED";
    FD1P3IX o_idl_word_i16 (.D(int_word[16]), .SP(dac_clk_p_c_enable_646), 
            .CD(n14199), .CK(dac_clk_p_c), .Q(idl_word[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i16.GSR = "DISABLED";
    FD1P3IX o_idl_word_i15 (.D(int_word[15]), .SP(dac_clk_p_c_enable_646), 
            .CD(n14199), .CK(dac_clk_p_c), .Q(idl_word[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i15.GSR = "DISABLED";
    FD1P3IX o_idl_word_i14 (.D(int_word[14]), .SP(dac_clk_p_c_enable_646), 
            .CD(n14199), .CK(dac_clk_p_c), .Q(idl_word[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i14.GSR = "DISABLED";
    FD1P3IX o_idl_word_i13 (.D(int_word[13]), .SP(dac_clk_p_c_enable_646), 
            .CD(n14199), .CK(dac_clk_p_c), .Q(idl_word[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i13.GSR = "DISABLED";
    FD1P3IX o_idl_word_i12 (.D(int_word[12]), .SP(dac_clk_p_c_enable_646), 
            .CD(n14199), .CK(dac_clk_p_c), .Q(idl_word[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i12.GSR = "DISABLED";
    FD1P3IX o_idl_word_i11 (.D(int_word[11]), .SP(dac_clk_p_c_enable_646), 
            .CD(n14199), .CK(dac_clk_p_c), .Q(idl_word[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=9, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i11.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module TSALL
// module not written out since it is a black-box. 
//

//
// Verilog Description of module efb_inst
//

module efb_inst (dac_clk_p_c, i_sw0_c, wb_cyc, wb_lo_data_7__N_34, wb_we, 
            \wb_addr[7] , \wb_addr[6] , \wb_addr[5] , \wb_addr[4] , 
            \wb_addr[3] , \wb_addr[2] , \wb_addr[1] , \wb_addr[0] , 
            \wb_odata[7] , \wb_odata[6] , \wb_odata[5] , \wb_odata[4] , 
            \wb_odata[3] , \wb_odata[2] , \wb_odata[1] , \wb_odata[0] , 
            pll_data_o, pll_ack, wb_lo_data, wb_lo_ack, pll_clk, pll_rst, 
            pll_stb, pll_we, pll_addr, pll_data_i, GND_net, VCC_net) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;
    input dac_clk_p_c;
    input i_sw0_c;
    input wb_cyc;
    input wb_lo_data_7__N_34;
    input wb_we;
    input \wb_addr[7] ;
    input \wb_addr[6] ;
    input \wb_addr[5] ;
    input \wb_addr[4] ;
    input \wb_addr[3] ;
    input \wb_addr[2] ;
    input \wb_addr[1] ;
    input \wb_addr[0] ;
    input \wb_odata[7] ;
    input \wb_odata[6] ;
    input \wb_odata[5] ;
    input \wb_odata[4] ;
    input \wb_odata[3] ;
    input \wb_odata[2] ;
    input \wb_odata[1] ;
    input \wb_odata[0] ;
    input [7:0]pll_data_o;
    input pll_ack;
    output [7:0]wb_lo_data;
    output wb_lo_ack;
    output pll_clk;
    output pll_rst;
    output pll_stb;
    output pll_we;
    output [4:0]pll_addr;
    output [7:0]pll_data_i;
    input GND_net;
    input VCC_net;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[29:38])
    
    EFB EFBInst_0 (.WBCLKI(dac_clk_p_c), .WBRSTI(i_sw0_c), .WBCYCI(wb_cyc), 
        .WBSTBI(wb_lo_data_7__N_34), .WBWEI(wb_we), .WBADRI0(\wb_addr[0] ), 
        .WBADRI1(\wb_addr[1] ), .WBADRI2(\wb_addr[2] ), .WBADRI3(\wb_addr[3] ), 
        .WBADRI4(\wb_addr[4] ), .WBADRI5(\wb_addr[5] ), .WBADRI6(\wb_addr[6] ), 
        .WBADRI7(\wb_addr[7] ), .WBDATI0(\wb_odata[0] ), .WBDATI1(\wb_odata[1] ), 
        .WBDATI2(\wb_odata[2] ), .WBDATI3(\wb_odata[3] ), .WBDATI4(\wb_odata[4] ), 
        .WBDATI5(\wb_odata[5] ), .WBDATI6(\wb_odata[6] ), .WBDATI7(\wb_odata[7] ), 
        .I2C1SCLI(GND_net), .I2C1SDAI(GND_net), .I2C2SCLI(GND_net), .I2C2SDAI(GND_net), 
        .SPISCKI(GND_net), .SPIMISOI(GND_net), .SPIMOSII(GND_net), .SPISCSN(GND_net), 
        .TCCLKI(GND_net), .TCRSTN(GND_net), .TCIC(GND_net), .UFMSN(VCC_net), 
        .PLL0DATI0(pll_data_o[0]), .PLL0DATI1(pll_data_o[1]), .PLL0DATI2(pll_data_o[2]), 
        .PLL0DATI3(pll_data_o[3]), .PLL0DATI4(pll_data_o[4]), .PLL0DATI5(pll_data_o[5]), 
        .PLL0DATI6(pll_data_o[6]), .PLL0DATI7(pll_data_o[7]), .PLL0ACKI(pll_ack), 
        .PLL1DATI0(GND_net), .PLL1DATI1(GND_net), .PLL1DATI2(GND_net), 
        .PLL1DATI3(GND_net), .PLL1DATI4(GND_net), .PLL1DATI5(GND_net), 
        .PLL1DATI6(GND_net), .PLL1DATI7(GND_net), .PLL1ACKI(GND_net), 
        .WBDATO0(wb_lo_data[0]), .WBDATO1(wb_lo_data[1]), .WBDATO2(wb_lo_data[2]), 
        .WBDATO3(wb_lo_data[3]), .WBDATO4(wb_lo_data[4]), .WBDATO5(wb_lo_data[5]), 
        .WBDATO6(wb_lo_data[6]), .WBDATO7(wb_lo_data[7]), .WBACKO(wb_lo_ack), 
        .PLLCLKO(pll_clk), .PLLRSTO(pll_rst), .PLL0STBO(pll_stb), .PLLWEO(pll_we), 
        .PLLADRO0(pll_addr[0]), .PLLADRO1(pll_addr[1]), .PLLADRO2(pll_addr[2]), 
        .PLLADRO3(pll_addr[3]), .PLLADRO4(pll_addr[4]), .PLLDATO0(pll_data_i[0]), 
        .PLLDATO1(pll_data_i[1]), .PLLDATO2(pll_data_i[2]), .PLLDATO3(pll_data_i[3]), 
        .PLLDATO4(pll_data_i[4]), .PLLDATO5(pll_data_i[5]), .PLLDATO6(pll_data_i[6]), 
        .PLLDATO7(pll_data_i[7])) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=7, LSE_LCOL=11, LSE_RCOL=4, LSE_LLINE=183, LSE_RLINE=195 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(183[11] 195[4])
    defparam EFBInst_0.EFB_I2C1 = "DISABLED";
    defparam EFBInst_0.EFB_I2C2 = "DISABLED";
    defparam EFBInst_0.EFB_SPI = "DISABLED";
    defparam EFBInst_0.EFB_TC = "DISABLED";
    defparam EFBInst_0.EFB_TC_PORTMODE = "WB";
    defparam EFBInst_0.EFB_UFM = "DISABLED";
    defparam EFBInst_0.EFB_WB_CLK_FREQ = "50.0";
    defparam EFBInst_0.DEV_DENSITY = "6900L";
    defparam EFBInst_0.UFM_INIT_PAGES = 0;
    defparam EFBInst_0.UFM_INIT_START_PAGE = 0;
    defparam EFBInst_0.UFM_INIT_ALL_ZEROS = "ENABLED";
    defparam EFBInst_0.UFM_INIT_FILE_NAME = "NONE";
    defparam EFBInst_0.UFM_INIT_FILE_FORMAT = "HEX";
    defparam EFBInst_0.I2C1_ADDRESSING = "7BIT";
    defparam EFBInst_0.I2C2_ADDRESSING = "7BIT";
    defparam EFBInst_0.I2C1_SLAVE_ADDR = "0b1000001";
    defparam EFBInst_0.I2C2_SLAVE_ADDR = "0b1000010";
    defparam EFBInst_0.I2C1_BUS_PERF = "100kHz";
    defparam EFBInst_0.I2C2_BUS_PERF = "100kHz";
    defparam EFBInst_0.I2C1_CLK_DIVIDER = 1;
    defparam EFBInst_0.I2C2_CLK_DIVIDER = 1;
    defparam EFBInst_0.I2C1_GEN_CALL = "DISABLED";
    defparam EFBInst_0.I2C2_GEN_CALL = "DISABLED";
    defparam EFBInst_0.I2C1_WAKEUP = "DISABLED";
    defparam EFBInst_0.I2C2_WAKEUP = "DISABLED";
    defparam EFBInst_0.SPI_MODE = "MASTER";
    defparam EFBInst_0.SPI_CLK_DIVIDER = 1;
    defparam EFBInst_0.SPI_LSB_FIRST = "DISABLED";
    defparam EFBInst_0.SPI_CLK_INV = "DISABLED";
    defparam EFBInst_0.SPI_PHASE_ADJ = "DISABLED";
    defparam EFBInst_0.SPI_SLAVE_HANDSHAKE = "DISABLED";
    defparam EFBInst_0.SPI_INTR_TXRDY = "DISABLED";
    defparam EFBInst_0.SPI_INTR_RXRDY = "DISABLED";
    defparam EFBInst_0.SPI_INTR_TXOVR = "DISABLED";
    defparam EFBInst_0.SPI_INTR_RXOVR = "DISABLED";
    defparam EFBInst_0.SPI_WAKEUP = "DISABLED";
    defparam EFBInst_0.TC_MODE = "CTCM";
    defparam EFBInst_0.TC_SCLK_SEL = "PCLOCK";
    defparam EFBInst_0.TC_CCLK_SEL = 1;
    defparam EFBInst_0.GSR = "ENABLED";
    defparam EFBInst_0.TC_TOP_SET = 65535;
    defparam EFBInst_0.TC_OCR_SET = 32767;
    defparam EFBInst_0.TC_OC_MODE = "TOGGLE";
    defparam EFBInst_0.TC_RESETN = "ENABLED";
    defparam EFBInst_0.TC_TOP_SEL = "OFF";
    defparam EFBInst_0.TC_OV_INT = "OFF";
    defparam EFBInst_0.TC_OCR_INT = "OFF";
    defparam EFBInst_0.TC_ICR_INT = "OFF";
    defparam EFBInst_0.TC_OVERFLOW = "DISABLED";
    defparam EFBInst_0.TC_ICAPTURE = "DISABLED";
    
endmodule
//
// Verilog Description of module sys_clk
//

module sys_clk (i_ref_clk_c, dac_clk_p_c, GND_net) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;
    input i_ref_clk_c;
    output dac_clk_p_c;
    input GND_net;
    
    wire i_ref_clk_c /* synthesis is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(26[12:21])
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[29:38])
    
    EHXPLLJ PLLInst_0 (.CLKI(i_ref_clk_c), .CLKFB(dac_clk_p_c), .PHASESEL0(GND_net), 
            .PHASESEL1(GND_net), .PHASEDIR(GND_net), .PHASESTEP(GND_net), 
            .LOADREG(GND_net), .STDBY(GND_net), .PLLWAKESYNC(GND_net), 
            .RST(GND_net), .RESETC(GND_net), .RESETD(GND_net), .RESETM(GND_net), 
            .ENCLKOP(GND_net), .ENCLKOS(GND_net), .ENCLKOS2(GND_net), 
            .ENCLKOS3(GND_net), .PLLCLK(GND_net), .PLLRST(GND_net), .PLLSTB(GND_net), 
            .PLLWE(GND_net), .PLLDATI0(GND_net), .PLLDATI1(GND_net), .PLLDATI2(GND_net), 
            .PLLDATI3(GND_net), .PLLDATI4(GND_net), .PLLDATI5(GND_net), 
            .PLLDATI6(GND_net), .PLLDATI7(GND_net), .PLLADDR0(GND_net), 
            .PLLADDR1(GND_net), .PLLADDR2(GND_net), .PLLADDR3(GND_net), 
            .PLLADDR4(GND_net), .CLKOP(dac_clk_p_c)) /* synthesis FREQUENCY_PIN_CLKOP="72.000000", FREQUENCY_PIN_CLKI="12.000000", ICP_CURRENT="9", LPF_RESISTOR="72", syn_instantiated=1, LSE_LINE_FILE_ID=7, LSE_LCOL=10, LSE_RCOL=54, LSE_LLINE=47, LSE_RLINE=47 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(47[10:54])
    defparam PLLInst_0.CLKI_DIV = 1;
    defparam PLLInst_0.CLKFB_DIV = 6;
    defparam PLLInst_0.CLKOP_DIV = 7;
    defparam PLLInst_0.CLKOS_DIV = 1;
    defparam PLLInst_0.CLKOS2_DIV = 1;
    defparam PLLInst_0.CLKOS3_DIV = 1;
    defparam PLLInst_0.CLKOP_ENABLE = "ENABLED";
    defparam PLLInst_0.CLKOS_ENABLE = "DISABLED";
    defparam PLLInst_0.CLKOS2_ENABLE = "DISABLED";
    defparam PLLInst_0.CLKOS3_ENABLE = "DISABLED";
    defparam PLLInst_0.VCO_BYPASS_A0 = "DISABLED";
    defparam PLLInst_0.VCO_BYPASS_B0 = "DISABLED";
    defparam PLLInst_0.VCO_BYPASS_C0 = "DISABLED";
    defparam PLLInst_0.VCO_BYPASS_D0 = "DISABLED";
    defparam PLLInst_0.CLKOP_CPHASE = 6;
    defparam PLLInst_0.CLKOS_CPHASE = 0;
    defparam PLLInst_0.CLKOS2_CPHASE = 0;
    defparam PLLInst_0.CLKOS3_CPHASE = 0;
    defparam PLLInst_0.CLKOP_FPHASE = 0;
    defparam PLLInst_0.CLKOS_FPHASE = 0;
    defparam PLLInst_0.CLKOS2_FPHASE = 0;
    defparam PLLInst_0.CLKOS3_FPHASE = 0;
    defparam PLLInst_0.FEEDBK_PATH = "CLKOP";
    defparam PLLInst_0.FRACN_ENABLE = "DISABLED";
    defparam PLLInst_0.FRACN_DIV = 0;
    defparam PLLInst_0.CLKOP_TRIM_POL = "RISING";
    defparam PLLInst_0.CLKOP_TRIM_DELAY = 0;
    defparam PLLInst_0.CLKOS_TRIM_POL = "FALLING";
    defparam PLLInst_0.CLKOS_TRIM_DELAY = 0;
    defparam PLLInst_0.PLL_USE_WB = "DISABLED";
    defparam PLLInst_0.PREDIVIDER_MUXA1 = 0;
    defparam PLLInst_0.PREDIVIDER_MUXB1 = 0;
    defparam PLLInst_0.PREDIVIDER_MUXC1 = 0;
    defparam PLLInst_0.PREDIVIDER_MUXD1 = 0;
    defparam PLLInst_0.OUTDIVIDER_MUXA2 = "DIVA";
    defparam PLLInst_0.OUTDIVIDER_MUXB2 = "DIVB";
    defparam PLLInst_0.OUTDIVIDER_MUXC2 = "DIVC";
    defparam PLLInst_0.OUTDIVIDER_MUXD2 = "DIVD";
    defparam PLLInst_0.PLL_LOCK_MODE = 0;
    defparam PLLInst_0.STDBY_ENABLE = "DISABLED";
    defparam PLLInst_0.DPHASE_SOURCE = "DISABLED";
    defparam PLLInst_0.PLLRST_ENA = "DISABLED";
    defparam PLLInst_0.MRST_ENA = "DISABLED";
    defparam PLLInst_0.DCRST_ENA = "DISABLED";
    defparam PLLInst_0.DDRST_ENA = "DISABLED";
    defparam PLLInst_0.INTFB_WAKE = "DISABLED";
    
endmodule
//
// Verilog Description of module dynamic_pll
//

module dynamic_pll (i_ref_clk_c, pll_clk, pll_rst, pll_stb, pll_we, 
            pll_data_i, pll_addr, lo_q, pll_data_o, pll_ack, GND_net, 
            lo_i_en, o_lo_i_c) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;
    input i_ref_clk_c;
    input pll_clk;
    input pll_rst;
    input pll_stb;
    input pll_we;
    input [7:0]pll_data_i;
    input [4:0]pll_addr;
    output lo_q;
    output [7:0]pll_data_o;
    output pll_ack;
    input GND_net;
    input lo_i_en;
    output o_lo_i_c;
    
    wire i_ref_clk_c /* synthesis is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(26[12:21])
    wire lo_i /* synthesis is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(159[18:22])
    wire lo_q /* synthesis is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(159[24:28])
    
    EHXPLLJ PLLInst_0 (.CLKI(i_ref_clk_c), .CLKFB(lo_i), .PHASESEL0(GND_net), 
            .PHASESEL1(GND_net), .PHASEDIR(GND_net), .PHASESTEP(GND_net), 
            .LOADREG(GND_net), .STDBY(GND_net), .PLLWAKESYNC(GND_net), 
            .RST(GND_net), .RESETC(GND_net), .RESETD(GND_net), .RESETM(GND_net), 
            .ENCLKOP(GND_net), .ENCLKOS(GND_net), .ENCLKOS2(GND_net), 
            .ENCLKOS3(GND_net), .PLLCLK(pll_clk), .PLLRST(pll_rst), .PLLSTB(pll_stb), 
            .PLLWE(pll_we), .PLLDATI0(pll_data_i[0]), .PLLDATI1(pll_data_i[1]), 
            .PLLDATI2(pll_data_i[2]), .PLLDATI3(pll_data_i[3]), .PLLDATI4(pll_data_i[4]), 
            .PLLDATI5(pll_data_i[5]), .PLLDATI6(pll_data_i[6]), .PLLDATI7(pll_data_i[7]), 
            .PLLADDR0(pll_addr[0]), .PLLADDR1(pll_addr[1]), .PLLADDR2(pll_addr[2]), 
            .PLLADDR3(pll_addr[3]), .PLLADDR4(pll_addr[4]), .CLKOP(lo_i), 
            .CLKOS(lo_q), .PLLDATO0(pll_data_o[0]), .PLLDATO1(pll_data_o[1]), 
            .PLLDATO2(pll_data_o[2]), .PLLDATO3(pll_data_o[3]), .PLLDATO4(pll_data_o[4]), 
            .PLLDATO5(pll_data_o[5]), .PLLDATO6(pll_data_o[6]), .PLLDATO7(pll_data_o[7]), 
            .PLLACK(pll_ack)) /* synthesis FREQUENCY_PIN_CLKOS="48.000000", FREQUENCY_PIN_CLKOP="48.000000", FREQUENCY_PIN_CLKI="12.000000", ICP_CURRENT="8", LPF_RESISTOR="8", syn_instantiated=1, LSE_LINE_FILE_ID=7, LSE_LCOL=14, LSE_RCOL=5, LSE_LLINE=169, LSE_RLINE=181 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(169[14] 181[5])
    defparam PLLInst_0.CLKI_DIV = 1;
    defparam PLLInst_0.CLKFB_DIV = 4;
    defparam PLLInst_0.CLKOP_DIV = 11;
    defparam PLLInst_0.CLKOS_DIV = 11;
    defparam PLLInst_0.CLKOS2_DIV = 1;
    defparam PLLInst_0.CLKOS3_DIV = 1;
    defparam PLLInst_0.CLKOP_ENABLE = "ENABLED";
    defparam PLLInst_0.CLKOS_ENABLE = "ENABLED";
    defparam PLLInst_0.CLKOS2_ENABLE = "DISABLED";
    defparam PLLInst_0.CLKOS3_ENABLE = "DISABLED";
    defparam PLLInst_0.VCO_BYPASS_A0 = "DISABLED";
    defparam PLLInst_0.VCO_BYPASS_B0 = "DISABLED";
    defparam PLLInst_0.VCO_BYPASS_C0 = "DISABLED";
    defparam PLLInst_0.VCO_BYPASS_D0 = "DISABLED";
    defparam PLLInst_0.CLKOP_CPHASE = 10;
    defparam PLLInst_0.CLKOS_CPHASE = 12;
    defparam PLLInst_0.CLKOS2_CPHASE = 0;
    defparam PLLInst_0.CLKOS3_CPHASE = 0;
    defparam PLLInst_0.CLKOP_FPHASE = 0;
    defparam PLLInst_0.CLKOS_FPHASE = 6;
    defparam PLLInst_0.CLKOS2_FPHASE = 0;
    defparam PLLInst_0.CLKOS3_FPHASE = 0;
    defparam PLLInst_0.FEEDBK_PATH = "CLKOP";
    defparam PLLInst_0.FRACN_ENABLE = "DISABLED";
    defparam PLLInst_0.FRACN_DIV = 0;
    defparam PLLInst_0.CLKOP_TRIM_POL = "RISING";
    defparam PLLInst_0.CLKOP_TRIM_DELAY = 0;
    defparam PLLInst_0.CLKOS_TRIM_POL = "RISING";
    defparam PLLInst_0.CLKOS_TRIM_DELAY = 0;
    defparam PLLInst_0.PLL_USE_WB = "ENABLED";
    defparam PLLInst_0.PREDIVIDER_MUXA1 = 0;
    defparam PLLInst_0.PREDIVIDER_MUXB1 = 0;
    defparam PLLInst_0.PREDIVIDER_MUXC1 = 0;
    defparam PLLInst_0.PREDIVIDER_MUXD1 = 0;
    defparam PLLInst_0.OUTDIVIDER_MUXA2 = "DIVA";
    defparam PLLInst_0.OUTDIVIDER_MUXB2 = "DIVB";
    defparam PLLInst_0.OUTDIVIDER_MUXC2 = "DIVC";
    defparam PLLInst_0.OUTDIVIDER_MUXD2 = "DIVD";
    defparam PLLInst_0.PLL_LOCK_MODE = 0;
    defparam PLLInst_0.STDBY_ENABLE = "DISABLED";
    defparam PLLInst_0.DPHASE_SOURCE = "DISABLED";
    defparam PLLInst_0.PLLRST_ENA = "DISABLED";
    defparam PLLInst_0.MRST_ENA = "DISABLED";
    defparam PLLInst_0.DCRST_ENA = "DISABLED";
    defparam PLLInst_0.DDRST_ENA = "DISABLED";
    defparam PLLInst_0.INTFB_WAKE = "DISABLED";
    LUT4 i1_2_lut (.A(lo_i), .B(lo_i_en), .Z(o_lo_i_c)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(169[14] 181[5])
    defparam i1_2_lut.init = 16'h8888;
    
endmodule
//
// Verilog Description of module fm_generator_wb_slave
//

module fm_generator_wb_slave (o_dac_b_c_0, dac_clk_p_c, wb_fm_data, i_sw0_c, 
            o_dac_a_c_0, GND_net, \wb_addr[0] , n29300, \wb_addr[2] , 
            \wb_addr[1] , wb_fm_ack, o_dac_a_9__N_1, dac_clk_p_c_enable_502, 
            wb_odata, n21641, n29065, n22458, dac_clk_p_c_enable_227, 
            o_dac_a_c_9, dac_clk_p_c_enable_241, dac_clk_p_c_enable_106, 
            o_dac_a_c_8, o_dac_a_c_7, o_dac_a_c_6, o_dac_a_c_5, o_dac_a_c_4, 
            o_dac_a_c_3, o_dac_a_c_2, o_dac_a_c_1, o_dac_b_c_9, o_dac_b_c_8, 
            o_dac_b_c_7, o_dac_b_c_6, o_dac_b_c_5, o_dac_b_c_4, o_dac_b_c_3, 
            o_dac_b_c_2, o_dac_b_c_1, dac_clk_p_c_enable_375, dac_clk_p_c_enable_407, 
            dac_clk_p_c_enable_439, dac_clk_p_c_enable_471, n21662, n29155, 
            n29197, n29199, o_dac_cw_b_c, n32067, n32066) /* synthesis syn_module_defined=1 */ ;
    output o_dac_b_c_0;
    input dac_clk_p_c;
    output [31:0]wb_fm_data;
    input i_sw0_c;
    output o_dac_a_c_0;
    input GND_net;
    input \wb_addr[0] ;
    output n29300;
    input \wb_addr[2] ;
    input \wb_addr[1] ;
    output wb_fm_ack;
    input o_dac_a_9__N_1;
    input dac_clk_p_c_enable_502;
    input [31:0]wb_odata;
    output n21641;
    input n29065;
    input n22458;
    output dac_clk_p_c_enable_227;
    output o_dac_a_c_9;
    output dac_clk_p_c_enable_241;
    output dac_clk_p_c_enable_106;
    output o_dac_a_c_8;
    output o_dac_a_c_7;
    output o_dac_a_c_6;
    output o_dac_a_c_5;
    output o_dac_a_c_4;
    output o_dac_a_c_3;
    output o_dac_a_c_2;
    output o_dac_a_c_1;
    output o_dac_b_c_9;
    output o_dac_b_c_8;
    output o_dac_b_c_7;
    output o_dac_b_c_6;
    output o_dac_b_c_5;
    output o_dac_b_c_4;
    output o_dac_b_c_3;
    output o_dac_b_c_2;
    output o_dac_b_c_1;
    input dac_clk_p_c_enable_375;
    input dac_clk_p_c_enable_407;
    input dac_clk_p_c_enable_439;
    input dac_clk_p_c_enable_471;
    output n21662;
    output n29155;
    output n29197;
    output n29199;
    output o_dac_cw_b_c;
    input n32067;
    input n32066;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[29:38])
    wire [15:0]o_sample_q /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(30[51:61])
    wire [15:0]modulation_output /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(86[39:56])
    wire [15:0]o_sample_i /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(30[39:49])
    wire [9:0]o_dac_b;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[40:47])
    wire [31:0]o_wb_data_31__N_1104;
    wire [30:0]carrier_increment;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(77[31:48])
    wire [30:0]carrier_increment_30__N_1296;
    
    wire cw_mux_dac_a_mux_sel;
    wire [16:0]o_sample_dc_offset_i;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(35[28:48])
    
    wire n19392;
    wire [31:0]\addr_space[0] ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(48[12:22])
    wire [29:0]carrier_center_increment_offset;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(112[20:51])
    
    wire n19393, n27179, n27178, n27180;
    wire [31:0]\addr_space[4] ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(48[12:22])
    wire [15:0]n694;
    wire [15:0]n34;
    
    wire n19391;
    wire [31:0]\addr_space[1] ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(48[12:22])
    wire [31:0]\addr_space[3] ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(48[12:22])
    
    wire n26951, n19390;
    wire [31:0]\addr_space[2] ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(48[12:22])
    
    wire n26952, n27104, n27103, n27105, n27204, n27203, n27086, 
        n27085, n27087, n27210, n27211, n27081, n27080, n27082, 
        n27225, n27226, n27238, n27237, n27076, n27075, n27077, 
        n27251, n27250, n27272, n27273, n27277, n27278, n27298, 
        n27297, n27068, n27067, n27069, n19389, n27063, n27062, 
        n27064, n19388, n27058, n27057, n27059, n27053, n27052, 
        n27054, n19387, n27048, n27047, n27049, n27043, n27042, 
        n27044, n27038, n27037, n27039, n27033, n27032, n27034, 
        n27028, n27027, n27029, n19386, n19385, n19384, n27023, 
        n27022, n27024, n27007, n27006, n27008;
    wire [15:0]n33;
    
    wire n27002, n27001, n27003, n26997, n26996, n26998, n26987, 
        n26986, n26988, n26982, n26981, n26983, n26972, n26971, 
        n26973, n26962, n26961, n26963, n26957, n26956, n26958, 
        n26953, n29455, n27299, n27279, n27274, n27252, n27239, 
        n27227, n27212, n27205, cw_N_1500, dac_clk_p_c_enable_595, 
        dac_clk_p_c_enable_598, n19398, n19397, dac_clk_p_c_enable_617, 
        n19396, cw, dac_clk_p_c_enable_630;
    wire [13:0]u_s;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(61[18:21])
    
    wire n9468;
    wire [13:0]u_s_adj_3684;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(61[18:21])
    
    wire n9444, n9446, n9448, n9450, n9452, n9454, n9458, n9460, 
        n9462, n9464, n9466;
    wire [13:0]u_s_adj_3685;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(61[18:21])
    
    wire n9490, n9492, n19395, n9494, n9496, n19394, n9498, n9504, 
        n9506, n9488, n9456;
    wire [15:0]quarter_wave_sample_register_i;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(22[24:54])
    
    FD1S3AX o_dac_b_registered_i1 (.D(o_dac_b[0]), .CK(dac_clk_p_c), .Q(o_dac_b_c_0)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(25[8] 28[4])
    defparam o_dac_b_registered_i1.GSR = "DISABLED";
    FD1S3AX o_wb_data_i0 (.D(o_wb_data_31__N_1104[0]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(64[8] 66[4])
    defparam o_wb_data_i0.GSR = "DISABLED";
    FD1S3DX carrier_increment_i0 (.D(carrier_increment_30__N_1296[0]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_increment[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(118[11] 120[5])
    defparam carrier_increment_i0.GSR = "DISABLED";
    FD1S3IX o_dac_a_registered_i1 (.D(o_sample_dc_offset_i[7]), .CK(dac_clk_p_c), 
            .CD(cw_mux_dac_a_mux_sel), .Q(o_dac_a_c_0)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(25[8] 28[4])
    defparam o_dac_a_registered_i1.GSR = "DISABLED";
    CCU2D addr_space_0__30__I_0_20 (.A0(\addr_space[0] [18]), .B0(carrier_center_increment_offset[18]), 
          .C0(GND_net), .D0(GND_net), .A1(\addr_space[0] [19]), .B1(carrier_center_increment_offset[19]), 
          .C1(GND_net), .D1(GND_net), .CIN(n19392), .COUT(n19393), .S0(carrier_increment_30__N_1296[18]), 
          .S1(carrier_increment_30__N_1296[19]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(119[24:82])
    defparam addr_space_0__30__I_0_20.INIT0 = 16'h5666;
    defparam addr_space_0__30__I_0_20.INIT1 = 16'h5666;
    defparam addr_space_0__30__I_0_20.INJECT1_0 = "NO";
    defparam addr_space_0__30__I_0_20.INJECT1_1 = "NO";
    PFUMX i25474 (.BLUT(n27179), .ALUT(n27178), .C0(\wb_addr[0] ), .Z(n27180));
    LUT4 n27180_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4] [9]), .C(\wb_addr[2] ), 
         .D(n27180), .Z(o_wb_data_31__N_1104[9])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n27180_bdd_3_lut_4_lut.init = 16'h8f80;
    FD1S3BX startup_timer_FSM_i0_i0 (.D(n34[0]), .CK(dac_clk_p_c), .PD(i_sw0_c), 
            .Q(n694[0]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(155[21:41])
    defparam startup_timer_FSM_i0_i0.GSR = "DISABLED";
    CCU2D addr_space_0__30__I_0_18 (.A0(\addr_space[0] [16]), .B0(carrier_center_increment_offset[16]), 
          .C0(GND_net), .D0(GND_net), .A1(\addr_space[0] [17]), .B1(carrier_center_increment_offset[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n19391), .COUT(n19392), .S0(carrier_increment_30__N_1296[16]), 
          .S1(carrier_increment_30__N_1296[17]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(119[24:82])
    defparam addr_space_0__30__I_0_18.INIT0 = 16'h5666;
    defparam addr_space_0__30__I_0_18.INIT1 = 16'h5666;
    defparam addr_space_0__30__I_0_18.INJECT1_0 = "NO";
    defparam addr_space_0__30__I_0_18.INJECT1_1 = "NO";
    LUT4 \addr_space_0[[31__bdd_3_lut_25271  (.A(\addr_space[1] [31]), .B(\addr_space[3] [31]), 
         .C(\wb_addr[1] ), .Z(n26951)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[31__bdd_3_lut_25271 .init = 16'hcaca;
    CCU2D addr_space_0__30__I_0_16 (.A0(\addr_space[0] [14]), .B0(carrier_center_increment_offset[14]), 
          .C0(GND_net), .D0(GND_net), .A1(\addr_space[0] [15]), .B1(carrier_center_increment_offset[15]), 
          .C1(GND_net), .D1(GND_net), .CIN(n19390), .COUT(n19391), .S0(carrier_increment_30__N_1296[14]), 
          .S1(carrier_increment_30__N_1296[15]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(119[24:82])
    defparam addr_space_0__30__I_0_16.INIT0 = 16'h5666;
    defparam addr_space_0__30__I_0_16.INIT1 = 16'h5666;
    defparam addr_space_0__30__I_0_16.INJECT1_0 = "NO";
    defparam addr_space_0__30__I_0_16.INJECT1_1 = "NO";
    FD1S3IX o_wb_ack_50 (.D(o_dac_a_9__N_1), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(wb_fm_ack)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(68[8] 73[4])
    defparam o_wb_ack_50.GSR = "DISABLED";
    FD1P3DX addr_space_4___i1 (.D(wb_odata[0]), .SP(dac_clk_p_c_enable_502), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[4] [0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i1.GSR = "DISABLED";
    LUT4 \addr_space_0[[31__bdd_3_lut_25642  (.A(\addr_space[0] [31]), .B(\addr_space[2] [31]), 
         .C(\wb_addr[1] ), .Z(n26952)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[31__bdd_3_lut_25642 .init = 16'hcaca;
    PFUMX i25396 (.BLUT(n27104), .ALUT(n27103), .C0(\wb_addr[0] ), .Z(n27105));
    LUT4 \addr_space_0[[8__bdd_3_lut_27067  (.A(\addr_space[0] [8]), .B(\addr_space[2] [8]), 
         .C(\wb_addr[1] ), .Z(n27204)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[8__bdd_3_lut_27067 .init = 16'hcaca;
    LUT4 \addr_space_0[[8__bdd_3_lut_25492  (.A(\addr_space[1] [8]), .B(\addr_space[3] [8]), 
         .C(\wb_addr[1] ), .Z(n27203)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[8__bdd_3_lut_25492 .init = 16'hcaca;
    PFUMX i25377 (.BLUT(n27086), .ALUT(n27085), .C0(\wb_addr[0] ), .Z(n27087));
    LUT4 i1_3_lut (.A(\wb_addr[0] ), .B(\wb_addr[1] ), .C(\wb_addr[2] ), 
         .Z(n21641)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(59[4:25])
    defparam i1_3_lut.init = 16'hfbfb;
    LUT4 \addr_space_0[[7__bdd_3_lut_25496  (.A(\addr_space[1] [7]), .B(\addr_space[3] [7]), 
         .C(\wb_addr[1] ), .Z(n27210)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[7__bdd_3_lut_25496 .init = 16'hcaca;
    LUT4 \addr_space_0[[7__bdd_3_lut_27063  (.A(\addr_space[0] [7]), .B(\addr_space[2] [7]), 
         .C(\wb_addr[1] ), .Z(n27211)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[7__bdd_3_lut_27063 .init = 16'hcaca;
    PFUMX i25373 (.BLUT(n27081), .ALUT(n27080), .C0(\wb_addr[0] ), .Z(n27082));
    LUT4 \addr_space_0[[6__bdd_3_lut_25510  (.A(\addr_space[1] [6]), .B(\addr_space[3] [6]), 
         .C(\wb_addr[1] ), .Z(n27225)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[6__bdd_3_lut_25510 .init = 16'hcaca;
    LUT4 \addr_space_0[[6__bdd_3_lut_27059  (.A(\addr_space[0] [6]), .B(\addr_space[2] [6]), 
         .C(\wb_addr[1] ), .Z(n27226)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[6__bdd_3_lut_27059 .init = 16'hcaca;
    LUT4 \addr_space_0[[5__bdd_3_lut_27053  (.A(\addr_space[0] [5]), .B(\addr_space[2] [5]), 
         .C(\wb_addr[1] ), .Z(n27238)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[5__bdd_3_lut_27053 .init = 16'hcaca;
    LUT4 \addr_space_0[[5__bdd_3_lut_25522  (.A(\addr_space[1] [5]), .B(\addr_space[3] [5]), 
         .C(\wb_addr[1] ), .Z(n27237)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[5__bdd_3_lut_25522 .init = 16'hcaca;
    PFUMX i25369 (.BLUT(n27076), .ALUT(n27075), .C0(\wb_addr[0] ), .Z(n27077));
    LUT4 \addr_space_0[[4__bdd_3_lut_27049  (.A(\addr_space[0] [4]), .B(\addr_space[2] [4]), 
         .C(\wb_addr[1] ), .Z(n27251)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[4__bdd_3_lut_27049 .init = 16'hcaca;
    LUT4 \addr_space_0[[4__bdd_3_lut_25532  (.A(\addr_space[1] [4]), .B(\addr_space[3] [4]), 
         .C(\wb_addr[1] ), .Z(n27250)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[4__bdd_3_lut_25532 .init = 16'hcaca;
    LUT4 \addr_space_0[[3__bdd_3_lut_25549  (.A(\addr_space[1] [3]), .B(\addr_space[3] [3]), 
         .C(\wb_addr[1] ), .Z(n27272)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[3__bdd_3_lut_25549 .init = 16'hcaca;
    LUT4 \addr_space_0[[3__bdd_3_lut_27045  (.A(\addr_space[0] [3]), .B(\addr_space[2] [3]), 
         .C(\wb_addr[1] ), .Z(n27273)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[3__bdd_3_lut_27045 .init = 16'hcaca;
    LUT4 \addr_space_0[[2__bdd_3_lut_25553  (.A(\addr_space[1] [2]), .B(\addr_space[3] [2]), 
         .C(\wb_addr[1] ), .Z(n27277)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[2__bdd_3_lut_25553 .init = 16'hcaca;
    LUT4 \addr_space_0[[2__bdd_3_lut_27041  (.A(\addr_space[0] [2]), .B(\addr_space[2] [2]), 
         .C(\wb_addr[1] ), .Z(n27278)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[2__bdd_3_lut_27041 .init = 16'hcaca;
    LUT4 \addr_space_0[[1__bdd_3_lut_27037  (.A(\addr_space[0] [1]), .B(\addr_space[2] [1]), 
         .C(\wb_addr[1] ), .Z(n27298)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[1__bdd_3_lut_27037 .init = 16'hcaca;
    LUT4 \addr_space_0[[1__bdd_3_lut_25571  (.A(\addr_space[1] [1]), .B(\addr_space[3] [1]), 
         .C(\wb_addr[1] ), .Z(n27297)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[1__bdd_3_lut_25571 .init = 16'hcaca;
    PFUMX i25363 (.BLUT(n27068), .ALUT(n27067), .C0(\wb_addr[0] ), .Z(n27069));
    CCU2D addr_space_0__30__I_0_14 (.A0(\addr_space[0] [12]), .B0(carrier_center_increment_offset[12]), 
          .C0(GND_net), .D0(GND_net), .A1(\addr_space[0] [13]), .B1(carrier_center_increment_offset[13]), 
          .C1(GND_net), .D1(GND_net), .CIN(n19389), .COUT(n19390), .S0(carrier_increment_30__N_1296[12]), 
          .S1(carrier_increment_30__N_1296[13]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(119[24:82])
    defparam addr_space_0__30__I_0_14.INIT0 = 16'h5666;
    defparam addr_space_0__30__I_0_14.INIT1 = 16'h5666;
    defparam addr_space_0__30__I_0_14.INJECT1_0 = "NO";
    defparam addr_space_0__30__I_0_14.INJECT1_1 = "NO";
    PFUMX i25359 (.BLUT(n27063), .ALUT(n27062), .C0(\wb_addr[0] ), .Z(n27064));
    CCU2D addr_space_0__30__I_0_12 (.A0(\addr_space[0] [10]), .B0(carrier_center_increment_offset[10]), 
          .C0(GND_net), .D0(GND_net), .A1(\addr_space[0] [11]), .B1(carrier_center_increment_offset[11]), 
          .C1(GND_net), .D1(GND_net), .CIN(n19388), .COUT(n19389), .S0(carrier_increment_30__N_1296[10]), 
          .S1(carrier_increment_30__N_1296[11]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(119[24:82])
    defparam addr_space_0__30__I_0_12.INIT0 = 16'h5666;
    defparam addr_space_0__30__I_0_12.INIT1 = 16'h5666;
    defparam addr_space_0__30__I_0_12.INJECT1_0 = "NO";
    defparam addr_space_0__30__I_0_12.INJECT1_1 = "NO";
    PFUMX i25355 (.BLUT(n27058), .ALUT(n27057), .C0(\wb_addr[0] ), .Z(n27059));
    PFUMX i25351 (.BLUT(n27053), .ALUT(n27052), .C0(\wb_addr[0] ), .Z(n27054));
    CCU2D addr_space_0__30__I_0_10 (.A0(\addr_space[0] [8]), .B0(carrier_center_increment_offset[8]), 
          .C0(GND_net), .D0(GND_net), .A1(\addr_space[0] [9]), .B1(carrier_center_increment_offset[9]), 
          .C1(GND_net), .D1(GND_net), .CIN(n19387), .COUT(n19388), .S0(carrier_increment_30__N_1296[8]), 
          .S1(carrier_increment_30__N_1296[9]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(119[24:82])
    defparam addr_space_0__30__I_0_10.INIT0 = 16'h5666;
    defparam addr_space_0__30__I_0_10.INIT1 = 16'h5666;
    defparam addr_space_0__30__I_0_10.INJECT1_0 = "NO";
    defparam addr_space_0__30__I_0_10.INJECT1_1 = "NO";
    PFUMX i25347 (.BLUT(n27048), .ALUT(n27047), .C0(\wb_addr[0] ), .Z(n27049));
    PFUMX i25343 (.BLUT(n27043), .ALUT(n27042), .C0(\wb_addr[0] ), .Z(n27044));
    PFUMX i25339 (.BLUT(n27038), .ALUT(n27037), .C0(\wb_addr[0] ), .Z(n27039));
    PFUMX i25335 (.BLUT(n27033), .ALUT(n27032), .C0(\wb_addr[0] ), .Z(n27034));
    PFUMX i25331 (.BLUT(n27028), .ALUT(n27027), .C0(\wb_addr[0] ), .Z(n27029));
    CCU2D addr_space_0__30__I_0_8 (.A0(\addr_space[0] [6]), .B0(carrier_center_increment_offset[6]), 
          .C0(GND_net), .D0(GND_net), .A1(\addr_space[0] [7]), .B1(carrier_center_increment_offset[7]), 
          .C1(GND_net), .D1(GND_net), .CIN(n19386), .COUT(n19387), .S0(carrier_increment_30__N_1296[6]), 
          .S1(carrier_increment_30__N_1296[7]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(119[24:82])
    defparam addr_space_0__30__I_0_8.INIT0 = 16'h5666;
    defparam addr_space_0__30__I_0_8.INIT1 = 16'h5666;
    defparam addr_space_0__30__I_0_8.INJECT1_0 = "NO";
    defparam addr_space_0__30__I_0_8.INJECT1_1 = "NO";
    CCU2D addr_space_0__30__I_0_6 (.A0(\addr_space[0] [4]), .B0(carrier_center_increment_offset[4]), 
          .C0(GND_net), .D0(GND_net), .A1(\addr_space[0] [5]), .B1(carrier_center_increment_offset[5]), 
          .C1(GND_net), .D1(GND_net), .CIN(n19385), .COUT(n19386), .S0(carrier_increment_30__N_1296[4]), 
          .S1(carrier_increment_30__N_1296[5]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(119[24:82])
    defparam addr_space_0__30__I_0_6.INIT0 = 16'h5666;
    defparam addr_space_0__30__I_0_6.INIT1 = 16'h5666;
    defparam addr_space_0__30__I_0_6.INJECT1_0 = "NO";
    defparam addr_space_0__30__I_0_6.INJECT1_1 = "NO";
    CCU2D addr_space_0__30__I_0_4 (.A0(\addr_space[0] [2]), .B0(carrier_center_increment_offset[2]), 
          .C0(GND_net), .D0(GND_net), .A1(\addr_space[0] [3]), .B1(carrier_center_increment_offset[3]), 
          .C1(GND_net), .D1(GND_net), .CIN(n19384), .COUT(n19385), .S0(carrier_increment_30__N_1296[2]), 
          .S1(carrier_increment_30__N_1296[3]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(119[24:82])
    defparam addr_space_0__30__I_0_4.INIT0 = 16'h5666;
    defparam addr_space_0__30__I_0_4.INIT1 = 16'h5666;
    defparam addr_space_0__30__I_0_4.INJECT1_0 = "NO";
    defparam addr_space_0__30__I_0_4.INJECT1_1 = "NO";
    CCU2D addr_space_0__30__I_0_2 (.A0(\addr_space[0] [0]), .B0(carrier_center_increment_offset[0]), 
          .C0(GND_net), .D0(GND_net), .A1(\addr_space[0] [1]), .B1(carrier_center_increment_offset[1]), 
          .C1(GND_net), .D1(GND_net), .COUT(n19384), .S1(carrier_increment_30__N_1296[1]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(119[24:82])
    defparam addr_space_0__30__I_0_2.INIT0 = 16'h7000;
    defparam addr_space_0__30__I_0_2.INIT1 = 16'h5666;
    defparam addr_space_0__30__I_0_2.INJECT1_0 = "NO";
    defparam addr_space_0__30__I_0_2.INJECT1_1 = "NO";
    PFUMX i25327 (.BLUT(n27023), .ALUT(n27022), .C0(\wb_addr[0] ), .Z(n27024));
    LUT4 i24714_3_lut_4_lut (.A(n29300), .B(\wb_addr[2] ), .C(n29065), 
         .D(n22458), .Z(dac_clk_p_c_enable_227)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(59[4:25])
    defparam i24714_3_lut_4_lut.init = 16'h0008;
    PFUMX i25313 (.BLUT(n27007), .ALUT(n27006), .C0(\wb_addr[0] ), .Z(n27008));
    LUT4 i17602_2_lut (.A(\addr_space[0] [0]), .B(carrier_center_increment_offset[0]), 
         .Z(carrier_increment_30__N_1296[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i17602_2_lut.init = 16'h6666;
    LUT4 i7125_2_lut (.A(n694[0]), .B(n33[15]), .Z(n34[0])) /* synthesis lut_function=(A (B)) */ ;
    defparam i7125_2_lut.init = 16'h8888;
    PFUMX i25309 (.BLUT(n27002), .ALUT(n27001), .C0(\wb_addr[0] ), .Z(n27003));
    PFUMX i25305 (.BLUT(n26997), .ALUT(n26996), .C0(\wb_addr[0] ), .Z(n26998));
    PFUMX i25298 (.BLUT(n26987), .ALUT(n26986), .C0(\wb_addr[0] ), .Z(n26988));
    PFUMX i25294 (.BLUT(n26982), .ALUT(n26981), .C0(\wb_addr[0] ), .Z(n26983));
    PFUMX i25287 (.BLUT(n26972), .ALUT(n26971), .C0(\wb_addr[0] ), .Z(n26973));
    PFUMX i25280 (.BLUT(n26962), .ALUT(n26961), .C0(\wb_addr[0] ), .Z(n26963));
    PFUMX i25276 (.BLUT(n26957), .ALUT(n26956), .C0(\wb_addr[0] ), .Z(n26958));
    PFUMX i25272 (.BLUT(n26952), .ALUT(n26951), .C0(\wb_addr[0] ), .Z(n26953));
    FD1S3IX o_dac_a_registered_i10 (.D(o_sample_dc_offset_i[16]), .CK(dac_clk_p_c), 
            .CD(cw_mux_dac_a_mux_sel), .Q(o_dac_a_c_9)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(25[8] 28[4])
    defparam o_dac_a_registered_i10.GSR = "DISABLED";
    LUT4 \addr_space_0[[9__bdd_3_lut  (.A(\addr_space[0] [9]), .B(\addr_space[2] [9]), 
         .C(\wb_addr[1] ), .Z(n27179)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[9__bdd_3_lut .init = 16'hcaca;
    LUT4 \addr_space_0[[9__bdd_3_lut_25473  (.A(\addr_space[1] [9]), .B(\addr_space[3] [9]), 
         .C(\wb_addr[1] ), .Z(n27178)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[9__bdd_3_lut_25473 .init = 16'hcaca;
    LUT4 i24646_2_lut_3_lut_4_lut (.A(\wb_addr[1] ), .B(n29455), .C(n29065), 
         .D(n22458), .Z(dac_clk_p_c_enable_241)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(59[4:25])
    defparam i24646_2_lut_3_lut_4_lut.init = 16'h0002;
    LUT4 i24650_2_lut_3_lut_4_lut (.A(\wb_addr[1] ), .B(n29455), .C(n29065), 
         .D(n22458), .Z(dac_clk_p_c_enable_106)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(59[4:25])
    defparam i24650_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 n27299_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4] [1]), .C(\wb_addr[2] ), 
         .D(n27299), .Z(o_wb_data_31__N_1104[1])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n27299_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 n27279_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4] [2]), .C(\wb_addr[2] ), 
         .D(n27279), .Z(o_wb_data_31__N_1104[2])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n27279_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 n27274_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4] [3]), .C(\wb_addr[2] ), 
         .D(n27274), .Z(o_wb_data_31__N_1104[3])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n27274_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 n27252_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4] [4]), .C(\wb_addr[2] ), 
         .D(n27252), .Z(o_wb_data_31__N_1104[4])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n27252_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 n27239_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4] [5]), .C(\wb_addr[2] ), 
         .D(n27239), .Z(o_wb_data_31__N_1104[5])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n27239_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 n27227_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4] [6]), .C(\wb_addr[2] ), 
         .D(n27227), .Z(o_wb_data_31__N_1104[6])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n27227_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 n27212_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4] [7]), .C(\wb_addr[2] ), 
         .D(n27212), .Z(o_wb_data_31__N_1104[7])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n27212_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 n27205_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4] [8]), .C(\wb_addr[2] ), 
         .D(n27205), .Z(o_wb_data_31__N_1104[8])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n27205_bdd_3_lut_4_lut.init = 16'h8f80;
    FD1S3JX o_dac_a_registered_i9 (.D(o_sample_dc_offset_i[15]), .CK(dac_clk_p_c), 
            .PD(cw_mux_dac_a_mux_sel), .Q(o_dac_a_c_8)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(25[8] 28[4])
    defparam o_dac_a_registered_i9.GSR = "DISABLED";
    FD1S3IX o_dac_a_registered_i8 (.D(o_sample_dc_offset_i[14]), .CK(dac_clk_p_c), 
            .CD(cw_mux_dac_a_mux_sel), .Q(o_dac_a_c_7)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(25[8] 28[4])
    defparam o_dac_a_registered_i8.GSR = "DISABLED";
    FD1S3IX o_dac_a_registered_i7 (.D(o_sample_dc_offset_i[13]), .CK(dac_clk_p_c), 
            .CD(cw_mux_dac_a_mux_sel), .Q(o_dac_a_c_6)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(25[8] 28[4])
    defparam o_dac_a_registered_i7.GSR = "DISABLED";
    FD1S3JX o_dac_a_registered_i6 (.D(o_sample_dc_offset_i[12]), .CK(dac_clk_p_c), 
            .PD(cw_mux_dac_a_mux_sel), .Q(o_dac_a_c_5)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(25[8] 28[4])
    defparam o_dac_a_registered_i6.GSR = "DISABLED";
    FD1S3IX o_dac_a_registered_i5 (.D(o_sample_dc_offset_i[11]), .CK(dac_clk_p_c), 
            .CD(cw_mux_dac_a_mux_sel), .Q(o_dac_a_c_4)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(25[8] 28[4])
    defparam o_dac_a_registered_i5.GSR = "DISABLED";
    FD1S3IX o_dac_a_registered_i4 (.D(o_sample_dc_offset_i[10]), .CK(dac_clk_p_c), 
            .CD(cw_mux_dac_a_mux_sel), .Q(o_dac_a_c_3)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(25[8] 28[4])
    defparam o_dac_a_registered_i4.GSR = "DISABLED";
    FD1S3IX o_dac_a_registered_i3 (.D(o_sample_dc_offset_i[9]), .CK(dac_clk_p_c), 
            .CD(cw_mux_dac_a_mux_sel), .Q(o_dac_a_c_2)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(25[8] 28[4])
    defparam o_dac_a_registered_i3.GSR = "DISABLED";
    FD1S3IX o_dac_a_registered_i2 (.D(o_sample_dc_offset_i[8]), .CK(dac_clk_p_c), 
            .CD(cw_mux_dac_a_mux_sel), .Q(o_dac_a_c_1)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(25[8] 28[4])
    defparam o_dac_a_registered_i2.GSR = "DISABLED";
    FD1S3DX carrier_increment_i30 (.D(carrier_increment_30__N_1296[30]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_increment[30])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(118[11] 120[5])
    defparam carrier_increment_i30.GSR = "DISABLED";
    FD1S3DX carrier_increment_i29 (.D(carrier_increment_30__N_1296[29]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_increment[29])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(118[11] 120[5])
    defparam carrier_increment_i29.GSR = "DISABLED";
    FD1S3DX carrier_increment_i28 (.D(carrier_increment_30__N_1296[28]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_increment[28])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(118[11] 120[5])
    defparam carrier_increment_i28.GSR = "DISABLED";
    FD1S3DX carrier_increment_i27 (.D(carrier_increment_30__N_1296[27]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_increment[27])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(118[11] 120[5])
    defparam carrier_increment_i27.GSR = "DISABLED";
    FD1S3DX carrier_increment_i26 (.D(carrier_increment_30__N_1296[26]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_increment[26])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(118[11] 120[5])
    defparam carrier_increment_i26.GSR = "DISABLED";
    FD1S3DX carrier_increment_i25 (.D(carrier_increment_30__N_1296[25]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_increment[25])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(118[11] 120[5])
    defparam carrier_increment_i25.GSR = "DISABLED";
    FD1S3DX carrier_increment_i24 (.D(carrier_increment_30__N_1296[24]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_increment[24])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(118[11] 120[5])
    defparam carrier_increment_i24.GSR = "DISABLED";
    FD1S3DX carrier_increment_i23 (.D(carrier_increment_30__N_1296[23]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_increment[23])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(118[11] 120[5])
    defparam carrier_increment_i23.GSR = "DISABLED";
    FD1S3DX carrier_increment_i22 (.D(carrier_increment_30__N_1296[22]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_increment[22])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(118[11] 120[5])
    defparam carrier_increment_i22.GSR = "DISABLED";
    FD1S3DX carrier_increment_i21 (.D(carrier_increment_30__N_1296[21]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_increment[21])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(118[11] 120[5])
    defparam carrier_increment_i21.GSR = "DISABLED";
    FD1S3DX carrier_increment_i20 (.D(carrier_increment_30__N_1296[20]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_increment[20])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(118[11] 120[5])
    defparam carrier_increment_i20.GSR = "DISABLED";
    FD1S3DX carrier_increment_i19 (.D(carrier_increment_30__N_1296[19]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_increment[19])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(118[11] 120[5])
    defparam carrier_increment_i19.GSR = "DISABLED";
    FD1S3DX carrier_increment_i18 (.D(carrier_increment_30__N_1296[18]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_increment[18])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(118[11] 120[5])
    defparam carrier_increment_i18.GSR = "DISABLED";
    FD1S3DX carrier_increment_i17 (.D(carrier_increment_30__N_1296[17]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_increment[17])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(118[11] 120[5])
    defparam carrier_increment_i17.GSR = "DISABLED";
    FD1S3DX carrier_increment_i16 (.D(carrier_increment_30__N_1296[16]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_increment[16])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(118[11] 120[5])
    defparam carrier_increment_i16.GSR = "DISABLED";
    FD1S3DX carrier_increment_i15 (.D(carrier_increment_30__N_1296[15]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_increment[15])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(118[11] 120[5])
    defparam carrier_increment_i15.GSR = "DISABLED";
    FD1S3DX carrier_increment_i14 (.D(carrier_increment_30__N_1296[14]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_increment[14])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(118[11] 120[5])
    defparam carrier_increment_i14.GSR = "DISABLED";
    FD1S3DX carrier_increment_i13 (.D(carrier_increment_30__N_1296[13]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_increment[13])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(118[11] 120[5])
    defparam carrier_increment_i13.GSR = "DISABLED";
    FD1S3DX carrier_increment_i12 (.D(carrier_increment_30__N_1296[12]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_increment[12])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(118[11] 120[5])
    defparam carrier_increment_i12.GSR = "DISABLED";
    FD1S3DX carrier_increment_i11 (.D(carrier_increment_30__N_1296[11]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_increment[11])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(118[11] 120[5])
    defparam carrier_increment_i11.GSR = "DISABLED";
    FD1S3DX carrier_increment_i10 (.D(carrier_increment_30__N_1296[10]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_increment[10])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(118[11] 120[5])
    defparam carrier_increment_i10.GSR = "DISABLED";
    FD1S3DX carrier_increment_i9 (.D(carrier_increment_30__N_1296[9]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_increment[9])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(118[11] 120[5])
    defparam carrier_increment_i9.GSR = "DISABLED";
    FD1S3DX carrier_increment_i8 (.D(carrier_increment_30__N_1296[8]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_increment[8])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(118[11] 120[5])
    defparam carrier_increment_i8.GSR = "DISABLED";
    FD1S3DX carrier_increment_i7 (.D(carrier_increment_30__N_1296[7]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_increment[7])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(118[11] 120[5])
    defparam carrier_increment_i7.GSR = "DISABLED";
    FD1S3DX carrier_increment_i6 (.D(carrier_increment_30__N_1296[6]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_increment[6])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(118[11] 120[5])
    defparam carrier_increment_i6.GSR = "DISABLED";
    FD1S3DX carrier_increment_i5 (.D(carrier_increment_30__N_1296[5]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_increment[5])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(118[11] 120[5])
    defparam carrier_increment_i5.GSR = "DISABLED";
    FD1S3DX carrier_increment_i4 (.D(carrier_increment_30__N_1296[4]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_increment[4])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(118[11] 120[5])
    defparam carrier_increment_i4.GSR = "DISABLED";
    FD1S3DX carrier_increment_i3 (.D(carrier_increment_30__N_1296[3]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_increment[3])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(118[11] 120[5])
    defparam carrier_increment_i3.GSR = "DISABLED";
    FD1S3DX carrier_increment_i2 (.D(carrier_increment_30__N_1296[2]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_increment[2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(118[11] 120[5])
    defparam carrier_increment_i2.GSR = "DISABLED";
    FD1S3DX carrier_increment_i1 (.D(carrier_increment_30__N_1296[1]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(carrier_increment[1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(118[11] 120[5])
    defparam carrier_increment_i1.GSR = "DISABLED";
    FD1S3AX o_wb_data_i31 (.D(o_wb_data_31__N_1104[31]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[31])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(64[8] 66[4])
    defparam o_wb_data_i31.GSR = "DISABLED";
    FD1S3AX o_wb_data_i30 (.D(o_wb_data_31__N_1104[30]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[30])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(64[8] 66[4])
    defparam o_wb_data_i30.GSR = "DISABLED";
    FD1S3AX o_wb_data_i29 (.D(o_wb_data_31__N_1104[29]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[29])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(64[8] 66[4])
    defparam o_wb_data_i29.GSR = "DISABLED";
    FD1S3AX o_wb_data_i28 (.D(o_wb_data_31__N_1104[28]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[28])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(64[8] 66[4])
    defparam o_wb_data_i28.GSR = "DISABLED";
    FD1S3AX o_wb_data_i27 (.D(o_wb_data_31__N_1104[27]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[27])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(64[8] 66[4])
    defparam o_wb_data_i27.GSR = "DISABLED";
    FD1S3AX o_wb_data_i26 (.D(o_wb_data_31__N_1104[26]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[26])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(64[8] 66[4])
    defparam o_wb_data_i26.GSR = "DISABLED";
    FD1S3AX o_wb_data_i25 (.D(o_wb_data_31__N_1104[25]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[25])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(64[8] 66[4])
    defparam o_wb_data_i25.GSR = "DISABLED";
    FD1S3AX o_wb_data_i24 (.D(o_wb_data_31__N_1104[24]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[24])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(64[8] 66[4])
    defparam o_wb_data_i24.GSR = "DISABLED";
    FD1S3AX o_wb_data_i23 (.D(o_wb_data_31__N_1104[23]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[23])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(64[8] 66[4])
    defparam o_wb_data_i23.GSR = "DISABLED";
    FD1S3AX o_wb_data_i22 (.D(o_wb_data_31__N_1104[22]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[22])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(64[8] 66[4])
    defparam o_wb_data_i22.GSR = "DISABLED";
    FD1S3AX o_wb_data_i21 (.D(o_wb_data_31__N_1104[21]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[21])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(64[8] 66[4])
    defparam o_wb_data_i21.GSR = "DISABLED";
    FD1S3AX o_wb_data_i20 (.D(o_wb_data_31__N_1104[20]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[20])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(64[8] 66[4])
    defparam o_wb_data_i20.GSR = "DISABLED";
    FD1S3AX o_wb_data_i19 (.D(o_wb_data_31__N_1104[19]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[19])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(64[8] 66[4])
    defparam o_wb_data_i19.GSR = "DISABLED";
    FD1S3AX o_wb_data_i18 (.D(o_wb_data_31__N_1104[18]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[18])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(64[8] 66[4])
    defparam o_wb_data_i18.GSR = "DISABLED";
    FD1S3AX o_wb_data_i17 (.D(o_wb_data_31__N_1104[17]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[17])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(64[8] 66[4])
    defparam o_wb_data_i17.GSR = "DISABLED";
    FD1S3AX o_wb_data_i16 (.D(o_wb_data_31__N_1104[16]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[16])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(64[8] 66[4])
    defparam o_wb_data_i16.GSR = "DISABLED";
    FD1S3AX o_wb_data_i15 (.D(o_wb_data_31__N_1104[15]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[15])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(64[8] 66[4])
    defparam o_wb_data_i15.GSR = "DISABLED";
    FD1S3AX o_wb_data_i14 (.D(o_wb_data_31__N_1104[14]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[14])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(64[8] 66[4])
    defparam o_wb_data_i14.GSR = "DISABLED";
    FD1S3AX o_wb_data_i13 (.D(o_wb_data_31__N_1104[13]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[13])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(64[8] 66[4])
    defparam o_wb_data_i13.GSR = "DISABLED";
    FD1S3AX o_wb_data_i12 (.D(o_wb_data_31__N_1104[12]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[12])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(64[8] 66[4])
    defparam o_wb_data_i12.GSR = "DISABLED";
    FD1S3AX o_wb_data_i11 (.D(o_wb_data_31__N_1104[11]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[11])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(64[8] 66[4])
    defparam o_wb_data_i11.GSR = "DISABLED";
    FD1S3AX o_wb_data_i10 (.D(o_wb_data_31__N_1104[10]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[10])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(64[8] 66[4])
    defparam o_wb_data_i10.GSR = "DISABLED";
    FD1S3AX o_wb_data_i9 (.D(o_wb_data_31__N_1104[9]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[9])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(64[8] 66[4])
    defparam o_wb_data_i9.GSR = "DISABLED";
    FD1S3AX o_wb_data_i8 (.D(o_wb_data_31__N_1104[8]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[8])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(64[8] 66[4])
    defparam o_wb_data_i8.GSR = "DISABLED";
    FD1S3AX o_wb_data_i7 (.D(o_wb_data_31__N_1104[7]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[7])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(64[8] 66[4])
    defparam o_wb_data_i7.GSR = "DISABLED";
    FD1S3AX o_wb_data_i6 (.D(o_wb_data_31__N_1104[6]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[6])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(64[8] 66[4])
    defparam o_wb_data_i6.GSR = "DISABLED";
    FD1S3AX o_wb_data_i5 (.D(o_wb_data_31__N_1104[5]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[5])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(64[8] 66[4])
    defparam o_wb_data_i5.GSR = "DISABLED";
    FD1S3AX o_wb_data_i4 (.D(o_wb_data_31__N_1104[4]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[4])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(64[8] 66[4])
    defparam o_wb_data_i4.GSR = "DISABLED";
    FD1S3AX o_wb_data_i3 (.D(o_wb_data_31__N_1104[3]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[3])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(64[8] 66[4])
    defparam o_wb_data_i3.GSR = "DISABLED";
    FD1S3AX o_wb_data_i2 (.D(o_wb_data_31__N_1104[2]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(64[8] 66[4])
    defparam o_wb_data_i2.GSR = "DISABLED";
    FD1S3AX o_wb_data_i1 (.D(o_wb_data_31__N_1104[1]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(64[8] 66[4])
    defparam o_wb_data_i1.GSR = "DISABLED";
    FD1S3AX o_dac_b_registered_i10 (.D(o_dac_b[9]), .CK(dac_clk_p_c), .Q(o_dac_b_c_9)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(25[8] 28[4])
    defparam o_dac_b_registered_i10.GSR = "DISABLED";
    LUT4 i1303_1_lut (.A(o_sample_dc_offset_i[15]), .Z(o_sample_dc_offset_i[16])) /* synthesis lut_function=(!(A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(37[31:77])
    defparam i1303_1_lut.init = 16'h5555;
    FD1S3AX o_dac_b_registered_i9 (.D(o_dac_b[8]), .CK(dac_clk_p_c), .Q(o_dac_b_c_8)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(25[8] 28[4])
    defparam o_dac_b_registered_i9.GSR = "DISABLED";
    FD1S3AX o_dac_b_registered_i8 (.D(o_dac_b[7]), .CK(dac_clk_p_c), .Q(o_dac_b_c_7)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(25[8] 28[4])
    defparam o_dac_b_registered_i8.GSR = "DISABLED";
    FD1S3AX o_dac_b_registered_i7 (.D(o_dac_b[6]), .CK(dac_clk_p_c), .Q(o_dac_b_c_6)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(25[8] 28[4])
    defparam o_dac_b_registered_i7.GSR = "DISABLED";
    FD1S3AX o_dac_b_registered_i6 (.D(o_dac_b[5]), .CK(dac_clk_p_c), .Q(o_dac_b_c_5)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(25[8] 28[4])
    defparam o_dac_b_registered_i6.GSR = "DISABLED";
    FD1S3AX o_dac_b_registered_i5 (.D(o_dac_b[4]), .CK(dac_clk_p_c), .Q(o_dac_b_c_4)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(25[8] 28[4])
    defparam o_dac_b_registered_i5.GSR = "DISABLED";
    FD1S3AX o_dac_b_registered_i4 (.D(o_dac_b[3]), .CK(dac_clk_p_c), .Q(o_dac_b_c_3)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(25[8] 28[4])
    defparam o_dac_b_registered_i4.GSR = "DISABLED";
    FD1S3AX o_dac_b_registered_i3 (.D(o_dac_b[2]), .CK(dac_clk_p_c), .Q(o_dac_b_c_2)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(25[8] 28[4])
    defparam o_dac_b_registered_i3.GSR = "DISABLED";
    FD1S3AX o_dac_b_registered_i2 (.D(o_dac_b[1]), .CK(dac_clk_p_c), .Q(o_dac_b_c_1)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(25[8] 28[4])
    defparam o_dac_b_registered_i2.GSR = "DISABLED";
    FD1P3DX addr_space_4___i160 (.D(wb_odata[31]), .SP(dac_clk_p_c_enable_375), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [31])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i160.GSR = "DISABLED";
    FD1P3DX addr_space_4___i159 (.D(wb_odata[30]), .SP(dac_clk_p_c_enable_375), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [30])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i159.GSR = "DISABLED";
    FD1P3DX addr_space_4___i158 (.D(wb_odata[29]), .SP(dac_clk_p_c_enable_375), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [29])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i158.GSR = "DISABLED";
    FD1P3DX addr_space_4___i157 (.D(wb_odata[28]), .SP(dac_clk_p_c_enable_375), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [28])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i157.GSR = "DISABLED";
    FD1P3DX addr_space_4___i156 (.D(wb_odata[27]), .SP(dac_clk_p_c_enable_375), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [27])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i156.GSR = "DISABLED";
    FD1P3DX addr_space_4___i155 (.D(wb_odata[26]), .SP(dac_clk_p_c_enable_375), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [26])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i155.GSR = "DISABLED";
    FD1P3DX addr_space_4___i154 (.D(wb_odata[25]), .SP(dac_clk_p_c_enable_375), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [25])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i154.GSR = "DISABLED";
    FD1P3DX addr_space_4___i153 (.D(wb_odata[24]), .SP(dac_clk_p_c_enable_375), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [24])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i153.GSR = "DISABLED";
    LUT4 n27105_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4] [10]), .C(\wb_addr[2] ), 
         .D(n27105), .Z(o_wb_data_31__N_1104[10])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n27105_bdd_3_lut_4_lut.init = 16'h8f80;
    FD1P3DX addr_space_4___i152 (.D(wb_odata[23]), .SP(dac_clk_p_c_enable_375), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [23])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i152.GSR = "DISABLED";
    FD1P3DX addr_space_4___i151 (.D(wb_odata[22]), .SP(dac_clk_p_c_enable_375), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [22])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i151.GSR = "DISABLED";
    FD1P3DX addr_space_4___i150 (.D(wb_odata[21]), .SP(dac_clk_p_c_enable_375), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [21])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i150.GSR = "DISABLED";
    FD1P3DX addr_space_4___i149 (.D(wb_odata[20]), .SP(dac_clk_p_c_enable_375), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [20])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i149.GSR = "DISABLED";
    FD1P3DX addr_space_4___i148 (.D(wb_odata[19]), .SP(dac_clk_p_c_enable_375), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [19])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i148.GSR = "DISABLED";
    FD1P3DX addr_space_4___i147 (.D(wb_odata[18]), .SP(dac_clk_p_c_enable_375), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [18])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i147.GSR = "DISABLED";
    FD1P3DX addr_space_4___i146 (.D(wb_odata[17]), .SP(dac_clk_p_c_enable_375), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [17])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i146.GSR = "DISABLED";
    FD1P3BX addr_space_4___i145 (.D(wb_odata[16]), .SP(dac_clk_p_c_enable_375), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(\addr_space[0] [16])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i145.GSR = "DISABLED";
    FD1P3BX addr_space_4___i144 (.D(wb_odata[15]), .SP(dac_clk_p_c_enable_375), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(\addr_space[0] [15])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i144.GSR = "DISABLED";
    FD1P3DX addr_space_4___i143 (.D(wb_odata[14]), .SP(dac_clk_p_c_enable_375), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [14])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i143.GSR = "DISABLED";
    FD1P3DX addr_space_4___i142 (.D(wb_odata[13]), .SP(dac_clk_p_c_enable_375), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [13])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i142.GSR = "DISABLED";
    FD1P3DX addr_space_4___i141 (.D(wb_odata[12]), .SP(dac_clk_p_c_enable_375), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [12])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i141.GSR = "DISABLED";
    FD1P3DX addr_space_4___i140 (.D(wb_odata[11]), .SP(dac_clk_p_c_enable_375), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [11])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i140.GSR = "DISABLED";
    FD1P3BX addr_space_4___i139 (.D(wb_odata[10]), .SP(dac_clk_p_c_enable_375), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(\addr_space[0] [10])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i139.GSR = "DISABLED";
    FD1P3BX addr_space_4___i138 (.D(wb_odata[9]), .SP(dac_clk_p_c_enable_375), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(\addr_space[0] [9])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i138.GSR = "DISABLED";
    FD1P3DX addr_space_4___i137 (.D(wb_odata[8]), .SP(dac_clk_p_c_enable_375), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [8])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i137.GSR = "DISABLED";
    FD1P3BX addr_space_4___i136 (.D(wb_odata[7]), .SP(dac_clk_p_c_enable_375), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(\addr_space[0] [7])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i136.GSR = "DISABLED";
    FD1P3DX addr_space_4___i135 (.D(wb_odata[6]), .SP(dac_clk_p_c_enable_375), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [6])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i135.GSR = "DISABLED";
    FD1P3BX addr_space_4___i134 (.D(wb_odata[5]), .SP(dac_clk_p_c_enable_375), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(\addr_space[0] [5])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i134.GSR = "DISABLED";
    FD1P3DX addr_space_4___i133 (.D(wb_odata[4]), .SP(dac_clk_p_c_enable_375), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [4])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i133.GSR = "DISABLED";
    FD1P3DX addr_space_4___i132 (.D(wb_odata[3]), .SP(dac_clk_p_c_enable_375), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [3])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i132.GSR = "DISABLED";
    FD1P3DX addr_space_4___i131 (.D(wb_odata[2]), .SP(dac_clk_p_c_enable_375), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i131.GSR = "DISABLED";
    FD1P3DX addr_space_4___i130 (.D(wb_odata[1]), .SP(dac_clk_p_c_enable_375), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i130.GSR = "DISABLED";
    FD1P3DX addr_space_4___i129 (.D(wb_odata[0]), .SP(dac_clk_p_c_enable_375), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[0] [0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i129.GSR = "DISABLED";
    FD1P3DX addr_space_4___i128 (.D(wb_odata[31]), .SP(dac_clk_p_c_enable_407), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[1] [31])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i128.GSR = "DISABLED";
    FD1P3DX addr_space_4___i127 (.D(wb_odata[30]), .SP(dac_clk_p_c_enable_407), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[1] [30])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i127.GSR = "DISABLED";
    FD1P3DX addr_space_4___i126 (.D(wb_odata[29]), .SP(dac_clk_p_c_enable_407), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[1] [29])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i126.GSR = "DISABLED";
    FD1P3DX addr_space_4___i125 (.D(wb_odata[28]), .SP(dac_clk_p_c_enable_407), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[1] [28])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i125.GSR = "DISABLED";
    FD1P3DX addr_space_4___i124 (.D(wb_odata[27]), .SP(dac_clk_p_c_enable_407), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[1] [27])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i124.GSR = "DISABLED";
    FD1P3DX addr_space_4___i123 (.D(wb_odata[26]), .SP(dac_clk_p_c_enable_407), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[1] [26])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i123.GSR = "DISABLED";
    FD1P3DX addr_space_4___i122 (.D(wb_odata[25]), .SP(dac_clk_p_c_enable_407), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[1] [25])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i122.GSR = "DISABLED";
    FD1P3DX addr_space_4___i121 (.D(wb_odata[24]), .SP(dac_clk_p_c_enable_407), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[1] [24])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i121.GSR = "DISABLED";
    FD1P3DX addr_space_4___i120 (.D(wb_odata[23]), .SP(dac_clk_p_c_enable_407), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[1] [23])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i120.GSR = "DISABLED";
    FD1P3DX addr_space_4___i119 (.D(wb_odata[22]), .SP(dac_clk_p_c_enable_407), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[1] [22])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i119.GSR = "DISABLED";
    FD1P3DX addr_space_4___i118 (.D(wb_odata[21]), .SP(dac_clk_p_c_enable_407), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[1] [21])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i118.GSR = "DISABLED";
    FD1P3DX addr_space_4___i117 (.D(wb_odata[20]), .SP(dac_clk_p_c_enable_407), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[1] [20])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i117.GSR = "DISABLED";
    FD1P3DX addr_space_4___i116 (.D(wb_odata[19]), .SP(dac_clk_p_c_enable_407), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[1] [19])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i116.GSR = "DISABLED";
    FD1P3DX addr_space_4___i115 (.D(wb_odata[18]), .SP(dac_clk_p_c_enable_407), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[1] [18])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i115.GSR = "DISABLED";
    FD1P3DX addr_space_4___i114 (.D(wb_odata[17]), .SP(dac_clk_p_c_enable_407), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[1] [17])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i114.GSR = "DISABLED";
    FD1P3BX addr_space_4___i113 (.D(wb_odata[16]), .SP(dac_clk_p_c_enable_407), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(\addr_space[1] [16])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i113.GSR = "DISABLED";
    FD1P3DX addr_space_4___i112 (.D(wb_odata[15]), .SP(dac_clk_p_c_enable_407), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[1] [15])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i112.GSR = "DISABLED";
    FD1P3BX addr_space_4___i111 (.D(wb_odata[14]), .SP(dac_clk_p_c_enable_407), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(\addr_space[1] [14])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i111.GSR = "DISABLED";
    FD1P3BX addr_space_4___i110 (.D(wb_odata[13]), .SP(dac_clk_p_c_enable_407), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(\addr_space[1] [13])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i110.GSR = "DISABLED";
    FD1P3BX addr_space_4___i109 (.D(wb_odata[12]), .SP(dac_clk_p_c_enable_407), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(\addr_space[1] [12])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i109.GSR = "DISABLED";
    FD1P3BX addr_space_4___i108 (.D(wb_odata[11]), .SP(dac_clk_p_c_enable_407), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(\addr_space[1] [11])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i108.GSR = "DISABLED";
    FD1P3DX addr_space_4___i107 (.D(wb_odata[10]), .SP(dac_clk_p_c_enable_407), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[1] [10])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i107.GSR = "DISABLED";
    FD1P3DX addr_space_4___i106 (.D(wb_odata[9]), .SP(dac_clk_p_c_enable_407), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[1] [9])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i106.GSR = "DISABLED";
    FD1P3BX addr_space_4___i105 (.D(wb_odata[8]), .SP(dac_clk_p_c_enable_407), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(\addr_space[1] [8])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i105.GSR = "DISABLED";
    FD1P3DX addr_space_4___i104 (.D(wb_odata[7]), .SP(dac_clk_p_c_enable_407), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[1] [7])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i104.GSR = "DISABLED";
    FD1P3DX addr_space_4___i103 (.D(wb_odata[6]), .SP(dac_clk_p_c_enable_407), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[1] [6])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i103.GSR = "DISABLED";
    FD1P3DX addr_space_4___i102 (.D(wb_odata[5]), .SP(dac_clk_p_c_enable_407), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[1] [5])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i102.GSR = "DISABLED";
    FD1P3DX addr_space_4___i101 (.D(wb_odata[4]), .SP(dac_clk_p_c_enable_407), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[1] [4])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i101.GSR = "DISABLED";
    FD1P3BX addr_space_4___i100 (.D(wb_odata[3]), .SP(dac_clk_p_c_enable_407), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(\addr_space[1] [3])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i100.GSR = "DISABLED";
    FD1P3DX addr_space_4___i99 (.D(wb_odata[2]), .SP(dac_clk_p_c_enable_407), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[1] [2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i99.GSR = "DISABLED";
    FD1P3BX addr_space_4___i98 (.D(wb_odata[1]), .SP(dac_clk_p_c_enable_407), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(\addr_space[1] [1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i98.GSR = "DISABLED";
    FD1P3BX addr_space_4___i97 (.D(wb_odata[0]), .SP(dac_clk_p_c_enable_407), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(\addr_space[1] [0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i97.GSR = "DISABLED";
    FD1P3DX addr_space_4___i96 (.D(wb_odata[31]), .SP(dac_clk_p_c_enable_439), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[2] [31])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i96.GSR = "DISABLED";
    FD1P3DX addr_space_4___i95 (.D(wb_odata[30]), .SP(dac_clk_p_c_enable_439), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[2] [30])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i95.GSR = "DISABLED";
    FD1P3DX addr_space_4___i94 (.D(wb_odata[29]), .SP(dac_clk_p_c_enable_439), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[2] [29])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i94.GSR = "DISABLED";
    FD1P3DX addr_space_4___i93 (.D(wb_odata[28]), .SP(dac_clk_p_c_enable_439), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[2] [28])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i93.GSR = "DISABLED";
    FD1P3DX addr_space_4___i92 (.D(wb_odata[27]), .SP(dac_clk_p_c_enable_439), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[2] [27])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i92.GSR = "DISABLED";
    FD1P3DX addr_space_4___i91 (.D(wb_odata[26]), .SP(dac_clk_p_c_enable_439), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[2] [26])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i91.GSR = "DISABLED";
    FD1P3DX addr_space_4___i90 (.D(wb_odata[25]), .SP(dac_clk_p_c_enable_439), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[2] [25])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i90.GSR = "DISABLED";
    FD1P3DX addr_space_4___i89 (.D(wb_odata[24]), .SP(dac_clk_p_c_enable_439), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[2] [24])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i89.GSR = "DISABLED";
    FD1P3DX addr_space_4___i88 (.D(wb_odata[23]), .SP(dac_clk_p_c_enable_439), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[2] [23])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i88.GSR = "DISABLED";
    FD1P3DX addr_space_4___i87 (.D(wb_odata[22]), .SP(dac_clk_p_c_enable_439), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[2] [22])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i87.GSR = "DISABLED";
    FD1P3DX addr_space_4___i86 (.D(wb_odata[21]), .SP(dac_clk_p_c_enable_439), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[2] [21])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i86.GSR = "DISABLED";
    FD1P3DX addr_space_4___i85 (.D(wb_odata[20]), .SP(dac_clk_p_c_enable_439), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[2] [20])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i85.GSR = "DISABLED";
    FD1P3DX addr_space_4___i84 (.D(wb_odata[19]), .SP(dac_clk_p_c_enable_439), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[2] [19])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i84.GSR = "DISABLED";
    FD1P3DX addr_space_4___i83 (.D(wb_odata[18]), .SP(dac_clk_p_c_enable_439), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[2] [18])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i83.GSR = "DISABLED";
    FD1P3DX addr_space_4___i82 (.D(wb_odata[17]), .SP(dac_clk_p_c_enable_439), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[2] [17])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i82.GSR = "DISABLED";
    FD1P3DX addr_space_4___i81 (.D(wb_odata[16]), .SP(dac_clk_p_c_enable_439), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[2] [16])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i81.GSR = "DISABLED";
    FD1P3DX addr_space_4___i80 (.D(wb_odata[15]), .SP(dac_clk_p_c_enable_439), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[2] [15])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i80.GSR = "DISABLED";
    FD1P3DX addr_space_4___i79 (.D(wb_odata[14]), .SP(dac_clk_p_c_enable_439), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[2] [14])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i79.GSR = "DISABLED";
    FD1P3DX addr_space_4___i78 (.D(wb_odata[13]), .SP(dac_clk_p_c_enable_439), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[2] [13])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i78.GSR = "DISABLED";
    FD1P3DX addr_space_4___i77 (.D(wb_odata[12]), .SP(dac_clk_p_c_enable_439), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[2] [12])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i77.GSR = "DISABLED";
    FD1P3DX addr_space_4___i76 (.D(wb_odata[11]), .SP(dac_clk_p_c_enable_439), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[2] [11])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i76.GSR = "DISABLED";
    FD1P3DX addr_space_4___i75 (.D(wb_odata[10]), .SP(dac_clk_p_c_enable_439), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[2] [10])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i75.GSR = "DISABLED";
    FD1P3DX addr_space_4___i74 (.D(wb_odata[9]), .SP(dac_clk_p_c_enable_439), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[2] [9])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i74.GSR = "DISABLED";
    FD1P3DX addr_space_4___i73 (.D(wb_odata[8]), .SP(dac_clk_p_c_enable_439), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[2] [8])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i73.GSR = "DISABLED";
    FD1P3DX addr_space_4___i72 (.D(wb_odata[7]), .SP(dac_clk_p_c_enable_439), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[2] [7])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i72.GSR = "DISABLED";
    FD1P3DX addr_space_4___i71 (.D(wb_odata[6]), .SP(dac_clk_p_c_enable_439), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[2] [6])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i71.GSR = "DISABLED";
    FD1P3DX addr_space_4___i70 (.D(wb_odata[5]), .SP(dac_clk_p_c_enable_439), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[2] [5])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i70.GSR = "DISABLED";
    FD1P3DX addr_space_4___i69 (.D(wb_odata[4]), .SP(dac_clk_p_c_enable_439), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[2] [4])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i69.GSR = "DISABLED";
    FD1P3DX addr_space_4___i68 (.D(wb_odata[3]), .SP(dac_clk_p_c_enable_439), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[2] [3])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i68.GSR = "DISABLED";
    FD1P3DX addr_space_4___i67 (.D(wb_odata[2]), .SP(dac_clk_p_c_enable_439), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[2] [2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i67.GSR = "DISABLED";
    FD1P3DX addr_space_4___i66 (.D(wb_odata[1]), .SP(dac_clk_p_c_enable_439), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[2] [1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i66.GSR = "DISABLED";
    FD1P3DX addr_space_4___i65 (.D(wb_odata[0]), .SP(dac_clk_p_c_enable_439), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[2] [0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i65.GSR = "DISABLED";
    FD1P3DX addr_space_4___i64 (.D(wb_odata[31]), .SP(dac_clk_p_c_enable_471), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[3] [31])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i64.GSR = "DISABLED";
    FD1P3DX addr_space_4___i63 (.D(wb_odata[30]), .SP(dac_clk_p_c_enable_471), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[3] [30])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i63.GSR = "DISABLED";
    FD1P3DX addr_space_4___i62 (.D(wb_odata[29]), .SP(dac_clk_p_c_enable_471), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[3] [29])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i62.GSR = "DISABLED";
    FD1P3DX addr_space_4___i61 (.D(wb_odata[28]), .SP(dac_clk_p_c_enable_471), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[3] [28])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i61.GSR = "DISABLED";
    FD1P3DX addr_space_4___i60 (.D(wb_odata[27]), .SP(dac_clk_p_c_enable_471), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[3] [27])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i60.GSR = "DISABLED";
    FD1P3DX addr_space_4___i59 (.D(wb_odata[26]), .SP(dac_clk_p_c_enable_471), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[3] [26])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i59.GSR = "DISABLED";
    FD1P3DX addr_space_4___i58 (.D(wb_odata[25]), .SP(dac_clk_p_c_enable_471), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[3] [25])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i58.GSR = "DISABLED";
    FD1P3DX addr_space_4___i57 (.D(wb_odata[24]), .SP(dac_clk_p_c_enable_471), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[3] [24])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i57.GSR = "DISABLED";
    FD1P3DX addr_space_4___i56 (.D(wb_odata[23]), .SP(dac_clk_p_c_enable_471), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[3] [23])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i56.GSR = "DISABLED";
    FD1P3DX addr_space_4___i55 (.D(wb_odata[22]), .SP(dac_clk_p_c_enable_471), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[3] [22])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i55.GSR = "DISABLED";
    FD1P3DX addr_space_4___i54 (.D(wb_odata[21]), .SP(dac_clk_p_c_enable_471), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[3] [21])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i54.GSR = "DISABLED";
    FD1P3DX addr_space_4___i53 (.D(wb_odata[20]), .SP(dac_clk_p_c_enable_471), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[3] [20])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i53.GSR = "DISABLED";
    FD1P3DX addr_space_4___i52 (.D(wb_odata[19]), .SP(dac_clk_p_c_enable_471), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[3] [19])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i52.GSR = "DISABLED";
    FD1P3DX addr_space_4___i51 (.D(wb_odata[18]), .SP(dac_clk_p_c_enable_471), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[3] [18])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i51.GSR = "DISABLED";
    FD1P3DX addr_space_4___i50 (.D(wb_odata[17]), .SP(dac_clk_p_c_enable_471), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[3] [17])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i50.GSR = "DISABLED";
    FD1P3DX addr_space_4___i49 (.D(wb_odata[16]), .SP(dac_clk_p_c_enable_471), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[3] [16])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i49.GSR = "DISABLED";
    FD1P3DX addr_space_4___i48 (.D(wb_odata[15]), .SP(dac_clk_p_c_enable_471), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[3] [15])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i48.GSR = "DISABLED";
    FD1P3DX addr_space_4___i47 (.D(wb_odata[14]), .SP(dac_clk_p_c_enable_471), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[3] [14])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i47.GSR = "DISABLED";
    FD1P3DX addr_space_4___i46 (.D(wb_odata[13]), .SP(dac_clk_p_c_enable_471), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[3] [13])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i46.GSR = "DISABLED";
    FD1P3BX addr_space_4___i45 (.D(wb_odata[12]), .SP(dac_clk_p_c_enable_471), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(\addr_space[3] [12])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i45.GSR = "DISABLED";
    FD1P3BX addr_space_4___i44 (.D(wb_odata[11]), .SP(dac_clk_p_c_enable_471), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(\addr_space[3] [11])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i44.GSR = "DISABLED";
    FD1P3BX addr_space_4___i43 (.D(wb_odata[10]), .SP(dac_clk_p_c_enable_471), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(\addr_space[3] [10])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i43.GSR = "DISABLED";
    FD1P3BX addr_space_4___i42 (.D(wb_odata[9]), .SP(dac_clk_p_c_enable_471), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(\addr_space[3] [9])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i42.GSR = "DISABLED";
    FD1P3BX addr_space_4___i41 (.D(wb_odata[8]), .SP(dac_clk_p_c_enable_471), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(\addr_space[3] [8])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i41.GSR = "DISABLED";
    FD1P3DX addr_space_4___i40 (.D(wb_odata[7]), .SP(dac_clk_p_c_enable_471), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[3] [7])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i40.GSR = "DISABLED";
    FD1P3BX addr_space_4___i39 (.D(wb_odata[6]), .SP(dac_clk_p_c_enable_471), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(\addr_space[3] [6])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i39.GSR = "DISABLED";
    FD1P3DX addr_space_4___i38 (.D(wb_odata[5]), .SP(dac_clk_p_c_enable_471), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[3] [5])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i38.GSR = "DISABLED";
    FD1P3DX addr_space_4___i37 (.D(wb_odata[4]), .SP(dac_clk_p_c_enable_471), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[3] [4])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i37.GSR = "DISABLED";
    FD1P3DX addr_space_4___i36 (.D(wb_odata[3]), .SP(dac_clk_p_c_enable_471), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[3] [3])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i36.GSR = "DISABLED";
    FD1P3DX addr_space_4___i35 (.D(wb_odata[2]), .SP(dac_clk_p_c_enable_471), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[3] [2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i35.GSR = "DISABLED";
    FD1P3DX addr_space_4___i34 (.D(wb_odata[1]), .SP(dac_clk_p_c_enable_471), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[3] [1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i34.GSR = "DISABLED";
    FD1P3DX addr_space_4___i33 (.D(wb_odata[0]), .SP(dac_clk_p_c_enable_471), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[3] [0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i33.GSR = "DISABLED";
    FD1P3DX addr_space_4___i32 (.D(wb_odata[31]), .SP(dac_clk_p_c_enable_502), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[4] [31])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i32.GSR = "DISABLED";
    FD1P3DX addr_space_4___i31 (.D(wb_odata[30]), .SP(dac_clk_p_c_enable_502), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[4] [30])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i31.GSR = "DISABLED";
    FD1P3DX addr_space_4___i30 (.D(wb_odata[29]), .SP(dac_clk_p_c_enable_502), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[4] [29])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i30.GSR = "DISABLED";
    FD1P3DX addr_space_4___i29 (.D(wb_odata[28]), .SP(dac_clk_p_c_enable_502), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[4] [28])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i29.GSR = "DISABLED";
    FD1P3DX addr_space_4___i28 (.D(wb_odata[27]), .SP(dac_clk_p_c_enable_502), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[4] [27])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i28.GSR = "DISABLED";
    FD1P3DX addr_space_4___i27 (.D(wb_odata[26]), .SP(dac_clk_p_c_enable_502), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[4] [26])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i27.GSR = "DISABLED";
    FD1P3DX addr_space_4___i26 (.D(wb_odata[25]), .SP(dac_clk_p_c_enable_502), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[4] [25])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i26.GSR = "DISABLED";
    FD1P3DX addr_space_4___i25 (.D(wb_odata[24]), .SP(dac_clk_p_c_enable_502), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[4] [24])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i25.GSR = "DISABLED";
    FD1P3DX addr_space_4___i24 (.D(wb_odata[23]), .SP(dac_clk_p_c_enable_502), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[4] [23])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i24.GSR = "DISABLED";
    FD1P3DX addr_space_4___i23 (.D(wb_odata[22]), .SP(dac_clk_p_c_enable_502), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[4] [22])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i23.GSR = "DISABLED";
    FD1P3DX addr_space_4___i22 (.D(wb_odata[21]), .SP(dac_clk_p_c_enable_502), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[4] [21])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i22.GSR = "DISABLED";
    FD1P3DX addr_space_4___i21 (.D(wb_odata[20]), .SP(dac_clk_p_c_enable_502), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[4] [20])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i21.GSR = "DISABLED";
    FD1P3DX addr_space_4___i20 (.D(wb_odata[19]), .SP(dac_clk_p_c_enable_502), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[4] [19])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i20.GSR = "DISABLED";
    FD1P3DX addr_space_4___i19 (.D(wb_odata[18]), .SP(dac_clk_p_c_enable_502), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[4] [18])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i19.GSR = "DISABLED";
    FD1P3DX addr_space_4___i18 (.D(wb_odata[17]), .SP(dac_clk_p_c_enable_502), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[4] [17])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i18.GSR = "DISABLED";
    FD1P3DX addr_space_4___i17 (.D(wb_odata[16]), .SP(dac_clk_p_c_enable_502), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[4] [16])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i17.GSR = "DISABLED";
    FD1P3DX addr_space_4___i16 (.D(wb_odata[15]), .SP(dac_clk_p_c_enable_502), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[4] [15])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i16.GSR = "DISABLED";
    FD1P3DX addr_space_4___i15 (.D(wb_odata[14]), .SP(dac_clk_p_c_enable_502), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[4] [14])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i15.GSR = "DISABLED";
    FD1P3DX addr_space_4___i14 (.D(wb_odata[13]), .SP(dac_clk_p_c_enable_502), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[4] [13])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i14.GSR = "DISABLED";
    FD1P3BX addr_space_4___i13 (.D(wb_odata[12]), .SP(dac_clk_p_c_enable_502), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(\addr_space[4] [12])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i13.GSR = "DISABLED";
    FD1P3BX addr_space_4___i12 (.D(wb_odata[11]), .SP(dac_clk_p_c_enable_502), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(\addr_space[4] [11])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i12.GSR = "DISABLED";
    FD1P3BX addr_space_4___i11 (.D(wb_odata[10]), .SP(dac_clk_p_c_enable_502), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(\addr_space[4] [10])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i11.GSR = "DISABLED";
    FD1P3BX addr_space_4___i10 (.D(wb_odata[9]), .SP(dac_clk_p_c_enable_502), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(\addr_space[4] [9])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i10.GSR = "DISABLED";
    FD1P3BX addr_space_4___i9 (.D(wb_odata[8]), .SP(dac_clk_p_c_enable_502), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(\addr_space[4] [8])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i9.GSR = "DISABLED";
    FD1P3DX addr_space_4___i8 (.D(wb_odata[7]), .SP(dac_clk_p_c_enable_502), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[4] [7])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i8.GSR = "DISABLED";
    FD1P3BX addr_space_4___i7 (.D(wb_odata[6]), .SP(dac_clk_p_c_enable_502), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(\addr_space[4] [6])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i7.GSR = "DISABLED";
    FD1P3DX addr_space_4___i6 (.D(wb_odata[5]), .SP(dac_clk_p_c_enable_502), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[4] [5])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i6.GSR = "DISABLED";
    FD1P3DX addr_space_4___i5 (.D(wb_odata[4]), .SP(dac_clk_p_c_enable_502), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[4] [4])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i5.GSR = "DISABLED";
    FD1P3DX addr_space_4___i4 (.D(wb_odata[3]), .SP(dac_clk_p_c_enable_502), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[4] [3])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i4.GSR = "DISABLED";
    FD1P3DX addr_space_4___i3 (.D(wb_odata[2]), .SP(dac_clk_p_c_enable_502), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[4] [2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i3.GSR = "DISABLED";
    FD1P3DX addr_space_4___i2 (.D(wb_odata[1]), .SP(dac_clk_p_c_enable_502), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(\addr_space[4] [1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(57[11] 61[5])
    defparam addr_space_4___i2.GSR = "DISABLED";
    LUT4 i24709_2_lut_rep_640 (.A(\wb_addr[0] ), .B(\wb_addr[1] ), .Z(n29300)) /* synthesis lut_function=(!(A+(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(59[4:25])
    defparam i24709_2_lut_rep_640.init = 16'h1111;
    LUT4 i1_2_lut_3_lut (.A(\wb_addr[0] ), .B(\wb_addr[1] ), .C(\wb_addr[2] ), 
         .Z(n21662)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(59[4:25])
    defparam i1_2_lut_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_rep_495_3_lut (.A(\wb_addr[0] ), .B(\wb_addr[1] ), .C(\wb_addr[2] ), 
         .Z(n29155)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(59[4:25])
    defparam i1_2_lut_rep_495_3_lut.init = 16'hefef;
    LUT4 i1295_1_lut (.A(o_dac_b[8]), .Z(o_dac_b[9])) /* synthesis lut_function=(!(A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(38[31:77])
    defparam i1295_1_lut.init = 16'h5555;
    LUT4 \addr_space_0[[30__bdd_3_lut_25275  (.A(\addr_space[1] [30]), .B(\addr_space[3] [30]), 
         .C(\wb_addr[1] ), .Z(n26956)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[30__bdd_3_lut_25275 .init = 16'hcaca;
    LUT4 \addr_space_0[[30__bdd_3_lut_25633  (.A(\addr_space[0] [30]), .B(\addr_space[2] [30]), 
         .C(\wb_addr[1] ), .Z(n26957)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[30__bdd_3_lut_25633 .init = 16'hcaca;
    LUT4 n27087_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4] [11]), .C(\wb_addr[2] ), 
         .D(n27087), .Z(o_wb_data_31__N_1104[11])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n27087_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 n27082_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4] [12]), .C(\wb_addr[2] ), 
         .D(n27082), .Z(o_wb_data_31__N_1104[12])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n27082_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 \addr_space_0[[29__bdd_3_lut_25279  (.A(\addr_space[1] [29]), .B(\addr_space[3] [29]), 
         .C(\wb_addr[1] ), .Z(n26961)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[29__bdd_3_lut_25279 .init = 16'hcaca;
    LUT4 \addr_space_0[[29__bdd_3_lut_25629  (.A(\addr_space[0] [29]), .B(\addr_space[2] [29]), 
         .C(\wb_addr[1] ), .Z(n26962)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[29__bdd_3_lut_25629 .init = 16'hcaca;
    LUT4 n27077_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4] [13]), .C(\wb_addr[2] ), 
         .D(n27077), .Z(o_wb_data_31__N_1104[13])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n27077_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 \addr_space_0[[28__bdd_3_lut_25621  (.A(\addr_space[0] [28]), .B(\addr_space[2] [28]), 
         .C(\wb_addr[1] ), .Z(n26972)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[28__bdd_3_lut_25621 .init = 16'hcaca;
    LUT4 \addr_space_0[[28__bdd_3_lut_25286  (.A(\addr_space[1] [28]), .B(\addr_space[3] [28]), 
         .C(\wb_addr[1] ), .Z(n26971)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[28__bdd_3_lut_25286 .init = 16'hcaca;
    LUT4 \addr_space_0[[27__bdd_3_lut_25617  (.A(\addr_space[0] [27]), .B(\addr_space[2] [27]), 
         .C(\wb_addr[1] ), .Z(n26982)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[27__bdd_3_lut_25617 .init = 16'hcaca;
    LUT4 \addr_space_0[[27__bdd_3_lut_25293  (.A(\addr_space[1] [27]), .B(\addr_space[3] [27]), 
         .C(\wb_addr[1] ), .Z(n26981)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[27__bdd_3_lut_25293 .init = 16'hcaca;
    LUT4 \addr_space_0[[26__bdd_3_lut_25297  (.A(\addr_space[1] [26]), .B(\addr_space[3] [26]), 
         .C(\wb_addr[1] ), .Z(n26986)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[26__bdd_3_lut_25297 .init = 16'hcaca;
    LUT4 \addr_space_0[[26__bdd_3_lut_25613  (.A(\addr_space[0] [26]), .B(\addr_space[2] [26]), 
         .C(\wb_addr[1] ), .Z(n26987)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[26__bdd_3_lut_25613 .init = 16'hcaca;
    LUT4 \addr_space_0[[25__bdd_3_lut_25609  (.A(\addr_space[0] [25]), .B(\addr_space[2] [25]), 
         .C(\wb_addr[1] ), .Z(n26997)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[25__bdd_3_lut_25609 .init = 16'hcaca;
    LUT4 \addr_space_0[[25__bdd_3_lut_25304  (.A(\addr_space[1] [25]), .B(\addr_space[3] [25]), 
         .C(\wb_addr[1] ), .Z(n26996)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[25__bdd_3_lut_25304 .init = 16'hcaca;
    LUT4 \addr_space_0[[0__bdd_3_lut_25308  (.A(\addr_space[1] [0]), .B(\addr_space[3] [0]), 
         .C(\wb_addr[1] ), .Z(n27001)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[0__bdd_3_lut_25308 .init = 16'hcaca;
    LUT4 \addr_space_0[[0__bdd_3_lut_25544  (.A(\addr_space[0] [0]), .B(\addr_space[2] [0]), 
         .C(\wb_addr[1] ), .Z(n27002)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[0__bdd_3_lut_25544 .init = 16'hcaca;
    LUT4 \addr_space_0[[24__bdd_3_lut_25312  (.A(\addr_space[1] [24]), .B(\addr_space[3] [24]), 
         .C(\wb_addr[1] ), .Z(n27006)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[24__bdd_3_lut_25312 .init = 16'hcaca;
    LUT4 n27069_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4] [14]), .C(\wb_addr[2] ), 
         .D(n27069), .Z(o_wb_data_31__N_1104[14])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n27069_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 n27064_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4] [15]), .C(\wb_addr[2] ), 
         .D(n27064), .Z(o_wb_data_31__N_1104[15])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n27064_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 n27059_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4] [16]), .C(\wb_addr[2] ), 
         .D(n27059), .Z(o_wb_data_31__N_1104[16])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n27059_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 \addr_space_0[[24__bdd_3_lut_25379  (.A(\addr_space[0] [24]), .B(\addr_space[2] [24]), 
         .C(\wb_addr[1] ), .Z(n27007)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[24__bdd_3_lut_25379 .init = 16'hcaca;
    LUT4 n27054_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4] [17]), .C(\wb_addr[2] ), 
         .D(n27054), .Z(o_wb_data_31__N_1104[17])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n27054_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 i1_2_lut_rep_795 (.A(\wb_addr[2] ), .B(\wb_addr[0] ), .Z(n29455)) /* synthesis lut_function=(A+!(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(59[4:25])
    defparam i1_2_lut_rep_795.init = 16'hbbbb;
    LUT4 n27049_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4] [18]), .C(\wb_addr[2] ), 
         .D(n27049), .Z(o_wb_data_31__N_1104[18])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n27049_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 n27044_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4] [19]), .C(\wb_addr[2] ), 
         .D(n27044), .Z(o_wb_data_31__N_1104[19])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n27044_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 n27039_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4] [20]), .C(\wb_addr[2] ), 
         .D(n27039), .Z(o_wb_data_31__N_1104[20])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n27039_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 n27034_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4] [21]), .C(\wb_addr[2] ), 
         .D(n27034), .Z(o_wb_data_31__N_1104[21])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n27034_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 n27029_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4] [22]), .C(\wb_addr[2] ), 
         .D(n27029), .Z(o_wb_data_31__N_1104[22])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n27029_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 i1_2_lut_rep_537_3_lut (.A(\wb_addr[2] ), .B(\wb_addr[0] ), .C(\wb_addr[1] ), 
         .Z(n29197)) /* synthesis lut_function=(A+!(B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(59[4:25])
    defparam i1_2_lut_rep_537_3_lut.init = 16'hbfbf;
    LUT4 n27024_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4] [23]), .C(\wb_addr[2] ), 
         .D(n27024), .Z(o_wb_data_31__N_1104[23])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n27024_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 i1_2_lut_rep_539_3_lut (.A(\wb_addr[2] ), .B(\wb_addr[0] ), .C(\wb_addr[1] ), 
         .Z(n29199)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(59[4:25])
    defparam i1_2_lut_rep_539_3_lut.init = 16'hfbfb;
    LUT4 n27008_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4] [24]), .C(\wb_addr[2] ), 
         .D(n27008), .Z(o_wb_data_31__N_1104[24])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n27008_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 n27003_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4] [0]), .C(\wb_addr[2] ), 
         .D(n27003), .Z(o_wb_data_31__N_1104[0])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n27003_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 n26998_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4] [25]), .C(\wb_addr[2] ), 
         .D(n26998), .Z(o_wb_data_31__N_1104[25])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n26998_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 n26988_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4] [26]), .C(\wb_addr[2] ), 
         .D(n26988), .Z(o_wb_data_31__N_1104[26])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n26988_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 n26983_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4] [27]), .C(\wb_addr[2] ), 
         .D(n26983), .Z(o_wb_data_31__N_1104[27])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n26983_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 n26973_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4] [28]), .C(\wb_addr[2] ), 
         .D(n26973), .Z(o_wb_data_31__N_1104[28])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n26973_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 n26963_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4] [29]), .C(\wb_addr[2] ), 
         .D(n26963), .Z(o_wb_data_31__N_1104[29])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n26963_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 i24576_4_lut (.A(n33[15]), .B(i_sw0_c), .C(cw_N_1500), .D(n33[10]), 
         .Z(dac_clk_p_c_enable_595)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C)))) */ ;
    defparam i24576_4_lut.init = 16'h3032;
    LUT4 i24574_3_lut (.A(n33[10]), .B(i_sw0_c), .C(cw_N_1500), .Z(dac_clk_p_c_enable_598)) /* synthesis lut_function=(!(A (B)+!A (B+!(C)))) */ ;
    defparam i24574_3_lut.init = 16'h3232;
    LUT4 \addr_space_0[[23__bdd_3_lut  (.A(\addr_space[0] [23]), .B(\addr_space[2] [23]), 
         .C(\wb_addr[1] ), .Z(n27023)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[23__bdd_3_lut .init = 16'hcaca;
    LUT4 \addr_space_0[[23__bdd_3_lut_25326  (.A(\addr_space[1] [23]), .B(\addr_space[3] [23]), 
         .C(\wb_addr[1] ), .Z(n27022)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[23__bdd_3_lut_25326 .init = 16'hcaca;
    CCU2D addr_space_0__30__I_0_32 (.A0(\addr_space[0] [30]), .B0(carrier_center_increment_offset[29]), 
          .C0(GND_net), .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n19398), .S0(carrier_increment_30__N_1296[30]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(119[24:82])
    defparam addr_space_0__30__I_0_32.INIT0 = 16'h5666;
    defparam addr_space_0__30__I_0_32.INIT1 = 16'h0000;
    defparam addr_space_0__30__I_0_32.INJECT1_0 = "NO";
    defparam addr_space_0__30__I_0_32.INJECT1_1 = "NO";
    LUT4 \addr_space_0[[22__bdd_3_lut_25330  (.A(\addr_space[1] [22]), .B(\addr_space[3] [22]), 
         .C(\wb_addr[1] ), .Z(n27027)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[22__bdd_3_lut_25330 .init = 16'hcaca;
    CCU2D addr_space_0__30__I_0_30 (.A0(\addr_space[0] [28]), .B0(carrier_center_increment_offset[28]), 
          .C0(GND_net), .D0(GND_net), .A1(\addr_space[0] [29]), .B1(carrier_center_increment_offset[29]), 
          .C1(GND_net), .D1(GND_net), .CIN(n19397), .COUT(n19398), .S0(carrier_increment_30__N_1296[28]), 
          .S1(carrier_increment_30__N_1296[29]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(119[24:82])
    defparam addr_space_0__30__I_0_30.INIT0 = 16'h5666;
    defparam addr_space_0__30__I_0_30.INIT1 = 16'h5666;
    defparam addr_space_0__30__I_0_30.INJECT1_0 = "NO";
    defparam addr_space_0__30__I_0_30.INJECT1_1 = "NO";
    LUT4 \addr_space_0[[22__bdd_3_lut  (.A(\addr_space[0] [22]), .B(\addr_space[2] [22]), 
         .C(\wb_addr[1] ), .Z(n27028)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[22__bdd_3_lut .init = 16'hcaca;
    LUT4 \addr_space_0[[21__bdd_3_lut_25334  (.A(\addr_space[1] [21]), .B(\addr_space[3] [21]), 
         .C(\wb_addr[1] ), .Z(n27032)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[21__bdd_3_lut_25334 .init = 16'hcaca;
    LUT4 \addr_space_0[[21__bdd_3_lut  (.A(\addr_space[0] [21]), .B(\addr_space[2] [21]), 
         .C(\wb_addr[1] ), .Z(n27033)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[21__bdd_3_lut .init = 16'hcaca;
    LUT4 \addr_space_0[[20__bdd_3_lut_25338  (.A(\addr_space[1] [20]), .B(\addr_space[3] [20]), 
         .C(\wb_addr[1] ), .Z(n27037)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[20__bdd_3_lut_25338 .init = 16'hcaca;
    LUT4 \addr_space_0[[20__bdd_3_lut  (.A(\addr_space[0] [20]), .B(\addr_space[2] [20]), 
         .C(\wb_addr[1] ), .Z(n27038)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[20__bdd_3_lut .init = 16'hcaca;
    LUT4 \addr_space_0[[19__bdd_3_lut_25342  (.A(\addr_space[1] [19]), .B(\addr_space[3] [19]), 
         .C(\wb_addr[1] ), .Z(n27042)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[19__bdd_3_lut_25342 .init = 16'hcaca;
    LUT4 \addr_space_0[[19__bdd_3_lut  (.A(\addr_space[0] [19]), .B(\addr_space[2] [19]), 
         .C(\wb_addr[1] ), .Z(n27043)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[19__bdd_3_lut .init = 16'hcaca;
    LUT4 \addr_space_0[[18__bdd_3_lut_25346  (.A(\addr_space[1] [18]), .B(\addr_space[3] [18]), 
         .C(\wb_addr[1] ), .Z(n27047)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[18__bdd_3_lut_25346 .init = 16'hcaca;
    LUT4 \addr_space_0[[18__bdd_3_lut  (.A(\addr_space[0] [18]), .B(\addr_space[2] [18]), 
         .C(\wb_addr[1] ), .Z(n27048)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[18__bdd_3_lut .init = 16'hcaca;
    LUT4 i11586_1_lut (.A(n33[15]), .Z(dac_clk_p_c_enable_617)) /* synthesis lut_function=(!(A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(155[21:41])
    defparam i11586_1_lut.init = 16'h5555;
    LUT4 \addr_space_0[[17__bdd_3_lut_25350  (.A(\addr_space[1] [17]), .B(\addr_space[3] [17]), 
         .C(\wb_addr[1] ), .Z(n27052)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[17__bdd_3_lut_25350 .init = 16'hcaca;
    LUT4 \addr_space_0[[17__bdd_3_lut  (.A(\addr_space[0] [17]), .B(\addr_space[2] [17]), 
         .C(\wb_addr[1] ), .Z(n27053)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[17__bdd_3_lut .init = 16'hcaca;
    CCU2D addr_space_0__30__I_0_28 (.A0(\addr_space[0] [26]), .B0(carrier_center_increment_offset[26]), 
          .C0(GND_net), .D0(GND_net), .A1(\addr_space[0] [27]), .B1(carrier_center_increment_offset[27]), 
          .C1(GND_net), .D1(GND_net), .CIN(n19396), .COUT(n19397), .S0(carrier_increment_30__N_1296[26]), 
          .S1(carrier_increment_30__N_1296[27]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(119[24:82])
    defparam addr_space_0__30__I_0_28.INIT0 = 16'h5666;
    defparam addr_space_0__30__I_0_28.INIT1 = 16'h5666;
    defparam addr_space_0__30__I_0_28.INJECT1_0 = "NO";
    defparam addr_space_0__30__I_0_28.INJECT1_1 = "NO";
    LUT4 \addr_space_0[[16__bdd_3_lut_25354  (.A(\addr_space[1] [16]), .B(\addr_space[3] [16]), 
         .C(\wb_addr[1] ), .Z(n27057)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[16__bdd_3_lut_25354 .init = 16'hcaca;
    LUT4 \addr_space_0[[16__bdd_3_lut  (.A(\addr_space[0] [16]), .B(\addr_space[2] [16]), 
         .C(\wb_addr[1] ), .Z(n27058)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[16__bdd_3_lut .init = 16'hcaca;
    LUT4 \addr_space_0[[15__bdd_3_lut_25358  (.A(\addr_space[1] [15]), .B(\addr_space[3] [15]), 
         .C(\wb_addr[1] ), .Z(n27062)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[15__bdd_3_lut_25358 .init = 16'hcaca;
    LUT4 \addr_space_0[[15__bdd_3_lut  (.A(\addr_space[0] [15]), .B(\addr_space[2] [15]), 
         .C(\wb_addr[1] ), .Z(n27063)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[15__bdd_3_lut .init = 16'hcaca;
    LUT4 n26958_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4] [30]), .C(\wb_addr[2] ), 
         .D(n26958), .Z(o_wb_data_31__N_1104[30])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n26958_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 \addr_space_0[[14__bdd_3_lut_25362  (.A(\addr_space[1] [14]), .B(\addr_space[3] [14]), 
         .C(\wb_addr[1] ), .Z(n27067)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[14__bdd_3_lut_25362 .init = 16'hcaca;
    LUT4 \addr_space_0[[14__bdd_3_lut  (.A(\addr_space[0] [14]), .B(\addr_space[2] [14]), 
         .C(\wb_addr[1] ), .Z(n27068)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[14__bdd_3_lut .init = 16'hcaca;
    LUT4 cw_I_0_1_lut (.A(cw), .Z(o_dac_cw_b_c)) /* synthesis lut_function=(!(A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(124[17:20])
    defparam cw_I_0_1_lut.init = 16'h5555;
    FD1P3AX cw_mux_dac_a_mux_sel_54 (.D(cw_N_1500), .SP(dac_clk_p_c_enable_595), 
            .CK(dac_clk_p_c), .Q(cw_mux_dac_a_mux_sel)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(145[11] 157[5])
    defparam cw_mux_dac_a_mux_sel_54.GSR = "DISABLED";
    FD1P3AX cw_53 (.D(cw_N_1500), .SP(dac_clk_p_c_enable_598), .CK(dac_clk_p_c), 
            .Q(cw)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=122, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(145[11] 157[5])
    defparam cw_53.GSR = "DISABLED";
    LUT4 i866_1_lut_rep_741 (.A(i_sw0_c), .Z(dac_clk_p_c_enable_630)) /* synthesis lut_function=(!(A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(31[12:17])
    defparam i866_1_lut_rep_741.init = 16'h5555;
    LUT4 i7237_2_lut_2_lut (.A(i_sw0_c), .B(u_s[2]), .Z(n9468)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(31[12:17])
    defparam i7237_2_lut_2_lut.init = 16'h4444;
    LUT4 i7213_2_lut_2_lut (.A(i_sw0_c), .B(u_s_adj_3684[12]), .Z(n9444)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(31[12:17])
    defparam i7213_2_lut_2_lut.init = 16'h4444;
    LUT4 i7215_2_lut_2_lut (.A(i_sw0_c), .B(u_s_adj_3684[10]), .Z(n9446)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(31[12:17])
    defparam i7215_2_lut_2_lut.init = 16'h4444;
    LUT4 i7217_2_lut_2_lut (.A(i_sw0_c), .B(u_s_adj_3684[8]), .Z(n9448)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(31[12:17])
    defparam i7217_2_lut_2_lut.init = 16'h4444;
    LUT4 i7219_2_lut_2_lut (.A(i_sw0_c), .B(u_s_adj_3684[6]), .Z(n9450)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(31[12:17])
    defparam i7219_2_lut_2_lut.init = 16'h4444;
    LUT4 n26953_bdd_3_lut_4_lut (.A(n29300), .B(\addr_space[4] [31]), .C(\wb_addr[2] ), 
         .D(n26953), .Z(o_wb_data_31__N_1104[31])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam n26953_bdd_3_lut_4_lut.init = 16'h8f80;
    LUT4 i7221_2_lut_2_lut (.A(i_sw0_c), .B(u_s_adj_3684[4]), .Z(n9452)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(31[12:17])
    defparam i7221_2_lut_2_lut.init = 16'h4444;
    LUT4 i7223_2_lut_2_lut (.A(i_sw0_c), .B(u_s_adj_3684[2]), .Z(n9454)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(31[12:17])
    defparam i7223_2_lut_2_lut.init = 16'h4444;
    LUT4 i7227_2_lut_2_lut (.A(i_sw0_c), .B(u_s[12]), .Z(n9458)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(31[12:17])
    defparam i7227_2_lut_2_lut.init = 16'h4444;
    LUT4 i7229_2_lut_2_lut (.A(i_sw0_c), .B(u_s[10]), .Z(n9460)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(31[12:17])
    defparam i7229_2_lut_2_lut.init = 16'h4444;
    LUT4 i7231_2_lut_2_lut (.A(i_sw0_c), .B(u_s[8]), .Z(n9462)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(31[12:17])
    defparam i7231_2_lut_2_lut.init = 16'h4444;
    LUT4 i7233_2_lut_2_lut (.A(i_sw0_c), .B(u_s[6]), .Z(n9464)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(31[12:17])
    defparam i7233_2_lut_2_lut.init = 16'h4444;
    LUT4 i7235_2_lut_2_lut (.A(i_sw0_c), .B(u_s[4]), .Z(n9466)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(31[12:17])
    defparam i7235_2_lut_2_lut.init = 16'h4444;
    LUT4 i7259_2_lut_2_lut (.A(i_sw0_c), .B(u_s_adj_3685[12]), .Z(n9490)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(31[12:17])
    defparam i7259_2_lut_2_lut.init = 16'h4444;
    LUT4 i7261_2_lut_2_lut (.A(i_sw0_c), .B(u_s_adj_3685[10]), .Z(n9492)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(31[12:17])
    defparam i7261_2_lut_2_lut.init = 16'h4444;
    CCU2D addr_space_0__30__I_0_26 (.A0(\addr_space[0] [24]), .B0(carrier_center_increment_offset[24]), 
          .C0(GND_net), .D0(GND_net), .A1(\addr_space[0] [25]), .B1(carrier_center_increment_offset[25]), 
          .C1(GND_net), .D1(GND_net), .CIN(n19395), .COUT(n19396), .S0(carrier_increment_30__N_1296[24]), 
          .S1(carrier_increment_30__N_1296[25]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(119[24:82])
    defparam addr_space_0__30__I_0_26.INIT0 = 16'h5666;
    defparam addr_space_0__30__I_0_26.INIT1 = 16'h5666;
    defparam addr_space_0__30__I_0_26.INJECT1_0 = "NO";
    defparam addr_space_0__30__I_0_26.INJECT1_1 = "NO";
    LUT4 i7263_2_lut_2_lut (.A(i_sw0_c), .B(u_s_adj_3685[8]), .Z(n9494)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(31[12:17])
    defparam i7263_2_lut_2_lut.init = 16'h4444;
    LUT4 i7265_2_lut_2_lut (.A(i_sw0_c), .B(u_s_adj_3685[6]), .Z(n9496)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(31[12:17])
    defparam i7265_2_lut_2_lut.init = 16'h4444;
    CCU2D addr_space_0__30__I_0_24 (.A0(\addr_space[0] [22]), .B0(carrier_center_increment_offset[22]), 
          .C0(GND_net), .D0(GND_net), .A1(\addr_space[0] [23]), .B1(carrier_center_increment_offset[23]), 
          .C1(GND_net), .D1(GND_net), .CIN(n19394), .COUT(n19395), .S0(carrier_increment_30__N_1296[22]), 
          .S1(carrier_increment_30__N_1296[23]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(119[24:82])
    defparam addr_space_0__30__I_0_24.INIT0 = 16'h5666;
    defparam addr_space_0__30__I_0_24.INIT1 = 16'h5666;
    defparam addr_space_0__30__I_0_24.INJECT1_0 = "NO";
    defparam addr_space_0__30__I_0_24.INJECT1_1 = "NO";
    LUT4 i7267_2_lut_2_lut (.A(i_sw0_c), .B(u_s_adj_3685[4]), .Z(n9498)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(31[12:17])
    defparam i7267_2_lut_2_lut.init = 16'h4444;
    LUT4 i7273_2_lut_2_lut (.A(i_sw0_c), .B(u_s_adj_3685[2]), .Z(n9504)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(31[12:17])
    defparam i7273_2_lut_2_lut.init = 16'h4444;
    LUT4 i7275_2_lut_2_lut (.A(i_sw0_c), .B(u_s_adj_3685[0]), .Z(n9506)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(31[12:17])
    defparam i7275_2_lut_2_lut.init = 16'h4444;
    LUT4 i7257_2_lut_2_lut (.A(i_sw0_c), .B(u_s[0]), .Z(n9488)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(31[12:17])
    defparam i7257_2_lut_2_lut.init = 16'h4444;
    LUT4 i7225_2_lut_2_lut (.A(i_sw0_c), .B(u_s_adj_3684[0]), .Z(n9456)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(31[12:17])
    defparam i7225_2_lut_2_lut.init = 16'h4444;
    LUT4 \addr_space_0[[13__bdd_3_lut_25368  (.A(\addr_space[1] [13]), .B(\addr_space[3] [13]), 
         .C(\wb_addr[1] ), .Z(n27075)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[13__bdd_3_lut_25368 .init = 16'hcaca;
    LUT4 \addr_space_0[[13__bdd_3_lut  (.A(\addr_space[0] [13]), .B(\addr_space[2] [13]), 
         .C(\wb_addr[1] ), .Z(n27076)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[13__bdd_3_lut .init = 16'hcaca;
    FD1P3DX startup_timer_FSM_i0_i15 (.D(n32067), .SP(n694[14]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(n33[15]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(155[21:41])
    defparam startup_timer_FSM_i0_i15.GSR = "DISABLED";
    FD1P3DX startup_timer_FSM_i0_i14 (.D(n694[13]), .SP(dac_clk_p_c_enable_617), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(n694[14]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(155[21:41])
    defparam startup_timer_FSM_i0_i14.GSR = "DISABLED";
    FD1P3DX startup_timer_FSM_i0_i13 (.D(n694[12]), .SP(dac_clk_p_c_enable_617), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(n694[13]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(155[21:41])
    defparam startup_timer_FSM_i0_i13.GSR = "DISABLED";
    LUT4 \addr_space_0[[12__bdd_3_lut_25372  (.A(\addr_space[1] [12]), .B(\addr_space[3] [12]), 
         .C(\wb_addr[1] ), .Z(n27080)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[12__bdd_3_lut_25372 .init = 16'hcaca;
    FD1P3DX startup_timer_FSM_i0_i12 (.D(n694[11]), .SP(dac_clk_p_c_enable_617), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(n694[12]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(155[21:41])
    defparam startup_timer_FSM_i0_i12.GSR = "DISABLED";
    FD1P3DX startup_timer_FSM_i0_i11 (.D(n33[10]), .SP(dac_clk_p_c_enable_617), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(n694[11]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(155[21:41])
    defparam startup_timer_FSM_i0_i11.GSR = "DISABLED";
    FD1P3DX startup_timer_FSM_i0_i10 (.D(n694[9]), .SP(dac_clk_p_c_enable_617), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(n33[10]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(155[21:41])
    defparam startup_timer_FSM_i0_i10.GSR = "DISABLED";
    FD1P3DX startup_timer_FSM_i0_i9 (.D(n694[8]), .SP(dac_clk_p_c_enable_617), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(n694[9]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(155[21:41])
    defparam startup_timer_FSM_i0_i9.GSR = "DISABLED";
    FD1P3DX startup_timer_FSM_i0_i8 (.D(n694[7]), .SP(dac_clk_p_c_enable_617), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(n694[8]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(155[21:41])
    defparam startup_timer_FSM_i0_i8.GSR = "DISABLED";
    LUT4 \addr_space_0[[12__bdd_3_lut  (.A(\addr_space[0] [12]), .B(\addr_space[2] [12]), 
         .C(\wb_addr[1] ), .Z(n27081)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[12__bdd_3_lut .init = 16'hcaca;
    FD1P3DX startup_timer_FSM_i0_i7 (.D(n694[6]), .SP(dac_clk_p_c_enable_617), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(n694[7]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(155[21:41])
    defparam startup_timer_FSM_i0_i7.GSR = "DISABLED";
    FD1P3DX startup_timer_FSM_i0_i6 (.D(n694[5]), .SP(dac_clk_p_c_enable_617), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(n694[6]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(155[21:41])
    defparam startup_timer_FSM_i0_i6.GSR = "DISABLED";
    FD1P3DX startup_timer_FSM_i0_i5 (.D(n694[4]), .SP(dac_clk_p_c_enable_617), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(n694[5]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(155[21:41])
    defparam startup_timer_FSM_i0_i5.GSR = "DISABLED";
    FD1P3DX startup_timer_FSM_i0_i4 (.D(cw_N_1500), .SP(dac_clk_p_c_enable_617), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(n694[4]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(155[21:41])
    defparam startup_timer_FSM_i0_i4.GSR = "DISABLED";
    FD1P3DX startup_timer_FSM_i0_i3 (.D(n694[2]), .SP(dac_clk_p_c_enable_617), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(cw_N_1500));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(155[21:41])
    defparam startup_timer_FSM_i0_i3.GSR = "DISABLED";
    FD1P3DX startup_timer_FSM_i0_i2 (.D(n694[1]), .SP(dac_clk_p_c_enable_617), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(n694[2]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(155[21:41])
    defparam startup_timer_FSM_i0_i2.GSR = "DISABLED";
    FD1P3DX startup_timer_FSM_i0_i1 (.D(n694[0]), .SP(dac_clk_p_c_enable_617), 
            .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(n694[1]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(155[21:41])
    defparam startup_timer_FSM_i0_i1.GSR = "DISABLED";
    CCU2D addr_space_0__30__I_0_22 (.A0(\addr_space[0] [20]), .B0(carrier_center_increment_offset[20]), 
          .C0(GND_net), .D0(GND_net), .A1(\addr_space[0] [21]), .B1(carrier_center_increment_offset[21]), 
          .C1(GND_net), .D1(GND_net), .CIN(n19393), .COUT(n19394), .S0(carrier_increment_30__N_1296[20]), 
          .S1(carrier_increment_30__N_1296[21]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(119[24:82])
    defparam addr_space_0__30__I_0_22.INIT0 = 16'h5666;
    defparam addr_space_0__30__I_0_22.INIT1 = 16'h5666;
    defparam addr_space_0__30__I_0_22.INJECT1_0 = "NO";
    defparam addr_space_0__30__I_0_22.INJECT1_1 = "NO";
    LUT4 \addr_space_0[[11__bdd_3_lut_25376  (.A(\addr_space[1] [11]), .B(\addr_space[3] [11]), 
         .C(\wb_addr[1] ), .Z(n27085)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[11__bdd_3_lut_25376 .init = 16'hcaca;
    LUT4 \addr_space_0[[11__bdd_3_lut  (.A(\addr_space[0] [11]), .B(\addr_space[2] [11]), 
         .C(\wb_addr[1] ), .Z(n27086)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[11__bdd_3_lut .init = 16'hcaca;
    LUT4 \addr_space_0[[10__bdd_3_lut  (.A(\addr_space[0] [10]), .B(\addr_space[2] [10]), 
         .C(\wb_addr[1] ), .Z(n27104)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[10__bdd_3_lut .init = 16'hcaca;
    LUT4 \addr_space_0[[10__bdd_3_lut_25395  (.A(\addr_space[1] [10]), .B(\addr_space[3] [10]), 
         .C(\wb_addr[1] ), .Z(n27103)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam \addr_space_0[[10__bdd_3_lut_25395 .init = 16'hcaca;
    PFUMX i25572 (.BLUT(n27298), .ALUT(n27297), .C0(\wb_addr[0] ), .Z(n27299));
    PFUMX i25554 (.BLUT(n27278), .ALUT(n27277), .C0(\wb_addr[0] ), .Z(n27279));
    PFUMX i25550 (.BLUT(n27273), .ALUT(n27272), .C0(\wb_addr[0] ), .Z(n27274));
    PFUMX i25533 (.BLUT(n27251), .ALUT(n27250), .C0(\wb_addr[0] ), .Z(n27252));
    PFUMX i25523 (.BLUT(n27238), .ALUT(n27237), .C0(\wb_addr[0] ), .Z(n27239));
    PFUMX i25511 (.BLUT(n27226), .ALUT(n27225), .C0(\wb_addr[0] ), .Z(n27227));
    PFUMX i25497 (.BLUT(n27211), .ALUT(n27210), .C0(\wb_addr[0] ), .Z(n27212));
    PFUMX i25493 (.BLUT(n27204), .ALUT(n27203), .C0(\wb_addr[0] ), .Z(n27205));
    sgnmpy_14x16 q_gain_multiplier (.u_s({Open_34, Open_35, Open_36, Open_37, 
            Open_38, Open_39, Open_40, Open_41, Open_42, Open_43, 
            Open_44, Open_45, Open_46, u_s[0]}), .dac_clk_p_c(dac_clk_p_c), 
            .i_sw0_c(i_sw0_c), .\o_dac_b[0] (o_dac_b[0]), .\addr_space[4][13] (\addr_space[4] [13]), 
            .o_sample_q({o_sample_q}), .GND_net(GND_net), .\addr_space[4][12] (\addr_space[4] [12]), 
            .\addr_space[4][10] (\addr_space[4] [10]), .\addr_space[4][11] (\addr_space[4] [11]), 
            .\addr_space[4][8] (\addr_space[4] [8]), .\addr_space[4][9] (\addr_space[4] [9]), 
            .\addr_space[4][6] (\addr_space[4] [6]), .\addr_space[4][7] (\addr_space[4] [7]), 
            .\addr_space[4][4] (\addr_space[4] [4]), .\addr_space[4][5] (\addr_space[4] [5]), 
            .\addr_space[4][2] (\addr_space[4] [2]), .\addr_space[4][3] (\addr_space[4] [3]), 
            .\addr_space[4][0] (\addr_space[4] [0]), .\addr_space[4][1] (\addr_space[4] [1]), 
            .\o_dac_b[8] (o_dac_b[8]), .\o_dac_b[7] (o_dac_b[7]), .\o_dac_b[6] (o_dac_b[6]), 
            .\o_dac_b[5] (o_dac_b[5]), .\o_dac_b[4] (o_dac_b[4]), .\o_dac_b[3] (o_dac_b[3]), 
            .\o_dac_b[2] (o_dac_b[2]), .\o_dac_b[1] (o_dac_b[1]), .\u_s[12] (u_s[12]), 
            .\u_s[10] (u_s[10]), .\u_s[8] (u_s[8]), .\u_s[6] (u_s[6]), 
            .\u_s[4] (u_s[4]), .\u_s[2] (u_s[2]), .n9458(n9458), .n9460(n9460), 
            .n9462(n9462), .n9464(n9464), .n9466(n9466), .n9468(n9468), 
            .n9488(n9488)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(109[14:99])
    sgnmpy_14x16_U24 modulation_amplitude_multiplier (.u_s({Open_47, Open_48, 
            Open_49, Open_50, Open_51, Open_52, Open_53, Open_54, 
            Open_55, Open_56, Open_57, Open_58, Open_59, u_s_adj_3684[0]}), 
            .dac_clk_p_c(dac_clk_p_c), .i_sw0_c(i_sw0_c), .carrier_center_increment_offset({carrier_center_increment_offset}), 
            .GND_net(GND_net), .\addr_space[2][13] (\addr_space[2] [13]), 
            .modulation_output({modulation_output}), .\addr_space[2][12] (\addr_space[2] [12]), 
            .\addr_space[2][10] (\addr_space[2] [10]), .\addr_space[2][11] (\addr_space[2] [11]), 
            .\addr_space[2][8] (\addr_space[2] [8]), .\addr_space[2][9] (\addr_space[2] [9]), 
            .\addr_space[2][6] (\addr_space[2] [6]), .\addr_space[2][7] (\addr_space[2] [7]), 
            .\addr_space[2][4] (\addr_space[2] [4]), .\addr_space[2][5] (\addr_space[2] [5]), 
            .\addr_space[2][2] (\addr_space[2] [2]), .\addr_space[2][3] (\addr_space[2] [3]), 
            .\addr_space[2][0] (\addr_space[2] [0]), .\addr_space[2][1] (\addr_space[2] [1]), 
            .\u_s[12] (u_s_adj_3684[12]), .\u_s[10] (u_s_adj_3684[10]), 
            .\u_s[8] (u_s_adj_3684[8]), .\u_s[6] (u_s_adj_3684[6]), .\u_s[4] (u_s_adj_3684[4]), 
            .\u_s[2] (u_s_adj_3684[2]), .n9444(n9444), .n9446(n9446), 
            .n9448(n9448), .n9450(n9450), .n9452(n9452), .n9454(n9454), 
            .n9456(n9456)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(113[14:154])
    dds modulation (.dac_clk_p_c(dac_clk_p_c), .i_sw0_c(i_sw0_c), .\addr_space[1][0] (\addr_space[1] [0]), 
        .\addr_space[1][30] (\addr_space[1] [30]), .\addr_space[1][29] (\addr_space[1] [29]), 
        .\addr_space[1][28] (\addr_space[1] [28]), .\addr_space[1][27] (\addr_space[1] [27]), 
        .\addr_space[1][26] (\addr_space[1] [26]), .\addr_space[1][25] (\addr_space[1] [25]), 
        .\addr_space[1][24] (\addr_space[1] [24]), .\addr_space[1][23] (\addr_space[1] [23]), 
        .\addr_space[1][22] (\addr_space[1] [22]), .\addr_space[1][21] (\addr_space[1] [21]), 
        .\addr_space[1][20] (\addr_space[1] [20]), .\addr_space[1][19] (\addr_space[1] [19]), 
        .\addr_space[1][18] (\addr_space[1] [18]), .\addr_space[1][17] (\addr_space[1] [17]), 
        .\addr_space[1][16] (\addr_space[1] [16]), .\addr_space[1][15] (\addr_space[1] [15]), 
        .\addr_space[1][14] (\addr_space[1] [14]), .\addr_space[1][13] (\addr_space[1] [13]), 
        .\addr_space[1][12] (\addr_space[1] [12]), .\addr_space[1][11] (\addr_space[1] [11]), 
        .\addr_space[1][10] (\addr_space[1] [10]), .\addr_space[1][9] (\addr_space[1] [9]), 
        .\addr_space[1][8] (\addr_space[1] [8]), .\addr_space[1][7] (\addr_space[1] [7]), 
        .\addr_space[1][6] (\addr_space[1] [6]), .\addr_space[1][5] (\addr_space[1] [5]), 
        .\addr_space[1][4] (\addr_space[1] [4]), .\addr_space[1][3] (\addr_space[1] [3]), 
        .\addr_space[1][2] (\addr_space[1] [2]), .\addr_space[1][1] (\addr_space[1] [1]), 
        .dac_clk_p_c_enable_630(dac_clk_p_c_enable_630), .modulation_output({modulation_output}), 
        .\quarter_wave_sample_register_i[15] (quarter_wave_sample_register_i[15]), 
        .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(96[4:161])
    sgnmpy_14x16_U25 i_gain_multiplier (.dac_clk_p_c(dac_clk_p_c), .i_sw0_c(i_sw0_c), 
            .\o_sample_dc_offset_i[7] (o_sample_dc_offset_i[7]), .u_s({Open_60, 
            Open_61, Open_62, Open_63, Open_64, Open_65, Open_66, 
            Open_67, Open_68, Open_69, Open_70, Open_71, Open_72, 
            u_s_adj_3685[0]}), .\addr_space[3][13] (\addr_space[3] [13]), 
            .o_sample_i({o_sample_i}), .GND_net(GND_net), .\u_s[12] (u_s_adj_3685[12]), 
            .\u_s[10] (u_s_adj_3685[10]), .\u_s[8] (u_s_adj_3685[8]), .\u_s[6] (u_s_adj_3685[6]), 
            .\u_s[4] (u_s_adj_3685[4]), .\u_s[2] (u_s_adj_3685[2]), .\addr_space[3][12] (\addr_space[3] [12]), 
            .\addr_space[3][10] (\addr_space[3] [10]), .\addr_space[3][11] (\addr_space[3] [11]), 
            .\addr_space[3][8] (\addr_space[3] [8]), .\addr_space[3][9] (\addr_space[3] [9]), 
            .\addr_space[3][6] (\addr_space[3] [6]), .\addr_space[3][7] (\addr_space[3] [7]), 
            .\addr_space[3][4] (\addr_space[3] [4]), .\addr_space[3][5] (\addr_space[3] [5]), 
            .\addr_space[3][2] (\addr_space[3] [2]), .\addr_space[3][3] (\addr_space[3] [3]), 
            .\addr_space[3][0] (\addr_space[3] [0]), .\addr_space[3][1] (\addr_space[3] [1]), 
            .\o_sample_dc_offset_i[15] (o_sample_dc_offset_i[15]), .\o_sample_dc_offset_i[14] (o_sample_dc_offset_i[14]), 
            .\o_sample_dc_offset_i[13] (o_sample_dc_offset_i[13]), .\o_sample_dc_offset_i[12] (o_sample_dc_offset_i[12]), 
            .\o_sample_dc_offset_i[11] (o_sample_dc_offset_i[11]), .\o_sample_dc_offset_i[10] (o_sample_dc_offset_i[10]), 
            .\o_sample_dc_offset_i[9] (o_sample_dc_offset_i[9]), .\o_sample_dc_offset_i[8] (o_sample_dc_offset_i[8]), 
            .n9490(n9490), .n9492(n9492), .n9494(n9494), .n9496(n9496), 
            .n9498(n9498), .n9504(n9504), .n9506(n9506)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(108[14:99])
    dds_U26 carrier (.dac_clk_p_c(dac_clk_p_c), .i_sw0_c(i_sw0_c), .carrier_increment({carrier_increment}), 
            .GND_net(GND_net), .dac_clk_p_c_enable_630(dac_clk_p_c_enable_630), 
            .o_sample_q({o_sample_q}), .o_sample_i({o_sample_i}), .\quarter_wave_sample_register_i[15] (quarter_wave_sample_register_i[15]), 
            .n32066(n32066)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(91[4:158])
    
endmodule
//
// Verilog Description of module sgnmpy_14x16
//

module sgnmpy_14x16 (u_s, dac_clk_p_c, i_sw0_c, \o_dac_b[0] , \addr_space[4][13] , 
            o_sample_q, GND_net, \addr_space[4][12] , \addr_space[4][10] , 
            \addr_space[4][11] , \addr_space[4][8] , \addr_space[4][9] , 
            \addr_space[4][6] , \addr_space[4][7] , \addr_space[4][4] , 
            \addr_space[4][5] , \addr_space[4][2] , \addr_space[4][3] , 
            \addr_space[4][0] , \addr_space[4][1] , \o_dac_b[8] , \o_dac_b[7] , 
            \o_dac_b[6] , \o_dac_b[5] , \o_dac_b[4] , \o_dac_b[3] , 
            \o_dac_b[2] , \o_dac_b[1] , \u_s[12] , \u_s[10] , \u_s[8] , 
            \u_s[6] , \u_s[4] , \u_s[2] , n9458, n9460, n9462, n9464, 
            n9466, n9468, n9488) /* synthesis syn_module_defined=1 */ ;
    output [13:0]u_s;
    input dac_clk_p_c;
    input i_sw0_c;
    output \o_dac_b[0] ;
    input \addr_space[4][13] ;
    input [15:0]o_sample_q;
    input GND_net;
    input \addr_space[4][12] ;
    input \addr_space[4][10] ;
    input \addr_space[4][11] ;
    input \addr_space[4][8] ;
    input \addr_space[4][9] ;
    input \addr_space[4][6] ;
    input \addr_space[4][7] ;
    input \addr_space[4][4] ;
    input \addr_space[4][5] ;
    input \addr_space[4][2] ;
    input \addr_space[4][3] ;
    input \addr_space[4][0] ;
    input \addr_space[4][1] ;
    output \o_dac_b[8] ;
    output \o_dac_b[7] ;
    output \o_dac_b[6] ;
    output \o_dac_b[5] ;
    output \o_dac_b[4] ;
    output \o_dac_b[3] ;
    output \o_dac_b[2] ;
    output \o_dac_b[1] ;
    output \u_s[12] ;
    output \u_s[10] ;
    output \u_s[8] ;
    output \u_s[6] ;
    output \u_s[4] ;
    output \u_s[2] ;
    input n9458;
    input n9460;
    input n9462;
    input n9464;
    input n9466;
    input n9468;
    input n9488;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[29:38])
    wire [15:0]o_sample_q_c /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(30[51:61])
    wire [13:0]u_s_13__N_1951;
    wire [15:0]u_l;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(62[18:21])
    wire [15:0]u_l_15__N_1965;
    wire [4:0]u_sgn;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(63[19:24])
    wire [4:0]u_sgn_4__N_1981;
    wire [29:0]o_p_29__N_1986;
    wire [29:0]u_r;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(93[21:24])
    wire [29:0]n215;
    
    wire n14230, n19801, n19800, n19799, n19798, n19797, n19796, 
        n19795, n19794, n19793, n19792, n19791, n19790, n19789, 
        n19788, n19623, n19622, n19621, n19620, n19619, n19618, 
        n19617, n19616, n19615, n19614, n19613, n19612, n19611, 
        n19610, n19609;
    wire [13:0]u_s_c;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(61[18:21])
    
    FD1S3IX u_s__i0 (.D(u_s_13__N_1951[0]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_s[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=109, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_s__i0.GSR = "DISABLED";
    FD1S3IX u_l__i0 (.D(u_l_15__N_1965[0]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_l[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=109, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_l__i0.GSR = "DISABLED";
    FD1S3IX u_sgn__i0 (.D(u_sgn_4__N_1981[0]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_sgn[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=109, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(87[9] 91[60])
    defparam u_sgn__i0.GSR = "DISABLED";
    FD1S3IX o_p__i1 (.D(o_p_29__N_1986[21]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_dac_b[0] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=109, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(98[9] 102[36])
    defparam o_p__i1.GSR = "DISABLED";
    LUT4 i17_2_lut (.A(\addr_space[4][13] ), .B(o_sample_q[15]), .Z(u_sgn_4__N_1981[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(91[32:57])
    defparam i17_2_lut.init = 16'h6666;
    LUT4 mux_644_i1_3_lut (.A(u_r[21]), .B(n215[21]), .C(u_sgn[4]), .Z(o_p_29__N_1986[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[10:35])
    defparam mux_644_i1_3_lut.init = 16'hcaca;
    LUT4 i11854_1_lut (.A(u_l[0]), .Z(n14230)) /* synthesis lut_function=(!(A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam i11854_1_lut.init = 16'h5555;
    CCU2D add_537_29 (.A0(u_r[28]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(u_r[29]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19801), 
          .S0(n215[28]), .S1(n215[29]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[25:31])
    defparam add_537_29.INIT0 = 16'hf555;
    defparam add_537_29.INIT1 = 16'hf555;
    defparam add_537_29.INJECT1_0 = "NO";
    defparam add_537_29.INJECT1_1 = "NO";
    CCU2D add_537_27 (.A0(u_r[26]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(u_r[27]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19800), 
          .COUT(n19801), .S0(n215[26]), .S1(n215[27]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[25:31])
    defparam add_537_27.INIT0 = 16'hf555;
    defparam add_537_27.INIT1 = 16'hf555;
    defparam add_537_27.INJECT1_0 = "NO";
    defparam add_537_27.INJECT1_1 = "NO";
    CCU2D add_537_25 (.A0(u_r[24]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(u_r[25]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19799), 
          .COUT(n19800), .S0(n215[24]), .S1(n215[25]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[25:31])
    defparam add_537_25.INIT0 = 16'hf555;
    defparam add_537_25.INIT1 = 16'hf555;
    defparam add_537_25.INJECT1_0 = "NO";
    defparam add_537_25.INJECT1_1 = "NO";
    CCU2D add_537_23 (.A0(u_r[22]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(u_r[23]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19798), 
          .COUT(n19799), .S0(n215[22]), .S1(n215[23]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[25:31])
    defparam add_537_23.INIT0 = 16'hf555;
    defparam add_537_23.INIT1 = 16'hf555;
    defparam add_537_23.INJECT1_0 = "NO";
    defparam add_537_23.INJECT1_1 = "NO";
    CCU2D add_537_21 (.A0(u_r[20]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(u_r[21]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19797), 
          .COUT(n19798), .S1(n215[21]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[25:31])
    defparam add_537_21.INIT0 = 16'hf555;
    defparam add_537_21.INIT1 = 16'hf555;
    defparam add_537_21.INJECT1_0 = "NO";
    defparam add_537_21.INJECT1_1 = "NO";
    CCU2D add_537_19 (.A0(u_r[18]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(u_r[19]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19796), 
          .COUT(n19797));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[25:31])
    defparam add_537_19.INIT0 = 16'hf555;
    defparam add_537_19.INIT1 = 16'hf555;
    defparam add_537_19.INJECT1_0 = "NO";
    defparam add_537_19.INJECT1_1 = "NO";
    CCU2D add_537_17 (.A0(u_r[16]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(u_r[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19795), 
          .COUT(n19796));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[25:31])
    defparam add_537_17.INIT0 = 16'hf555;
    defparam add_537_17.INIT1 = 16'hf555;
    defparam add_537_17.INJECT1_0 = "NO";
    defparam add_537_17.INJECT1_1 = "NO";
    CCU2D add_537_15 (.A0(u_r[14]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(u_r[15]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19794), 
          .COUT(n19795));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[25:31])
    defparam add_537_15.INIT0 = 16'hf555;
    defparam add_537_15.INIT1 = 16'hf555;
    defparam add_537_15.INJECT1_0 = "NO";
    defparam add_537_15.INJECT1_1 = "NO";
    CCU2D add_537_13 (.A0(u_r[12]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(u_r[13]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19793), 
          .COUT(n19794));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[25:31])
    defparam add_537_13.INIT0 = 16'hf555;
    defparam add_537_13.INIT1 = 16'hf555;
    defparam add_537_13.INJECT1_0 = "NO";
    defparam add_537_13.INJECT1_1 = "NO";
    CCU2D add_537_11 (.A0(u_r[10]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(u_r[11]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19792), 
          .COUT(n19793));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[25:31])
    defparam add_537_11.INIT0 = 16'hf555;
    defparam add_537_11.INIT1 = 16'hf555;
    defparam add_537_11.INJECT1_0 = "NO";
    defparam add_537_11.INJECT1_1 = "NO";
    CCU2D add_537_9 (.A0(u_r[8]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(u_r[9]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19791), 
          .COUT(n19792));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[25:31])
    defparam add_537_9.INIT0 = 16'hf555;
    defparam add_537_9.INIT1 = 16'hf555;
    defparam add_537_9.INJECT1_0 = "NO";
    defparam add_537_9.INJECT1_1 = "NO";
    CCU2D add_537_7 (.A0(u_r[6]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(u_r[7]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19790), 
          .COUT(n19791));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[25:31])
    defparam add_537_7.INIT0 = 16'hf555;
    defparam add_537_7.INIT1 = 16'hf555;
    defparam add_537_7.INJECT1_0 = "NO";
    defparam add_537_7.INJECT1_1 = "NO";
    CCU2D add_537_5 (.A0(u_r[4]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(u_r[5]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19789), 
          .COUT(n19790));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[25:31])
    defparam add_537_5.INIT0 = 16'hf555;
    defparam add_537_5.INIT1 = 16'hf555;
    defparam add_537_5.INJECT1_0 = "NO";
    defparam add_537_5.INJECT1_1 = "NO";
    CCU2D add_537_3 (.A0(u_r[2]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(u_r[3]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19788), 
          .COUT(n19789));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[25:31])
    defparam add_537_3.INIT0 = 16'hf555;
    defparam add_537_3.INIT1 = 16'hf555;
    defparam add_537_3.INJECT1_0 = "NO";
    defparam add_537_3.INJECT1_1 = "NO";
    CCU2D add_537_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(u_r[0]), .B1(u_r[1]), .C1(GND_net), .D1(GND_net), .COUT(n19788));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[25:31])
    defparam add_537_1.INIT0 = 16'hF000;
    defparam add_537_1.INIT1 = 16'ha666;
    defparam add_537_1.INJECT1_0 = "NO";
    defparam add_537_1.INJECT1_1 = "NO";
    CCU2D unary_minus_8_add_3_17 (.A0(o_sample_q[14]), .B0(o_sample_q[15]), 
          .C0(GND_net), .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n19623), .S0(u_l_15__N_1965[15]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(83[22:28])
    defparam unary_minus_8_add_3_17.INIT0 = 16'hd111;
    defparam unary_minus_8_add_3_17.INIT1 = 16'h0000;
    defparam unary_minus_8_add_3_17.INJECT1_0 = "NO";
    defparam unary_minus_8_add_3_17.INJECT1_1 = "NO";
    CCU2D unary_minus_8_add_3_15 (.A0(o_sample_q[12]), .B0(o_sample_q[15]), 
          .C0(o_sample_q[13]), .D0(GND_net), .A1(o_sample_q[13]), .B1(o_sample_q[15]), 
          .C1(o_sample_q[14]), .D1(GND_net), .CIN(n19622), .COUT(n19623), 
          .S0(u_l_15__N_1965[13]), .S1(u_l_15__N_1965[14]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(83[22:28])
    defparam unary_minus_8_add_3_15.INIT0 = 16'hdd2d;
    defparam unary_minus_8_add_3_15.INIT1 = 16'hdd2d;
    defparam unary_minus_8_add_3_15.INJECT1_0 = "NO";
    defparam unary_minus_8_add_3_15.INJECT1_1 = "NO";
    CCU2D unary_minus_8_add_3_13 (.A0(o_sample_q[10]), .B0(o_sample_q[15]), 
          .C0(o_sample_q[11]), .D0(GND_net), .A1(o_sample_q[11]), .B1(o_sample_q[15]), 
          .C1(o_sample_q[12]), .D1(GND_net), .CIN(n19621), .COUT(n19622), 
          .S0(u_l_15__N_1965[11]), .S1(u_l_15__N_1965[12]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(83[22:28])
    defparam unary_minus_8_add_3_13.INIT0 = 16'hdd2d;
    defparam unary_minus_8_add_3_13.INIT1 = 16'hdd2d;
    defparam unary_minus_8_add_3_13.INJECT1_0 = "NO";
    defparam unary_minus_8_add_3_13.INJECT1_1 = "NO";
    CCU2D unary_minus_8_add_3_11 (.A0(o_sample_q[8]), .B0(o_sample_q[15]), 
          .C0(o_sample_q[9]), .D0(GND_net), .A1(o_sample_q[9]), .B1(o_sample_q[15]), 
          .C1(o_sample_q[10]), .D1(GND_net), .CIN(n19620), .COUT(n19621), 
          .S0(u_l_15__N_1965[9]), .S1(u_l_15__N_1965[10]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(83[22:28])
    defparam unary_minus_8_add_3_11.INIT0 = 16'hdd2d;
    defparam unary_minus_8_add_3_11.INIT1 = 16'hdd2d;
    defparam unary_minus_8_add_3_11.INJECT1_0 = "NO";
    defparam unary_minus_8_add_3_11.INJECT1_1 = "NO";
    CCU2D unary_minus_8_add_3_9 (.A0(o_sample_q[6]), .B0(o_sample_q[15]), 
          .C0(o_sample_q[7]), .D0(GND_net), .A1(o_sample_q[7]), .B1(o_sample_q[15]), 
          .C1(o_sample_q[8]), .D1(GND_net), .CIN(n19619), .COUT(n19620), 
          .S0(u_l_15__N_1965[7]), .S1(u_l_15__N_1965[8]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(83[22:28])
    defparam unary_minus_8_add_3_9.INIT0 = 16'hdd2d;
    defparam unary_minus_8_add_3_9.INIT1 = 16'hdd2d;
    defparam unary_minus_8_add_3_9.INJECT1_0 = "NO";
    defparam unary_minus_8_add_3_9.INJECT1_1 = "NO";
    CCU2D unary_minus_8_add_3_7 (.A0(o_sample_q[4]), .B0(o_sample_q[15]), 
          .C0(o_sample_q[5]), .D0(GND_net), .A1(o_sample_q[5]), .B1(o_sample_q[15]), 
          .C1(o_sample_q[6]), .D1(GND_net), .CIN(n19618), .COUT(n19619), 
          .S0(u_l_15__N_1965[5]), .S1(u_l_15__N_1965[6]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(83[22:28])
    defparam unary_minus_8_add_3_7.INIT0 = 16'hdd2d;
    defparam unary_minus_8_add_3_7.INIT1 = 16'hdd2d;
    defparam unary_minus_8_add_3_7.INJECT1_0 = "NO";
    defparam unary_minus_8_add_3_7.INJECT1_1 = "NO";
    CCU2D unary_minus_8_add_3_5 (.A0(o_sample_q[2]), .B0(o_sample_q[15]), 
          .C0(o_sample_q[3]), .D0(GND_net), .A1(o_sample_q[3]), .B1(o_sample_q[15]), 
          .C1(o_sample_q[4]), .D1(GND_net), .CIN(n19617), .COUT(n19618), 
          .S0(u_l_15__N_1965[3]), .S1(u_l_15__N_1965[4]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(83[22:28])
    defparam unary_minus_8_add_3_5.INIT0 = 16'hdd2d;
    defparam unary_minus_8_add_3_5.INIT1 = 16'hdd2d;
    defparam unary_minus_8_add_3_5.INJECT1_0 = "NO";
    defparam unary_minus_8_add_3_5.INJECT1_1 = "NO";
    CCU2D unary_minus_8_add_3_3 (.A0(o_sample_q[0]), .B0(o_sample_q[15]), 
          .C0(o_sample_q[1]), .D0(GND_net), .A1(o_sample_q[1]), .B1(o_sample_q[15]), 
          .C1(o_sample_q[2]), .D1(GND_net), .CIN(n19616), .COUT(n19617), 
          .S0(u_l_15__N_1965[1]), .S1(u_l_15__N_1965[2]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(83[22:28])
    defparam unary_minus_8_add_3_3.INIT0 = 16'hdd2d;
    defparam unary_minus_8_add_3_3.INIT1 = 16'hdd2d;
    defparam unary_minus_8_add_3_3.INJECT1_0 = "NO";
    defparam unary_minus_8_add_3_3.INJECT1_1 = "NO";
    CCU2D unary_minus_8_add_3_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(o_sample_q[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n19616), .S1(u_l_15__N_1965[0]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(83[22:28])
    defparam unary_minus_8_add_3_1.INIT0 = 16'hF000;
    defparam unary_minus_8_add_3_1.INIT1 = 16'h0aaa;
    defparam unary_minus_8_add_3_1.INJECT1_0 = "NO";
    defparam unary_minus_8_add_3_1.INJECT1_1 = "NO";
    CCU2D unary_minus_6_add_3_15 (.A0(\addr_space[4][12] ), .B0(\addr_space[4][13] ), 
          .C0(GND_net), .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n19615), .S0(u_s_13__N_1951[13]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(82[22:28])
    defparam unary_minus_6_add_3_15.INIT0 = 16'hd111;
    defparam unary_minus_6_add_3_15.INIT1 = 16'h0000;
    defparam unary_minus_6_add_3_15.INJECT1_0 = "NO";
    defparam unary_minus_6_add_3_15.INJECT1_1 = "NO";
    CCU2D unary_minus_6_add_3_13 (.A0(\addr_space[4][10] ), .B0(\addr_space[4][13] ), 
          .C0(\addr_space[4][11] ), .D0(GND_net), .A1(\addr_space[4][11] ), 
          .B1(\addr_space[4][13] ), .C1(\addr_space[4][12] ), .D1(GND_net), 
          .CIN(n19614), .COUT(n19615), .S0(u_s_13__N_1951[11]), .S1(u_s_13__N_1951[12]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(82[22:28])
    defparam unary_minus_6_add_3_13.INIT0 = 16'hdd2d;
    defparam unary_minus_6_add_3_13.INIT1 = 16'hdd2d;
    defparam unary_minus_6_add_3_13.INJECT1_0 = "NO";
    defparam unary_minus_6_add_3_13.INJECT1_1 = "NO";
    CCU2D unary_minus_6_add_3_11 (.A0(\addr_space[4][8] ), .B0(\addr_space[4][13] ), 
          .C0(\addr_space[4][9] ), .D0(GND_net), .A1(\addr_space[4][9] ), 
          .B1(\addr_space[4][13] ), .C1(\addr_space[4][10] ), .D1(GND_net), 
          .CIN(n19613), .COUT(n19614), .S0(u_s_13__N_1951[9]), .S1(u_s_13__N_1951[10]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(82[22:28])
    defparam unary_minus_6_add_3_11.INIT0 = 16'hdd2d;
    defparam unary_minus_6_add_3_11.INIT1 = 16'hdd2d;
    defparam unary_minus_6_add_3_11.INJECT1_0 = "NO";
    defparam unary_minus_6_add_3_11.INJECT1_1 = "NO";
    CCU2D unary_minus_6_add_3_9 (.A0(\addr_space[4][6] ), .B0(\addr_space[4][13] ), 
          .C0(\addr_space[4][7] ), .D0(GND_net), .A1(\addr_space[4][7] ), 
          .B1(\addr_space[4][13] ), .C1(\addr_space[4][8] ), .D1(GND_net), 
          .CIN(n19612), .COUT(n19613), .S0(u_s_13__N_1951[7]), .S1(u_s_13__N_1951[8]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(82[22:28])
    defparam unary_minus_6_add_3_9.INIT0 = 16'hdd2d;
    defparam unary_minus_6_add_3_9.INIT1 = 16'hdd2d;
    defparam unary_minus_6_add_3_9.INJECT1_0 = "NO";
    defparam unary_minus_6_add_3_9.INJECT1_1 = "NO";
    CCU2D unary_minus_6_add_3_7 (.A0(\addr_space[4][4] ), .B0(\addr_space[4][13] ), 
          .C0(\addr_space[4][5] ), .D0(GND_net), .A1(\addr_space[4][5] ), 
          .B1(\addr_space[4][13] ), .C1(\addr_space[4][6] ), .D1(GND_net), 
          .CIN(n19611), .COUT(n19612), .S0(u_s_13__N_1951[5]), .S1(u_s_13__N_1951[6]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(82[22:28])
    defparam unary_minus_6_add_3_7.INIT0 = 16'hdd2d;
    defparam unary_minus_6_add_3_7.INIT1 = 16'hdd2d;
    defparam unary_minus_6_add_3_7.INJECT1_0 = "NO";
    defparam unary_minus_6_add_3_7.INJECT1_1 = "NO";
    CCU2D unary_minus_6_add_3_5 (.A0(\addr_space[4][2] ), .B0(\addr_space[4][13] ), 
          .C0(\addr_space[4][3] ), .D0(GND_net), .A1(\addr_space[4][3] ), 
          .B1(\addr_space[4][13] ), .C1(\addr_space[4][4] ), .D1(GND_net), 
          .CIN(n19610), .COUT(n19611), .S0(u_s_13__N_1951[3]), .S1(u_s_13__N_1951[4]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(82[22:28])
    defparam unary_minus_6_add_3_5.INIT0 = 16'hdd2d;
    defparam unary_minus_6_add_3_5.INIT1 = 16'hdd2d;
    defparam unary_minus_6_add_3_5.INJECT1_0 = "NO";
    defparam unary_minus_6_add_3_5.INJECT1_1 = "NO";
    CCU2D unary_minus_6_add_3_3 (.A0(\addr_space[4][0] ), .B0(\addr_space[4][13] ), 
          .C0(\addr_space[4][1] ), .D0(GND_net), .A1(\addr_space[4][1] ), 
          .B1(\addr_space[4][13] ), .C1(\addr_space[4][2] ), .D1(GND_net), 
          .CIN(n19609), .COUT(n19610), .S0(u_s_13__N_1951[1]), .S1(u_s_13__N_1951[2]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(82[22:28])
    defparam unary_minus_6_add_3_3.INIT0 = 16'hdd2d;
    defparam unary_minus_6_add_3_3.INIT1 = 16'hdd2d;
    defparam unary_minus_6_add_3_3.INJECT1_0 = "NO";
    defparam unary_minus_6_add_3_3.INJECT1_1 = "NO";
    CCU2D unary_minus_6_add_3_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\addr_space[4][0] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n19609), .S1(u_s_13__N_1951[0]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(82[22:28])
    defparam unary_minus_6_add_3_1.INIT0 = 16'hF000;
    defparam unary_minus_6_add_3_1.INIT1 = 16'h0aaa;
    defparam unary_minus_6_add_3_1.INJECT1_0 = "NO";
    defparam unary_minus_6_add_3_1.INJECT1_1 = "NO";
    LUT4 mux_644_i9_3_lut (.A(u_r[29]), .B(n215[29]), .C(u_sgn[4]), .Z(o_p_29__N_1986[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[10:35])
    defparam mux_644_i9_3_lut.init = 16'hcaca;
    LUT4 mux_644_i8_3_lut (.A(u_r[28]), .B(n215[28]), .C(u_sgn[4]), .Z(o_p_29__N_1986[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[10:35])
    defparam mux_644_i8_3_lut.init = 16'hcaca;
    LUT4 mux_644_i7_3_lut (.A(u_r[27]), .B(n215[27]), .C(u_sgn[4]), .Z(o_p_29__N_1986[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[10:35])
    defparam mux_644_i7_3_lut.init = 16'hcaca;
    LUT4 mux_644_i6_3_lut (.A(u_r[26]), .B(n215[26]), .C(u_sgn[4]), .Z(o_p_29__N_1986[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[10:35])
    defparam mux_644_i6_3_lut.init = 16'hcaca;
    LUT4 mux_644_i5_3_lut (.A(u_r[25]), .B(n215[25]), .C(u_sgn[4]), .Z(o_p_29__N_1986[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[10:35])
    defparam mux_644_i5_3_lut.init = 16'hcaca;
    LUT4 mux_644_i4_3_lut (.A(u_r[24]), .B(n215[24]), .C(u_sgn[4]), .Z(o_p_29__N_1986[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[10:35])
    defparam mux_644_i4_3_lut.init = 16'hcaca;
    LUT4 mux_644_i3_3_lut (.A(u_r[23]), .B(n215[23]), .C(u_sgn[4]), .Z(o_p_29__N_1986[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[10:35])
    defparam mux_644_i3_3_lut.init = 16'hcaca;
    LUT4 mux_644_i2_3_lut (.A(u_r[22]), .B(n215[22]), .C(u_sgn[4]), .Z(o_p_29__N_1986[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[10:35])
    defparam mux_644_i2_3_lut.init = 16'hcaca;
    FD1S3IX o_p__i9 (.D(o_p_29__N_1986[29]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_dac_b[8] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=109, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(98[9] 102[36])
    defparam o_p__i9.GSR = "DISABLED";
    FD1S3IX o_p__i8 (.D(o_p_29__N_1986[28]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_dac_b[7] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=109, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(98[9] 102[36])
    defparam o_p__i8.GSR = "DISABLED";
    FD1S3IX o_p__i7 (.D(o_p_29__N_1986[27]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_dac_b[6] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=109, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(98[9] 102[36])
    defparam o_p__i7.GSR = "DISABLED";
    FD1S3IX o_p__i6 (.D(o_p_29__N_1986[26]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_dac_b[5] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=109, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(98[9] 102[36])
    defparam o_p__i6.GSR = "DISABLED";
    FD1S3IX o_p__i5 (.D(o_p_29__N_1986[25]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_dac_b[4] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=109, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(98[9] 102[36])
    defparam o_p__i5.GSR = "DISABLED";
    FD1S3IX o_p__i4 (.D(o_p_29__N_1986[24]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_dac_b[3] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=109, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(98[9] 102[36])
    defparam o_p__i4.GSR = "DISABLED";
    FD1S3IX o_p__i3 (.D(o_p_29__N_1986[23]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_dac_b[2] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=109, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(98[9] 102[36])
    defparam o_p__i3.GSR = "DISABLED";
    FD1S3IX o_p__i2 (.D(o_p_29__N_1986[22]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_dac_b[1] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=109, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(98[9] 102[36])
    defparam o_p__i2.GSR = "DISABLED";
    FD1S3IX u_sgn__i4 (.D(u_sgn[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(u_sgn[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=109, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(87[9] 91[60])
    defparam u_sgn__i4.GSR = "DISABLED";
    FD1S3IX u_sgn__i3 (.D(u_sgn[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(u_sgn[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=109, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(87[9] 91[60])
    defparam u_sgn__i3.GSR = "DISABLED";
    FD1S3IX u_sgn__i2 (.D(u_sgn[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(u_sgn[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=109, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(87[9] 91[60])
    defparam u_sgn__i2.GSR = "DISABLED";
    FD1S3IX u_sgn__i1 (.D(u_sgn[0]), .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(u_sgn[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=109, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(87[9] 91[60])
    defparam u_sgn__i1.GSR = "DISABLED";
    FD1S3IX u_l__i15 (.D(u_l_15__N_1965[15]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_l[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=109, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_l__i15.GSR = "DISABLED";
    FD1S3IX u_l__i14 (.D(u_l_15__N_1965[14]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_l[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=109, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_l__i14.GSR = "DISABLED";
    FD1S3IX u_l__i13 (.D(u_l_15__N_1965[13]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_l[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=109, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_l__i13.GSR = "DISABLED";
    FD1S3IX u_l__i12 (.D(u_l_15__N_1965[12]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_l[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=109, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_l__i12.GSR = "DISABLED";
    FD1S3IX u_l__i11 (.D(u_l_15__N_1965[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_l[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=109, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_l__i11.GSR = "DISABLED";
    FD1S3IX u_l__i10 (.D(u_l_15__N_1965[10]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_l[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=109, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_l__i10.GSR = "DISABLED";
    FD1S3IX u_l__i9 (.D(u_l_15__N_1965[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_l[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=109, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_l__i9.GSR = "DISABLED";
    FD1S3IX u_l__i8 (.D(u_l_15__N_1965[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_l[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=109, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_l__i8.GSR = "DISABLED";
    FD1S3IX u_l__i7 (.D(u_l_15__N_1965[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_l[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=109, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_l__i7.GSR = "DISABLED";
    FD1S3IX u_l__i6 (.D(u_l_15__N_1965[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_l[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=109, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_l__i6.GSR = "DISABLED";
    FD1S3IX u_l__i5 (.D(u_l_15__N_1965[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_l[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=109, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_l__i5.GSR = "DISABLED";
    FD1S3IX u_l__i4 (.D(u_l_15__N_1965[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_l[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=109, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_l__i4.GSR = "DISABLED";
    FD1S3IX u_l__i3 (.D(u_l_15__N_1965[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_l[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=109, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_l__i3.GSR = "DISABLED";
    FD1S3IX u_l__i2 (.D(u_l_15__N_1965[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_l[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=109, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_l__i2.GSR = "DISABLED";
    FD1S3IX u_l__i1 (.D(u_l_15__N_1965[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_l[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=109, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_l__i1.GSR = "DISABLED";
    FD1S3IX u_s__i13 (.D(u_s_13__N_1951[13]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_s_c[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=109, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_s__i13.GSR = "DISABLED";
    FD1S3IX u_s__i12 (.D(u_s_13__N_1951[12]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\u_s[12] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=109, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_s__i12.GSR = "DISABLED";
    FD1S3IX u_s__i11 (.D(u_s_13__N_1951[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_s_c[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=109, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_s__i11.GSR = "DISABLED";
    FD1S3IX u_s__i10 (.D(u_s_13__N_1951[10]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\u_s[10] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=109, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_s__i10.GSR = "DISABLED";
    FD1S3IX u_s__i9 (.D(u_s_13__N_1951[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_s_c[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=109, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_s__i9.GSR = "DISABLED";
    FD1S3IX u_s__i8 (.D(u_s_13__N_1951[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\u_s[8] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=109, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_s__i8.GSR = "DISABLED";
    FD1S3IX u_s__i7 (.D(u_s_13__N_1951[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_s_c[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=109, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_s__i7.GSR = "DISABLED";
    FD1S3IX u_s__i6 (.D(u_s_13__N_1951[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\u_s[6] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=109, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_s__i6.GSR = "DISABLED";
    FD1S3IX u_s__i5 (.D(u_s_13__N_1951[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_s_c[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=109, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_s__i5.GSR = "DISABLED";
    FD1S3IX u_s__i4 (.D(u_s_13__N_1951[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\u_s[4] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=109, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_s__i4.GSR = "DISABLED";
    FD1S3IX u_s__i3 (.D(u_s_13__N_1951[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_s_c[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=109, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_s__i3.GSR = "DISABLED";
    FD1S3IX u_s__i2 (.D(u_s_13__N_1951[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\u_s[2] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=109, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_s__i2.GSR = "DISABLED";
    FD1S3IX u_s__i1 (.D(u_s_13__N_1951[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_s_c[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=109, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_s__i1.GSR = "DISABLED";
    umpy_14x16 umpy (.dac_clk_p_c(dac_clk_p_c), .i_sw0_c(i_sw0_c), .u_r({u_r}), 
            .GND_net(GND_net), .n14230(n14230), .n9458(n9458), .u_l({u_l}), 
            .u_s({u_s_c[13], \u_s[12] , u_s_c[11], \u_s[10] , u_s_c[9], 
            \u_s[8] , u_s_c[7], \u_s[6] , u_s_c[5], \u_s[4] , u_s_c[3], 
            \u_s[2] , u_s_c[1], u_s[0]}), .n9460(n9460), .n9462(n9462), 
            .n9464(n9464), .n9466(n9466), .n9468(n9468), .n9488(n9488)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(95[13:68])
    
endmodule
//
// Verilog Description of module umpy_14x16
//

module umpy_14x16 (dac_clk_p_c, i_sw0_c, u_r, GND_net, n14230, n9458, 
            u_l, u_s, n9460, n9462, n9464, n9466, n9468, n9488) /* synthesis syn_module_defined=1 */ ;
    input dac_clk_p_c;
    input i_sw0_c;
    output [29:0]u_r;
    input GND_net;
    input n14230;
    input n9458;
    input [15:0]u_l;
    input [13:0]u_s;
    input n9460;
    input n9462;
    input n9464;
    input n9466;
    input n9468;
    input n9488;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[29:38])
    wire [20:0]S_1_00;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(103[17:23])
    wire [17:0]S_0_00;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(71[14:20])
    wire [20:0]S_1_01;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(104[17:23])
    wire [17:0]S_0_02;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(77[14:20])
    wire [25:0]S_2_01_25__N_2294;
    wire [17:0]S_0_04;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(83[14:20])
    wire [20:0]S_1_03;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(106[17:23])
    wire [17:0]S_0_06;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(89[14:20])
    wire [29:0]o_p_29__N_2320;
    wire [25:0]S_2_01;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(140[17:23])
    
    wire n19864;
    wire [20:0]S_1_02_20__N_2226;
    
    wire n19863;
    wire [17:0]S_0_05;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(86[14:20])
    
    wire n19862, n19861, n19860, n19859, n19858, n19857, n19856, 
        n19854;
    wire [25:0]S_2_00_25__N_2268;
    
    wire n19853, n19852, n19851, n19850, n19849, n19848, n19847, 
        n19846, n19845, n19843;
    wire [20:0]S_1_00_20__N_2184;
    
    wire n19842;
    wire [17:0]S_0_01;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(74[14:20])
    
    wire n19841, n19840, n19839, n19838, n19837, n19836, n19835, 
        n19645;
    wire [20:0]S_1_01_20__N_2205;
    
    wire n19644;
    wire [17:0]S_0_03;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(80[14:20])
    
    wire n19643, n19642, n19641, n19640, n19639, n19638, n19637, 
        n19634, n19633, n19632;
    wire [25:0]S_2_00;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(139[17:23])
    
    wire n19631, n19630, n19629, n19628, n19627, n19626, n19625;
    wire [20:0]S_1_02;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(105[17:23])
    
    wire n19570, n19569, n19568, n19567, n19566, n19565, n19564, 
        n19563;
    
    FD1S3IX S_1_00__i0 (.D(S_0_00[0]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_00[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i0.GSR = "DISABLED";
    FD1S3IX S_1_01__i0 (.D(S_0_02[0]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i0.GSR = "DISABLED";
    FD1S3IX S_1_02__i1 (.D(S_0_04[0]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01_25__N_2294[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i1.GSR = "DISABLED";
    FD1S3IX S_1_03__i1 (.D(S_0_06[0]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_03[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_03__i1.GSR = "DISABLED";
    FD1S3IX S_2_00__i1 (.D(S_1_00[0]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_p_29__N_2320[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i1.GSR = "DISABLED";
    FD1S3IX S_2_01__i1 (.D(S_2_01_25__N_2294[0]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i1.GSR = "DISABLED";
    FD1S3IX S_3_00__i0 (.D(o_p_29__N_2320[0]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i0.GSR = "DISABLED";
    CCU2D add_848_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19864), 
          .S0(S_1_02_20__N_2226[20]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(124[13:48])
    defparam add_848_cout.INIT0 = 16'h0000;
    defparam add_848_cout.INIT1 = 16'h0000;
    defparam add_848_cout.INJECT1_0 = "NO";
    defparam add_848_cout.INJECT1_1 = "NO";
    CCU2D add_848_18 (.A0(S_0_05[16]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(S_0_05[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n19863), .COUT(n19864), .S0(S_1_02_20__N_2226[18]), .S1(S_1_02_20__N_2226[19]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(124[13:48])
    defparam add_848_18.INIT0 = 16'hfaaa;
    defparam add_848_18.INIT1 = 16'hfaaa;
    defparam add_848_18.INJECT1_0 = "NO";
    defparam add_848_18.INJECT1_1 = "NO";
    CCU2D add_848_16 (.A0(S_0_04[16]), .B0(S_0_05[14]), .C0(GND_net), 
          .D0(GND_net), .A1(S_0_04[17]), .B1(S_0_05[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n19862), .COUT(n19863), .S0(S_1_02_20__N_2226[16]), 
          .S1(S_1_02_20__N_2226[17]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(124[13:48])
    defparam add_848_16.INIT0 = 16'h5666;
    defparam add_848_16.INIT1 = 16'h5666;
    defparam add_848_16.INJECT1_0 = "NO";
    defparam add_848_16.INJECT1_1 = "NO";
    CCU2D add_848_14 (.A0(S_0_04[14]), .B0(S_0_05[12]), .C0(GND_net), 
          .D0(GND_net), .A1(S_0_04[15]), .B1(S_0_05[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n19861), .COUT(n19862), .S0(S_1_02_20__N_2226[14]), 
          .S1(S_1_02_20__N_2226[15]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(124[13:48])
    defparam add_848_14.INIT0 = 16'h5666;
    defparam add_848_14.INIT1 = 16'h5666;
    defparam add_848_14.INJECT1_0 = "NO";
    defparam add_848_14.INJECT1_1 = "NO";
    CCU2D add_848_12 (.A0(S_0_04[12]), .B0(S_0_05[10]), .C0(GND_net), 
          .D0(GND_net), .A1(S_0_04[13]), .B1(S_0_05[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n19860), .COUT(n19861), .S0(S_1_02_20__N_2226[12]), 
          .S1(S_1_02_20__N_2226[13]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(124[13:48])
    defparam add_848_12.INIT0 = 16'h5666;
    defparam add_848_12.INIT1 = 16'h5666;
    defparam add_848_12.INJECT1_0 = "NO";
    defparam add_848_12.INJECT1_1 = "NO";
    CCU2D add_848_10 (.A0(S_0_04[10]), .B0(S_0_05[8]), .C0(GND_net), .D0(GND_net), 
          .A1(S_0_04[11]), .B1(S_0_05[9]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19859), .COUT(n19860), .S0(S_1_02_20__N_2226[10]), .S1(S_1_02_20__N_2226[11]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(124[13:48])
    defparam add_848_10.INIT0 = 16'h5666;
    defparam add_848_10.INIT1 = 16'h5666;
    defparam add_848_10.INJECT1_0 = "NO";
    defparam add_848_10.INJECT1_1 = "NO";
    CCU2D add_848_8 (.A0(S_0_04[8]), .B0(S_0_05[6]), .C0(GND_net), .D0(GND_net), 
          .A1(S_0_04[9]), .B1(S_0_05[7]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19858), .COUT(n19859), .S0(S_1_02_20__N_2226[8]), .S1(S_1_02_20__N_2226[9]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(124[13:48])
    defparam add_848_8.INIT0 = 16'h5666;
    defparam add_848_8.INIT1 = 16'h5666;
    defparam add_848_8.INJECT1_0 = "NO";
    defparam add_848_8.INJECT1_1 = "NO";
    CCU2D add_848_6 (.A0(S_0_04[6]), .B0(S_0_05[4]), .C0(GND_net), .D0(GND_net), 
          .A1(S_0_04[7]), .B1(S_0_05[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19857), .COUT(n19858), .S0(S_1_02_20__N_2226[6]), .S1(S_1_02_20__N_2226[7]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(124[13:48])
    defparam add_848_6.INIT0 = 16'h5666;
    defparam add_848_6.INIT1 = 16'h5666;
    defparam add_848_6.INJECT1_0 = "NO";
    defparam add_848_6.INJECT1_1 = "NO";
    CCU2D add_848_4 (.A0(S_0_04[4]), .B0(S_0_05[2]), .C0(GND_net), .D0(GND_net), 
          .A1(S_0_04[5]), .B1(S_0_05[3]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19856), .COUT(n19857), .S0(S_1_02_20__N_2226[4]), .S1(S_1_02_20__N_2226[5]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(124[13:48])
    defparam add_848_4.INIT0 = 16'h5666;
    defparam add_848_4.INIT1 = 16'h5666;
    defparam add_848_4.INJECT1_0 = "NO";
    defparam add_848_4.INJECT1_1 = "NO";
    CCU2D add_848_2 (.A0(S_0_04[2]), .B0(S_0_05[0]), .C0(GND_net), .D0(GND_net), 
          .A1(S_0_04[3]), .B1(S_0_05[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n19856), .S1(S_1_02_20__N_2226[3]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(124[13:48])
    defparam add_848_2.INIT0 = 16'h7000;
    defparam add_848_2.INIT1 = 16'h5666;
    defparam add_848_2.INJECT1_0 = "NO";
    defparam add_848_2.INJECT1_1 = "NO";
    CCU2D add_847_22 (.A0(S_1_01[20]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19854), 
          .S0(S_2_00_25__N_2268[24]), .S1(S_2_00_25__N_2268[25]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(152[13:48])
    defparam add_847_22.INIT0 = 16'hfaaa;
    defparam add_847_22.INIT1 = 16'h0000;
    defparam add_847_22.INJECT1_0 = "NO";
    defparam add_847_22.INJECT1_1 = "NO";
    CCU2D add_847_20 (.A0(S_1_01[18]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(S_1_01[19]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n19853), .COUT(n19854), .S0(S_2_00_25__N_2268[22]), .S1(S_2_00_25__N_2268[23]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(152[13:48])
    defparam add_847_20.INIT0 = 16'hfaaa;
    defparam add_847_20.INIT1 = 16'hfaaa;
    defparam add_847_20.INJECT1_0 = "NO";
    defparam add_847_20.INJECT1_1 = "NO";
    CCU2D add_847_18 (.A0(S_1_00[20]), .B0(S_1_01[16]), .C0(GND_net), 
          .D0(GND_net), .A1(S_1_01[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n19852), .COUT(n19853), .S0(S_2_00_25__N_2268[20]), 
          .S1(S_2_00_25__N_2268[21]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(152[13:48])
    defparam add_847_18.INIT0 = 16'h5666;
    defparam add_847_18.INIT1 = 16'hfaaa;
    defparam add_847_18.INJECT1_0 = "NO";
    defparam add_847_18.INJECT1_1 = "NO";
    CCU2D add_847_16 (.A0(S_1_00[18]), .B0(S_1_01[14]), .C0(GND_net), 
          .D0(GND_net), .A1(S_1_00[19]), .B1(S_1_01[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n19851), .COUT(n19852), .S0(S_2_00_25__N_2268[18]), 
          .S1(S_2_00_25__N_2268[19]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(152[13:48])
    defparam add_847_16.INIT0 = 16'h5666;
    defparam add_847_16.INIT1 = 16'h5666;
    defparam add_847_16.INJECT1_0 = "NO";
    defparam add_847_16.INJECT1_1 = "NO";
    CCU2D add_847_14 (.A0(S_1_00[16]), .B0(S_1_01[12]), .C0(GND_net), 
          .D0(GND_net), .A1(S_1_00[17]), .B1(S_1_01[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n19850), .COUT(n19851), .S0(S_2_00_25__N_2268[16]), 
          .S1(S_2_00_25__N_2268[17]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(152[13:48])
    defparam add_847_14.INIT0 = 16'h5666;
    defparam add_847_14.INIT1 = 16'h5666;
    defparam add_847_14.INJECT1_0 = "NO";
    defparam add_847_14.INJECT1_1 = "NO";
    CCU2D add_847_12 (.A0(S_1_00[14]), .B0(S_1_01[10]), .C0(GND_net), 
          .D0(GND_net), .A1(S_1_00[15]), .B1(S_1_01[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n19849), .COUT(n19850), .S0(S_2_00_25__N_2268[14]), 
          .S1(S_2_00_25__N_2268[15]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(152[13:48])
    defparam add_847_12.INIT0 = 16'h5666;
    defparam add_847_12.INIT1 = 16'h5666;
    defparam add_847_12.INJECT1_0 = "NO";
    defparam add_847_12.INJECT1_1 = "NO";
    CCU2D add_847_10 (.A0(S_1_00[12]), .B0(S_1_01[8]), .C0(GND_net), .D0(GND_net), 
          .A1(S_1_00[13]), .B1(S_1_01[9]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19848), .COUT(n19849), .S0(S_2_00_25__N_2268[12]), .S1(S_2_00_25__N_2268[13]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(152[13:48])
    defparam add_847_10.INIT0 = 16'h5666;
    defparam add_847_10.INIT1 = 16'h5666;
    defparam add_847_10.INJECT1_0 = "NO";
    defparam add_847_10.INJECT1_1 = "NO";
    CCU2D add_847_8 (.A0(S_1_00[10]), .B0(S_1_01[6]), .C0(GND_net), .D0(GND_net), 
          .A1(S_1_00[11]), .B1(S_1_01[7]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19847), .COUT(n19848), .S0(S_2_00_25__N_2268[10]), .S1(S_2_00_25__N_2268[11]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(152[13:48])
    defparam add_847_8.INIT0 = 16'h5666;
    defparam add_847_8.INIT1 = 16'h5666;
    defparam add_847_8.INJECT1_0 = "NO";
    defparam add_847_8.INJECT1_1 = "NO";
    CCU2D add_847_6 (.A0(S_1_00[8]), .B0(S_1_01[4]), .C0(GND_net), .D0(GND_net), 
          .A1(S_1_00[9]), .B1(S_1_01[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19846), .COUT(n19847), .S0(S_2_00_25__N_2268[8]), .S1(S_2_00_25__N_2268[9]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(152[13:48])
    defparam add_847_6.INIT0 = 16'h5666;
    defparam add_847_6.INIT1 = 16'h5666;
    defparam add_847_6.INJECT1_0 = "NO";
    defparam add_847_6.INJECT1_1 = "NO";
    CCU2D add_847_4 (.A0(S_1_00[6]), .B0(S_1_01[2]), .C0(GND_net), .D0(GND_net), 
          .A1(S_1_00[7]), .B1(S_1_01[3]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19845), .COUT(n19846), .S0(S_2_00_25__N_2268[6]), .S1(S_2_00_25__N_2268[7]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(152[13:48])
    defparam add_847_4.INIT0 = 16'h5666;
    defparam add_847_4.INIT1 = 16'h5666;
    defparam add_847_4.INJECT1_0 = "NO";
    defparam add_847_4.INJECT1_1 = "NO";
    CCU2D add_847_2 (.A0(S_1_00[4]), .B0(S_1_01[0]), .C0(GND_net), .D0(GND_net), 
          .A1(S_1_00[5]), .B1(S_1_01[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n19845), .S1(S_2_00_25__N_2268[5]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(152[13:48])
    defparam add_847_2.INIT0 = 16'h7000;
    defparam add_847_2.INIT1 = 16'h5666;
    defparam add_847_2.INJECT1_0 = "NO";
    defparam add_847_2.INJECT1_1 = "NO";
    CCU2D add_846_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19843), 
          .S0(S_1_00_20__N_2184[20]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(122[13:48])
    defparam add_846_cout.INIT0 = 16'h0000;
    defparam add_846_cout.INIT1 = 16'h0000;
    defparam add_846_cout.INJECT1_0 = "NO";
    defparam add_846_cout.INJECT1_1 = "NO";
    CCU2D add_846_18 (.A0(S_0_01[16]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(S_0_01[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n19842), .COUT(n19843), .S0(S_1_00_20__N_2184[18]), .S1(S_1_00_20__N_2184[19]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(122[13:48])
    defparam add_846_18.INIT0 = 16'hfaaa;
    defparam add_846_18.INIT1 = 16'hfaaa;
    defparam add_846_18.INJECT1_0 = "NO";
    defparam add_846_18.INJECT1_1 = "NO";
    CCU2D add_846_16 (.A0(S_0_00[16]), .B0(S_0_01[14]), .C0(GND_net), 
          .D0(GND_net), .A1(S_0_00[17]), .B1(S_0_01[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n19841), .COUT(n19842), .S0(S_1_00_20__N_2184[16]), 
          .S1(S_1_00_20__N_2184[17]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(122[13:48])
    defparam add_846_16.INIT0 = 16'h5666;
    defparam add_846_16.INIT1 = 16'h5666;
    defparam add_846_16.INJECT1_0 = "NO";
    defparam add_846_16.INJECT1_1 = "NO";
    CCU2D add_846_14 (.A0(S_0_00[14]), .B0(S_0_01[12]), .C0(GND_net), 
          .D0(GND_net), .A1(S_0_00[15]), .B1(S_0_01[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n19840), .COUT(n19841), .S0(S_1_00_20__N_2184[14]), 
          .S1(S_1_00_20__N_2184[15]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(122[13:48])
    defparam add_846_14.INIT0 = 16'h5666;
    defparam add_846_14.INIT1 = 16'h5666;
    defparam add_846_14.INJECT1_0 = "NO";
    defparam add_846_14.INJECT1_1 = "NO";
    CCU2D add_846_12 (.A0(S_0_00[12]), .B0(S_0_01[10]), .C0(GND_net), 
          .D0(GND_net), .A1(S_0_00[13]), .B1(S_0_01[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n19839), .COUT(n19840), .S0(S_1_00_20__N_2184[12]), 
          .S1(S_1_00_20__N_2184[13]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(122[13:48])
    defparam add_846_12.INIT0 = 16'h5666;
    defparam add_846_12.INIT1 = 16'h5666;
    defparam add_846_12.INJECT1_0 = "NO";
    defparam add_846_12.INJECT1_1 = "NO";
    CCU2D add_846_10 (.A0(S_0_00[10]), .B0(S_0_01[8]), .C0(GND_net), .D0(GND_net), 
          .A1(S_0_00[11]), .B1(S_0_01[9]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19838), .COUT(n19839), .S0(S_1_00_20__N_2184[10]), .S1(S_1_00_20__N_2184[11]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(122[13:48])
    defparam add_846_10.INIT0 = 16'h5666;
    defparam add_846_10.INIT1 = 16'h5666;
    defparam add_846_10.INJECT1_0 = "NO";
    defparam add_846_10.INJECT1_1 = "NO";
    CCU2D add_846_8 (.A0(S_0_00[8]), .B0(S_0_01[6]), .C0(GND_net), .D0(GND_net), 
          .A1(S_0_00[9]), .B1(S_0_01[7]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19837), .COUT(n19838), .S0(S_1_00_20__N_2184[8]), .S1(S_1_00_20__N_2184[9]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(122[13:48])
    defparam add_846_8.INIT0 = 16'h5666;
    defparam add_846_8.INIT1 = 16'h5666;
    defparam add_846_8.INJECT1_0 = "NO";
    defparam add_846_8.INJECT1_1 = "NO";
    CCU2D add_846_6 (.A0(S_0_00[6]), .B0(S_0_01[4]), .C0(GND_net), .D0(GND_net), 
          .A1(S_0_00[7]), .B1(S_0_01[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19836), .COUT(n19837), .S0(S_1_00_20__N_2184[6]), .S1(S_1_00_20__N_2184[7]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(122[13:48])
    defparam add_846_6.INIT0 = 16'h5666;
    defparam add_846_6.INIT1 = 16'h5666;
    defparam add_846_6.INJECT1_0 = "NO";
    defparam add_846_6.INJECT1_1 = "NO";
    CCU2D add_846_4 (.A0(S_0_00[4]), .B0(S_0_01[2]), .C0(GND_net), .D0(GND_net), 
          .A1(S_0_00[5]), .B1(S_0_01[3]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19835), .COUT(n19836), .S0(S_1_00_20__N_2184[4]), .S1(S_1_00_20__N_2184[5]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(122[13:48])
    defparam add_846_4.INIT0 = 16'h5666;
    defparam add_846_4.INIT1 = 16'h5666;
    defparam add_846_4.INJECT1_0 = "NO";
    defparam add_846_4.INJECT1_1 = "NO";
    CCU2D add_846_2 (.A0(S_0_00[2]), .B0(S_0_01[0]), .C0(GND_net), .D0(GND_net), 
          .A1(S_0_00[3]), .B1(S_0_01[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n19835), .S1(S_1_00_20__N_2184[3]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(122[13:48])
    defparam add_846_2.INIT0 = 16'h7000;
    defparam add_846_2.INIT1 = 16'h5666;
    defparam add_846_2.INJECT1_0 = "NO";
    defparam add_846_2.INJECT1_1 = "NO";
    CCU2D add_836_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19645), 
          .S0(S_1_01_20__N_2205[20]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(123[13:48])
    defparam add_836_cout.INIT0 = 16'h0000;
    defparam add_836_cout.INIT1 = 16'h0000;
    defparam add_836_cout.INJECT1_0 = "NO";
    defparam add_836_cout.INJECT1_1 = "NO";
    CCU2D add_836_18 (.A0(S_0_03[16]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(S_0_03[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n19644), .COUT(n19645), .S0(S_1_01_20__N_2205[18]), .S1(S_1_01_20__N_2205[19]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(123[13:48])
    defparam add_836_18.INIT0 = 16'hfaaa;
    defparam add_836_18.INIT1 = 16'hfaaa;
    defparam add_836_18.INJECT1_0 = "NO";
    defparam add_836_18.INJECT1_1 = "NO";
    CCU2D add_836_16 (.A0(S_0_02[16]), .B0(S_0_03[14]), .C0(GND_net), 
          .D0(GND_net), .A1(S_0_02[17]), .B1(S_0_03[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n19643), .COUT(n19644), .S0(S_1_01_20__N_2205[16]), 
          .S1(S_1_01_20__N_2205[17]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(123[13:48])
    defparam add_836_16.INIT0 = 16'h5666;
    defparam add_836_16.INIT1 = 16'h5666;
    defparam add_836_16.INJECT1_0 = "NO";
    defparam add_836_16.INJECT1_1 = "NO";
    CCU2D add_836_14 (.A0(S_0_02[14]), .B0(S_0_03[12]), .C0(GND_net), 
          .D0(GND_net), .A1(S_0_02[15]), .B1(S_0_03[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n19642), .COUT(n19643), .S0(S_1_01_20__N_2205[14]), 
          .S1(S_1_01_20__N_2205[15]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(123[13:48])
    defparam add_836_14.INIT0 = 16'h5666;
    defparam add_836_14.INIT1 = 16'h5666;
    defparam add_836_14.INJECT1_0 = "NO";
    defparam add_836_14.INJECT1_1 = "NO";
    CCU2D add_836_12 (.A0(S_0_02[12]), .B0(S_0_03[10]), .C0(GND_net), 
          .D0(GND_net), .A1(S_0_02[13]), .B1(S_0_03[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n19641), .COUT(n19642), .S0(S_1_01_20__N_2205[12]), 
          .S1(S_1_01_20__N_2205[13]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(123[13:48])
    defparam add_836_12.INIT0 = 16'h5666;
    defparam add_836_12.INIT1 = 16'h5666;
    defparam add_836_12.INJECT1_0 = "NO";
    defparam add_836_12.INJECT1_1 = "NO";
    CCU2D add_836_10 (.A0(S_0_02[10]), .B0(S_0_03[8]), .C0(GND_net), .D0(GND_net), 
          .A1(S_0_02[11]), .B1(S_0_03[9]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19640), .COUT(n19641), .S0(S_1_01_20__N_2205[10]), .S1(S_1_01_20__N_2205[11]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(123[13:48])
    defparam add_836_10.INIT0 = 16'h5666;
    defparam add_836_10.INIT1 = 16'h5666;
    defparam add_836_10.INJECT1_0 = "NO";
    defparam add_836_10.INJECT1_1 = "NO";
    CCU2D add_836_8 (.A0(S_0_02[8]), .B0(S_0_03[6]), .C0(GND_net), .D0(GND_net), 
          .A1(S_0_02[9]), .B1(S_0_03[7]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19639), .COUT(n19640), .S0(S_1_01_20__N_2205[8]), .S1(S_1_01_20__N_2205[9]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(123[13:48])
    defparam add_836_8.INIT0 = 16'h5666;
    defparam add_836_8.INIT1 = 16'h5666;
    defparam add_836_8.INJECT1_0 = "NO";
    defparam add_836_8.INJECT1_1 = "NO";
    CCU2D add_836_6 (.A0(S_0_02[6]), .B0(S_0_03[4]), .C0(GND_net), .D0(GND_net), 
          .A1(S_0_02[7]), .B1(S_0_03[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19638), .COUT(n19639), .S0(S_1_01_20__N_2205[6]), .S1(S_1_01_20__N_2205[7]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(123[13:48])
    defparam add_836_6.INIT0 = 16'h5666;
    defparam add_836_6.INIT1 = 16'h5666;
    defparam add_836_6.INJECT1_0 = "NO";
    defparam add_836_6.INJECT1_1 = "NO";
    CCU2D add_836_4 (.A0(S_0_02[4]), .B0(S_0_03[2]), .C0(GND_net), .D0(GND_net), 
          .A1(S_0_02[5]), .B1(S_0_03[3]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19637), .COUT(n19638), .S0(S_1_01_20__N_2205[4]), .S1(S_1_01_20__N_2205[5]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(123[13:48])
    defparam add_836_4.INIT0 = 16'h5666;
    defparam add_836_4.INIT1 = 16'h5666;
    defparam add_836_4.INJECT1_0 = "NO";
    defparam add_836_4.INJECT1_1 = "NO";
    CCU2D add_836_2 (.A0(S_0_02[2]), .B0(S_0_03[0]), .C0(GND_net), .D0(GND_net), 
          .A1(S_0_02[3]), .B1(S_0_03[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n19637), .S1(S_1_01_20__N_2205[3]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(123[13:48])
    defparam add_836_2.INIT0 = 16'h7000;
    defparam add_836_2.INIT1 = 16'h5666;
    defparam add_836_2.INJECT1_0 = "NO";
    defparam add_836_2.INJECT1_1 = "NO";
    CCU2D add_35_22 (.A0(S_2_01[20]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(S_2_01[21]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n19634), .S0(o_p_29__N_2320[28]), .S1(o_p_29__N_2320[29]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(177[13] 178[15])
    defparam add_35_22.INIT0 = 16'hfaaa;
    defparam add_35_22.INIT1 = 16'hfaaa;
    defparam add_35_22.INJECT1_0 = "NO";
    defparam add_35_22.INJECT1_1 = "NO";
    CCU2D add_35_20 (.A0(S_2_01[18]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(S_2_01[19]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n19633), .COUT(n19634), .S0(o_p_29__N_2320[26]), .S1(o_p_29__N_2320[27]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(177[13] 178[15])
    defparam add_35_20.INIT0 = 16'hfaaa;
    defparam add_35_20.INIT1 = 16'hfaaa;
    defparam add_35_20.INJECT1_0 = "NO";
    defparam add_35_20.INJECT1_1 = "NO";
    CCU2D add_35_18 (.A0(S_2_00[24]), .B0(S_2_01[16]), .C0(GND_net), .D0(GND_net), 
          .A1(S_2_00[25]), .B1(S_2_01[17]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19632), .COUT(n19633), .S0(o_p_29__N_2320[24]), .S1(o_p_29__N_2320[25]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(177[13] 178[15])
    defparam add_35_18.INIT0 = 16'h5666;
    defparam add_35_18.INIT1 = 16'h5666;
    defparam add_35_18.INJECT1_0 = "NO";
    defparam add_35_18.INJECT1_1 = "NO";
    CCU2D add_35_16 (.A0(S_2_00[22]), .B0(S_2_01[14]), .C0(GND_net), .D0(GND_net), 
          .A1(S_2_00[23]), .B1(S_2_01[15]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19631), .COUT(n19632), .S0(o_p_29__N_2320[22]), .S1(o_p_29__N_2320[23]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(177[13] 178[15])
    defparam add_35_16.INIT0 = 16'h5666;
    defparam add_35_16.INIT1 = 16'h5666;
    defparam add_35_16.INJECT1_0 = "NO";
    defparam add_35_16.INJECT1_1 = "NO";
    CCU2D add_35_14 (.A0(S_2_00[20]), .B0(S_2_01[12]), .C0(GND_net), .D0(GND_net), 
          .A1(S_2_00[21]), .B1(S_2_01[13]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19630), .COUT(n19631), .S0(o_p_29__N_2320[20]), .S1(o_p_29__N_2320[21]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(177[13] 178[15])
    defparam add_35_14.INIT0 = 16'h5666;
    defparam add_35_14.INIT1 = 16'h5666;
    defparam add_35_14.INJECT1_0 = "NO";
    defparam add_35_14.INJECT1_1 = "NO";
    CCU2D add_35_12 (.A0(S_2_00[18]), .B0(S_2_01[10]), .C0(GND_net), .D0(GND_net), 
          .A1(S_2_00[19]), .B1(S_2_01[11]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19629), .COUT(n19630), .S0(o_p_29__N_2320[18]), .S1(o_p_29__N_2320[19]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(177[13] 178[15])
    defparam add_35_12.INIT0 = 16'h5666;
    defparam add_35_12.INIT1 = 16'h5666;
    defparam add_35_12.INJECT1_0 = "NO";
    defparam add_35_12.INJECT1_1 = "NO";
    CCU2D add_35_10 (.A0(S_2_00[16]), .B0(S_2_01[8]), .C0(GND_net), .D0(GND_net), 
          .A1(S_2_00[17]), .B1(S_2_01[9]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19628), .COUT(n19629), .S0(o_p_29__N_2320[16]), .S1(o_p_29__N_2320[17]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(177[13] 178[15])
    defparam add_35_10.INIT0 = 16'h5666;
    defparam add_35_10.INIT1 = 16'h5666;
    defparam add_35_10.INJECT1_0 = "NO";
    defparam add_35_10.INJECT1_1 = "NO";
    CCU2D add_35_8 (.A0(S_2_00[14]), .B0(S_2_01[6]), .C0(GND_net), .D0(GND_net), 
          .A1(S_2_00[15]), .B1(S_2_01[7]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19627), .COUT(n19628), .S0(o_p_29__N_2320[14]), .S1(o_p_29__N_2320[15]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(177[13] 178[15])
    defparam add_35_8.INIT0 = 16'h5666;
    defparam add_35_8.INIT1 = 16'h5666;
    defparam add_35_8.INJECT1_0 = "NO";
    defparam add_35_8.INJECT1_1 = "NO";
    CCU2D add_35_6 (.A0(S_2_00[12]), .B0(S_2_01[4]), .C0(GND_net), .D0(GND_net), 
          .A1(S_2_00[13]), .B1(S_2_01[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19626), .COUT(n19627), .S0(o_p_29__N_2320[12]), .S1(o_p_29__N_2320[13]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(177[13] 178[15])
    defparam add_35_6.INIT0 = 16'h5666;
    defparam add_35_6.INIT1 = 16'h5666;
    defparam add_35_6.INJECT1_0 = "NO";
    defparam add_35_6.INJECT1_1 = "NO";
    CCU2D add_35_4 (.A0(S_2_00[10]), .B0(S_2_01[2]), .C0(GND_net), .D0(GND_net), 
          .A1(S_2_00[11]), .B1(S_2_01[3]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19625), .COUT(n19626), .S0(o_p_29__N_2320[10]), .S1(o_p_29__N_2320[11]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(177[13] 178[15])
    defparam add_35_4.INIT0 = 16'h5666;
    defparam add_35_4.INIT1 = 16'h5666;
    defparam add_35_4.INJECT1_0 = "NO";
    defparam add_35_4.INJECT1_1 = "NO";
    CCU2D add_35_2 (.A0(S_2_00[8]), .B0(S_2_01[0]), .C0(GND_net), .D0(GND_net), 
          .A1(S_2_00[9]), .B1(S_2_01[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n19625), .S1(o_p_29__N_2320[9]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(177[13] 178[15])
    defparam add_35_2.INIT0 = 16'h7000;
    defparam add_35_2.INIT1 = 16'h5666;
    defparam add_35_2.INJECT1_0 = "NO";
    defparam add_35_2.INJECT1_1 = "NO";
    LUT4 i17608_2_lut (.A(S_2_00[8]), .B(S_2_01[0]), .Z(o_p_29__N_2320[8])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i17608_2_lut.init = 16'h6666;
    LUT4 i17605_2_lut (.A(S_1_02[4]), .B(S_1_03[0]), .Z(S_2_01_25__N_2294[4])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i17605_2_lut.init = 16'h6666;
    LUT4 i17617_2_lut (.A(S_1_00[4]), .B(S_1_01[0]), .Z(S_2_00_25__N_2268[4])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i17617_2_lut.init = 16'h6666;
    LUT4 i17618_2_lut (.A(S_0_04[2]), .B(S_0_05[0]), .Z(S_1_02_20__N_2226[2])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i17618_2_lut.init = 16'h6666;
    LUT4 i17609_2_lut (.A(S_0_02[2]), .B(S_0_03[0]), .Z(S_1_01_20__N_2205[2])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i17609_2_lut.init = 16'h6666;
    LUT4 i17616_2_lut (.A(S_0_00[2]), .B(S_0_01[0]), .Z(S_1_00_20__N_2184[2])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i17616_2_lut.init = 16'h6666;
    FD1S3IX S_3_00__i29 (.D(o_p_29__N_2320[29]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i29.GSR = "DISABLED";
    FD1S3IX S_3_00__i28 (.D(o_p_29__N_2320[28]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i28.GSR = "DISABLED";
    FD1S3IX S_3_00__i27 (.D(o_p_29__N_2320[27]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i27.GSR = "DISABLED";
    FD1S3IX S_3_00__i26 (.D(o_p_29__N_2320[26]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i26.GSR = "DISABLED";
    FD1S3IX S_3_00__i25 (.D(o_p_29__N_2320[25]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i25.GSR = "DISABLED";
    FD1S3IX S_3_00__i24 (.D(o_p_29__N_2320[24]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i24.GSR = "DISABLED";
    FD1S3IX S_3_00__i23 (.D(o_p_29__N_2320[23]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i23.GSR = "DISABLED";
    FD1S3IX S_3_00__i22 (.D(o_p_29__N_2320[22]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i22.GSR = "DISABLED";
    FD1S3IX S_3_00__i21 (.D(o_p_29__N_2320[21]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i21.GSR = "DISABLED";
    FD1S3IX S_3_00__i20 (.D(o_p_29__N_2320[20]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i20.GSR = "DISABLED";
    FD1S3IX S_3_00__i19 (.D(o_p_29__N_2320[19]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i19.GSR = "DISABLED";
    FD1S3IX S_3_00__i18 (.D(o_p_29__N_2320[18]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i18.GSR = "DISABLED";
    FD1S3IX S_3_00__i17 (.D(o_p_29__N_2320[17]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i17.GSR = "DISABLED";
    FD1S3IX S_3_00__i16 (.D(o_p_29__N_2320[16]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i16.GSR = "DISABLED";
    FD1S3IX S_3_00__i15 (.D(o_p_29__N_2320[15]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i15.GSR = "DISABLED";
    FD1S3IX S_3_00__i14 (.D(o_p_29__N_2320[14]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i14.GSR = "DISABLED";
    FD1S3IX S_3_00__i13 (.D(o_p_29__N_2320[13]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i13.GSR = "DISABLED";
    FD1S3IX S_3_00__i12 (.D(o_p_29__N_2320[12]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i12.GSR = "DISABLED";
    FD1S3IX S_3_00__i11 (.D(o_p_29__N_2320[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i11.GSR = "DISABLED";
    FD1S3IX S_3_00__i10 (.D(o_p_29__N_2320[10]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i10.GSR = "DISABLED";
    FD1S3IX S_3_00__i9 (.D(o_p_29__N_2320[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i9.GSR = "DISABLED";
    FD1S3IX S_3_00__i8 (.D(o_p_29__N_2320[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i8.GSR = "DISABLED";
    FD1S3IX S_3_00__i7 (.D(o_p_29__N_2320[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i7.GSR = "DISABLED";
    FD1S3IX S_3_00__i6 (.D(o_p_29__N_2320[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i6.GSR = "DISABLED";
    FD1S3IX S_3_00__i5 (.D(o_p_29__N_2320[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i5.GSR = "DISABLED";
    FD1S3IX S_3_00__i4 (.D(o_p_29__N_2320[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i4.GSR = "DISABLED";
    FD1S3IX S_3_00__i3 (.D(o_p_29__N_2320[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i3.GSR = "DISABLED";
    FD1S3IX S_3_00__i2 (.D(o_p_29__N_2320[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i2.GSR = "DISABLED";
    FD1S3IX S_3_00__i1 (.D(o_p_29__N_2320[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i1.GSR = "DISABLED";
    FD1S3IX S_2_01__i22 (.D(S_2_01_25__N_2294[21]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i22.GSR = "DISABLED";
    FD1S3IX S_2_01__i21 (.D(S_2_01_25__N_2294[20]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i21.GSR = "DISABLED";
    FD1S3IX S_2_01__i20 (.D(S_2_01_25__N_2294[19]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i20.GSR = "DISABLED";
    FD1S3IX S_2_01__i19 (.D(S_2_01_25__N_2294[18]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i19.GSR = "DISABLED";
    FD1S3IX S_2_01__i18 (.D(S_2_01_25__N_2294[17]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i18.GSR = "DISABLED";
    FD1S3IX S_2_01__i17 (.D(S_2_01_25__N_2294[16]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i17.GSR = "DISABLED";
    FD1S3IX S_2_01__i16 (.D(S_2_01_25__N_2294[15]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i16.GSR = "DISABLED";
    FD1S3IX S_2_01__i15 (.D(S_2_01_25__N_2294[14]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i15.GSR = "DISABLED";
    FD1S3IX S_2_01__i14 (.D(S_2_01_25__N_2294[13]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i14.GSR = "DISABLED";
    FD1S3IX S_2_01__i13 (.D(S_2_01_25__N_2294[12]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i13.GSR = "DISABLED";
    FD1S3IX S_2_01__i12 (.D(S_2_01_25__N_2294[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i12.GSR = "DISABLED";
    FD1S3IX S_2_01__i11 (.D(S_2_01_25__N_2294[10]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i11.GSR = "DISABLED";
    FD1S3IX S_2_01__i10 (.D(S_2_01_25__N_2294[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i10.GSR = "DISABLED";
    FD1S3IX S_2_01__i9 (.D(S_2_01_25__N_2294[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i9.GSR = "DISABLED";
    FD1S3IX S_2_01__i8 (.D(S_2_01_25__N_2294[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i8.GSR = "DISABLED";
    FD1S3IX S_2_01__i7 (.D(S_2_01_25__N_2294[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i7.GSR = "DISABLED";
    FD1S3IX S_2_01__i6 (.D(S_2_01_25__N_2294[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i6.GSR = "DISABLED";
    FD1S3IX S_2_01__i5 (.D(S_2_01_25__N_2294[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i5.GSR = "DISABLED";
    FD1S3IX S_2_01__i4 (.D(S_2_01_25__N_2294[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i4.GSR = "DISABLED";
    FD1S3IX S_2_01__i3 (.D(S_2_01_25__N_2294[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i3.GSR = "DISABLED";
    FD1S3IX S_2_01__i2 (.D(S_2_01_25__N_2294[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i2.GSR = "DISABLED";
    FD1S3IX S_2_00__i26 (.D(S_2_00_25__N_2268[25]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i26.GSR = "DISABLED";
    FD1S3IX S_2_00__i25 (.D(S_2_00_25__N_2268[24]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i25.GSR = "DISABLED";
    FD1S3IX S_2_00__i24 (.D(S_2_00_25__N_2268[23]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i24.GSR = "DISABLED";
    FD1S3IX S_2_00__i23 (.D(S_2_00_25__N_2268[22]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i23.GSR = "DISABLED";
    FD1S3IX S_2_00__i22 (.D(S_2_00_25__N_2268[21]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i22.GSR = "DISABLED";
    FD1S3IX S_2_00__i21 (.D(S_2_00_25__N_2268[20]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i21.GSR = "DISABLED";
    FD1S3IX S_2_00__i20 (.D(S_2_00_25__N_2268[19]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i20.GSR = "DISABLED";
    FD1S3IX S_2_00__i19 (.D(S_2_00_25__N_2268[18]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i19.GSR = "DISABLED";
    FD1S3IX S_2_00__i18 (.D(S_2_00_25__N_2268[17]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i18.GSR = "DISABLED";
    FD1S3IX S_2_00__i17 (.D(S_2_00_25__N_2268[16]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i17.GSR = "DISABLED";
    FD1S3IX S_2_00__i16 (.D(S_2_00_25__N_2268[15]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i16.GSR = "DISABLED";
    FD1S3IX S_2_00__i15 (.D(S_2_00_25__N_2268[14]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i15.GSR = "DISABLED";
    FD1S3IX S_2_00__i14 (.D(S_2_00_25__N_2268[13]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i14.GSR = "DISABLED";
    FD1S3IX S_2_00__i13 (.D(S_2_00_25__N_2268[12]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i13.GSR = "DISABLED";
    FD1S3IX S_2_00__i12 (.D(S_2_00_25__N_2268[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i12.GSR = "DISABLED";
    FD1S3IX S_2_00__i11 (.D(S_2_00_25__N_2268[10]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i11.GSR = "DISABLED";
    FD1S3IX S_2_00__i10 (.D(S_2_00_25__N_2268[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i10.GSR = "DISABLED";
    FD1S3IX S_2_00__i9 (.D(S_2_00_25__N_2268[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i9.GSR = "DISABLED";
    FD1S3IX S_2_00__i8 (.D(S_2_00_25__N_2268[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_p_29__N_2320[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i8.GSR = "DISABLED";
    FD1S3IX S_2_00__i7 (.D(S_2_00_25__N_2268[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_p_29__N_2320[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i7.GSR = "DISABLED";
    FD1S3IX S_2_00__i6 (.D(S_2_00_25__N_2268[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_p_29__N_2320[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i6.GSR = "DISABLED";
    FD1S3IX S_2_00__i5 (.D(S_2_00_25__N_2268[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_p_29__N_2320[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i5.GSR = "DISABLED";
    FD1S3IX S_2_00__i4 (.D(S_2_00_25__N_2268[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_p_29__N_2320[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i4.GSR = "DISABLED";
    FD1S3IX S_2_00__i3 (.D(S_2_00_25__N_2268[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_p_29__N_2320[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i3.GSR = "DISABLED";
    FD1S3IX S_2_00__i2 (.D(S_2_00_25__N_2268[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_p_29__N_2320[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i2.GSR = "DISABLED";
    FD1S3IX S_1_03__i18 (.D(S_0_06[17]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_03[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_03__i18.GSR = "DISABLED";
    FD1S3IX S_1_03__i17 (.D(S_0_06[16]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_03[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_03__i17.GSR = "DISABLED";
    FD1S3IX S_1_03__i16 (.D(S_0_06[15]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_03[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_03__i16.GSR = "DISABLED";
    FD1S3IX S_1_03__i15 (.D(S_0_06[14]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_03[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_03__i15.GSR = "DISABLED";
    FD1S3IX S_1_03__i14 (.D(S_0_06[13]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_03[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_03__i14.GSR = "DISABLED";
    FD1S3IX S_1_03__i13 (.D(S_0_06[12]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_03[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_03__i13.GSR = "DISABLED";
    FD1S3IX S_1_03__i12 (.D(S_0_06[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_03[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_03__i12.GSR = "DISABLED";
    FD1S3IX S_1_03__i11 (.D(S_0_06[10]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_03[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_03__i11.GSR = "DISABLED";
    FD1S3IX S_1_03__i10 (.D(S_0_06[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_03[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_03__i10.GSR = "DISABLED";
    FD1S3IX S_1_03__i9 (.D(S_0_06[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_03[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_03__i9.GSR = "DISABLED";
    FD1S3IX S_1_03__i8 (.D(S_0_06[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_03[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_03__i8.GSR = "DISABLED";
    FD1S3IX S_1_03__i7 (.D(S_0_06[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_03[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_03__i7.GSR = "DISABLED";
    FD1S3IX S_1_03__i6 (.D(S_0_06[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_03[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_03__i6.GSR = "DISABLED";
    FD1S3IX S_1_03__i5 (.D(S_0_06[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_03[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_03__i5.GSR = "DISABLED";
    FD1S3IX S_1_03__i4 (.D(S_0_06[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_03[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_03__i4.GSR = "DISABLED";
    FD1S3IX S_1_03__i3 (.D(S_0_06[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_03[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_03__i3.GSR = "DISABLED";
    FD1S3IX S_1_03__i2 (.D(S_0_06[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_03[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_03__i2.GSR = "DISABLED";
    FD1S3IX S_1_02__i21 (.D(S_1_02_20__N_2226[20]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_02[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i21.GSR = "DISABLED";
    FD1S3IX S_1_02__i20 (.D(S_1_02_20__N_2226[19]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_02[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i20.GSR = "DISABLED";
    FD1S3IX S_1_02__i19 (.D(S_1_02_20__N_2226[18]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_02[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i19.GSR = "DISABLED";
    FD1S3IX S_1_02__i18 (.D(S_1_02_20__N_2226[17]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_02[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i18.GSR = "DISABLED";
    FD1S3IX S_1_02__i17 (.D(S_1_02_20__N_2226[16]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_02[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i17.GSR = "DISABLED";
    FD1S3IX S_1_02__i16 (.D(S_1_02_20__N_2226[15]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_02[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i16.GSR = "DISABLED";
    FD1S3IX S_1_02__i15 (.D(S_1_02_20__N_2226[14]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_02[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i15.GSR = "DISABLED";
    FD1S3IX S_1_02__i14 (.D(S_1_02_20__N_2226[13]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_02[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i14.GSR = "DISABLED";
    FD1S3IX S_1_02__i13 (.D(S_1_02_20__N_2226[12]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_02[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i13.GSR = "DISABLED";
    FD1S3IX S_1_02__i12 (.D(S_1_02_20__N_2226[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_02[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i12.GSR = "DISABLED";
    FD1S3IX S_1_02__i11 (.D(S_1_02_20__N_2226[10]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_02[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i11.GSR = "DISABLED";
    FD1S3IX S_1_02__i10 (.D(S_1_02_20__N_2226[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_02[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i10.GSR = "DISABLED";
    FD1S3IX S_1_02__i9 (.D(S_1_02_20__N_2226[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_02[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i9.GSR = "DISABLED";
    FD1S3IX S_1_02__i8 (.D(S_1_02_20__N_2226[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_02[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i8.GSR = "DISABLED";
    FD1S3IX S_1_02__i7 (.D(S_1_02_20__N_2226[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_02[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i7.GSR = "DISABLED";
    FD1S3IX S_1_02__i6 (.D(S_1_02_20__N_2226[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_02[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i6.GSR = "DISABLED";
    FD1S3IX S_1_02__i5 (.D(S_1_02_20__N_2226[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_02[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i5.GSR = "DISABLED";
    FD1S3IX S_1_02__i4 (.D(S_1_02_20__N_2226[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01_25__N_2294[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i4.GSR = "DISABLED";
    FD1S3IX S_1_02__i3 (.D(S_1_02_20__N_2226[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01_25__N_2294[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i3.GSR = "DISABLED";
    FD1S3IX S_1_02__i2 (.D(S_1_02_20__N_2226[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01_25__N_2294[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i2.GSR = "DISABLED";
    FD1S3IX S_1_01__i20 (.D(S_1_01_20__N_2205[20]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i20.GSR = "DISABLED";
    FD1S3IX S_1_01__i19 (.D(S_1_01_20__N_2205[19]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i19.GSR = "DISABLED";
    FD1S3IX S_1_01__i18 (.D(S_1_01_20__N_2205[18]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i18.GSR = "DISABLED";
    FD1S3IX S_1_01__i17 (.D(S_1_01_20__N_2205[17]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i17.GSR = "DISABLED";
    FD1S3IX S_1_01__i16 (.D(S_1_01_20__N_2205[16]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i16.GSR = "DISABLED";
    FD1S3IX S_1_01__i15 (.D(S_1_01_20__N_2205[15]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i15.GSR = "DISABLED";
    FD1S3IX S_1_01__i14 (.D(S_1_01_20__N_2205[14]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i14.GSR = "DISABLED";
    FD1S3IX S_1_01__i13 (.D(S_1_01_20__N_2205[13]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i13.GSR = "DISABLED";
    FD1S3IX S_1_01__i12 (.D(S_1_01_20__N_2205[12]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i12.GSR = "DISABLED";
    FD1S3IX S_1_01__i11 (.D(S_1_01_20__N_2205[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i11.GSR = "DISABLED";
    FD1S3IX S_1_01__i10 (.D(S_1_01_20__N_2205[10]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i10.GSR = "DISABLED";
    FD1S3IX S_1_01__i9 (.D(S_1_01_20__N_2205[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i9.GSR = "DISABLED";
    FD1S3IX S_1_01__i8 (.D(S_1_01_20__N_2205[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i8.GSR = "DISABLED";
    FD1S3IX S_1_01__i7 (.D(S_1_01_20__N_2205[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i7.GSR = "DISABLED";
    FD1S3IX S_1_01__i6 (.D(S_1_01_20__N_2205[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i6.GSR = "DISABLED";
    FD1S3IX S_1_01__i5 (.D(S_1_01_20__N_2205[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i5.GSR = "DISABLED";
    FD1S3IX S_1_01__i4 (.D(S_1_01_20__N_2205[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i4.GSR = "DISABLED";
    FD1S3IX S_1_01__i3 (.D(S_1_01_20__N_2205[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i3.GSR = "DISABLED";
    FD1S3IX S_1_01__i2 (.D(S_1_01_20__N_2205[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i2.GSR = "DISABLED";
    FD1S3IX S_1_01__i1 (.D(S_1_01_20__N_2205[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i1.GSR = "DISABLED";
    FD1S3IX S_1_00__i20 (.D(S_1_00_20__N_2184[20]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_00[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i20.GSR = "DISABLED";
    FD1S3IX S_1_00__i19 (.D(S_1_00_20__N_2184[19]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_00[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i19.GSR = "DISABLED";
    FD1S3IX S_1_00__i18 (.D(S_1_00_20__N_2184[18]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_00[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i18.GSR = "DISABLED";
    FD1S3IX S_1_00__i17 (.D(S_1_00_20__N_2184[17]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_00[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i17.GSR = "DISABLED";
    FD1S3IX S_1_00__i16 (.D(S_1_00_20__N_2184[16]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_00[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i16.GSR = "DISABLED";
    FD1S3IX S_1_00__i15 (.D(S_1_00_20__N_2184[15]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_00[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i15.GSR = "DISABLED";
    FD1S3IX S_1_00__i14 (.D(S_1_00_20__N_2184[14]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_00[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i14.GSR = "DISABLED";
    FD1S3IX S_1_00__i13 (.D(S_1_00_20__N_2184[13]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_00[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i13.GSR = "DISABLED";
    FD1S3IX S_1_00__i12 (.D(S_1_00_20__N_2184[12]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_00[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i12.GSR = "DISABLED";
    FD1S3IX S_1_00__i11 (.D(S_1_00_20__N_2184[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_00[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i11.GSR = "DISABLED";
    FD1S3IX S_1_00__i10 (.D(S_1_00_20__N_2184[10]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_00[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i10.GSR = "DISABLED";
    FD1S3IX S_1_00__i9 (.D(S_1_00_20__N_2184[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_00[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i9.GSR = "DISABLED";
    FD1S3IX S_1_00__i8 (.D(S_1_00_20__N_2184[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_00[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i8.GSR = "DISABLED";
    FD1S3IX S_1_00__i7 (.D(S_1_00_20__N_2184[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_00[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i7.GSR = "DISABLED";
    FD1S3IX S_1_00__i6 (.D(S_1_00_20__N_2184[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_00[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i6.GSR = "DISABLED";
    FD1S3IX S_1_00__i5 (.D(S_1_00_20__N_2184[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_00[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i5.GSR = "DISABLED";
    FD1S3IX S_1_00__i4 (.D(S_1_00_20__N_2184[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_00[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i4.GSR = "DISABLED";
    FD1S3IX S_1_00__i3 (.D(S_1_00_20__N_2184[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00_25__N_2268[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i3.GSR = "DISABLED";
    FD1S3IX S_1_00__i2 (.D(S_1_00_20__N_2184[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00_25__N_2268[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i2.GSR = "DISABLED";
    FD1S3IX S_1_00__i1 (.D(S_1_00_20__N_2184[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00_25__N_2268[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i1.GSR = "DISABLED";
    CCU2D add_411_18 (.A0(S_1_02[20]), .B0(S_1_03[16]), .C0(GND_net), 
          .D0(GND_net), .A1(S_1_03[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n19570), .S0(S_2_01_25__N_2294[20]), .S1(S_2_01_25__N_2294[21]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(153[13:48])
    defparam add_411_18.INIT0 = 16'h5666;
    defparam add_411_18.INIT1 = 16'hfaaa;
    defparam add_411_18.INJECT1_0 = "NO";
    defparam add_411_18.INJECT1_1 = "NO";
    CCU2D add_411_16 (.A0(S_1_02[18]), .B0(S_1_03[14]), .C0(GND_net), 
          .D0(GND_net), .A1(S_1_02[19]), .B1(S_1_03[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n19569), .COUT(n19570), .S0(S_2_01_25__N_2294[18]), 
          .S1(S_2_01_25__N_2294[19]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(153[13:48])
    defparam add_411_16.INIT0 = 16'h5666;
    defparam add_411_16.INIT1 = 16'h5666;
    defparam add_411_16.INJECT1_0 = "NO";
    defparam add_411_16.INJECT1_1 = "NO";
    CCU2D add_411_14 (.A0(S_1_02[16]), .B0(S_1_03[12]), .C0(GND_net), 
          .D0(GND_net), .A1(S_1_02[17]), .B1(S_1_03[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n19568), .COUT(n19569), .S0(S_2_01_25__N_2294[16]), 
          .S1(S_2_01_25__N_2294[17]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(153[13:48])
    defparam add_411_14.INIT0 = 16'h5666;
    defparam add_411_14.INIT1 = 16'h5666;
    defparam add_411_14.INJECT1_0 = "NO";
    defparam add_411_14.INJECT1_1 = "NO";
    CCU2D add_411_12 (.A0(S_1_02[14]), .B0(S_1_03[10]), .C0(GND_net), 
          .D0(GND_net), .A1(S_1_02[15]), .B1(S_1_03[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n19567), .COUT(n19568), .S0(S_2_01_25__N_2294[14]), 
          .S1(S_2_01_25__N_2294[15]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(153[13:48])
    defparam add_411_12.INIT0 = 16'h5666;
    defparam add_411_12.INIT1 = 16'h5666;
    defparam add_411_12.INJECT1_0 = "NO";
    defparam add_411_12.INJECT1_1 = "NO";
    CCU2D add_411_10 (.A0(S_1_02[12]), .B0(S_1_03[8]), .C0(GND_net), .D0(GND_net), 
          .A1(S_1_02[13]), .B1(S_1_03[9]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19566), .COUT(n19567), .S0(S_2_01_25__N_2294[12]), .S1(S_2_01_25__N_2294[13]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(153[13:48])
    defparam add_411_10.INIT0 = 16'h5666;
    defparam add_411_10.INIT1 = 16'h5666;
    defparam add_411_10.INJECT1_0 = "NO";
    defparam add_411_10.INJECT1_1 = "NO";
    CCU2D add_411_8 (.A0(S_1_02[10]), .B0(S_1_03[6]), .C0(GND_net), .D0(GND_net), 
          .A1(S_1_02[11]), .B1(S_1_03[7]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19565), .COUT(n19566), .S0(S_2_01_25__N_2294[10]), .S1(S_2_01_25__N_2294[11]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(153[13:48])
    defparam add_411_8.INIT0 = 16'h5666;
    defparam add_411_8.INIT1 = 16'h5666;
    defparam add_411_8.INJECT1_0 = "NO";
    defparam add_411_8.INJECT1_1 = "NO";
    CCU2D add_411_6 (.A0(S_1_02[8]), .B0(S_1_03[4]), .C0(GND_net), .D0(GND_net), 
          .A1(S_1_02[9]), .B1(S_1_03[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19564), .COUT(n19565), .S0(S_2_01_25__N_2294[8]), .S1(S_2_01_25__N_2294[9]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(153[13:48])
    defparam add_411_6.INIT0 = 16'h5666;
    defparam add_411_6.INIT1 = 16'h5666;
    defparam add_411_6.INJECT1_0 = "NO";
    defparam add_411_6.INJECT1_1 = "NO";
    CCU2D add_411_4 (.A0(S_1_02[6]), .B0(S_1_03[2]), .C0(GND_net), .D0(GND_net), 
          .A1(S_1_02[7]), .B1(S_1_03[3]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19563), .COUT(n19564), .S0(S_2_01_25__N_2294[6]), .S1(S_2_01_25__N_2294[7]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(153[13:48])
    defparam add_411_4.INIT0 = 16'h5666;
    defparam add_411_4.INIT1 = 16'h5666;
    defparam add_411_4.INJECT1_0 = "NO";
    defparam add_411_4.INJECT1_1 = "NO";
    CCU2D add_411_2 (.A0(S_1_02[4]), .B0(S_1_03[0]), .C0(GND_net), .D0(GND_net), 
          .A1(S_1_02[5]), .B1(S_1_03[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n19563), .S1(S_2_01_25__N_2294[5]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(153[13:48])
    defparam add_411_2.INIT0 = 16'h7000;
    defparam add_411_2.INIT1 = 16'h5666;
    defparam add_411_2.INJECT1_0 = "NO";
    defparam add_411_2.INJECT1_1 = "NO";
    \bimpy(BW=16)  initialmpy_6_0 (.S_0_06({S_0_06}), .dac_clk_p_c(dac_clk_p_c), 
            .n14230(n14230), .n9458(n9458), .GND_net(GND_net), .u_l({u_l}), 
            .\u_s[13] (u_s[13]), .\u_s[12] (u_s[12]), .i_sw0_c(i_sw0_c)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(90[14:75])
    \bimpy(BW=16)_U0  initialmpy_5_0 (.S_0_05({S_0_05}), .dac_clk_p_c(dac_clk_p_c), 
            .n14230(n14230), .n9460(n9460), .GND_net(GND_net), .u_l({u_l}), 
            .\u_s[11] (u_s[11]), .\u_s[10] (u_s[10]), .i_sw0_c(i_sw0_c)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(87[14:75])
    \bimpy(BW=16)_U1  initialmpy_4_0 (.\S_0_04[0] (S_0_04[0]), .dac_clk_p_c(dac_clk_p_c), 
            .n14230(n14230), .n9462(n9462), .GND_net(GND_net), .u_l({u_l}), 
            .\u_s[9] (u_s[9]), .\u_s[8] (u_s[8]), .\S_0_04[17] (S_0_04[17]), 
            .i_sw0_c(i_sw0_c), .\S_0_04[16] (S_0_04[16]), .\S_0_04[15] (S_0_04[15]), 
            .\S_0_04[14] (S_0_04[14]), .\S_0_04[13] (S_0_04[13]), .\S_0_04[12] (S_0_04[12]), 
            .\S_0_04[11] (S_0_04[11]), .\S_0_04[10] (S_0_04[10]), .\S_0_04[9] (S_0_04[9]), 
            .\S_0_04[8] (S_0_04[8]), .\S_0_04[7] (S_0_04[7]), .\S_0_04[6] (S_0_04[6]), 
            .\S_0_04[5] (S_0_04[5]), .\S_0_04[4] (S_0_04[4]), .\S_0_04[3] (S_0_04[3]), 
            .\S_0_04[2] (S_0_04[2]), .\S_1_02_20__N_2226[1] (S_1_02_20__N_2226[1])) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(84[14:73])
    \bimpy(BW=16)_U2  initialmpy_3_0 (.u_l({u_l}), .\u_s[6] (u_s[6]), .\u_s[7] (u_s[7]), 
            .S_0_03({S_0_03}), .dac_clk_p_c(dac_clk_p_c), .n14230(n14230), 
            .n9464(n9464), .GND_net(GND_net), .i_sw0_c(i_sw0_c)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(81[14:73])
    \bimpy(BW=16)_U3  initialmpy_2_0 (.\S_0_02[0] (S_0_02[0]), .dac_clk_p_c(dac_clk_p_c), 
            .n14230(n14230), .n9466(n9466), .u_l({u_l}), .\u_s[4] (u_s[4]), 
            .\u_s[5] (u_s[5]), .GND_net(GND_net), .\S_0_02[17] (S_0_02[17]), 
            .i_sw0_c(i_sw0_c), .\S_0_02[16] (S_0_02[16]), .\S_0_02[15] (S_0_02[15]), 
            .\S_0_02[14] (S_0_02[14]), .\S_0_02[13] (S_0_02[13]), .\S_0_02[12] (S_0_02[12]), 
            .\S_0_02[11] (S_0_02[11]), .\S_0_02[10] (S_0_02[10]), .\S_0_02[9] (S_0_02[9]), 
            .\S_0_02[8] (S_0_02[8]), .\S_0_02[7] (S_0_02[7]), .\S_0_02[6] (S_0_02[6]), 
            .\S_0_02[5] (S_0_02[5]), .\S_0_02[4] (S_0_02[4]), .\S_0_02[3] (S_0_02[3]), 
            .\S_0_02[2] (S_0_02[2]), .\S_1_01_20__N_2205[1] (S_1_01_20__N_2205[1])) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(78[14:73])
    \bimpy(BW=16)_U4  initialmpy_1_0 (.S_0_01({S_0_01}), .dac_clk_p_c(dac_clk_p_c), 
            .n14230(n14230), .n9468(n9468), .GND_net(GND_net), .u_l({u_l}), 
            .\u_s[3] (u_s[3]), .\u_s[2] (u_s[2]), .i_sw0_c(i_sw0_c)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(75[14:73])
    \bimpy(BW=16)_U5  initialmpy_0_0 (.\S_0_00[0] (S_0_00[0]), .dac_clk_p_c(dac_clk_p_c), 
            .n14230(n14230), .n9488(n9488), .GND_net(GND_net), .u_l({u_l}), 
            .\u_s[1] (u_s[1]), .\u_s[0] (u_s[0]), .\S_0_00[17] (S_0_00[17]), 
            .i_sw0_c(i_sw0_c), .\S_0_00[16] (S_0_00[16]), .\S_0_00[15] (S_0_00[15]), 
            .\S_0_00[14] (S_0_00[14]), .\S_0_00[13] (S_0_00[13]), .\S_0_00[12] (S_0_00[12]), 
            .\S_0_00[11] (S_0_00[11]), .\S_0_00[10] (S_0_00[10]), .\S_0_00[9] (S_0_00[9]), 
            .\S_0_00[8] (S_0_00[8]), .\S_0_00[7] (S_0_00[7]), .\S_0_00[6] (S_0_00[6]), 
            .\S_0_00[5] (S_0_00[5]), .\S_0_00[4] (S_0_00[4]), .\S_0_00[3] (S_0_00[3]), 
            .\S_0_00[2] (S_0_00[2]), .\S_1_00_20__N_2184[1] (S_1_00_20__N_2184[1])) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(72[14:73])
    
endmodule
//
// Verilog Description of module \bimpy(BW=16) 
//

module \bimpy(BW=16)  (S_0_06, dac_clk_p_c, n14230, n9458, GND_net, 
            u_l, \u_s[13] , \u_s[12] , i_sw0_c) /* synthesis syn_module_defined=1 */ ;
    output [17:0]S_0_06;
    input dac_clk_p_c;
    input n14230;
    input n9458;
    input GND_net;
    input [15:0]u_l;
    input \u_s[13] ;
    input \u_s[12] ;
    input i_sw0_c;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[29:38])
    
    wire n19382;
    wire [17:0]o_r_17__N_2438;
    
    wire n19381;
    wire [14:0]c_15__N_2408;
    wire [14:0]c_15__N_2423;
    
    wire n19380, n19379, n19378, n19377, n19376, n19375, n29289, 
        n29288;
    
    FD1S3IX o_r__i0 (.D(n9458), .CK(dac_clk_p_c), .CD(n14230), .Q(S_0_06[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=90, LSE_RLINE=90 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i0.GSR = "DISABLED";
    CCU2D add_818_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19382), 
          .S0(o_r_17__N_2438[17]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_818_cout.INIT0 = 16'h0000;
    defparam add_818_cout.INIT1 = 16'h0000;
    defparam add_818_cout.INJECT1_0 = "NO";
    defparam add_818_cout.INJECT1_1 = "NO";
    CCU2D add_818_15 (.A0(c_15__N_2408[14]), .B0(c_15__N_2423[14]), .C0(c_15__N_2408[13]), 
          .D0(c_15__N_2423[13]), .A1(u_l[15]), .B1(\u_s[13] ), .C1(c_15__N_2408[14]), 
          .D1(c_15__N_2423[14]), .CIN(n19381), .COUT(n19382), .S0(o_r_17__N_2438[15]), 
          .S1(o_r_17__N_2438[16]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_818_15.INIT0 = 16'h9666;
    defparam add_818_15.INIT1 = 16'h7888;
    defparam add_818_15.INJECT1_0 = "NO";
    defparam add_818_15.INJECT1_1 = "NO";
    CCU2D add_818_13 (.A0(c_15__N_2408[12]), .B0(c_15__N_2423[12]), .C0(c_15__N_2408[11]), 
          .D0(c_15__N_2423[11]), .A1(c_15__N_2408[13]), .B1(c_15__N_2423[13]), 
          .C1(c_15__N_2408[12]), .D1(c_15__N_2423[12]), .CIN(n19380), 
          .COUT(n19381), .S0(o_r_17__N_2438[13]), .S1(o_r_17__N_2438[14]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_818_13.INIT0 = 16'h9666;
    defparam add_818_13.INIT1 = 16'h9666;
    defparam add_818_13.INJECT1_0 = "NO";
    defparam add_818_13.INJECT1_1 = "NO";
    CCU2D add_818_11 (.A0(c_15__N_2408[10]), .B0(c_15__N_2423[10]), .C0(c_15__N_2408[9]), 
          .D0(c_15__N_2423[9]), .A1(c_15__N_2408[11]), .B1(c_15__N_2423[11]), 
          .C1(c_15__N_2408[10]), .D1(c_15__N_2423[10]), .CIN(n19379), 
          .COUT(n19380), .S0(o_r_17__N_2438[11]), .S1(o_r_17__N_2438[12]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_818_11.INIT0 = 16'h9666;
    defparam add_818_11.INIT1 = 16'h9666;
    defparam add_818_11.INJECT1_0 = "NO";
    defparam add_818_11.INJECT1_1 = "NO";
    CCU2D add_818_9 (.A0(c_15__N_2408[8]), .B0(c_15__N_2423[8]), .C0(c_15__N_2408[7]), 
          .D0(c_15__N_2423[7]), .A1(c_15__N_2408[9]), .B1(c_15__N_2423[9]), 
          .C1(c_15__N_2408[8]), .D1(c_15__N_2423[8]), .CIN(n19378), .COUT(n19379), 
          .S0(o_r_17__N_2438[9]), .S1(o_r_17__N_2438[10]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_818_9.INIT0 = 16'h9666;
    defparam add_818_9.INIT1 = 16'h9666;
    defparam add_818_9.INJECT1_0 = "NO";
    defparam add_818_9.INJECT1_1 = "NO";
    CCU2D add_818_7 (.A0(c_15__N_2408[6]), .B0(c_15__N_2423[6]), .C0(c_15__N_2408[5]), 
          .D0(c_15__N_2423[5]), .A1(c_15__N_2408[7]), .B1(c_15__N_2423[7]), 
          .C1(c_15__N_2408[6]), .D1(c_15__N_2423[6]), .CIN(n19377), .COUT(n19378), 
          .S0(o_r_17__N_2438[7]), .S1(o_r_17__N_2438[8]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_818_7.INIT0 = 16'h9666;
    defparam add_818_7.INIT1 = 16'h9666;
    defparam add_818_7.INJECT1_0 = "NO";
    defparam add_818_7.INJECT1_1 = "NO";
    CCU2D add_818_5 (.A0(c_15__N_2408[4]), .B0(c_15__N_2423[4]), .C0(c_15__N_2408[3]), 
          .D0(c_15__N_2423[3]), .A1(c_15__N_2408[5]), .B1(c_15__N_2423[5]), 
          .C1(c_15__N_2408[4]), .D1(c_15__N_2423[4]), .CIN(n19376), .COUT(n19377), 
          .S0(o_r_17__N_2438[5]), .S1(o_r_17__N_2438[6]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_818_5.INIT0 = 16'h9666;
    defparam add_818_5.INIT1 = 16'h9666;
    defparam add_818_5.INJECT1_0 = "NO";
    defparam add_818_5.INJECT1_1 = "NO";
    CCU2D add_818_3 (.A0(c_15__N_2408[2]), .B0(c_15__N_2423[2]), .C0(c_15__N_2408[1]), 
          .D0(c_15__N_2423[1]), .A1(c_15__N_2408[3]), .B1(c_15__N_2423[3]), 
          .C1(c_15__N_2408[2]), .D1(c_15__N_2423[2]), .CIN(n19375), .COUT(n19376), 
          .S0(o_r_17__N_2438[3]), .S1(o_r_17__N_2438[4]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_818_3.INIT0 = 16'h9666;
    defparam add_818_3.INIT1 = 16'h9666;
    defparam add_818_3.INJECT1_0 = "NO";
    defparam add_818_3.INJECT1_1 = "NO";
    CCU2D add_818_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(c_15__N_2408[1]), .B1(c_15__N_2423[1]), .C1(n29289), .D1(n29288), 
          .COUT(n19375), .S1(o_r_17__N_2438[2]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_818_1.INIT0 = 16'hF000;
    defparam add_818_1.INIT1 = 16'h9666;
    defparam add_818_1.INJECT1_0 = "NO";
    defparam add_818_1.INJECT1_1 = "NO";
    LUT4 i13418_2_lut (.A(u_l[14]), .B(\u_s[13] ), .Z(c_15__N_2408[14])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13418_2_lut.init = 16'h8888;
    LUT4 i13404_2_lut (.A(u_l[15]), .B(\u_s[12] ), .Z(c_15__N_2423[14])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13404_2_lut.init = 16'h8888;
    LUT4 i13419_2_lut (.A(u_l[13]), .B(\u_s[13] ), .Z(c_15__N_2408[13])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13419_2_lut.init = 16'h8888;
    LUT4 i13405_2_lut (.A(u_l[14]), .B(\u_s[12] ), .Z(c_15__N_2423[13])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13405_2_lut.init = 16'h8888;
    LUT4 i13420_2_lut (.A(u_l[12]), .B(\u_s[13] ), .Z(c_15__N_2408[12])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13420_2_lut.init = 16'h8888;
    LUT4 i13406_2_lut (.A(u_l[13]), .B(\u_s[12] ), .Z(c_15__N_2423[12])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13406_2_lut.init = 16'h8888;
    LUT4 i13421_2_lut (.A(u_l[11]), .B(\u_s[13] ), .Z(c_15__N_2408[11])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13421_2_lut.init = 16'h8888;
    LUT4 i13407_2_lut (.A(u_l[12]), .B(\u_s[12] ), .Z(c_15__N_2423[11])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13407_2_lut.init = 16'h8888;
    LUT4 i13422_2_lut (.A(u_l[10]), .B(\u_s[13] ), .Z(c_15__N_2408[10])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13422_2_lut.init = 16'h8888;
    LUT4 i13408_2_lut (.A(u_l[11]), .B(\u_s[12] ), .Z(c_15__N_2423[10])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13408_2_lut.init = 16'h8888;
    LUT4 i13423_2_lut (.A(u_l[9]), .B(\u_s[13] ), .Z(c_15__N_2408[9])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13423_2_lut.init = 16'h8888;
    LUT4 i13409_2_lut (.A(u_l[10]), .B(\u_s[12] ), .Z(c_15__N_2423[9])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13409_2_lut.init = 16'h8888;
    LUT4 i13424_2_lut (.A(u_l[8]), .B(\u_s[13] ), .Z(c_15__N_2408[8])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13424_2_lut.init = 16'h8888;
    LUT4 i13410_2_lut (.A(u_l[9]), .B(\u_s[12] ), .Z(c_15__N_2423[8])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13410_2_lut.init = 16'h8888;
    LUT4 i13425_2_lut (.A(u_l[7]), .B(\u_s[13] ), .Z(c_15__N_2408[7])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13425_2_lut.init = 16'h8888;
    LUT4 i13411_2_lut (.A(u_l[8]), .B(\u_s[12] ), .Z(c_15__N_2423[7])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13411_2_lut.init = 16'h8888;
    LUT4 i13426_2_lut (.A(u_l[6]), .B(\u_s[13] ), .Z(c_15__N_2408[6])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13426_2_lut.init = 16'h8888;
    LUT4 i13412_2_lut (.A(u_l[7]), .B(\u_s[12] ), .Z(c_15__N_2423[6])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13412_2_lut.init = 16'h8888;
    LUT4 i13427_2_lut (.A(u_l[5]), .B(\u_s[13] ), .Z(c_15__N_2408[5])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13427_2_lut.init = 16'h8888;
    LUT4 i13413_2_lut (.A(u_l[6]), .B(\u_s[12] ), .Z(c_15__N_2423[5])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13413_2_lut.init = 16'h8888;
    LUT4 i13428_2_lut (.A(u_l[4]), .B(\u_s[13] ), .Z(c_15__N_2408[4])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13428_2_lut.init = 16'h8888;
    LUT4 i13414_2_lut (.A(u_l[5]), .B(\u_s[12] ), .Z(c_15__N_2423[4])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13414_2_lut.init = 16'h8888;
    LUT4 i13429_2_lut (.A(u_l[3]), .B(\u_s[13] ), .Z(c_15__N_2408[3])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13429_2_lut.init = 16'h8888;
    LUT4 i13415_2_lut (.A(u_l[4]), .B(\u_s[12] ), .Z(c_15__N_2423[3])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13415_2_lut.init = 16'h8888;
    LUT4 i13430_2_lut (.A(u_l[2]), .B(\u_s[13] ), .Z(c_15__N_2408[2])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13430_2_lut.init = 16'h8888;
    LUT4 i13416_2_lut (.A(u_l[3]), .B(\u_s[12] ), .Z(c_15__N_2423[2])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13416_2_lut.init = 16'h8888;
    LUT4 i13431_2_lut (.A(u_l[1]), .B(\u_s[13] ), .Z(c_15__N_2408[1])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13431_2_lut.init = 16'h8888;
    LUT4 i13417_2_lut (.A(u_l[2]), .B(\u_s[12] ), .Z(c_15__N_2423[1])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13417_2_lut.init = 16'h8888;
    LUT4 i12501_2_lut_rep_628 (.A(u_l[1]), .B(\u_s[12] ), .Z(n29288)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i12501_2_lut_rep_628.init = 16'h8888;
    LUT4 i12500_2_lut_rep_629 (.A(u_l[0]), .B(\u_s[13] ), .Z(n29289)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(51[18:45])
    defparam i12500_2_lut_rep_629.init = 16'h8888;
    LUT4 w_r_16__I_0_i2_2_lut_3_lut_4_lut (.A(u_l[0]), .B(\u_s[13] ), .C(\u_s[12] ), 
         .D(u_l[1]), .Z(o_r_17__N_2438[1])) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(51[18:45])
    defparam w_r_16__I_0_i2_2_lut_3_lut_4_lut.init = 16'h7888;
    FD1S3IX o_r__i17 (.D(o_r_17__N_2438[17]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_06[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=90, LSE_RLINE=90 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i17.GSR = "DISABLED";
    FD1S3IX o_r__i16 (.D(o_r_17__N_2438[16]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_06[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=90, LSE_RLINE=90 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i16.GSR = "DISABLED";
    FD1S3IX o_r__i15 (.D(o_r_17__N_2438[15]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_06[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=90, LSE_RLINE=90 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i15.GSR = "DISABLED";
    FD1S3IX o_r__i14 (.D(o_r_17__N_2438[14]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_06[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=90, LSE_RLINE=90 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i14.GSR = "DISABLED";
    FD1S3IX o_r__i13 (.D(o_r_17__N_2438[13]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_06[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=90, LSE_RLINE=90 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i13.GSR = "DISABLED";
    FD1S3IX o_r__i12 (.D(o_r_17__N_2438[12]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_06[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=90, LSE_RLINE=90 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i12.GSR = "DISABLED";
    FD1S3IX o_r__i11 (.D(o_r_17__N_2438[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_06[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=90, LSE_RLINE=90 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i11.GSR = "DISABLED";
    FD1S3IX o_r__i10 (.D(o_r_17__N_2438[10]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_06[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=90, LSE_RLINE=90 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i10.GSR = "DISABLED";
    FD1S3IX o_r__i9 (.D(o_r_17__N_2438[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_06[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=90, LSE_RLINE=90 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i9.GSR = "DISABLED";
    FD1S3IX o_r__i8 (.D(o_r_17__N_2438[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_06[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=90, LSE_RLINE=90 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i8.GSR = "DISABLED";
    FD1S3IX o_r__i7 (.D(o_r_17__N_2438[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_06[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=90, LSE_RLINE=90 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i7.GSR = "DISABLED";
    FD1S3IX o_r__i6 (.D(o_r_17__N_2438[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_06[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=90, LSE_RLINE=90 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i6.GSR = "DISABLED";
    FD1S3IX o_r__i5 (.D(o_r_17__N_2438[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_06[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=90, LSE_RLINE=90 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i5.GSR = "DISABLED";
    FD1S3IX o_r__i4 (.D(o_r_17__N_2438[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_06[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=90, LSE_RLINE=90 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i4.GSR = "DISABLED";
    FD1S3IX o_r__i3 (.D(o_r_17__N_2438[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_06[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=90, LSE_RLINE=90 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i3.GSR = "DISABLED";
    FD1S3IX o_r__i2 (.D(o_r_17__N_2438[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_06[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=90, LSE_RLINE=90 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i2.GSR = "DISABLED";
    FD1S3IX o_r__i1 (.D(o_r_17__N_2438[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_06[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=90, LSE_RLINE=90 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i1.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module \bimpy(BW=16)_U0 
//

module \bimpy(BW=16)_U0  (S_0_05, dac_clk_p_c, n14230, n9460, GND_net, 
            u_l, \u_s[11] , \u_s[10] , i_sw0_c) /* synthesis syn_module_defined=1 */ ;
    output [17:0]S_0_05;
    input dac_clk_p_c;
    input n14230;
    input n9460;
    input GND_net;
    input [15:0]u_l;
    input \u_s[11] ;
    input \u_s[10] ;
    input i_sw0_c;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[29:38])
    
    wire n19487;
    wire [17:0]o_r_17__N_2438;
    
    wire n19486;
    wire [14:0]c_15__N_2408;
    wire [14:0]c_15__N_2423;
    
    wire n19485, n19484, n19483, n19482, n19481, n19480, n29270, 
        n29269;
    
    FD1S3IX o_r__i0 (.D(n9460), .CK(dac_clk_p_c), .CD(n14230), .Q(S_0_05[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=87, LSE_RLINE=87 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i0.GSR = "DISABLED";
    CCU2D add_826_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19487), 
          .S0(o_r_17__N_2438[17]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_826_cout.INIT0 = 16'h0000;
    defparam add_826_cout.INIT1 = 16'h0000;
    defparam add_826_cout.INJECT1_0 = "NO";
    defparam add_826_cout.INJECT1_1 = "NO";
    CCU2D add_826_15 (.A0(c_15__N_2408[14]), .B0(c_15__N_2423[14]), .C0(c_15__N_2408[13]), 
          .D0(c_15__N_2423[13]), .A1(u_l[15]), .B1(\u_s[11] ), .C1(c_15__N_2408[14]), 
          .D1(c_15__N_2423[14]), .CIN(n19486), .COUT(n19487), .S0(o_r_17__N_2438[15]), 
          .S1(o_r_17__N_2438[16]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_826_15.INIT0 = 16'h9666;
    defparam add_826_15.INIT1 = 16'h7888;
    defparam add_826_15.INJECT1_0 = "NO";
    defparam add_826_15.INJECT1_1 = "NO";
    CCU2D add_826_13 (.A0(c_15__N_2408[12]), .B0(c_15__N_2423[12]), .C0(c_15__N_2408[11]), 
          .D0(c_15__N_2423[11]), .A1(c_15__N_2408[13]), .B1(c_15__N_2423[13]), 
          .C1(c_15__N_2408[12]), .D1(c_15__N_2423[12]), .CIN(n19485), 
          .COUT(n19486), .S0(o_r_17__N_2438[13]), .S1(o_r_17__N_2438[14]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_826_13.INIT0 = 16'h9666;
    defparam add_826_13.INIT1 = 16'h9666;
    defparam add_826_13.INJECT1_0 = "NO";
    defparam add_826_13.INJECT1_1 = "NO";
    CCU2D add_826_11 (.A0(c_15__N_2408[10]), .B0(c_15__N_2423[10]), .C0(c_15__N_2408[9]), 
          .D0(c_15__N_2423[9]), .A1(c_15__N_2408[11]), .B1(c_15__N_2423[11]), 
          .C1(c_15__N_2408[10]), .D1(c_15__N_2423[10]), .CIN(n19484), 
          .COUT(n19485), .S0(o_r_17__N_2438[11]), .S1(o_r_17__N_2438[12]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_826_11.INIT0 = 16'h9666;
    defparam add_826_11.INIT1 = 16'h9666;
    defparam add_826_11.INJECT1_0 = "NO";
    defparam add_826_11.INJECT1_1 = "NO";
    CCU2D add_826_9 (.A0(c_15__N_2408[8]), .B0(c_15__N_2423[8]), .C0(c_15__N_2408[7]), 
          .D0(c_15__N_2423[7]), .A1(c_15__N_2408[9]), .B1(c_15__N_2423[9]), 
          .C1(c_15__N_2408[8]), .D1(c_15__N_2423[8]), .CIN(n19483), .COUT(n19484), 
          .S0(o_r_17__N_2438[9]), .S1(o_r_17__N_2438[10]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_826_9.INIT0 = 16'h9666;
    defparam add_826_9.INIT1 = 16'h9666;
    defparam add_826_9.INJECT1_0 = "NO";
    defparam add_826_9.INJECT1_1 = "NO";
    CCU2D add_826_7 (.A0(c_15__N_2408[6]), .B0(c_15__N_2423[6]), .C0(c_15__N_2408[5]), 
          .D0(c_15__N_2423[5]), .A1(c_15__N_2408[7]), .B1(c_15__N_2423[7]), 
          .C1(c_15__N_2408[6]), .D1(c_15__N_2423[6]), .CIN(n19482), .COUT(n19483), 
          .S0(o_r_17__N_2438[7]), .S1(o_r_17__N_2438[8]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_826_7.INIT0 = 16'h9666;
    defparam add_826_7.INIT1 = 16'h9666;
    defparam add_826_7.INJECT1_0 = "NO";
    defparam add_826_7.INJECT1_1 = "NO";
    CCU2D add_826_5 (.A0(c_15__N_2408[4]), .B0(c_15__N_2423[4]), .C0(c_15__N_2408[3]), 
          .D0(c_15__N_2423[3]), .A1(c_15__N_2408[5]), .B1(c_15__N_2423[5]), 
          .C1(c_15__N_2408[4]), .D1(c_15__N_2423[4]), .CIN(n19481), .COUT(n19482), 
          .S0(o_r_17__N_2438[5]), .S1(o_r_17__N_2438[6]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_826_5.INIT0 = 16'h9666;
    defparam add_826_5.INIT1 = 16'h9666;
    defparam add_826_5.INJECT1_0 = "NO";
    defparam add_826_5.INJECT1_1 = "NO";
    CCU2D add_826_3 (.A0(c_15__N_2408[2]), .B0(c_15__N_2423[2]), .C0(c_15__N_2408[1]), 
          .D0(c_15__N_2423[1]), .A1(c_15__N_2408[3]), .B1(c_15__N_2423[3]), 
          .C1(c_15__N_2408[2]), .D1(c_15__N_2423[2]), .CIN(n19480), .COUT(n19481), 
          .S0(o_r_17__N_2438[3]), .S1(o_r_17__N_2438[4]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_826_3.INIT0 = 16'h9666;
    defparam add_826_3.INIT1 = 16'h9666;
    defparam add_826_3.INJECT1_0 = "NO";
    defparam add_826_3.INJECT1_1 = "NO";
    CCU2D add_826_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(c_15__N_2408[1]), .B1(c_15__N_2423[1]), .C1(n29270), .D1(n29269), 
          .COUT(n19480), .S1(o_r_17__N_2438[2]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_826_1.INIT0 = 16'hF000;
    defparam add_826_1.INIT1 = 16'h9666;
    defparam add_826_1.INJECT1_0 = "NO";
    defparam add_826_1.INJECT1_1 = "NO";
    LUT4 i13450_2_lut (.A(u_l[14]), .B(\u_s[11] ), .Z(c_15__N_2408[14])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13450_2_lut.init = 16'h8888;
    LUT4 i13435_2_lut (.A(u_l[15]), .B(\u_s[10] ), .Z(c_15__N_2423[14])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13435_2_lut.init = 16'h8888;
    LUT4 i13451_2_lut (.A(u_l[13]), .B(\u_s[11] ), .Z(c_15__N_2408[13])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13451_2_lut.init = 16'h8888;
    LUT4 i13436_2_lut (.A(u_l[14]), .B(\u_s[10] ), .Z(c_15__N_2423[13])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13436_2_lut.init = 16'h8888;
    LUT4 i13452_2_lut (.A(u_l[12]), .B(\u_s[11] ), .Z(c_15__N_2408[12])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13452_2_lut.init = 16'h8888;
    LUT4 i13437_2_lut (.A(u_l[13]), .B(\u_s[10] ), .Z(c_15__N_2423[12])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13437_2_lut.init = 16'h8888;
    LUT4 i13453_2_lut (.A(u_l[11]), .B(\u_s[11] ), .Z(c_15__N_2408[11])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13453_2_lut.init = 16'h8888;
    LUT4 i13438_2_lut (.A(u_l[12]), .B(\u_s[10] ), .Z(c_15__N_2423[11])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13438_2_lut.init = 16'h8888;
    LUT4 i13454_2_lut (.A(u_l[10]), .B(\u_s[11] ), .Z(c_15__N_2408[10])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13454_2_lut.init = 16'h8888;
    LUT4 i13439_2_lut (.A(u_l[11]), .B(\u_s[10] ), .Z(c_15__N_2423[10])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13439_2_lut.init = 16'h8888;
    LUT4 i13455_2_lut (.A(u_l[9]), .B(\u_s[11] ), .Z(c_15__N_2408[9])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13455_2_lut.init = 16'h8888;
    LUT4 i13440_2_lut (.A(u_l[10]), .B(\u_s[10] ), .Z(c_15__N_2423[9])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13440_2_lut.init = 16'h8888;
    LUT4 i13456_2_lut (.A(u_l[8]), .B(\u_s[11] ), .Z(c_15__N_2408[8])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13456_2_lut.init = 16'h8888;
    LUT4 i13441_2_lut (.A(u_l[9]), .B(\u_s[10] ), .Z(c_15__N_2423[8])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13441_2_lut.init = 16'h8888;
    LUT4 i13457_2_lut (.A(u_l[7]), .B(\u_s[11] ), .Z(c_15__N_2408[7])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13457_2_lut.init = 16'h8888;
    LUT4 i13442_2_lut (.A(u_l[8]), .B(\u_s[10] ), .Z(c_15__N_2423[7])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13442_2_lut.init = 16'h8888;
    LUT4 i13458_2_lut (.A(u_l[6]), .B(\u_s[11] ), .Z(c_15__N_2408[6])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13458_2_lut.init = 16'h8888;
    LUT4 i13443_2_lut (.A(u_l[7]), .B(\u_s[10] ), .Z(c_15__N_2423[6])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13443_2_lut.init = 16'h8888;
    LUT4 i13459_2_lut (.A(u_l[5]), .B(\u_s[11] ), .Z(c_15__N_2408[5])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13459_2_lut.init = 16'h8888;
    LUT4 i13444_2_lut (.A(u_l[6]), .B(\u_s[10] ), .Z(c_15__N_2423[5])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13444_2_lut.init = 16'h8888;
    LUT4 i13460_2_lut (.A(u_l[4]), .B(\u_s[11] ), .Z(c_15__N_2408[4])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13460_2_lut.init = 16'h8888;
    LUT4 i13445_2_lut (.A(u_l[5]), .B(\u_s[10] ), .Z(c_15__N_2423[4])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13445_2_lut.init = 16'h8888;
    LUT4 i13461_2_lut (.A(u_l[3]), .B(\u_s[11] ), .Z(c_15__N_2408[3])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13461_2_lut.init = 16'h8888;
    LUT4 i13446_2_lut (.A(u_l[4]), .B(\u_s[10] ), .Z(c_15__N_2423[3])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13446_2_lut.init = 16'h8888;
    LUT4 i13462_2_lut (.A(u_l[2]), .B(\u_s[11] ), .Z(c_15__N_2408[2])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13462_2_lut.init = 16'h8888;
    LUT4 i13448_2_lut (.A(u_l[3]), .B(\u_s[10] ), .Z(c_15__N_2423[2])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13448_2_lut.init = 16'h8888;
    LUT4 i13463_2_lut (.A(u_l[1]), .B(\u_s[11] ), .Z(c_15__N_2408[1])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13463_2_lut.init = 16'h8888;
    LUT4 i13449_2_lut (.A(u_l[2]), .B(\u_s[10] ), .Z(c_15__N_2423[1])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13449_2_lut.init = 16'h8888;
    FD1S3IX o_r__i17 (.D(o_r_17__N_2438[17]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_05[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=87, LSE_RLINE=87 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i17.GSR = "DISABLED";
    FD1S3IX o_r__i16 (.D(o_r_17__N_2438[16]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_05[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=87, LSE_RLINE=87 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i16.GSR = "DISABLED";
    FD1S3IX o_r__i15 (.D(o_r_17__N_2438[15]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_05[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=87, LSE_RLINE=87 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i15.GSR = "DISABLED";
    FD1S3IX o_r__i14 (.D(o_r_17__N_2438[14]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_05[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=87, LSE_RLINE=87 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i14.GSR = "DISABLED";
    FD1S3IX o_r__i13 (.D(o_r_17__N_2438[13]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_05[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=87, LSE_RLINE=87 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i13.GSR = "DISABLED";
    FD1S3IX o_r__i12 (.D(o_r_17__N_2438[12]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_05[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=87, LSE_RLINE=87 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i12.GSR = "DISABLED";
    FD1S3IX o_r__i11 (.D(o_r_17__N_2438[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_05[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=87, LSE_RLINE=87 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i11.GSR = "DISABLED";
    FD1S3IX o_r__i10 (.D(o_r_17__N_2438[10]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_05[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=87, LSE_RLINE=87 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i10.GSR = "DISABLED";
    FD1S3IX o_r__i9 (.D(o_r_17__N_2438[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_05[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=87, LSE_RLINE=87 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i9.GSR = "DISABLED";
    FD1S3IX o_r__i8 (.D(o_r_17__N_2438[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_05[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=87, LSE_RLINE=87 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i8.GSR = "DISABLED";
    FD1S3IX o_r__i7 (.D(o_r_17__N_2438[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_05[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=87, LSE_RLINE=87 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i7.GSR = "DISABLED";
    FD1S3IX o_r__i6 (.D(o_r_17__N_2438[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_05[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=87, LSE_RLINE=87 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i6.GSR = "DISABLED";
    FD1S3IX o_r__i5 (.D(o_r_17__N_2438[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_05[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=87, LSE_RLINE=87 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i5.GSR = "DISABLED";
    FD1S3IX o_r__i4 (.D(o_r_17__N_2438[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_05[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=87, LSE_RLINE=87 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i4.GSR = "DISABLED";
    FD1S3IX o_r__i3 (.D(o_r_17__N_2438[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_05[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=87, LSE_RLINE=87 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i3.GSR = "DISABLED";
    FD1S3IX o_r__i2 (.D(o_r_17__N_2438[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_05[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=87, LSE_RLINE=87 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i2.GSR = "DISABLED";
    FD1S3IX o_r__i1 (.D(o_r_17__N_2438[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_05[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=87, LSE_RLINE=87 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i1.GSR = "DISABLED";
    LUT4 i12499_2_lut_rep_609 (.A(u_l[1]), .B(\u_s[10] ), .Z(n29269)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i12499_2_lut_rep_609.init = 16'h8888;
    LUT4 i12498_2_lut_rep_610 (.A(u_l[0]), .B(\u_s[11] ), .Z(n29270)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(51[18:45])
    defparam i12498_2_lut_rep_610.init = 16'h8888;
    LUT4 w_r_16__I_0_i2_2_lut_3_lut_4_lut (.A(u_l[0]), .B(\u_s[11] ), .C(\u_s[10] ), 
         .D(u_l[1]), .Z(o_r_17__N_2438[1])) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(51[18:45])
    defparam w_r_16__I_0_i2_2_lut_3_lut_4_lut.init = 16'h7888;
    
endmodule
//
// Verilog Description of module \bimpy(BW=16)_U1 
//

module \bimpy(BW=16)_U1  (\S_0_04[0] , dac_clk_p_c, n14230, n9462, GND_net, 
            u_l, \u_s[9] , \u_s[8] , \S_0_04[17] , i_sw0_c, \S_0_04[16] , 
            \S_0_04[15] , \S_0_04[14] , \S_0_04[13] , \S_0_04[12] , 
            \S_0_04[11] , \S_0_04[10] , \S_0_04[9] , \S_0_04[8] , \S_0_04[7] , 
            \S_0_04[6] , \S_0_04[5] , \S_0_04[4] , \S_0_04[3] , \S_0_04[2] , 
            \S_1_02_20__N_2226[1] ) /* synthesis syn_module_defined=1 */ ;
    output \S_0_04[0] ;
    input dac_clk_p_c;
    input n14230;
    input n9462;
    input GND_net;
    input [15:0]u_l;
    input \u_s[9] ;
    input \u_s[8] ;
    output \S_0_04[17] ;
    input i_sw0_c;
    output \S_0_04[16] ;
    output \S_0_04[15] ;
    output \S_0_04[14] ;
    output \S_0_04[13] ;
    output \S_0_04[12] ;
    output \S_0_04[11] ;
    output \S_0_04[10] ;
    output \S_0_04[9] ;
    output \S_0_04[8] ;
    output \S_0_04[7] ;
    output \S_0_04[6] ;
    output \S_0_04[5] ;
    output \S_0_04[4] ;
    output \S_0_04[3] ;
    output \S_0_04[2] ;
    output \S_1_02_20__N_2226[1] ;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[29:38])
    
    wire n19495;
    wire [17:0]o_r_17__N_2438;
    
    wire n19494;
    wire [14:0]c_15__N_2408;
    wire [14:0]c_15__N_2423;
    
    wire n19493, n19492, n19491, n19490, n19489, n19488, n29273, 
        n29272;
    
    FD1S3IX o_r__i0 (.D(n9462), .CK(dac_clk_p_c), .CD(n14230), .Q(\S_0_04[0] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=84, LSE_RLINE=84 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i0.GSR = "DISABLED";
    CCU2D add_827_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19495), 
          .S0(o_r_17__N_2438[17]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_827_cout.INIT0 = 16'h0000;
    defparam add_827_cout.INIT1 = 16'h0000;
    defparam add_827_cout.INJECT1_0 = "NO";
    defparam add_827_cout.INJECT1_1 = "NO";
    CCU2D add_827_15 (.A0(c_15__N_2408[14]), .B0(c_15__N_2423[14]), .C0(c_15__N_2408[13]), 
          .D0(c_15__N_2423[13]), .A1(u_l[15]), .B1(\u_s[9] ), .C1(c_15__N_2408[14]), 
          .D1(c_15__N_2423[14]), .CIN(n19494), .COUT(n19495), .S0(o_r_17__N_2438[15]), 
          .S1(o_r_17__N_2438[16]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_827_15.INIT0 = 16'h9666;
    defparam add_827_15.INIT1 = 16'h7888;
    defparam add_827_15.INJECT1_0 = "NO";
    defparam add_827_15.INJECT1_1 = "NO";
    CCU2D add_827_13 (.A0(c_15__N_2408[12]), .B0(c_15__N_2423[12]), .C0(c_15__N_2408[11]), 
          .D0(c_15__N_2423[11]), .A1(c_15__N_2408[13]), .B1(c_15__N_2423[13]), 
          .C1(c_15__N_2408[12]), .D1(c_15__N_2423[12]), .CIN(n19493), 
          .COUT(n19494), .S0(o_r_17__N_2438[13]), .S1(o_r_17__N_2438[14]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_827_13.INIT0 = 16'h9666;
    defparam add_827_13.INIT1 = 16'h9666;
    defparam add_827_13.INJECT1_0 = "NO";
    defparam add_827_13.INJECT1_1 = "NO";
    CCU2D add_827_11 (.A0(c_15__N_2408[10]), .B0(c_15__N_2423[10]), .C0(c_15__N_2408[9]), 
          .D0(c_15__N_2423[9]), .A1(c_15__N_2408[11]), .B1(c_15__N_2423[11]), 
          .C1(c_15__N_2408[10]), .D1(c_15__N_2423[10]), .CIN(n19492), 
          .COUT(n19493), .S0(o_r_17__N_2438[11]), .S1(o_r_17__N_2438[12]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_827_11.INIT0 = 16'h9666;
    defparam add_827_11.INIT1 = 16'h9666;
    defparam add_827_11.INJECT1_0 = "NO";
    defparam add_827_11.INJECT1_1 = "NO";
    CCU2D add_827_9 (.A0(c_15__N_2408[8]), .B0(c_15__N_2423[8]), .C0(c_15__N_2408[7]), 
          .D0(c_15__N_2423[7]), .A1(c_15__N_2408[9]), .B1(c_15__N_2423[9]), 
          .C1(c_15__N_2408[8]), .D1(c_15__N_2423[8]), .CIN(n19491), .COUT(n19492), 
          .S0(o_r_17__N_2438[9]), .S1(o_r_17__N_2438[10]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_827_9.INIT0 = 16'h9666;
    defparam add_827_9.INIT1 = 16'h9666;
    defparam add_827_9.INJECT1_0 = "NO";
    defparam add_827_9.INJECT1_1 = "NO";
    CCU2D add_827_7 (.A0(c_15__N_2408[6]), .B0(c_15__N_2423[6]), .C0(c_15__N_2408[5]), 
          .D0(c_15__N_2423[5]), .A1(c_15__N_2408[7]), .B1(c_15__N_2423[7]), 
          .C1(c_15__N_2408[6]), .D1(c_15__N_2423[6]), .CIN(n19490), .COUT(n19491), 
          .S0(o_r_17__N_2438[7]), .S1(o_r_17__N_2438[8]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_827_7.INIT0 = 16'h9666;
    defparam add_827_7.INIT1 = 16'h9666;
    defparam add_827_7.INJECT1_0 = "NO";
    defparam add_827_7.INJECT1_1 = "NO";
    CCU2D add_827_5 (.A0(c_15__N_2408[4]), .B0(c_15__N_2423[4]), .C0(c_15__N_2408[3]), 
          .D0(c_15__N_2423[3]), .A1(c_15__N_2408[5]), .B1(c_15__N_2423[5]), 
          .C1(c_15__N_2408[4]), .D1(c_15__N_2423[4]), .CIN(n19489), .COUT(n19490), 
          .S0(o_r_17__N_2438[5]), .S1(o_r_17__N_2438[6]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_827_5.INIT0 = 16'h9666;
    defparam add_827_5.INIT1 = 16'h9666;
    defparam add_827_5.INJECT1_0 = "NO";
    defparam add_827_5.INJECT1_1 = "NO";
    CCU2D add_827_3 (.A0(c_15__N_2408[2]), .B0(c_15__N_2423[2]), .C0(c_15__N_2408[1]), 
          .D0(c_15__N_2423[1]), .A1(c_15__N_2408[3]), .B1(c_15__N_2423[3]), 
          .C1(c_15__N_2408[2]), .D1(c_15__N_2423[2]), .CIN(n19488), .COUT(n19489), 
          .S0(o_r_17__N_2438[3]), .S1(o_r_17__N_2438[4]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_827_3.INIT0 = 16'h9666;
    defparam add_827_3.INIT1 = 16'h9666;
    defparam add_827_3.INJECT1_0 = "NO";
    defparam add_827_3.INJECT1_1 = "NO";
    CCU2D add_827_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(c_15__N_2408[1]), .B1(c_15__N_2423[1]), .C1(n29273), .D1(n29272), 
          .COUT(n19488), .S1(o_r_17__N_2438[2]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_827_1.INIT0 = 16'hF000;
    defparam add_827_1.INIT1 = 16'h9666;
    defparam add_827_1.INJECT1_0 = "NO";
    defparam add_827_1.INJECT1_1 = "NO";
    LUT4 i13481_2_lut (.A(u_l[14]), .B(\u_s[9] ), .Z(c_15__N_2408[14])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13481_2_lut.init = 16'h8888;
    LUT4 i13467_2_lut (.A(u_l[15]), .B(\u_s[8] ), .Z(c_15__N_2423[14])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13467_2_lut.init = 16'h8888;
    LUT4 i13482_2_lut (.A(u_l[13]), .B(\u_s[9] ), .Z(c_15__N_2408[13])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13482_2_lut.init = 16'h8888;
    LUT4 i13468_2_lut (.A(u_l[14]), .B(\u_s[8] ), .Z(c_15__N_2423[13])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13468_2_lut.init = 16'h8888;
    LUT4 i13483_2_lut (.A(u_l[12]), .B(\u_s[9] ), .Z(c_15__N_2408[12])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13483_2_lut.init = 16'h8888;
    LUT4 i13469_2_lut (.A(u_l[13]), .B(\u_s[8] ), .Z(c_15__N_2423[12])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13469_2_lut.init = 16'h8888;
    LUT4 i13484_2_lut (.A(u_l[11]), .B(\u_s[9] ), .Z(c_15__N_2408[11])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13484_2_lut.init = 16'h8888;
    LUT4 i13470_2_lut (.A(u_l[12]), .B(\u_s[8] ), .Z(c_15__N_2423[11])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13470_2_lut.init = 16'h8888;
    LUT4 i13485_2_lut (.A(u_l[10]), .B(\u_s[9] ), .Z(c_15__N_2408[10])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13485_2_lut.init = 16'h8888;
    LUT4 i13471_2_lut (.A(u_l[11]), .B(\u_s[8] ), .Z(c_15__N_2423[10])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13471_2_lut.init = 16'h8888;
    LUT4 i13486_2_lut (.A(u_l[9]), .B(\u_s[9] ), .Z(c_15__N_2408[9])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13486_2_lut.init = 16'h8888;
    LUT4 i13472_2_lut (.A(u_l[10]), .B(\u_s[8] ), .Z(c_15__N_2423[9])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13472_2_lut.init = 16'h8888;
    LUT4 i13487_2_lut (.A(u_l[8]), .B(\u_s[9] ), .Z(c_15__N_2408[8])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13487_2_lut.init = 16'h8888;
    LUT4 i13473_2_lut (.A(u_l[9]), .B(\u_s[8] ), .Z(c_15__N_2423[8])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13473_2_lut.init = 16'h8888;
    LUT4 i13488_2_lut (.A(u_l[7]), .B(\u_s[9] ), .Z(c_15__N_2408[7])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13488_2_lut.init = 16'h8888;
    LUT4 i13474_2_lut (.A(u_l[8]), .B(\u_s[8] ), .Z(c_15__N_2423[7])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13474_2_lut.init = 16'h8888;
    LUT4 i13489_2_lut (.A(u_l[6]), .B(\u_s[9] ), .Z(c_15__N_2408[6])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13489_2_lut.init = 16'h8888;
    LUT4 i13475_2_lut (.A(u_l[7]), .B(\u_s[8] ), .Z(c_15__N_2423[6])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13475_2_lut.init = 16'h8888;
    LUT4 i13490_2_lut (.A(u_l[5]), .B(\u_s[9] ), .Z(c_15__N_2408[5])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13490_2_lut.init = 16'h8888;
    LUT4 i13476_2_lut (.A(u_l[6]), .B(\u_s[8] ), .Z(c_15__N_2423[5])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13476_2_lut.init = 16'h8888;
    LUT4 i13491_2_lut (.A(u_l[4]), .B(\u_s[9] ), .Z(c_15__N_2408[4])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13491_2_lut.init = 16'h8888;
    LUT4 i13477_2_lut (.A(u_l[5]), .B(\u_s[8] ), .Z(c_15__N_2423[4])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13477_2_lut.init = 16'h8888;
    LUT4 i13492_2_lut (.A(u_l[3]), .B(\u_s[9] ), .Z(c_15__N_2408[3])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13492_2_lut.init = 16'h8888;
    LUT4 i13478_2_lut (.A(u_l[4]), .B(\u_s[8] ), .Z(c_15__N_2423[3])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13478_2_lut.init = 16'h8888;
    LUT4 i13493_2_lut (.A(u_l[2]), .B(\u_s[9] ), .Z(c_15__N_2408[2])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13493_2_lut.init = 16'h8888;
    LUT4 i13479_2_lut (.A(u_l[3]), .B(\u_s[8] ), .Z(c_15__N_2423[2])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13479_2_lut.init = 16'h8888;
    LUT4 i13494_2_lut (.A(u_l[1]), .B(\u_s[9] ), .Z(c_15__N_2408[1])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13494_2_lut.init = 16'h8888;
    LUT4 i13480_2_lut (.A(u_l[2]), .B(\u_s[8] ), .Z(c_15__N_2423[1])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13480_2_lut.init = 16'h8888;
    FD1S3IX o_r__i17 (.D(o_r_17__N_2438[17]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_04[17] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=84, LSE_RLINE=84 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i17.GSR = "DISABLED";
    FD1S3IX o_r__i16 (.D(o_r_17__N_2438[16]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_04[16] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=84, LSE_RLINE=84 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i16.GSR = "DISABLED";
    FD1S3IX o_r__i15 (.D(o_r_17__N_2438[15]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_04[15] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=84, LSE_RLINE=84 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i15.GSR = "DISABLED";
    FD1S3IX o_r__i14 (.D(o_r_17__N_2438[14]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_04[14] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=84, LSE_RLINE=84 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i14.GSR = "DISABLED";
    FD1S3IX o_r__i13 (.D(o_r_17__N_2438[13]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_04[13] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=84, LSE_RLINE=84 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i13.GSR = "DISABLED";
    FD1S3IX o_r__i12 (.D(o_r_17__N_2438[12]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_04[12] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=84, LSE_RLINE=84 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i12.GSR = "DISABLED";
    FD1S3IX o_r__i11 (.D(o_r_17__N_2438[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_04[11] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=84, LSE_RLINE=84 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i11.GSR = "DISABLED";
    FD1S3IX o_r__i10 (.D(o_r_17__N_2438[10]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_04[10] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=84, LSE_RLINE=84 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i10.GSR = "DISABLED";
    FD1S3IX o_r__i9 (.D(o_r_17__N_2438[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_04[9] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=84, LSE_RLINE=84 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i9.GSR = "DISABLED";
    FD1S3IX o_r__i8 (.D(o_r_17__N_2438[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_04[8] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=84, LSE_RLINE=84 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i8.GSR = "DISABLED";
    FD1S3IX o_r__i7 (.D(o_r_17__N_2438[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_04[7] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=84, LSE_RLINE=84 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i7.GSR = "DISABLED";
    FD1S3IX o_r__i6 (.D(o_r_17__N_2438[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_04[6] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=84, LSE_RLINE=84 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i6.GSR = "DISABLED";
    FD1S3IX o_r__i5 (.D(o_r_17__N_2438[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_04[5] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=84, LSE_RLINE=84 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i5.GSR = "DISABLED";
    FD1S3IX o_r__i4 (.D(o_r_17__N_2438[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_04[4] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=84, LSE_RLINE=84 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i4.GSR = "DISABLED";
    FD1S3IX o_r__i3 (.D(o_r_17__N_2438[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_04[3] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=84, LSE_RLINE=84 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i3.GSR = "DISABLED";
    FD1S3IX o_r__i2 (.D(o_r_17__N_2438[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_04[2] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=84, LSE_RLINE=84 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i2.GSR = "DISABLED";
    FD1S3IX o_r__i1 (.D(o_r_17__N_2438[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_1_02_20__N_2226[1] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=84, LSE_RLINE=84 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i1.GSR = "DISABLED";
    LUT4 i12497_2_lut_rep_612 (.A(u_l[1]), .B(\u_s[8] ), .Z(n29272)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i12497_2_lut_rep_612.init = 16'h8888;
    LUT4 i12496_2_lut_rep_613 (.A(u_l[0]), .B(\u_s[9] ), .Z(n29273)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(51[18:45])
    defparam i12496_2_lut_rep_613.init = 16'h8888;
    LUT4 w_r_16__I_0_i2_2_lut_3_lut_4_lut (.A(u_l[0]), .B(\u_s[9] ), .C(\u_s[8] ), 
         .D(u_l[1]), .Z(o_r_17__N_2438[1])) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(51[18:45])
    defparam w_r_16__I_0_i2_2_lut_3_lut_4_lut.init = 16'h7888;
    
endmodule
//
// Verilog Description of module \bimpy(BW=16)_U2 
//

module \bimpy(BW=16)_U2  (u_l, \u_s[6] , \u_s[7] , S_0_03, dac_clk_p_c, 
            n14230, n9464, GND_net, i_sw0_c) /* synthesis syn_module_defined=1 */ ;
    input [15:0]u_l;
    input \u_s[6] ;
    input \u_s[7] ;
    output [17:0]S_0_03;
    input dac_clk_p_c;
    input n14230;
    input n9464;
    input GND_net;
    input i_sw0_c;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[29:38])
    
    wire n29277, n29278;
    wire [17:0]o_r_17__N_2438;
    
    wire n19503, n19502;
    wire [14:0]c_15__N_2408;
    wire [14:0]c_15__N_2423;
    
    wire n19501, n19500, n19499, n19498, n19497, n19496;
    
    LUT4 i12495_2_lut_rep_617 (.A(u_l[1]), .B(\u_s[6] ), .Z(n29277)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i12495_2_lut_rep_617.init = 16'h8888;
    LUT4 i12494_2_lut_rep_618 (.A(u_l[0]), .B(\u_s[7] ), .Z(n29278)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(51[18:45])
    defparam i12494_2_lut_rep_618.init = 16'h8888;
    LUT4 w_r_16__I_0_i2_2_lut_3_lut_4_lut (.A(u_l[0]), .B(\u_s[7] ), .C(\u_s[6] ), 
         .D(u_l[1]), .Z(o_r_17__N_2438[1])) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(51[18:45])
    defparam w_r_16__I_0_i2_2_lut_3_lut_4_lut.init = 16'h7888;
    FD1S3IX o_r__i0 (.D(n9464), .CK(dac_clk_p_c), .CD(n14230), .Q(S_0_03[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=81, LSE_RLINE=81 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i0.GSR = "DISABLED";
    CCU2D add_828_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19503), 
          .S0(o_r_17__N_2438[17]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_828_cout.INIT0 = 16'h0000;
    defparam add_828_cout.INIT1 = 16'h0000;
    defparam add_828_cout.INJECT1_0 = "NO";
    defparam add_828_cout.INJECT1_1 = "NO";
    CCU2D add_828_15 (.A0(c_15__N_2408[14]), .B0(c_15__N_2423[14]), .C0(c_15__N_2408[13]), 
          .D0(c_15__N_2423[13]), .A1(u_l[15]), .B1(\u_s[7] ), .C1(c_15__N_2408[14]), 
          .D1(c_15__N_2423[14]), .CIN(n19502), .COUT(n19503), .S0(o_r_17__N_2438[15]), 
          .S1(o_r_17__N_2438[16]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_828_15.INIT0 = 16'h9666;
    defparam add_828_15.INIT1 = 16'h7888;
    defparam add_828_15.INJECT1_0 = "NO";
    defparam add_828_15.INJECT1_1 = "NO";
    CCU2D add_828_13 (.A0(c_15__N_2408[12]), .B0(c_15__N_2423[12]), .C0(c_15__N_2408[11]), 
          .D0(c_15__N_2423[11]), .A1(c_15__N_2408[13]), .B1(c_15__N_2423[13]), 
          .C1(c_15__N_2408[12]), .D1(c_15__N_2423[12]), .CIN(n19501), 
          .COUT(n19502), .S0(o_r_17__N_2438[13]), .S1(o_r_17__N_2438[14]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_828_13.INIT0 = 16'h9666;
    defparam add_828_13.INIT1 = 16'h9666;
    defparam add_828_13.INJECT1_0 = "NO";
    defparam add_828_13.INJECT1_1 = "NO";
    CCU2D add_828_11 (.A0(c_15__N_2408[10]), .B0(c_15__N_2423[10]), .C0(c_15__N_2408[9]), 
          .D0(c_15__N_2423[9]), .A1(c_15__N_2408[11]), .B1(c_15__N_2423[11]), 
          .C1(c_15__N_2408[10]), .D1(c_15__N_2423[10]), .CIN(n19500), 
          .COUT(n19501), .S0(o_r_17__N_2438[11]), .S1(o_r_17__N_2438[12]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_828_11.INIT0 = 16'h9666;
    defparam add_828_11.INIT1 = 16'h9666;
    defparam add_828_11.INJECT1_0 = "NO";
    defparam add_828_11.INJECT1_1 = "NO";
    CCU2D add_828_9 (.A0(c_15__N_2408[8]), .B0(c_15__N_2423[8]), .C0(c_15__N_2408[7]), 
          .D0(c_15__N_2423[7]), .A1(c_15__N_2408[9]), .B1(c_15__N_2423[9]), 
          .C1(c_15__N_2408[8]), .D1(c_15__N_2423[8]), .CIN(n19499), .COUT(n19500), 
          .S0(o_r_17__N_2438[9]), .S1(o_r_17__N_2438[10]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_828_9.INIT0 = 16'h9666;
    defparam add_828_9.INIT1 = 16'h9666;
    defparam add_828_9.INJECT1_0 = "NO";
    defparam add_828_9.INJECT1_1 = "NO";
    CCU2D add_828_7 (.A0(c_15__N_2408[6]), .B0(c_15__N_2423[6]), .C0(c_15__N_2408[5]), 
          .D0(c_15__N_2423[5]), .A1(c_15__N_2408[7]), .B1(c_15__N_2423[7]), 
          .C1(c_15__N_2408[6]), .D1(c_15__N_2423[6]), .CIN(n19498), .COUT(n19499), 
          .S0(o_r_17__N_2438[7]), .S1(o_r_17__N_2438[8]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_828_7.INIT0 = 16'h9666;
    defparam add_828_7.INIT1 = 16'h9666;
    defparam add_828_7.INJECT1_0 = "NO";
    defparam add_828_7.INJECT1_1 = "NO";
    CCU2D add_828_5 (.A0(c_15__N_2408[4]), .B0(c_15__N_2423[4]), .C0(c_15__N_2408[3]), 
          .D0(c_15__N_2423[3]), .A1(c_15__N_2408[5]), .B1(c_15__N_2423[5]), 
          .C1(c_15__N_2408[4]), .D1(c_15__N_2423[4]), .CIN(n19497), .COUT(n19498), 
          .S0(o_r_17__N_2438[5]), .S1(o_r_17__N_2438[6]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_828_5.INIT0 = 16'h9666;
    defparam add_828_5.INIT1 = 16'h9666;
    defparam add_828_5.INJECT1_0 = "NO";
    defparam add_828_5.INJECT1_1 = "NO";
    CCU2D add_828_3 (.A0(c_15__N_2408[2]), .B0(c_15__N_2423[2]), .C0(c_15__N_2408[1]), 
          .D0(c_15__N_2423[1]), .A1(c_15__N_2408[3]), .B1(c_15__N_2423[3]), 
          .C1(c_15__N_2408[2]), .D1(c_15__N_2423[2]), .CIN(n19496), .COUT(n19497), 
          .S0(o_r_17__N_2438[3]), .S1(o_r_17__N_2438[4]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_828_3.INIT0 = 16'h9666;
    defparam add_828_3.INIT1 = 16'h9666;
    defparam add_828_3.INJECT1_0 = "NO";
    defparam add_828_3.INJECT1_1 = "NO";
    CCU2D add_828_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(c_15__N_2408[1]), .B1(c_15__N_2423[1]), .C1(n29278), .D1(n29277), 
          .COUT(n19496), .S1(o_r_17__N_2438[2]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_828_1.INIT0 = 16'hF000;
    defparam add_828_1.INIT1 = 16'h9666;
    defparam add_828_1.INJECT1_0 = "NO";
    defparam add_828_1.INJECT1_1 = "NO";
    LUT4 i13510_2_lut (.A(u_l[14]), .B(\u_s[7] ), .Z(c_15__N_2408[14])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13510_2_lut.init = 16'h8888;
    LUT4 i13496_2_lut (.A(u_l[15]), .B(\u_s[6] ), .Z(c_15__N_2423[14])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13496_2_lut.init = 16'h8888;
    LUT4 i13511_2_lut (.A(u_l[13]), .B(\u_s[7] ), .Z(c_15__N_2408[13])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13511_2_lut.init = 16'h8888;
    LUT4 i13497_2_lut (.A(u_l[14]), .B(\u_s[6] ), .Z(c_15__N_2423[13])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13497_2_lut.init = 16'h8888;
    LUT4 i13512_2_lut (.A(u_l[12]), .B(\u_s[7] ), .Z(c_15__N_2408[12])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13512_2_lut.init = 16'h8888;
    LUT4 i13498_2_lut (.A(u_l[13]), .B(\u_s[6] ), .Z(c_15__N_2423[12])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13498_2_lut.init = 16'h8888;
    LUT4 i13513_2_lut (.A(u_l[11]), .B(\u_s[7] ), .Z(c_15__N_2408[11])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13513_2_lut.init = 16'h8888;
    LUT4 i13499_2_lut (.A(u_l[12]), .B(\u_s[6] ), .Z(c_15__N_2423[11])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13499_2_lut.init = 16'h8888;
    LUT4 i13514_2_lut (.A(u_l[10]), .B(\u_s[7] ), .Z(c_15__N_2408[10])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13514_2_lut.init = 16'h8888;
    LUT4 i13500_2_lut (.A(u_l[11]), .B(\u_s[6] ), .Z(c_15__N_2423[10])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13500_2_lut.init = 16'h8888;
    LUT4 i13515_2_lut (.A(u_l[9]), .B(\u_s[7] ), .Z(c_15__N_2408[9])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13515_2_lut.init = 16'h8888;
    LUT4 i13501_2_lut (.A(u_l[10]), .B(\u_s[6] ), .Z(c_15__N_2423[9])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13501_2_lut.init = 16'h8888;
    LUT4 i13516_2_lut (.A(u_l[8]), .B(\u_s[7] ), .Z(c_15__N_2408[8])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13516_2_lut.init = 16'h8888;
    LUT4 i13502_2_lut (.A(u_l[9]), .B(\u_s[6] ), .Z(c_15__N_2423[8])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13502_2_lut.init = 16'h8888;
    LUT4 i13517_2_lut (.A(u_l[7]), .B(\u_s[7] ), .Z(c_15__N_2408[7])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13517_2_lut.init = 16'h8888;
    LUT4 i13503_2_lut (.A(u_l[8]), .B(\u_s[6] ), .Z(c_15__N_2423[7])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13503_2_lut.init = 16'h8888;
    LUT4 i13518_2_lut (.A(u_l[6]), .B(\u_s[7] ), .Z(c_15__N_2408[6])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13518_2_lut.init = 16'h8888;
    LUT4 i13504_2_lut (.A(u_l[7]), .B(\u_s[6] ), .Z(c_15__N_2423[6])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13504_2_lut.init = 16'h8888;
    LUT4 i13519_2_lut (.A(u_l[5]), .B(\u_s[7] ), .Z(c_15__N_2408[5])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13519_2_lut.init = 16'h8888;
    LUT4 i13505_2_lut (.A(u_l[6]), .B(\u_s[6] ), .Z(c_15__N_2423[5])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13505_2_lut.init = 16'h8888;
    LUT4 i13520_2_lut (.A(u_l[4]), .B(\u_s[7] ), .Z(c_15__N_2408[4])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13520_2_lut.init = 16'h8888;
    LUT4 i13506_2_lut (.A(u_l[5]), .B(\u_s[6] ), .Z(c_15__N_2423[4])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13506_2_lut.init = 16'h8888;
    LUT4 i13521_2_lut (.A(u_l[3]), .B(\u_s[7] ), .Z(c_15__N_2408[3])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13521_2_lut.init = 16'h8888;
    LUT4 i13507_2_lut (.A(u_l[4]), .B(\u_s[6] ), .Z(c_15__N_2423[3])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13507_2_lut.init = 16'h8888;
    LUT4 i13522_2_lut (.A(u_l[2]), .B(\u_s[7] ), .Z(c_15__N_2408[2])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13522_2_lut.init = 16'h8888;
    LUT4 i13508_2_lut (.A(u_l[3]), .B(\u_s[6] ), .Z(c_15__N_2423[2])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13508_2_lut.init = 16'h8888;
    LUT4 i13523_2_lut (.A(u_l[1]), .B(\u_s[7] ), .Z(c_15__N_2408[1])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13523_2_lut.init = 16'h8888;
    LUT4 i13509_2_lut (.A(u_l[2]), .B(\u_s[6] ), .Z(c_15__N_2423[1])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13509_2_lut.init = 16'h8888;
    FD1S3IX o_r__i17 (.D(o_r_17__N_2438[17]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_03[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=81, LSE_RLINE=81 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i17.GSR = "DISABLED";
    FD1S3IX o_r__i16 (.D(o_r_17__N_2438[16]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_03[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=81, LSE_RLINE=81 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i16.GSR = "DISABLED";
    FD1S3IX o_r__i15 (.D(o_r_17__N_2438[15]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_03[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=81, LSE_RLINE=81 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i15.GSR = "DISABLED";
    FD1S3IX o_r__i14 (.D(o_r_17__N_2438[14]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_03[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=81, LSE_RLINE=81 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i14.GSR = "DISABLED";
    FD1S3IX o_r__i13 (.D(o_r_17__N_2438[13]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_03[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=81, LSE_RLINE=81 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i13.GSR = "DISABLED";
    FD1S3IX o_r__i12 (.D(o_r_17__N_2438[12]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_03[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=81, LSE_RLINE=81 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i12.GSR = "DISABLED";
    FD1S3IX o_r__i11 (.D(o_r_17__N_2438[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_03[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=81, LSE_RLINE=81 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i11.GSR = "DISABLED";
    FD1S3IX o_r__i10 (.D(o_r_17__N_2438[10]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_03[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=81, LSE_RLINE=81 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i10.GSR = "DISABLED";
    FD1S3IX o_r__i9 (.D(o_r_17__N_2438[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_03[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=81, LSE_RLINE=81 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i9.GSR = "DISABLED";
    FD1S3IX o_r__i8 (.D(o_r_17__N_2438[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_03[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=81, LSE_RLINE=81 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i8.GSR = "DISABLED";
    FD1S3IX o_r__i7 (.D(o_r_17__N_2438[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_03[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=81, LSE_RLINE=81 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i7.GSR = "DISABLED";
    FD1S3IX o_r__i6 (.D(o_r_17__N_2438[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_03[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=81, LSE_RLINE=81 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i6.GSR = "DISABLED";
    FD1S3IX o_r__i5 (.D(o_r_17__N_2438[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_03[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=81, LSE_RLINE=81 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i5.GSR = "DISABLED";
    FD1S3IX o_r__i4 (.D(o_r_17__N_2438[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_03[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=81, LSE_RLINE=81 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i4.GSR = "DISABLED";
    FD1S3IX o_r__i3 (.D(o_r_17__N_2438[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_03[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=81, LSE_RLINE=81 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i3.GSR = "DISABLED";
    FD1S3IX o_r__i2 (.D(o_r_17__N_2438[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_03[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=81, LSE_RLINE=81 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i2.GSR = "DISABLED";
    FD1S3IX o_r__i1 (.D(o_r_17__N_2438[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_03[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=81, LSE_RLINE=81 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i1.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module \bimpy(BW=16)_U3 
//

module \bimpy(BW=16)_U3  (\S_0_02[0] , dac_clk_p_c, n14230, n9466, u_l, 
            \u_s[4] , \u_s[5] , GND_net, \S_0_02[17] , i_sw0_c, \S_0_02[16] , 
            \S_0_02[15] , \S_0_02[14] , \S_0_02[13] , \S_0_02[12] , 
            \S_0_02[11] , \S_0_02[10] , \S_0_02[9] , \S_0_02[8] , \S_0_02[7] , 
            \S_0_02[6] , \S_0_02[5] , \S_0_02[4] , \S_0_02[3] , \S_0_02[2] , 
            \S_1_01_20__N_2205[1] ) /* synthesis syn_module_defined=1 */ ;
    output \S_0_02[0] ;
    input dac_clk_p_c;
    input n14230;
    input n9466;
    input [15:0]u_l;
    input \u_s[4] ;
    input \u_s[5] ;
    input GND_net;
    output \S_0_02[17] ;
    input i_sw0_c;
    output \S_0_02[16] ;
    output \S_0_02[15] ;
    output \S_0_02[14] ;
    output \S_0_02[13] ;
    output \S_0_02[12] ;
    output \S_0_02[11] ;
    output \S_0_02[10] ;
    output \S_0_02[9] ;
    output \S_0_02[8] ;
    output \S_0_02[7] ;
    output \S_0_02[6] ;
    output \S_0_02[5] ;
    output \S_0_02[4] ;
    output \S_0_02[3] ;
    output \S_0_02[2] ;
    output \S_1_01_20__N_2205[1] ;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[29:38])
    
    wire n29279, n29280;
    wire [17:0]o_r_17__N_2438;
    
    wire n19511, n19510;
    wire [14:0]c_15__N_2408;
    wire [14:0]c_15__N_2423;
    
    wire n19509, n19508, n19507, n19506, n19505, n19504;
    
    FD1S3IX o_r__i0 (.D(n9466), .CK(dac_clk_p_c), .CD(n14230), .Q(\S_0_02[0] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i0.GSR = "DISABLED";
    LUT4 i12493_2_lut_rep_619 (.A(u_l[1]), .B(\u_s[4] ), .Z(n29279)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i12493_2_lut_rep_619.init = 16'h8888;
    LUT4 i12492_2_lut_rep_620 (.A(u_l[0]), .B(\u_s[5] ), .Z(n29280)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(51[18:45])
    defparam i12492_2_lut_rep_620.init = 16'h8888;
    LUT4 w_r_16__I_0_i2_2_lut_3_lut_4_lut (.A(u_l[0]), .B(\u_s[5] ), .C(\u_s[4] ), 
         .D(u_l[1]), .Z(o_r_17__N_2438[1])) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(51[18:45])
    defparam w_r_16__I_0_i2_2_lut_3_lut_4_lut.init = 16'h7888;
    CCU2D add_829_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19511), 
          .S0(o_r_17__N_2438[17]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_829_cout.INIT0 = 16'h0000;
    defparam add_829_cout.INIT1 = 16'h0000;
    defparam add_829_cout.INJECT1_0 = "NO";
    defparam add_829_cout.INJECT1_1 = "NO";
    CCU2D add_829_15 (.A0(c_15__N_2408[14]), .B0(c_15__N_2423[14]), .C0(c_15__N_2408[13]), 
          .D0(c_15__N_2423[13]), .A1(u_l[15]), .B1(\u_s[5] ), .C1(c_15__N_2408[14]), 
          .D1(c_15__N_2423[14]), .CIN(n19510), .COUT(n19511), .S0(o_r_17__N_2438[15]), 
          .S1(o_r_17__N_2438[16]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_829_15.INIT0 = 16'h9666;
    defparam add_829_15.INIT1 = 16'h7888;
    defparam add_829_15.INJECT1_0 = "NO";
    defparam add_829_15.INJECT1_1 = "NO";
    CCU2D add_829_13 (.A0(c_15__N_2408[12]), .B0(c_15__N_2423[12]), .C0(c_15__N_2408[11]), 
          .D0(c_15__N_2423[11]), .A1(c_15__N_2408[13]), .B1(c_15__N_2423[13]), 
          .C1(c_15__N_2408[12]), .D1(c_15__N_2423[12]), .CIN(n19509), 
          .COUT(n19510), .S0(o_r_17__N_2438[13]), .S1(o_r_17__N_2438[14]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_829_13.INIT0 = 16'h9666;
    defparam add_829_13.INIT1 = 16'h9666;
    defparam add_829_13.INJECT1_0 = "NO";
    defparam add_829_13.INJECT1_1 = "NO";
    CCU2D add_829_11 (.A0(c_15__N_2408[10]), .B0(c_15__N_2423[10]), .C0(c_15__N_2408[9]), 
          .D0(c_15__N_2423[9]), .A1(c_15__N_2408[11]), .B1(c_15__N_2423[11]), 
          .C1(c_15__N_2408[10]), .D1(c_15__N_2423[10]), .CIN(n19508), 
          .COUT(n19509), .S0(o_r_17__N_2438[11]), .S1(o_r_17__N_2438[12]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_829_11.INIT0 = 16'h9666;
    defparam add_829_11.INIT1 = 16'h9666;
    defparam add_829_11.INJECT1_0 = "NO";
    defparam add_829_11.INJECT1_1 = "NO";
    CCU2D add_829_9 (.A0(c_15__N_2408[8]), .B0(c_15__N_2423[8]), .C0(c_15__N_2408[7]), 
          .D0(c_15__N_2423[7]), .A1(c_15__N_2408[9]), .B1(c_15__N_2423[9]), 
          .C1(c_15__N_2408[8]), .D1(c_15__N_2423[8]), .CIN(n19507), .COUT(n19508), 
          .S0(o_r_17__N_2438[9]), .S1(o_r_17__N_2438[10]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_829_9.INIT0 = 16'h9666;
    defparam add_829_9.INIT1 = 16'h9666;
    defparam add_829_9.INJECT1_0 = "NO";
    defparam add_829_9.INJECT1_1 = "NO";
    CCU2D add_829_7 (.A0(c_15__N_2408[6]), .B0(c_15__N_2423[6]), .C0(c_15__N_2408[5]), 
          .D0(c_15__N_2423[5]), .A1(c_15__N_2408[7]), .B1(c_15__N_2423[7]), 
          .C1(c_15__N_2408[6]), .D1(c_15__N_2423[6]), .CIN(n19506), .COUT(n19507), 
          .S0(o_r_17__N_2438[7]), .S1(o_r_17__N_2438[8]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_829_7.INIT0 = 16'h9666;
    defparam add_829_7.INIT1 = 16'h9666;
    defparam add_829_7.INJECT1_0 = "NO";
    defparam add_829_7.INJECT1_1 = "NO";
    CCU2D add_829_5 (.A0(c_15__N_2408[4]), .B0(c_15__N_2423[4]), .C0(c_15__N_2408[3]), 
          .D0(c_15__N_2423[3]), .A1(c_15__N_2408[5]), .B1(c_15__N_2423[5]), 
          .C1(c_15__N_2408[4]), .D1(c_15__N_2423[4]), .CIN(n19505), .COUT(n19506), 
          .S0(o_r_17__N_2438[5]), .S1(o_r_17__N_2438[6]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_829_5.INIT0 = 16'h9666;
    defparam add_829_5.INIT1 = 16'h9666;
    defparam add_829_5.INJECT1_0 = "NO";
    defparam add_829_5.INJECT1_1 = "NO";
    CCU2D add_829_3 (.A0(c_15__N_2408[2]), .B0(c_15__N_2423[2]), .C0(c_15__N_2408[1]), 
          .D0(c_15__N_2423[1]), .A1(c_15__N_2408[3]), .B1(c_15__N_2423[3]), 
          .C1(c_15__N_2408[2]), .D1(c_15__N_2423[2]), .CIN(n19504), .COUT(n19505), 
          .S0(o_r_17__N_2438[3]), .S1(o_r_17__N_2438[4]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_829_3.INIT0 = 16'h9666;
    defparam add_829_3.INIT1 = 16'h9666;
    defparam add_829_3.INJECT1_0 = "NO";
    defparam add_829_3.INJECT1_1 = "NO";
    CCU2D add_829_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(c_15__N_2408[1]), .B1(c_15__N_2423[1]), .C1(n29280), .D1(n29279), 
          .COUT(n19504), .S1(o_r_17__N_2438[2]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_829_1.INIT0 = 16'hF000;
    defparam add_829_1.INIT1 = 16'h9666;
    defparam add_829_1.INJECT1_0 = "NO";
    defparam add_829_1.INJECT1_1 = "NO";
    LUT4 i13539_2_lut (.A(u_l[14]), .B(\u_s[5] ), .Z(c_15__N_2408[14])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13539_2_lut.init = 16'h8888;
    LUT4 i13525_2_lut (.A(u_l[15]), .B(\u_s[4] ), .Z(c_15__N_2423[14])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13525_2_lut.init = 16'h8888;
    LUT4 i13540_2_lut (.A(u_l[13]), .B(\u_s[5] ), .Z(c_15__N_2408[13])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13540_2_lut.init = 16'h8888;
    LUT4 i13526_2_lut (.A(u_l[14]), .B(\u_s[4] ), .Z(c_15__N_2423[13])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13526_2_lut.init = 16'h8888;
    LUT4 i13541_2_lut (.A(u_l[12]), .B(\u_s[5] ), .Z(c_15__N_2408[12])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13541_2_lut.init = 16'h8888;
    LUT4 i13527_2_lut (.A(u_l[13]), .B(\u_s[4] ), .Z(c_15__N_2423[12])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13527_2_lut.init = 16'h8888;
    LUT4 i13542_2_lut (.A(u_l[11]), .B(\u_s[5] ), .Z(c_15__N_2408[11])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13542_2_lut.init = 16'h8888;
    LUT4 i13528_2_lut (.A(u_l[12]), .B(\u_s[4] ), .Z(c_15__N_2423[11])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13528_2_lut.init = 16'h8888;
    LUT4 i13543_2_lut (.A(u_l[10]), .B(\u_s[5] ), .Z(c_15__N_2408[10])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13543_2_lut.init = 16'h8888;
    LUT4 i13529_2_lut (.A(u_l[11]), .B(\u_s[4] ), .Z(c_15__N_2423[10])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13529_2_lut.init = 16'h8888;
    LUT4 i13544_2_lut (.A(u_l[9]), .B(\u_s[5] ), .Z(c_15__N_2408[9])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13544_2_lut.init = 16'h8888;
    LUT4 i13530_2_lut (.A(u_l[10]), .B(\u_s[4] ), .Z(c_15__N_2423[9])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13530_2_lut.init = 16'h8888;
    LUT4 i13545_2_lut (.A(u_l[8]), .B(\u_s[5] ), .Z(c_15__N_2408[8])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13545_2_lut.init = 16'h8888;
    LUT4 i13531_2_lut (.A(u_l[9]), .B(\u_s[4] ), .Z(c_15__N_2423[8])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13531_2_lut.init = 16'h8888;
    LUT4 i13546_2_lut (.A(u_l[7]), .B(\u_s[5] ), .Z(c_15__N_2408[7])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13546_2_lut.init = 16'h8888;
    LUT4 i13532_2_lut (.A(u_l[8]), .B(\u_s[4] ), .Z(c_15__N_2423[7])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13532_2_lut.init = 16'h8888;
    LUT4 i13547_2_lut (.A(u_l[6]), .B(\u_s[5] ), .Z(c_15__N_2408[6])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13547_2_lut.init = 16'h8888;
    LUT4 i13533_2_lut (.A(u_l[7]), .B(\u_s[4] ), .Z(c_15__N_2423[6])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13533_2_lut.init = 16'h8888;
    LUT4 i13548_2_lut (.A(u_l[5]), .B(\u_s[5] ), .Z(c_15__N_2408[5])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13548_2_lut.init = 16'h8888;
    LUT4 i13534_2_lut (.A(u_l[6]), .B(\u_s[4] ), .Z(c_15__N_2423[5])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13534_2_lut.init = 16'h8888;
    LUT4 i13549_2_lut (.A(u_l[4]), .B(\u_s[5] ), .Z(c_15__N_2408[4])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13549_2_lut.init = 16'h8888;
    LUT4 i13535_2_lut (.A(u_l[5]), .B(\u_s[4] ), .Z(c_15__N_2423[4])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13535_2_lut.init = 16'h8888;
    LUT4 i13550_2_lut (.A(u_l[3]), .B(\u_s[5] ), .Z(c_15__N_2408[3])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13550_2_lut.init = 16'h8888;
    LUT4 i13536_2_lut (.A(u_l[4]), .B(\u_s[4] ), .Z(c_15__N_2423[3])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13536_2_lut.init = 16'h8888;
    LUT4 i13551_2_lut (.A(u_l[2]), .B(\u_s[5] ), .Z(c_15__N_2408[2])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13551_2_lut.init = 16'h8888;
    LUT4 i13537_2_lut (.A(u_l[3]), .B(\u_s[4] ), .Z(c_15__N_2423[2])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13537_2_lut.init = 16'h8888;
    LUT4 i13552_2_lut (.A(u_l[1]), .B(\u_s[5] ), .Z(c_15__N_2408[1])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13552_2_lut.init = 16'h8888;
    LUT4 i13538_2_lut (.A(u_l[2]), .B(\u_s[4] ), .Z(c_15__N_2423[1])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13538_2_lut.init = 16'h8888;
    FD1S3IX o_r__i17 (.D(o_r_17__N_2438[17]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_02[17] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i17.GSR = "DISABLED";
    FD1S3IX o_r__i16 (.D(o_r_17__N_2438[16]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_02[16] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i16.GSR = "DISABLED";
    FD1S3IX o_r__i15 (.D(o_r_17__N_2438[15]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_02[15] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i15.GSR = "DISABLED";
    FD1S3IX o_r__i14 (.D(o_r_17__N_2438[14]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_02[14] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i14.GSR = "DISABLED";
    FD1S3IX o_r__i13 (.D(o_r_17__N_2438[13]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_02[13] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i13.GSR = "DISABLED";
    FD1S3IX o_r__i12 (.D(o_r_17__N_2438[12]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_02[12] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i12.GSR = "DISABLED";
    FD1S3IX o_r__i11 (.D(o_r_17__N_2438[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_02[11] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i11.GSR = "DISABLED";
    FD1S3IX o_r__i10 (.D(o_r_17__N_2438[10]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_02[10] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i10.GSR = "DISABLED";
    FD1S3IX o_r__i9 (.D(o_r_17__N_2438[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_02[9] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i9.GSR = "DISABLED";
    FD1S3IX o_r__i8 (.D(o_r_17__N_2438[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_02[8] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i8.GSR = "DISABLED";
    FD1S3IX o_r__i7 (.D(o_r_17__N_2438[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_02[7] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i7.GSR = "DISABLED";
    FD1S3IX o_r__i6 (.D(o_r_17__N_2438[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_02[6] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i6.GSR = "DISABLED";
    FD1S3IX o_r__i5 (.D(o_r_17__N_2438[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_02[5] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i5.GSR = "DISABLED";
    FD1S3IX o_r__i4 (.D(o_r_17__N_2438[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_02[4] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i4.GSR = "DISABLED";
    FD1S3IX o_r__i3 (.D(o_r_17__N_2438[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_02[3] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i3.GSR = "DISABLED";
    FD1S3IX o_r__i2 (.D(o_r_17__N_2438[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_02[2] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i2.GSR = "DISABLED";
    FD1S3IX o_r__i1 (.D(o_r_17__N_2438[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_1_01_20__N_2205[1] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i1.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module \bimpy(BW=16)_U4 
//

module \bimpy(BW=16)_U4  (S_0_01, dac_clk_p_c, n14230, n9468, GND_net, 
            u_l, \u_s[3] , \u_s[2] , i_sw0_c) /* synthesis syn_module_defined=1 */ ;
    output [17:0]S_0_01;
    input dac_clk_p_c;
    input n14230;
    input n9468;
    input GND_net;
    input [15:0]u_l;
    input \u_s[3] ;
    input \u_s[2] ;
    input i_sw0_c;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[29:38])
    
    wire n19519;
    wire [17:0]o_r_17__N_2438;
    
    wire n19518;
    wire [14:0]c_15__N_2408;
    wire [14:0]c_15__N_2423;
    
    wire n19517, n19516, n19515, n19514, n19513, n19512, n29287, 
        n29286;
    
    FD1S3IX o_r__i0 (.D(n9468), .CK(dac_clk_p_c), .CD(n14230), .Q(S_0_01[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=75, LSE_RLINE=75 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i0.GSR = "DISABLED";
    CCU2D add_830_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19519), 
          .S0(o_r_17__N_2438[17]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_830_cout.INIT0 = 16'h0000;
    defparam add_830_cout.INIT1 = 16'h0000;
    defparam add_830_cout.INJECT1_0 = "NO";
    defparam add_830_cout.INJECT1_1 = "NO";
    CCU2D add_830_15 (.A0(c_15__N_2408[14]), .B0(c_15__N_2423[14]), .C0(c_15__N_2408[13]), 
          .D0(c_15__N_2423[13]), .A1(u_l[15]), .B1(\u_s[3] ), .C1(c_15__N_2408[14]), 
          .D1(c_15__N_2423[14]), .CIN(n19518), .COUT(n19519), .S0(o_r_17__N_2438[15]), 
          .S1(o_r_17__N_2438[16]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_830_15.INIT0 = 16'h9666;
    defparam add_830_15.INIT1 = 16'h7888;
    defparam add_830_15.INJECT1_0 = "NO";
    defparam add_830_15.INJECT1_1 = "NO";
    CCU2D add_830_13 (.A0(c_15__N_2408[12]), .B0(c_15__N_2423[12]), .C0(c_15__N_2408[11]), 
          .D0(c_15__N_2423[11]), .A1(c_15__N_2408[13]), .B1(c_15__N_2423[13]), 
          .C1(c_15__N_2408[12]), .D1(c_15__N_2423[12]), .CIN(n19517), 
          .COUT(n19518), .S0(o_r_17__N_2438[13]), .S1(o_r_17__N_2438[14]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_830_13.INIT0 = 16'h9666;
    defparam add_830_13.INIT1 = 16'h9666;
    defparam add_830_13.INJECT1_0 = "NO";
    defparam add_830_13.INJECT1_1 = "NO";
    CCU2D add_830_11 (.A0(c_15__N_2408[10]), .B0(c_15__N_2423[10]), .C0(c_15__N_2408[9]), 
          .D0(c_15__N_2423[9]), .A1(c_15__N_2408[11]), .B1(c_15__N_2423[11]), 
          .C1(c_15__N_2408[10]), .D1(c_15__N_2423[10]), .CIN(n19516), 
          .COUT(n19517), .S0(o_r_17__N_2438[11]), .S1(o_r_17__N_2438[12]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_830_11.INIT0 = 16'h9666;
    defparam add_830_11.INIT1 = 16'h9666;
    defparam add_830_11.INJECT1_0 = "NO";
    defparam add_830_11.INJECT1_1 = "NO";
    CCU2D add_830_9 (.A0(c_15__N_2408[8]), .B0(c_15__N_2423[8]), .C0(c_15__N_2408[7]), 
          .D0(c_15__N_2423[7]), .A1(c_15__N_2408[9]), .B1(c_15__N_2423[9]), 
          .C1(c_15__N_2408[8]), .D1(c_15__N_2423[8]), .CIN(n19515), .COUT(n19516), 
          .S0(o_r_17__N_2438[9]), .S1(o_r_17__N_2438[10]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_830_9.INIT0 = 16'h9666;
    defparam add_830_9.INIT1 = 16'h9666;
    defparam add_830_9.INJECT1_0 = "NO";
    defparam add_830_9.INJECT1_1 = "NO";
    CCU2D add_830_7 (.A0(c_15__N_2408[6]), .B0(c_15__N_2423[6]), .C0(c_15__N_2408[5]), 
          .D0(c_15__N_2423[5]), .A1(c_15__N_2408[7]), .B1(c_15__N_2423[7]), 
          .C1(c_15__N_2408[6]), .D1(c_15__N_2423[6]), .CIN(n19514), .COUT(n19515), 
          .S0(o_r_17__N_2438[7]), .S1(o_r_17__N_2438[8]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_830_7.INIT0 = 16'h9666;
    defparam add_830_7.INIT1 = 16'h9666;
    defparam add_830_7.INJECT1_0 = "NO";
    defparam add_830_7.INJECT1_1 = "NO";
    CCU2D add_830_5 (.A0(c_15__N_2408[4]), .B0(c_15__N_2423[4]), .C0(c_15__N_2408[3]), 
          .D0(c_15__N_2423[3]), .A1(c_15__N_2408[5]), .B1(c_15__N_2423[5]), 
          .C1(c_15__N_2408[4]), .D1(c_15__N_2423[4]), .CIN(n19513), .COUT(n19514), 
          .S0(o_r_17__N_2438[5]), .S1(o_r_17__N_2438[6]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_830_5.INIT0 = 16'h9666;
    defparam add_830_5.INIT1 = 16'h9666;
    defparam add_830_5.INJECT1_0 = "NO";
    defparam add_830_5.INJECT1_1 = "NO";
    CCU2D add_830_3 (.A0(c_15__N_2408[2]), .B0(c_15__N_2423[2]), .C0(c_15__N_2408[1]), 
          .D0(c_15__N_2423[1]), .A1(c_15__N_2408[3]), .B1(c_15__N_2423[3]), 
          .C1(c_15__N_2408[2]), .D1(c_15__N_2423[2]), .CIN(n19512), .COUT(n19513), 
          .S0(o_r_17__N_2438[3]), .S1(o_r_17__N_2438[4]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_830_3.INIT0 = 16'h9666;
    defparam add_830_3.INIT1 = 16'h9666;
    defparam add_830_3.INJECT1_0 = "NO";
    defparam add_830_3.INJECT1_1 = "NO";
    CCU2D add_830_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(c_15__N_2408[1]), .B1(c_15__N_2423[1]), .C1(n29287), .D1(n29286), 
          .COUT(n19512), .S1(o_r_17__N_2438[2]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_830_1.INIT0 = 16'hF000;
    defparam add_830_1.INIT1 = 16'h9666;
    defparam add_830_1.INJECT1_0 = "NO";
    defparam add_830_1.INJECT1_1 = "NO";
    LUT4 i13568_2_lut (.A(u_l[14]), .B(\u_s[3] ), .Z(c_15__N_2408[14])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13568_2_lut.init = 16'h8888;
    LUT4 i13554_2_lut (.A(u_l[15]), .B(\u_s[2] ), .Z(c_15__N_2423[14])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13554_2_lut.init = 16'h8888;
    LUT4 i13569_2_lut (.A(u_l[13]), .B(\u_s[3] ), .Z(c_15__N_2408[13])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13569_2_lut.init = 16'h8888;
    LUT4 i13555_2_lut (.A(u_l[14]), .B(\u_s[2] ), .Z(c_15__N_2423[13])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13555_2_lut.init = 16'h8888;
    LUT4 i13570_2_lut (.A(u_l[12]), .B(\u_s[3] ), .Z(c_15__N_2408[12])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13570_2_lut.init = 16'h8888;
    LUT4 i13556_2_lut (.A(u_l[13]), .B(\u_s[2] ), .Z(c_15__N_2423[12])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13556_2_lut.init = 16'h8888;
    LUT4 i13571_2_lut (.A(u_l[11]), .B(\u_s[3] ), .Z(c_15__N_2408[11])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13571_2_lut.init = 16'h8888;
    LUT4 i13557_2_lut (.A(u_l[12]), .B(\u_s[2] ), .Z(c_15__N_2423[11])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13557_2_lut.init = 16'h8888;
    LUT4 i13572_2_lut (.A(u_l[10]), .B(\u_s[3] ), .Z(c_15__N_2408[10])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13572_2_lut.init = 16'h8888;
    LUT4 i13558_2_lut (.A(u_l[11]), .B(\u_s[2] ), .Z(c_15__N_2423[10])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13558_2_lut.init = 16'h8888;
    LUT4 i13573_2_lut (.A(u_l[9]), .B(\u_s[3] ), .Z(c_15__N_2408[9])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13573_2_lut.init = 16'h8888;
    LUT4 i13559_2_lut (.A(u_l[10]), .B(\u_s[2] ), .Z(c_15__N_2423[9])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13559_2_lut.init = 16'h8888;
    LUT4 i13574_2_lut (.A(u_l[8]), .B(\u_s[3] ), .Z(c_15__N_2408[8])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13574_2_lut.init = 16'h8888;
    LUT4 i13560_2_lut (.A(u_l[9]), .B(\u_s[2] ), .Z(c_15__N_2423[8])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13560_2_lut.init = 16'h8888;
    LUT4 i13575_2_lut (.A(u_l[7]), .B(\u_s[3] ), .Z(c_15__N_2408[7])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13575_2_lut.init = 16'h8888;
    LUT4 i13561_2_lut (.A(u_l[8]), .B(\u_s[2] ), .Z(c_15__N_2423[7])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13561_2_lut.init = 16'h8888;
    LUT4 i13576_2_lut (.A(u_l[6]), .B(\u_s[3] ), .Z(c_15__N_2408[6])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13576_2_lut.init = 16'h8888;
    LUT4 i13562_2_lut (.A(u_l[7]), .B(\u_s[2] ), .Z(c_15__N_2423[6])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13562_2_lut.init = 16'h8888;
    LUT4 i13577_2_lut (.A(u_l[5]), .B(\u_s[3] ), .Z(c_15__N_2408[5])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13577_2_lut.init = 16'h8888;
    LUT4 i13563_2_lut (.A(u_l[6]), .B(\u_s[2] ), .Z(c_15__N_2423[5])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13563_2_lut.init = 16'h8888;
    LUT4 i13578_2_lut (.A(u_l[4]), .B(\u_s[3] ), .Z(c_15__N_2408[4])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13578_2_lut.init = 16'h8888;
    LUT4 i13564_2_lut (.A(u_l[5]), .B(\u_s[2] ), .Z(c_15__N_2423[4])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13564_2_lut.init = 16'h8888;
    LUT4 i13579_2_lut (.A(u_l[3]), .B(\u_s[3] ), .Z(c_15__N_2408[3])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13579_2_lut.init = 16'h8888;
    LUT4 i13565_2_lut (.A(u_l[4]), .B(\u_s[2] ), .Z(c_15__N_2423[3])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13565_2_lut.init = 16'h8888;
    LUT4 i13580_2_lut (.A(u_l[2]), .B(\u_s[3] ), .Z(c_15__N_2408[2])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13580_2_lut.init = 16'h8888;
    LUT4 i13566_2_lut (.A(u_l[3]), .B(\u_s[2] ), .Z(c_15__N_2423[2])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13566_2_lut.init = 16'h8888;
    LUT4 i13581_2_lut (.A(u_l[1]), .B(\u_s[3] ), .Z(c_15__N_2408[1])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13581_2_lut.init = 16'h8888;
    LUT4 i13567_2_lut (.A(u_l[2]), .B(\u_s[2] ), .Z(c_15__N_2423[1])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13567_2_lut.init = 16'h8888;
    LUT4 i12491_2_lut_rep_626 (.A(u_l[1]), .B(\u_s[2] ), .Z(n29286)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i12491_2_lut_rep_626.init = 16'h8888;
    LUT4 i12490_2_lut_rep_627 (.A(u_l[0]), .B(\u_s[3] ), .Z(n29287)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(51[18:45])
    defparam i12490_2_lut_rep_627.init = 16'h8888;
    LUT4 w_r_16__I_0_i2_2_lut_3_lut_4_lut (.A(u_l[0]), .B(\u_s[3] ), .C(\u_s[2] ), 
         .D(u_l[1]), .Z(o_r_17__N_2438[1])) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(51[18:45])
    defparam w_r_16__I_0_i2_2_lut_3_lut_4_lut.init = 16'h7888;
    FD1S3IX o_r__i17 (.D(o_r_17__N_2438[17]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_01[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=75, LSE_RLINE=75 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i17.GSR = "DISABLED";
    FD1S3IX o_r__i16 (.D(o_r_17__N_2438[16]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_01[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=75, LSE_RLINE=75 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i16.GSR = "DISABLED";
    FD1S3IX o_r__i15 (.D(o_r_17__N_2438[15]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_01[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=75, LSE_RLINE=75 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i15.GSR = "DISABLED";
    FD1S3IX o_r__i14 (.D(o_r_17__N_2438[14]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_01[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=75, LSE_RLINE=75 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i14.GSR = "DISABLED";
    FD1S3IX o_r__i13 (.D(o_r_17__N_2438[13]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_01[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=75, LSE_RLINE=75 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i13.GSR = "DISABLED";
    FD1S3IX o_r__i12 (.D(o_r_17__N_2438[12]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_01[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=75, LSE_RLINE=75 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i12.GSR = "DISABLED";
    FD1S3IX o_r__i11 (.D(o_r_17__N_2438[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_01[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=75, LSE_RLINE=75 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i11.GSR = "DISABLED";
    FD1S3IX o_r__i10 (.D(o_r_17__N_2438[10]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_01[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=75, LSE_RLINE=75 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i10.GSR = "DISABLED";
    FD1S3IX o_r__i9 (.D(o_r_17__N_2438[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_01[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=75, LSE_RLINE=75 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i9.GSR = "DISABLED";
    FD1S3IX o_r__i8 (.D(o_r_17__N_2438[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_01[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=75, LSE_RLINE=75 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i8.GSR = "DISABLED";
    FD1S3IX o_r__i7 (.D(o_r_17__N_2438[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_01[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=75, LSE_RLINE=75 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i7.GSR = "DISABLED";
    FD1S3IX o_r__i6 (.D(o_r_17__N_2438[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_01[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=75, LSE_RLINE=75 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i6.GSR = "DISABLED";
    FD1S3IX o_r__i5 (.D(o_r_17__N_2438[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_01[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=75, LSE_RLINE=75 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i5.GSR = "DISABLED";
    FD1S3IX o_r__i4 (.D(o_r_17__N_2438[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_01[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=75, LSE_RLINE=75 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i4.GSR = "DISABLED";
    FD1S3IX o_r__i3 (.D(o_r_17__N_2438[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_01[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=75, LSE_RLINE=75 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i3.GSR = "DISABLED";
    FD1S3IX o_r__i2 (.D(o_r_17__N_2438[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_01[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=75, LSE_RLINE=75 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i2.GSR = "DISABLED";
    FD1S3IX o_r__i1 (.D(o_r_17__N_2438[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_01[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=75, LSE_RLINE=75 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i1.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module \bimpy(BW=16)_U5 
//

module \bimpy(BW=16)_U5  (\S_0_00[0] , dac_clk_p_c, n14230, n9488, GND_net, 
            u_l, \u_s[1] , \u_s[0] , \S_0_00[17] , i_sw0_c, \S_0_00[16] , 
            \S_0_00[15] , \S_0_00[14] , \S_0_00[13] , \S_0_00[12] , 
            \S_0_00[11] , \S_0_00[10] , \S_0_00[9] , \S_0_00[8] , \S_0_00[7] , 
            \S_0_00[6] , \S_0_00[5] , \S_0_00[4] , \S_0_00[3] , \S_0_00[2] , 
            \S_1_00_20__N_2184[1] ) /* synthesis syn_module_defined=1 */ ;
    output \S_0_00[0] ;
    input dac_clk_p_c;
    input n14230;
    input n9488;
    input GND_net;
    input [15:0]u_l;
    input \u_s[1] ;
    input \u_s[0] ;
    output \S_0_00[17] ;
    input i_sw0_c;
    output \S_0_00[16] ;
    output \S_0_00[15] ;
    output \S_0_00[14] ;
    output \S_0_00[13] ;
    output \S_0_00[12] ;
    output \S_0_00[11] ;
    output \S_0_00[10] ;
    output \S_0_00[9] ;
    output \S_0_00[8] ;
    output \S_0_00[7] ;
    output \S_0_00[6] ;
    output \S_0_00[5] ;
    output \S_0_00[4] ;
    output \S_0_00[3] ;
    output \S_0_00[2] ;
    output \S_1_00_20__N_2184[1] ;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[29:38])
    
    wire n19527;
    wire [17:0]o_r_17__N_2438;
    
    wire n19526;
    wire [14:0]c_15__N_2408;
    wire [14:0]c_15__N_2423;
    
    wire n19525, n19524, n19523, n19522, n19521, n19520, n29293, 
        n29292;
    
    FD1S3IX o_r__i0 (.D(n9488), .CK(dac_clk_p_c), .CD(n14230), .Q(\S_0_00[0] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i0.GSR = "DISABLED";
    CCU2D add_831_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19527), 
          .S0(o_r_17__N_2438[17]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_831_cout.INIT0 = 16'h0000;
    defparam add_831_cout.INIT1 = 16'h0000;
    defparam add_831_cout.INJECT1_0 = "NO";
    defparam add_831_cout.INJECT1_1 = "NO";
    CCU2D add_831_15 (.A0(c_15__N_2408[14]), .B0(c_15__N_2423[14]), .C0(c_15__N_2408[13]), 
          .D0(c_15__N_2423[13]), .A1(u_l[15]), .B1(\u_s[1] ), .C1(c_15__N_2408[14]), 
          .D1(c_15__N_2423[14]), .CIN(n19526), .COUT(n19527), .S0(o_r_17__N_2438[15]), 
          .S1(o_r_17__N_2438[16]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_831_15.INIT0 = 16'h9666;
    defparam add_831_15.INIT1 = 16'h7888;
    defparam add_831_15.INJECT1_0 = "NO";
    defparam add_831_15.INJECT1_1 = "NO";
    CCU2D add_831_13 (.A0(c_15__N_2408[12]), .B0(c_15__N_2423[12]), .C0(c_15__N_2408[11]), 
          .D0(c_15__N_2423[11]), .A1(c_15__N_2408[13]), .B1(c_15__N_2423[13]), 
          .C1(c_15__N_2408[12]), .D1(c_15__N_2423[12]), .CIN(n19525), 
          .COUT(n19526), .S0(o_r_17__N_2438[13]), .S1(o_r_17__N_2438[14]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_831_13.INIT0 = 16'h9666;
    defparam add_831_13.INIT1 = 16'h9666;
    defparam add_831_13.INJECT1_0 = "NO";
    defparam add_831_13.INJECT1_1 = "NO";
    CCU2D add_831_11 (.A0(c_15__N_2408[10]), .B0(c_15__N_2423[10]), .C0(c_15__N_2408[9]), 
          .D0(c_15__N_2423[9]), .A1(c_15__N_2408[11]), .B1(c_15__N_2423[11]), 
          .C1(c_15__N_2408[10]), .D1(c_15__N_2423[10]), .CIN(n19524), 
          .COUT(n19525), .S0(o_r_17__N_2438[11]), .S1(o_r_17__N_2438[12]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_831_11.INIT0 = 16'h9666;
    defparam add_831_11.INIT1 = 16'h9666;
    defparam add_831_11.INJECT1_0 = "NO";
    defparam add_831_11.INJECT1_1 = "NO";
    CCU2D add_831_9 (.A0(c_15__N_2408[8]), .B0(c_15__N_2423[8]), .C0(c_15__N_2408[7]), 
          .D0(c_15__N_2423[7]), .A1(c_15__N_2408[9]), .B1(c_15__N_2423[9]), 
          .C1(c_15__N_2408[8]), .D1(c_15__N_2423[8]), .CIN(n19523), .COUT(n19524), 
          .S0(o_r_17__N_2438[9]), .S1(o_r_17__N_2438[10]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_831_9.INIT0 = 16'h9666;
    defparam add_831_9.INIT1 = 16'h9666;
    defparam add_831_9.INJECT1_0 = "NO";
    defparam add_831_9.INJECT1_1 = "NO";
    CCU2D add_831_7 (.A0(c_15__N_2408[6]), .B0(c_15__N_2423[6]), .C0(c_15__N_2408[5]), 
          .D0(c_15__N_2423[5]), .A1(c_15__N_2408[7]), .B1(c_15__N_2423[7]), 
          .C1(c_15__N_2408[6]), .D1(c_15__N_2423[6]), .CIN(n19522), .COUT(n19523), 
          .S0(o_r_17__N_2438[7]), .S1(o_r_17__N_2438[8]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_831_7.INIT0 = 16'h9666;
    defparam add_831_7.INIT1 = 16'h9666;
    defparam add_831_7.INJECT1_0 = "NO";
    defparam add_831_7.INJECT1_1 = "NO";
    CCU2D add_831_5 (.A0(c_15__N_2408[4]), .B0(c_15__N_2423[4]), .C0(c_15__N_2408[3]), 
          .D0(c_15__N_2423[3]), .A1(c_15__N_2408[5]), .B1(c_15__N_2423[5]), 
          .C1(c_15__N_2408[4]), .D1(c_15__N_2423[4]), .CIN(n19521), .COUT(n19522), 
          .S0(o_r_17__N_2438[5]), .S1(o_r_17__N_2438[6]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_831_5.INIT0 = 16'h9666;
    defparam add_831_5.INIT1 = 16'h9666;
    defparam add_831_5.INJECT1_0 = "NO";
    defparam add_831_5.INJECT1_1 = "NO";
    CCU2D add_831_3 (.A0(c_15__N_2408[2]), .B0(c_15__N_2423[2]), .C0(c_15__N_2408[1]), 
          .D0(c_15__N_2423[1]), .A1(c_15__N_2408[3]), .B1(c_15__N_2423[3]), 
          .C1(c_15__N_2408[2]), .D1(c_15__N_2423[2]), .CIN(n19520), .COUT(n19521), 
          .S0(o_r_17__N_2438[3]), .S1(o_r_17__N_2438[4]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_831_3.INIT0 = 16'h9666;
    defparam add_831_3.INIT1 = 16'h9666;
    defparam add_831_3.INJECT1_0 = "NO";
    defparam add_831_3.INJECT1_1 = "NO";
    CCU2D add_831_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(c_15__N_2408[1]), .B1(c_15__N_2423[1]), .C1(n29293), .D1(n29292), 
          .COUT(n19520), .S1(o_r_17__N_2438[2]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_831_1.INIT0 = 16'hF000;
    defparam add_831_1.INIT1 = 16'h9666;
    defparam add_831_1.INJECT1_0 = "NO";
    defparam add_831_1.INJECT1_1 = "NO";
    LUT4 i13598_2_lut (.A(u_l[14]), .B(\u_s[1] ), .Z(c_15__N_2408[14])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13598_2_lut.init = 16'h8888;
    LUT4 i13584_2_lut (.A(u_l[15]), .B(\u_s[0] ), .Z(c_15__N_2423[14])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13584_2_lut.init = 16'h8888;
    LUT4 i13599_2_lut (.A(u_l[13]), .B(\u_s[1] ), .Z(c_15__N_2408[13])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13599_2_lut.init = 16'h8888;
    LUT4 i13585_2_lut (.A(u_l[14]), .B(\u_s[0] ), .Z(c_15__N_2423[13])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13585_2_lut.init = 16'h8888;
    LUT4 i13600_2_lut (.A(u_l[12]), .B(\u_s[1] ), .Z(c_15__N_2408[12])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13600_2_lut.init = 16'h8888;
    LUT4 i13586_2_lut (.A(u_l[13]), .B(\u_s[0] ), .Z(c_15__N_2423[12])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13586_2_lut.init = 16'h8888;
    LUT4 i13601_2_lut (.A(u_l[11]), .B(\u_s[1] ), .Z(c_15__N_2408[11])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13601_2_lut.init = 16'h8888;
    LUT4 i13587_2_lut (.A(u_l[12]), .B(\u_s[0] ), .Z(c_15__N_2423[11])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13587_2_lut.init = 16'h8888;
    LUT4 i13602_2_lut (.A(u_l[10]), .B(\u_s[1] ), .Z(c_15__N_2408[10])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13602_2_lut.init = 16'h8888;
    LUT4 i13588_2_lut (.A(u_l[11]), .B(\u_s[0] ), .Z(c_15__N_2423[10])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13588_2_lut.init = 16'h8888;
    LUT4 i13603_2_lut (.A(u_l[9]), .B(\u_s[1] ), .Z(c_15__N_2408[9])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13603_2_lut.init = 16'h8888;
    LUT4 i13589_2_lut (.A(u_l[10]), .B(\u_s[0] ), .Z(c_15__N_2423[9])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13589_2_lut.init = 16'h8888;
    LUT4 i13604_2_lut (.A(u_l[8]), .B(\u_s[1] ), .Z(c_15__N_2408[8])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13604_2_lut.init = 16'h8888;
    LUT4 i13590_2_lut (.A(u_l[9]), .B(\u_s[0] ), .Z(c_15__N_2423[8])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13590_2_lut.init = 16'h8888;
    LUT4 i13605_2_lut (.A(u_l[7]), .B(\u_s[1] ), .Z(c_15__N_2408[7])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13605_2_lut.init = 16'h8888;
    LUT4 i13591_2_lut (.A(u_l[8]), .B(\u_s[0] ), .Z(c_15__N_2423[7])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13591_2_lut.init = 16'h8888;
    LUT4 i13606_2_lut (.A(u_l[6]), .B(\u_s[1] ), .Z(c_15__N_2408[6])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13606_2_lut.init = 16'h8888;
    LUT4 i13592_2_lut (.A(u_l[7]), .B(\u_s[0] ), .Z(c_15__N_2423[6])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13592_2_lut.init = 16'h8888;
    LUT4 i13607_2_lut (.A(u_l[5]), .B(\u_s[1] ), .Z(c_15__N_2408[5])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13607_2_lut.init = 16'h8888;
    LUT4 i13593_2_lut (.A(u_l[6]), .B(\u_s[0] ), .Z(c_15__N_2423[5])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13593_2_lut.init = 16'h8888;
    LUT4 i13608_2_lut (.A(u_l[4]), .B(\u_s[1] ), .Z(c_15__N_2408[4])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13608_2_lut.init = 16'h8888;
    LUT4 i13594_2_lut (.A(u_l[5]), .B(\u_s[0] ), .Z(c_15__N_2423[4])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13594_2_lut.init = 16'h8888;
    LUT4 i13609_2_lut (.A(u_l[3]), .B(\u_s[1] ), .Z(c_15__N_2408[3])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13609_2_lut.init = 16'h8888;
    LUT4 i13595_2_lut (.A(u_l[4]), .B(\u_s[0] ), .Z(c_15__N_2423[3])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13595_2_lut.init = 16'h8888;
    LUT4 i13610_2_lut (.A(u_l[2]), .B(\u_s[1] ), .Z(c_15__N_2408[2])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13610_2_lut.init = 16'h8888;
    LUT4 i13596_2_lut (.A(u_l[3]), .B(\u_s[0] ), .Z(c_15__N_2423[2])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13596_2_lut.init = 16'h8888;
    LUT4 i13611_2_lut (.A(u_l[1]), .B(\u_s[1] ), .Z(c_15__N_2408[1])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13611_2_lut.init = 16'h8888;
    LUT4 i13597_2_lut (.A(u_l[2]), .B(\u_s[0] ), .Z(c_15__N_2423[1])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13597_2_lut.init = 16'h8888;
    LUT4 i12489_2_lut_rep_632 (.A(u_l[1]), .B(\u_s[0] ), .Z(n29292)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i12489_2_lut_rep_632.init = 16'h8888;
    LUT4 i12484_2_lut_rep_633 (.A(u_l[0]), .B(\u_s[1] ), .Z(n29293)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(51[18:45])
    defparam i12484_2_lut_rep_633.init = 16'h8888;
    LUT4 w_r_16__I_0_i2_2_lut_3_lut_4_lut (.A(u_l[0]), .B(\u_s[1] ), .C(\u_s[0] ), 
         .D(u_l[1]), .Z(o_r_17__N_2438[1])) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(51[18:45])
    defparam w_r_16__I_0_i2_2_lut_3_lut_4_lut.init = 16'h7888;
    FD1S3IX o_r__i17 (.D(o_r_17__N_2438[17]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_00[17] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i17.GSR = "DISABLED";
    FD1S3IX o_r__i16 (.D(o_r_17__N_2438[16]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_00[16] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i16.GSR = "DISABLED";
    FD1S3IX o_r__i15 (.D(o_r_17__N_2438[15]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_00[15] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i15.GSR = "DISABLED";
    FD1S3IX o_r__i14 (.D(o_r_17__N_2438[14]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_00[14] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i14.GSR = "DISABLED";
    FD1S3IX o_r__i13 (.D(o_r_17__N_2438[13]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_00[13] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i13.GSR = "DISABLED";
    FD1S3IX o_r__i12 (.D(o_r_17__N_2438[12]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_00[12] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i12.GSR = "DISABLED";
    FD1S3IX o_r__i11 (.D(o_r_17__N_2438[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_00[11] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i11.GSR = "DISABLED";
    FD1S3IX o_r__i10 (.D(o_r_17__N_2438[10]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_00[10] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i10.GSR = "DISABLED";
    FD1S3IX o_r__i9 (.D(o_r_17__N_2438[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_00[9] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i9.GSR = "DISABLED";
    FD1S3IX o_r__i8 (.D(o_r_17__N_2438[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_00[8] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i8.GSR = "DISABLED";
    FD1S3IX o_r__i7 (.D(o_r_17__N_2438[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_00[7] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i7.GSR = "DISABLED";
    FD1S3IX o_r__i6 (.D(o_r_17__N_2438[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_00[6] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i6.GSR = "DISABLED";
    FD1S3IX o_r__i5 (.D(o_r_17__N_2438[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_00[5] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i5.GSR = "DISABLED";
    FD1S3IX o_r__i4 (.D(o_r_17__N_2438[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_00[4] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i4.GSR = "DISABLED";
    FD1S3IX o_r__i3 (.D(o_r_17__N_2438[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_00[3] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i3.GSR = "DISABLED";
    FD1S3IX o_r__i2 (.D(o_r_17__N_2438[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_00[2] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i2.GSR = "DISABLED";
    FD1S3IX o_r__i1 (.D(o_r_17__N_2438[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_1_00_20__N_2184[1] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i1.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module sgnmpy_14x16_U24
//

module sgnmpy_14x16_U24 (u_s, dac_clk_p_c, i_sw0_c, carrier_center_increment_offset, 
            GND_net, \addr_space[2][13] , modulation_output, \addr_space[2][12] , 
            \addr_space[2][10] , \addr_space[2][11] , \addr_space[2][8] , 
            \addr_space[2][9] , \addr_space[2][6] , \addr_space[2][7] , 
            \addr_space[2][4] , \addr_space[2][5] , \addr_space[2][2] , 
            \addr_space[2][3] , \addr_space[2][0] , \addr_space[2][1] , 
            \u_s[12] , \u_s[10] , \u_s[8] , \u_s[6] , \u_s[4] , \u_s[2] , 
            n9444, n9446, n9448, n9450, n9452, n9454, n9456) /* synthesis syn_module_defined=1 */ ;
    output [13:0]u_s;
    input dac_clk_p_c;
    input i_sw0_c;
    output [29:0]carrier_center_increment_offset;
    input GND_net;
    input \addr_space[2][13] ;
    input [15:0]modulation_output;
    input \addr_space[2][12] ;
    input \addr_space[2][10] ;
    input \addr_space[2][11] ;
    input \addr_space[2][8] ;
    input \addr_space[2][9] ;
    input \addr_space[2][6] ;
    input \addr_space[2][7] ;
    input \addr_space[2][4] ;
    input \addr_space[2][5] ;
    input \addr_space[2][2] ;
    input \addr_space[2][3] ;
    input \addr_space[2][0] ;
    input \addr_space[2][1] ;
    output \u_s[12] ;
    output \u_s[10] ;
    output \u_s[8] ;
    output \u_s[6] ;
    output \u_s[4] ;
    output \u_s[2] ;
    input n9444;
    input n9446;
    input n9448;
    input n9450;
    input n9452;
    input n9454;
    input n9456;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[29:38])
    wire [15:0]modulation_output_c /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(86[39:56])
    wire [13:0]u_s_13__N_1951;
    wire [15:0]u_l;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(62[18:21])
    wire [15:0]u_l_15__N_1965;
    wire [4:0]u_sgn;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(63[19:24])
    wire [4:0]u_sgn_4__N_1981;
    wire [29:0]o_p_29__N_1986;
    
    wire n19697;
    wire [29:0]u_r;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(93[21:24])
    wire [29:0]n215;
    
    wire n19696, n19695, n19694, n19693, n19692, n19691, n19690, 
        n19689, n19688, n19687, n19686, n19685, n19684, n19683, 
        n19660, n19659, n19658, n19657, n19656, n19655, n19654, 
        n19653, n19652, n14231, n19651, n19650, n19649, n19648, 
        n19647, n19646;
    wire [13:0]u_s_c;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(61[18:21])
    
    FD1S3IX u_s__i0 (.D(u_s_13__N_1951[0]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_s[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_s__i0.GSR = "DISABLED";
    FD1S3IX u_l__i0 (.D(u_l_15__N_1965[0]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_l[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_l__i0.GSR = "DISABLED";
    FD1S3IX u_sgn__i0 (.D(u_sgn_4__N_1981[0]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_sgn[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(87[9] 91[60])
    defparam u_sgn__i0.GSR = "DISABLED";
    FD1S3IX o_p__i0 (.D(o_p_29__N_1986[0]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(carrier_center_increment_offset[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(98[9] 102[36])
    defparam o_p__i0.GSR = "DISABLED";
    CCU2D unary_minus_20_add_3_31 (.A0(u_r[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n19697), .S0(n215[29]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[25:31])
    defparam unary_minus_20_add_3_31.INIT0 = 16'hf555;
    defparam unary_minus_20_add_3_31.INIT1 = 16'h0000;
    defparam unary_minus_20_add_3_31.INJECT1_0 = "NO";
    defparam unary_minus_20_add_3_31.INJECT1_1 = "NO";
    CCU2D unary_minus_20_add_3_29 (.A0(u_r[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(u_r[28]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n19696), .COUT(n19697), .S0(n215[27]), .S1(n215[28]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[25:31])
    defparam unary_minus_20_add_3_29.INIT0 = 16'hf555;
    defparam unary_minus_20_add_3_29.INIT1 = 16'hf555;
    defparam unary_minus_20_add_3_29.INJECT1_0 = "NO";
    defparam unary_minus_20_add_3_29.INJECT1_1 = "NO";
    CCU2D unary_minus_20_add_3_27 (.A0(u_r[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(u_r[26]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n19695), .COUT(n19696), .S0(n215[25]), .S1(n215[26]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[25:31])
    defparam unary_minus_20_add_3_27.INIT0 = 16'hf555;
    defparam unary_minus_20_add_3_27.INIT1 = 16'hf555;
    defparam unary_minus_20_add_3_27.INJECT1_0 = "NO";
    defparam unary_minus_20_add_3_27.INJECT1_1 = "NO";
    CCU2D unary_minus_20_add_3_25 (.A0(u_r[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(u_r[24]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n19694), .COUT(n19695), .S0(n215[23]), .S1(n215[24]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[25:31])
    defparam unary_minus_20_add_3_25.INIT0 = 16'hf555;
    defparam unary_minus_20_add_3_25.INIT1 = 16'hf555;
    defparam unary_minus_20_add_3_25.INJECT1_0 = "NO";
    defparam unary_minus_20_add_3_25.INJECT1_1 = "NO";
    CCU2D unary_minus_20_add_3_23 (.A0(u_r[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(u_r[22]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n19693), .COUT(n19694), .S0(n215[21]), .S1(n215[22]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[25:31])
    defparam unary_minus_20_add_3_23.INIT0 = 16'hf555;
    defparam unary_minus_20_add_3_23.INIT1 = 16'hf555;
    defparam unary_minus_20_add_3_23.INJECT1_0 = "NO";
    defparam unary_minus_20_add_3_23.INJECT1_1 = "NO";
    CCU2D unary_minus_20_add_3_21 (.A0(u_r[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(u_r[20]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n19692), .COUT(n19693), .S0(n215[19]), .S1(n215[20]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[25:31])
    defparam unary_minus_20_add_3_21.INIT0 = 16'hf555;
    defparam unary_minus_20_add_3_21.INIT1 = 16'hf555;
    defparam unary_minus_20_add_3_21.INJECT1_0 = "NO";
    defparam unary_minus_20_add_3_21.INJECT1_1 = "NO";
    CCU2D unary_minus_20_add_3_19 (.A0(u_r[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(u_r[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n19691), .COUT(n19692), .S0(n215[17]), .S1(n215[18]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[25:31])
    defparam unary_minus_20_add_3_19.INIT0 = 16'hf555;
    defparam unary_minus_20_add_3_19.INIT1 = 16'hf555;
    defparam unary_minus_20_add_3_19.INJECT1_0 = "NO";
    defparam unary_minus_20_add_3_19.INJECT1_1 = "NO";
    CCU2D unary_minus_20_add_3_17 (.A0(u_r[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(u_r[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n19690), .COUT(n19691), .S0(n215[15]), .S1(n215[16]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[25:31])
    defparam unary_minus_20_add_3_17.INIT0 = 16'hf555;
    defparam unary_minus_20_add_3_17.INIT1 = 16'hf555;
    defparam unary_minus_20_add_3_17.INJECT1_0 = "NO";
    defparam unary_minus_20_add_3_17.INJECT1_1 = "NO";
    CCU2D unary_minus_20_add_3_15 (.A0(u_r[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(u_r[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n19689), .COUT(n19690), .S0(n215[13]), .S1(n215[14]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[25:31])
    defparam unary_minus_20_add_3_15.INIT0 = 16'hf555;
    defparam unary_minus_20_add_3_15.INIT1 = 16'hf555;
    defparam unary_minus_20_add_3_15.INJECT1_0 = "NO";
    defparam unary_minus_20_add_3_15.INJECT1_1 = "NO";
    CCU2D unary_minus_20_add_3_13 (.A0(u_r[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(u_r[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n19688), .COUT(n19689), .S0(n215[11]), .S1(n215[12]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[25:31])
    defparam unary_minus_20_add_3_13.INIT0 = 16'hf555;
    defparam unary_minus_20_add_3_13.INIT1 = 16'hf555;
    defparam unary_minus_20_add_3_13.INJECT1_0 = "NO";
    defparam unary_minus_20_add_3_13.INJECT1_1 = "NO";
    CCU2D unary_minus_20_add_3_11 (.A0(u_r[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(u_r[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n19687), .COUT(n19688), .S0(n215[9]), .S1(n215[10]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[25:31])
    defparam unary_minus_20_add_3_11.INIT0 = 16'hf555;
    defparam unary_minus_20_add_3_11.INIT1 = 16'hf555;
    defparam unary_minus_20_add_3_11.INJECT1_0 = "NO";
    defparam unary_minus_20_add_3_11.INJECT1_1 = "NO";
    CCU2D unary_minus_20_add_3_9 (.A0(u_r[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(u_r[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n19686), .COUT(n19687), .S0(n215[7]), .S1(n215[8]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[25:31])
    defparam unary_minus_20_add_3_9.INIT0 = 16'hf555;
    defparam unary_minus_20_add_3_9.INIT1 = 16'hf555;
    defparam unary_minus_20_add_3_9.INJECT1_0 = "NO";
    defparam unary_minus_20_add_3_9.INJECT1_1 = "NO";
    CCU2D unary_minus_20_add_3_7 (.A0(u_r[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(u_r[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n19685), .COUT(n19686), .S0(n215[5]), .S1(n215[6]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[25:31])
    defparam unary_minus_20_add_3_7.INIT0 = 16'hf555;
    defparam unary_minus_20_add_3_7.INIT1 = 16'hf555;
    defparam unary_minus_20_add_3_7.INJECT1_0 = "NO";
    defparam unary_minus_20_add_3_7.INJECT1_1 = "NO";
    CCU2D unary_minus_20_add_3_5 (.A0(u_r[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(u_r[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n19684), .COUT(n19685), .S0(n215[3]), .S1(n215[4]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[25:31])
    defparam unary_minus_20_add_3_5.INIT0 = 16'hf555;
    defparam unary_minus_20_add_3_5.INIT1 = 16'hf555;
    defparam unary_minus_20_add_3_5.INJECT1_0 = "NO";
    defparam unary_minus_20_add_3_5.INJECT1_1 = "NO";
    CCU2D unary_minus_20_add_3_3 (.A0(u_r[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(u_r[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n19683), .COUT(n19684), .S0(n215[1]), .S1(n215[2]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[25:31])
    defparam unary_minus_20_add_3_3.INIT0 = 16'hf555;
    defparam unary_minus_20_add_3_3.INIT1 = 16'hf555;
    defparam unary_minus_20_add_3_3.INJECT1_0 = "NO";
    defparam unary_minus_20_add_3_3.INJECT1_1 = "NO";
    CCU2D unary_minus_20_add_3_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(u_r[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n19683), .S1(n215[0]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[25:31])
    defparam unary_minus_20_add_3_1.INIT0 = 16'hF000;
    defparam unary_minus_20_add_3_1.INIT1 = 16'h0aaa;
    defparam unary_minus_20_add_3_1.INJECT1_0 = "NO";
    defparam unary_minus_20_add_3_1.INJECT1_1 = "NO";
    LUT4 i17_2_lut (.A(\addr_space[2][13] ), .B(modulation_output[15]), 
         .Z(u_sgn_4__N_1981[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(91[32:57])
    defparam i17_2_lut.init = 16'h6666;
    LUT4 mux_21_i1_3_lut (.A(u_r[0]), .B(n215[0]), .C(u_sgn[4]), .Z(o_p_29__N_1986[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[10:35])
    defparam mux_21_i1_3_lut.init = 16'hcaca;
    CCU2D unary_minus_8_add_3_17 (.A0(modulation_output[14]), .B0(modulation_output[15]), 
          .C0(GND_net), .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n19660), .S0(u_l_15__N_1965[15]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(83[22:28])
    defparam unary_minus_8_add_3_17.INIT0 = 16'hd111;
    defparam unary_minus_8_add_3_17.INIT1 = 16'h0000;
    defparam unary_minus_8_add_3_17.INJECT1_0 = "NO";
    defparam unary_minus_8_add_3_17.INJECT1_1 = "NO";
    CCU2D unary_minus_8_add_3_15 (.A0(modulation_output[12]), .B0(modulation_output[15]), 
          .C0(modulation_output[13]), .D0(GND_net), .A1(modulation_output[13]), 
          .B1(modulation_output[15]), .C1(modulation_output[14]), .D1(GND_net), 
          .CIN(n19659), .COUT(n19660), .S0(u_l_15__N_1965[13]), .S1(u_l_15__N_1965[14]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(83[22:28])
    defparam unary_minus_8_add_3_15.INIT0 = 16'hdd2d;
    defparam unary_minus_8_add_3_15.INIT1 = 16'hdd2d;
    defparam unary_minus_8_add_3_15.INJECT1_0 = "NO";
    defparam unary_minus_8_add_3_15.INJECT1_1 = "NO";
    CCU2D unary_minus_8_add_3_13 (.A0(modulation_output[10]), .B0(modulation_output[15]), 
          .C0(modulation_output[11]), .D0(GND_net), .A1(modulation_output[11]), 
          .B1(modulation_output[15]), .C1(modulation_output[12]), .D1(GND_net), 
          .CIN(n19658), .COUT(n19659), .S0(u_l_15__N_1965[11]), .S1(u_l_15__N_1965[12]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(83[22:28])
    defparam unary_minus_8_add_3_13.INIT0 = 16'hdd2d;
    defparam unary_minus_8_add_3_13.INIT1 = 16'hdd2d;
    defparam unary_minus_8_add_3_13.INJECT1_0 = "NO";
    defparam unary_minus_8_add_3_13.INJECT1_1 = "NO";
    CCU2D unary_minus_8_add_3_11 (.A0(modulation_output[8]), .B0(modulation_output[15]), 
          .C0(modulation_output[9]), .D0(GND_net), .A1(modulation_output[9]), 
          .B1(modulation_output[15]), .C1(modulation_output[10]), .D1(GND_net), 
          .CIN(n19657), .COUT(n19658), .S0(u_l_15__N_1965[9]), .S1(u_l_15__N_1965[10]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(83[22:28])
    defparam unary_minus_8_add_3_11.INIT0 = 16'hdd2d;
    defparam unary_minus_8_add_3_11.INIT1 = 16'hdd2d;
    defparam unary_minus_8_add_3_11.INJECT1_0 = "NO";
    defparam unary_minus_8_add_3_11.INJECT1_1 = "NO";
    CCU2D unary_minus_8_add_3_9 (.A0(modulation_output[6]), .B0(modulation_output[15]), 
          .C0(modulation_output[7]), .D0(GND_net), .A1(modulation_output[7]), 
          .B1(modulation_output[15]), .C1(modulation_output[8]), .D1(GND_net), 
          .CIN(n19656), .COUT(n19657), .S0(u_l_15__N_1965[7]), .S1(u_l_15__N_1965[8]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(83[22:28])
    defparam unary_minus_8_add_3_9.INIT0 = 16'hdd2d;
    defparam unary_minus_8_add_3_9.INIT1 = 16'hdd2d;
    defparam unary_minus_8_add_3_9.INJECT1_0 = "NO";
    defparam unary_minus_8_add_3_9.INJECT1_1 = "NO";
    CCU2D unary_minus_8_add_3_7 (.A0(modulation_output[4]), .B0(modulation_output[15]), 
          .C0(modulation_output[5]), .D0(GND_net), .A1(modulation_output[5]), 
          .B1(modulation_output[15]), .C1(modulation_output[6]), .D1(GND_net), 
          .CIN(n19655), .COUT(n19656), .S0(u_l_15__N_1965[5]), .S1(u_l_15__N_1965[6]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(83[22:28])
    defparam unary_minus_8_add_3_7.INIT0 = 16'hdd2d;
    defparam unary_minus_8_add_3_7.INIT1 = 16'hdd2d;
    defparam unary_minus_8_add_3_7.INJECT1_0 = "NO";
    defparam unary_minus_8_add_3_7.INJECT1_1 = "NO";
    CCU2D unary_minus_8_add_3_5 (.A0(modulation_output[2]), .B0(modulation_output[15]), 
          .C0(modulation_output[3]), .D0(GND_net), .A1(modulation_output[3]), 
          .B1(modulation_output[15]), .C1(modulation_output[4]), .D1(GND_net), 
          .CIN(n19654), .COUT(n19655), .S0(u_l_15__N_1965[3]), .S1(u_l_15__N_1965[4]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(83[22:28])
    defparam unary_minus_8_add_3_5.INIT0 = 16'hdd2d;
    defparam unary_minus_8_add_3_5.INIT1 = 16'hdd2d;
    defparam unary_minus_8_add_3_5.INJECT1_0 = "NO";
    defparam unary_minus_8_add_3_5.INJECT1_1 = "NO";
    CCU2D unary_minus_8_add_3_3 (.A0(modulation_output[0]), .B0(modulation_output[15]), 
          .C0(modulation_output[1]), .D0(GND_net), .A1(modulation_output[1]), 
          .B1(modulation_output[15]), .C1(modulation_output[2]), .D1(GND_net), 
          .CIN(n19653), .COUT(n19654), .S0(u_l_15__N_1965[1]), .S1(u_l_15__N_1965[2]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(83[22:28])
    defparam unary_minus_8_add_3_3.INIT0 = 16'hdd2d;
    defparam unary_minus_8_add_3_3.INIT1 = 16'hdd2d;
    defparam unary_minus_8_add_3_3.INJECT1_0 = "NO";
    defparam unary_minus_8_add_3_3.INJECT1_1 = "NO";
    CCU2D unary_minus_8_add_3_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(modulation_output[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n19653), .S1(u_l_15__N_1965[0]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(83[22:28])
    defparam unary_minus_8_add_3_1.INIT0 = 16'hF000;
    defparam unary_minus_8_add_3_1.INIT1 = 16'h0aaa;
    defparam unary_minus_8_add_3_1.INJECT1_0 = "NO";
    defparam unary_minus_8_add_3_1.INJECT1_1 = "NO";
    CCU2D unary_minus_6_add_3_15 (.A0(\addr_space[2][12] ), .B0(\addr_space[2][13] ), 
          .C0(GND_net), .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n19652), .S0(u_s_13__N_1951[13]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(82[22:28])
    defparam unary_minus_6_add_3_15.INIT0 = 16'hd111;
    defparam unary_minus_6_add_3_15.INIT1 = 16'h0000;
    defparam unary_minus_6_add_3_15.INJECT1_0 = "NO";
    defparam unary_minus_6_add_3_15.INJECT1_1 = "NO";
    LUT4 i11855_1_lut (.A(u_l[0]), .Z(n14231)) /* synthesis lut_function=(!(A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam i11855_1_lut.init = 16'h5555;
    CCU2D unary_minus_6_add_3_13 (.A0(\addr_space[2][10] ), .B0(\addr_space[2][13] ), 
          .C0(\addr_space[2][11] ), .D0(GND_net), .A1(\addr_space[2][11] ), 
          .B1(\addr_space[2][13] ), .C1(\addr_space[2][12] ), .D1(GND_net), 
          .CIN(n19651), .COUT(n19652), .S0(u_s_13__N_1951[11]), .S1(u_s_13__N_1951[12]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(82[22:28])
    defparam unary_minus_6_add_3_13.INIT0 = 16'hdd2d;
    defparam unary_minus_6_add_3_13.INIT1 = 16'hdd2d;
    defparam unary_minus_6_add_3_13.INJECT1_0 = "NO";
    defparam unary_minus_6_add_3_13.INJECT1_1 = "NO";
    CCU2D unary_minus_6_add_3_11 (.A0(\addr_space[2][8] ), .B0(\addr_space[2][13] ), 
          .C0(\addr_space[2][9] ), .D0(GND_net), .A1(\addr_space[2][9] ), 
          .B1(\addr_space[2][13] ), .C1(\addr_space[2][10] ), .D1(GND_net), 
          .CIN(n19650), .COUT(n19651), .S0(u_s_13__N_1951[9]), .S1(u_s_13__N_1951[10]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(82[22:28])
    defparam unary_minus_6_add_3_11.INIT0 = 16'hdd2d;
    defparam unary_minus_6_add_3_11.INIT1 = 16'hdd2d;
    defparam unary_minus_6_add_3_11.INJECT1_0 = "NO";
    defparam unary_minus_6_add_3_11.INJECT1_1 = "NO";
    CCU2D unary_minus_6_add_3_9 (.A0(\addr_space[2][6] ), .B0(\addr_space[2][13] ), 
          .C0(\addr_space[2][7] ), .D0(GND_net), .A1(\addr_space[2][7] ), 
          .B1(\addr_space[2][13] ), .C1(\addr_space[2][8] ), .D1(GND_net), 
          .CIN(n19649), .COUT(n19650), .S0(u_s_13__N_1951[7]), .S1(u_s_13__N_1951[8]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(82[22:28])
    defparam unary_minus_6_add_3_9.INIT0 = 16'hdd2d;
    defparam unary_minus_6_add_3_9.INIT1 = 16'hdd2d;
    defparam unary_minus_6_add_3_9.INJECT1_0 = "NO";
    defparam unary_minus_6_add_3_9.INJECT1_1 = "NO";
    CCU2D unary_minus_6_add_3_7 (.A0(\addr_space[2][4] ), .B0(\addr_space[2][13] ), 
          .C0(\addr_space[2][5] ), .D0(GND_net), .A1(\addr_space[2][5] ), 
          .B1(\addr_space[2][13] ), .C1(\addr_space[2][6] ), .D1(GND_net), 
          .CIN(n19648), .COUT(n19649), .S0(u_s_13__N_1951[5]), .S1(u_s_13__N_1951[6]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(82[22:28])
    defparam unary_minus_6_add_3_7.INIT0 = 16'hdd2d;
    defparam unary_minus_6_add_3_7.INIT1 = 16'hdd2d;
    defparam unary_minus_6_add_3_7.INJECT1_0 = "NO";
    defparam unary_minus_6_add_3_7.INJECT1_1 = "NO";
    CCU2D unary_minus_6_add_3_5 (.A0(\addr_space[2][2] ), .B0(\addr_space[2][13] ), 
          .C0(\addr_space[2][3] ), .D0(GND_net), .A1(\addr_space[2][3] ), 
          .B1(\addr_space[2][13] ), .C1(\addr_space[2][4] ), .D1(GND_net), 
          .CIN(n19647), .COUT(n19648), .S0(u_s_13__N_1951[3]), .S1(u_s_13__N_1951[4]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(82[22:28])
    defparam unary_minus_6_add_3_5.INIT0 = 16'hdd2d;
    defparam unary_minus_6_add_3_5.INIT1 = 16'hdd2d;
    defparam unary_minus_6_add_3_5.INJECT1_0 = "NO";
    defparam unary_minus_6_add_3_5.INJECT1_1 = "NO";
    CCU2D unary_minus_6_add_3_3 (.A0(\addr_space[2][0] ), .B0(\addr_space[2][13] ), 
          .C0(\addr_space[2][1] ), .D0(GND_net), .A1(\addr_space[2][1] ), 
          .B1(\addr_space[2][13] ), .C1(\addr_space[2][2] ), .D1(GND_net), 
          .CIN(n19646), .COUT(n19647), .S0(u_s_13__N_1951[1]), .S1(u_s_13__N_1951[2]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(82[22:28])
    defparam unary_minus_6_add_3_3.INIT0 = 16'hdd2d;
    defparam unary_minus_6_add_3_3.INIT1 = 16'hdd2d;
    defparam unary_minus_6_add_3_3.INJECT1_0 = "NO";
    defparam unary_minus_6_add_3_3.INJECT1_1 = "NO";
    CCU2D unary_minus_6_add_3_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\addr_space[2][0] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n19646), .S1(u_s_13__N_1951[0]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(82[22:28])
    defparam unary_minus_6_add_3_1.INIT0 = 16'hF000;
    defparam unary_minus_6_add_3_1.INIT1 = 16'h0aaa;
    defparam unary_minus_6_add_3_1.INJECT1_0 = "NO";
    defparam unary_minus_6_add_3_1.INJECT1_1 = "NO";
    LUT4 mux_21_i30_3_lut (.A(u_r[29]), .B(n215[29]), .C(u_sgn[4]), .Z(o_p_29__N_1986[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[10:35])
    defparam mux_21_i30_3_lut.init = 16'hcaca;
    LUT4 mux_21_i29_3_lut (.A(u_r[28]), .B(n215[28]), .C(u_sgn[4]), .Z(o_p_29__N_1986[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[10:35])
    defparam mux_21_i29_3_lut.init = 16'hcaca;
    LUT4 mux_21_i28_3_lut (.A(u_r[27]), .B(n215[27]), .C(u_sgn[4]), .Z(o_p_29__N_1986[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[10:35])
    defparam mux_21_i28_3_lut.init = 16'hcaca;
    LUT4 mux_21_i27_3_lut (.A(u_r[26]), .B(n215[26]), .C(u_sgn[4]), .Z(o_p_29__N_1986[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[10:35])
    defparam mux_21_i27_3_lut.init = 16'hcaca;
    LUT4 mux_21_i26_3_lut (.A(u_r[25]), .B(n215[25]), .C(u_sgn[4]), .Z(o_p_29__N_1986[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[10:35])
    defparam mux_21_i26_3_lut.init = 16'hcaca;
    LUT4 mux_21_i25_3_lut (.A(u_r[24]), .B(n215[24]), .C(u_sgn[4]), .Z(o_p_29__N_1986[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[10:35])
    defparam mux_21_i25_3_lut.init = 16'hcaca;
    LUT4 mux_21_i24_3_lut (.A(u_r[23]), .B(n215[23]), .C(u_sgn[4]), .Z(o_p_29__N_1986[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[10:35])
    defparam mux_21_i24_3_lut.init = 16'hcaca;
    LUT4 mux_21_i23_3_lut (.A(u_r[22]), .B(n215[22]), .C(u_sgn[4]), .Z(o_p_29__N_1986[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[10:35])
    defparam mux_21_i23_3_lut.init = 16'hcaca;
    LUT4 mux_21_i22_3_lut (.A(u_r[21]), .B(n215[21]), .C(u_sgn[4]), .Z(o_p_29__N_1986[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[10:35])
    defparam mux_21_i22_3_lut.init = 16'hcaca;
    LUT4 mux_21_i21_3_lut (.A(u_r[20]), .B(n215[20]), .C(u_sgn[4]), .Z(o_p_29__N_1986[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[10:35])
    defparam mux_21_i21_3_lut.init = 16'hcaca;
    LUT4 mux_21_i20_3_lut (.A(u_r[19]), .B(n215[19]), .C(u_sgn[4]), .Z(o_p_29__N_1986[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[10:35])
    defparam mux_21_i20_3_lut.init = 16'hcaca;
    LUT4 mux_21_i19_3_lut (.A(u_r[18]), .B(n215[18]), .C(u_sgn[4]), .Z(o_p_29__N_1986[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[10:35])
    defparam mux_21_i19_3_lut.init = 16'hcaca;
    LUT4 mux_21_i18_3_lut (.A(u_r[17]), .B(n215[17]), .C(u_sgn[4]), .Z(o_p_29__N_1986[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[10:35])
    defparam mux_21_i18_3_lut.init = 16'hcaca;
    LUT4 mux_21_i17_3_lut (.A(u_r[16]), .B(n215[16]), .C(u_sgn[4]), .Z(o_p_29__N_1986[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[10:35])
    defparam mux_21_i17_3_lut.init = 16'hcaca;
    LUT4 mux_21_i16_3_lut (.A(u_r[15]), .B(n215[15]), .C(u_sgn[4]), .Z(o_p_29__N_1986[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[10:35])
    defparam mux_21_i16_3_lut.init = 16'hcaca;
    LUT4 mux_21_i15_3_lut (.A(u_r[14]), .B(n215[14]), .C(u_sgn[4]), .Z(o_p_29__N_1986[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[10:35])
    defparam mux_21_i15_3_lut.init = 16'hcaca;
    LUT4 mux_21_i14_3_lut (.A(u_r[13]), .B(n215[13]), .C(u_sgn[4]), .Z(o_p_29__N_1986[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[10:35])
    defparam mux_21_i14_3_lut.init = 16'hcaca;
    LUT4 mux_21_i13_3_lut (.A(u_r[12]), .B(n215[12]), .C(u_sgn[4]), .Z(o_p_29__N_1986[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[10:35])
    defparam mux_21_i13_3_lut.init = 16'hcaca;
    LUT4 mux_21_i12_3_lut (.A(u_r[11]), .B(n215[11]), .C(u_sgn[4]), .Z(o_p_29__N_1986[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[10:35])
    defparam mux_21_i12_3_lut.init = 16'hcaca;
    LUT4 mux_21_i11_3_lut (.A(u_r[10]), .B(n215[10]), .C(u_sgn[4]), .Z(o_p_29__N_1986[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[10:35])
    defparam mux_21_i11_3_lut.init = 16'hcaca;
    LUT4 mux_21_i10_3_lut (.A(u_r[9]), .B(n215[9]), .C(u_sgn[4]), .Z(o_p_29__N_1986[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[10:35])
    defparam mux_21_i10_3_lut.init = 16'hcaca;
    LUT4 mux_21_i9_3_lut (.A(u_r[8]), .B(n215[8]), .C(u_sgn[4]), .Z(o_p_29__N_1986[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[10:35])
    defparam mux_21_i9_3_lut.init = 16'hcaca;
    LUT4 mux_21_i8_3_lut (.A(u_r[7]), .B(n215[7]), .C(u_sgn[4]), .Z(o_p_29__N_1986[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[10:35])
    defparam mux_21_i8_3_lut.init = 16'hcaca;
    LUT4 mux_21_i7_3_lut (.A(u_r[6]), .B(n215[6]), .C(u_sgn[4]), .Z(o_p_29__N_1986[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[10:35])
    defparam mux_21_i7_3_lut.init = 16'hcaca;
    LUT4 mux_21_i6_3_lut (.A(u_r[5]), .B(n215[5]), .C(u_sgn[4]), .Z(o_p_29__N_1986[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[10:35])
    defparam mux_21_i6_3_lut.init = 16'hcaca;
    LUT4 mux_21_i5_3_lut (.A(u_r[4]), .B(n215[4]), .C(u_sgn[4]), .Z(o_p_29__N_1986[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[10:35])
    defparam mux_21_i5_3_lut.init = 16'hcaca;
    LUT4 mux_21_i4_3_lut (.A(u_r[3]), .B(n215[3]), .C(u_sgn[4]), .Z(o_p_29__N_1986[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[10:35])
    defparam mux_21_i4_3_lut.init = 16'hcaca;
    LUT4 mux_21_i3_3_lut (.A(u_r[2]), .B(n215[2]), .C(u_sgn[4]), .Z(o_p_29__N_1986[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[10:35])
    defparam mux_21_i3_3_lut.init = 16'hcaca;
    LUT4 mux_21_i2_3_lut (.A(u_r[1]), .B(n215[1]), .C(u_sgn[4]), .Z(o_p_29__N_1986[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[10:35])
    defparam mux_21_i2_3_lut.init = 16'hcaca;
    FD1S3IX o_p__i29 (.D(o_p_29__N_1986[29]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(carrier_center_increment_offset[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(98[9] 102[36])
    defparam o_p__i29.GSR = "DISABLED";
    FD1S3IX o_p__i28 (.D(o_p_29__N_1986[28]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(carrier_center_increment_offset[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(98[9] 102[36])
    defparam o_p__i28.GSR = "DISABLED";
    FD1S3IX o_p__i27 (.D(o_p_29__N_1986[27]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(carrier_center_increment_offset[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(98[9] 102[36])
    defparam o_p__i27.GSR = "DISABLED";
    FD1S3IX o_p__i26 (.D(o_p_29__N_1986[26]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(carrier_center_increment_offset[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(98[9] 102[36])
    defparam o_p__i26.GSR = "DISABLED";
    FD1S3IX o_p__i25 (.D(o_p_29__N_1986[25]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(carrier_center_increment_offset[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(98[9] 102[36])
    defparam o_p__i25.GSR = "DISABLED";
    FD1S3IX o_p__i24 (.D(o_p_29__N_1986[24]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(carrier_center_increment_offset[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(98[9] 102[36])
    defparam o_p__i24.GSR = "DISABLED";
    FD1S3IX o_p__i23 (.D(o_p_29__N_1986[23]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(carrier_center_increment_offset[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(98[9] 102[36])
    defparam o_p__i23.GSR = "DISABLED";
    FD1S3IX o_p__i22 (.D(o_p_29__N_1986[22]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(carrier_center_increment_offset[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(98[9] 102[36])
    defparam o_p__i22.GSR = "DISABLED";
    FD1S3IX o_p__i21 (.D(o_p_29__N_1986[21]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(carrier_center_increment_offset[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(98[9] 102[36])
    defparam o_p__i21.GSR = "DISABLED";
    FD1S3IX o_p__i20 (.D(o_p_29__N_1986[20]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(carrier_center_increment_offset[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(98[9] 102[36])
    defparam o_p__i20.GSR = "DISABLED";
    FD1S3IX o_p__i19 (.D(o_p_29__N_1986[19]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(carrier_center_increment_offset[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(98[9] 102[36])
    defparam o_p__i19.GSR = "DISABLED";
    FD1S3IX o_p__i18 (.D(o_p_29__N_1986[18]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(carrier_center_increment_offset[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(98[9] 102[36])
    defparam o_p__i18.GSR = "DISABLED";
    FD1S3IX o_p__i17 (.D(o_p_29__N_1986[17]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(carrier_center_increment_offset[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(98[9] 102[36])
    defparam o_p__i17.GSR = "DISABLED";
    FD1S3IX o_p__i16 (.D(o_p_29__N_1986[16]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(carrier_center_increment_offset[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(98[9] 102[36])
    defparam o_p__i16.GSR = "DISABLED";
    FD1S3IX o_p__i15 (.D(o_p_29__N_1986[15]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(carrier_center_increment_offset[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(98[9] 102[36])
    defparam o_p__i15.GSR = "DISABLED";
    FD1S3IX o_p__i14 (.D(o_p_29__N_1986[14]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(carrier_center_increment_offset[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(98[9] 102[36])
    defparam o_p__i14.GSR = "DISABLED";
    FD1S3IX o_p__i13 (.D(o_p_29__N_1986[13]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(carrier_center_increment_offset[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(98[9] 102[36])
    defparam o_p__i13.GSR = "DISABLED";
    FD1S3IX o_p__i12 (.D(o_p_29__N_1986[12]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(carrier_center_increment_offset[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(98[9] 102[36])
    defparam o_p__i12.GSR = "DISABLED";
    FD1S3IX o_p__i11 (.D(o_p_29__N_1986[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(carrier_center_increment_offset[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(98[9] 102[36])
    defparam o_p__i11.GSR = "DISABLED";
    FD1S3IX o_p__i10 (.D(o_p_29__N_1986[10]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(carrier_center_increment_offset[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(98[9] 102[36])
    defparam o_p__i10.GSR = "DISABLED";
    FD1S3IX o_p__i9 (.D(o_p_29__N_1986[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(carrier_center_increment_offset[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(98[9] 102[36])
    defparam o_p__i9.GSR = "DISABLED";
    FD1S3IX o_p__i8 (.D(o_p_29__N_1986[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(carrier_center_increment_offset[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(98[9] 102[36])
    defparam o_p__i8.GSR = "DISABLED";
    FD1S3IX o_p__i7 (.D(o_p_29__N_1986[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(carrier_center_increment_offset[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(98[9] 102[36])
    defparam o_p__i7.GSR = "DISABLED";
    FD1S3IX o_p__i6 (.D(o_p_29__N_1986[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(carrier_center_increment_offset[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(98[9] 102[36])
    defparam o_p__i6.GSR = "DISABLED";
    FD1S3IX o_p__i5 (.D(o_p_29__N_1986[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(carrier_center_increment_offset[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(98[9] 102[36])
    defparam o_p__i5.GSR = "DISABLED";
    FD1S3IX o_p__i4 (.D(o_p_29__N_1986[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(carrier_center_increment_offset[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(98[9] 102[36])
    defparam o_p__i4.GSR = "DISABLED";
    FD1S3IX o_p__i3 (.D(o_p_29__N_1986[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(carrier_center_increment_offset[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(98[9] 102[36])
    defparam o_p__i3.GSR = "DISABLED";
    FD1S3IX o_p__i2 (.D(o_p_29__N_1986[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(carrier_center_increment_offset[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(98[9] 102[36])
    defparam o_p__i2.GSR = "DISABLED";
    FD1S3IX o_p__i1 (.D(o_p_29__N_1986[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(carrier_center_increment_offset[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(98[9] 102[36])
    defparam o_p__i1.GSR = "DISABLED";
    FD1S3IX u_sgn__i4 (.D(u_sgn[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(u_sgn[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(87[9] 91[60])
    defparam u_sgn__i4.GSR = "DISABLED";
    FD1S3IX u_sgn__i3 (.D(u_sgn[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(u_sgn[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(87[9] 91[60])
    defparam u_sgn__i3.GSR = "DISABLED";
    FD1S3IX u_sgn__i2 (.D(u_sgn[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(u_sgn[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(87[9] 91[60])
    defparam u_sgn__i2.GSR = "DISABLED";
    FD1S3IX u_sgn__i1 (.D(u_sgn[0]), .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(u_sgn[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(87[9] 91[60])
    defparam u_sgn__i1.GSR = "DISABLED";
    FD1S3IX u_l__i15 (.D(u_l_15__N_1965[15]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_l[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_l__i15.GSR = "DISABLED";
    FD1S3IX u_l__i14 (.D(u_l_15__N_1965[14]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_l[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_l__i14.GSR = "DISABLED";
    FD1S3IX u_l__i13 (.D(u_l_15__N_1965[13]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_l[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_l__i13.GSR = "DISABLED";
    FD1S3IX u_l__i12 (.D(u_l_15__N_1965[12]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_l[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_l__i12.GSR = "DISABLED";
    FD1S3IX u_l__i11 (.D(u_l_15__N_1965[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_l[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_l__i11.GSR = "DISABLED";
    FD1S3IX u_l__i10 (.D(u_l_15__N_1965[10]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_l[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_l__i10.GSR = "DISABLED";
    FD1S3IX u_l__i9 (.D(u_l_15__N_1965[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_l[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_l__i9.GSR = "DISABLED";
    FD1S3IX u_l__i8 (.D(u_l_15__N_1965[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_l[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_l__i8.GSR = "DISABLED";
    FD1S3IX u_l__i7 (.D(u_l_15__N_1965[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_l[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_l__i7.GSR = "DISABLED";
    FD1S3IX u_l__i6 (.D(u_l_15__N_1965[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_l[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_l__i6.GSR = "DISABLED";
    FD1S3IX u_l__i5 (.D(u_l_15__N_1965[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_l[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_l__i5.GSR = "DISABLED";
    FD1S3IX u_l__i4 (.D(u_l_15__N_1965[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_l[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_l__i4.GSR = "DISABLED";
    FD1S3IX u_l__i3 (.D(u_l_15__N_1965[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_l[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_l__i3.GSR = "DISABLED";
    FD1S3IX u_l__i2 (.D(u_l_15__N_1965[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_l[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_l__i2.GSR = "DISABLED";
    FD1S3IX u_l__i1 (.D(u_l_15__N_1965[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_l[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_l__i1.GSR = "DISABLED";
    FD1S3IX u_s__i13 (.D(u_s_13__N_1951[13]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_s_c[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_s__i13.GSR = "DISABLED";
    FD1S3IX u_s__i12 (.D(u_s_13__N_1951[12]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\u_s[12] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_s__i12.GSR = "DISABLED";
    FD1S3IX u_s__i11 (.D(u_s_13__N_1951[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_s_c[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_s__i11.GSR = "DISABLED";
    FD1S3IX u_s__i10 (.D(u_s_13__N_1951[10]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\u_s[10] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_s__i10.GSR = "DISABLED";
    FD1S3IX u_s__i9 (.D(u_s_13__N_1951[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_s_c[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_s__i9.GSR = "DISABLED";
    FD1S3IX u_s__i8 (.D(u_s_13__N_1951[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\u_s[8] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_s__i8.GSR = "DISABLED";
    FD1S3IX u_s__i7 (.D(u_s_13__N_1951[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_s_c[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_s__i7.GSR = "DISABLED";
    FD1S3IX u_s__i6 (.D(u_s_13__N_1951[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\u_s[6] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_s__i6.GSR = "DISABLED";
    FD1S3IX u_s__i5 (.D(u_s_13__N_1951[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_s_c[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_s__i5.GSR = "DISABLED";
    FD1S3IX u_s__i4 (.D(u_s_13__N_1951[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\u_s[4] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_s__i4.GSR = "DISABLED";
    FD1S3IX u_s__i3 (.D(u_s_13__N_1951[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_s_c[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_s__i3.GSR = "DISABLED";
    FD1S3IX u_s__i2 (.D(u_s_13__N_1951[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\u_s[2] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_s__i2.GSR = "DISABLED";
    FD1S3IX u_s__i1 (.D(u_s_13__N_1951[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_s_c[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=154, LSE_LLINE=113, LSE_RLINE=113 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_s__i1.GSR = "DISABLED";
    umpy_14x16_U20 umpy (.dac_clk_p_c(dac_clk_p_c), .i_sw0_c(i_sw0_c), .u_r({u_r}), 
            .GND_net(GND_net), .u_l({u_l}), .u_s({u_s_c[13], \u_s[12] , 
            u_s_c[11], \u_s[10] , u_s_c[9], \u_s[8] , u_s_c[7], \u_s[6] , 
            u_s_c[5], \u_s[4] , u_s_c[3], \u_s[2] , u_s_c[1], u_s[0]}), 
            .n14231(n14231), .n9444(n9444), .n9446(n9446), .n9448(n9448), 
            .n9450(n9450), .n9452(n9452), .n9454(n9454), .n9456(n9456)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(95[13:68])
    
endmodule
//
// Verilog Description of module umpy_14x16_U20
//

module umpy_14x16_U20 (dac_clk_p_c, i_sw0_c, u_r, GND_net, u_l, u_s, 
            n14231, n9444, n9446, n9448, n9450, n9452, n9454, 
            n9456) /* synthesis syn_module_defined=1 */ ;
    input dac_clk_p_c;
    input i_sw0_c;
    output [29:0]u_r;
    input GND_net;
    input [15:0]u_l;
    input [13:0]u_s;
    input n14231;
    input n9444;
    input n9446;
    input n9448;
    input n9450;
    input n9452;
    input n9454;
    input n9456;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[29:38])
    wire [20:0]S_1_00;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(103[17:23])
    wire [17:0]S_0_00;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(71[14:20])
    wire [20:0]S_1_01;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(104[17:23])
    wire [17:0]S_0_02;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(77[14:20])
    wire [25:0]S_2_01_25__N_2294;
    wire [17:0]S_0_04;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(83[14:20])
    wire [20:0]S_1_03;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(106[17:23])
    wire [17:0]S_0_06;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(89[14:20])
    wire [29:0]o_p_29__N_2320;
    wire [25:0]S_2_01;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(140[17:23])
    
    wire n19671, n19670, n19669;
    wire [25:0]S_2_00;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(139[17:23])
    
    wire n19833;
    wire [20:0]S_1_01_20__N_2205;
    
    wire n19832;
    wire [17:0]S_0_03;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(80[14:20])
    
    wire n19668, n19667, n19666, n19665, n19831, n19830, n19664, 
        n19663, n19829, n19662, n19828, n19827, n19826, n19825, 
        n19823;
    wire [20:0]S_1_02_20__N_2226;
    
    wire n19822;
    wire [17:0]S_0_05;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(86[14:20])
    
    wire n19821, n19820, n19819, n19818, n19817, n19816, n19815, 
        n19813;
    wire [25:0]S_2_00_25__N_2268;
    
    wire n19812, n19811, n19810, n19809, n19808, n19807, n19806, 
        n19805, n19804, n19763;
    wire [20:0]S_1_00_20__N_2184;
    
    wire n19762;
    wire [17:0]S_0_01;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(74[14:20])
    
    wire n19761, n19607;
    wire [20:0]S_1_02;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(105[17:23])
    
    wire n19606, n19605, n19760, n19759, n19758, n19757, n19604, 
        n19756, n19603, n19602, n19755, n19601, n19600;
    
    FD1S3IX S_1_00__i0 (.D(S_0_00[0]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_00[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i0.GSR = "DISABLED";
    FD1S3IX S_1_01__i0 (.D(S_0_02[0]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i0.GSR = "DISABLED";
    FD1S3IX S_1_02__i1 (.D(S_0_04[0]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01_25__N_2294[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i1.GSR = "DISABLED";
    FD1S3IX S_1_03__i1 (.D(S_0_06[0]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_03[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_03__i1.GSR = "DISABLED";
    FD1S3IX S_2_00__i1 (.D(S_1_00[0]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_p_29__N_2320[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i1.GSR = "DISABLED";
    FD1S3IX S_2_01__i1 (.D(S_2_01_25__N_2294[0]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i1.GSR = "DISABLED";
    FD1S3IX S_3_00__i0 (.D(o_p_29__N_2320[0]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i0.GSR = "DISABLED";
    CCU2D add_35_22 (.A0(S_2_01[20]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(S_2_01[21]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n19671), .S0(o_p_29__N_2320[28]), .S1(o_p_29__N_2320[29]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(177[13] 178[15])
    defparam add_35_22.INIT0 = 16'hfaaa;
    defparam add_35_22.INIT1 = 16'hfaaa;
    defparam add_35_22.INJECT1_0 = "NO";
    defparam add_35_22.INJECT1_1 = "NO";
    CCU2D add_35_20 (.A0(S_2_01[18]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(S_2_01[19]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n19670), .COUT(n19671), .S0(o_p_29__N_2320[26]), .S1(o_p_29__N_2320[27]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(177[13] 178[15])
    defparam add_35_20.INIT0 = 16'hfaaa;
    defparam add_35_20.INIT1 = 16'hfaaa;
    defparam add_35_20.INJECT1_0 = "NO";
    defparam add_35_20.INJECT1_1 = "NO";
    CCU2D add_35_18 (.A0(S_2_00[24]), .B0(S_2_01[16]), .C0(GND_net), .D0(GND_net), 
          .A1(S_2_00[25]), .B1(S_2_01[17]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19669), .COUT(n19670), .S0(o_p_29__N_2320[24]), .S1(o_p_29__N_2320[25]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(177[13] 178[15])
    defparam add_35_18.INIT0 = 16'h5666;
    defparam add_35_18.INIT1 = 16'h5666;
    defparam add_35_18.INJECT1_0 = "NO";
    defparam add_35_18.INJECT1_1 = "NO";
    CCU2D add_845_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19833), 
          .S0(S_1_01_20__N_2205[20]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(123[13:48])
    defparam add_845_cout.INIT0 = 16'h0000;
    defparam add_845_cout.INIT1 = 16'h0000;
    defparam add_845_cout.INJECT1_0 = "NO";
    defparam add_845_cout.INJECT1_1 = "NO";
    CCU2D add_845_18 (.A0(S_0_03[16]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(S_0_03[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n19832), .COUT(n19833), .S0(S_1_01_20__N_2205[18]), .S1(S_1_01_20__N_2205[19]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(123[13:48])
    defparam add_845_18.INIT0 = 16'hfaaa;
    defparam add_845_18.INIT1 = 16'hfaaa;
    defparam add_845_18.INJECT1_0 = "NO";
    defparam add_845_18.INJECT1_1 = "NO";
    CCU2D add_35_16 (.A0(S_2_00[22]), .B0(S_2_01[14]), .C0(GND_net), .D0(GND_net), 
          .A1(S_2_00[23]), .B1(S_2_01[15]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19668), .COUT(n19669), .S0(o_p_29__N_2320[22]), .S1(o_p_29__N_2320[23]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(177[13] 178[15])
    defparam add_35_16.INIT0 = 16'h5666;
    defparam add_35_16.INIT1 = 16'h5666;
    defparam add_35_16.INJECT1_0 = "NO";
    defparam add_35_16.INJECT1_1 = "NO";
    CCU2D add_35_14 (.A0(S_2_00[20]), .B0(S_2_01[12]), .C0(GND_net), .D0(GND_net), 
          .A1(S_2_00[21]), .B1(S_2_01[13]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19667), .COUT(n19668), .S0(o_p_29__N_2320[20]), .S1(o_p_29__N_2320[21]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(177[13] 178[15])
    defparam add_35_14.INIT0 = 16'h5666;
    defparam add_35_14.INIT1 = 16'h5666;
    defparam add_35_14.INJECT1_0 = "NO";
    defparam add_35_14.INJECT1_1 = "NO";
    CCU2D add_35_12 (.A0(S_2_00[18]), .B0(S_2_01[10]), .C0(GND_net), .D0(GND_net), 
          .A1(S_2_00[19]), .B1(S_2_01[11]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19666), .COUT(n19667), .S0(o_p_29__N_2320[18]), .S1(o_p_29__N_2320[19]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(177[13] 178[15])
    defparam add_35_12.INIT0 = 16'h5666;
    defparam add_35_12.INIT1 = 16'h5666;
    defparam add_35_12.INJECT1_0 = "NO";
    defparam add_35_12.INJECT1_1 = "NO";
    CCU2D add_35_10 (.A0(S_2_00[16]), .B0(S_2_01[8]), .C0(GND_net), .D0(GND_net), 
          .A1(S_2_00[17]), .B1(S_2_01[9]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19665), .COUT(n19666), .S0(o_p_29__N_2320[16]), .S1(o_p_29__N_2320[17]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(177[13] 178[15])
    defparam add_35_10.INIT0 = 16'h5666;
    defparam add_35_10.INIT1 = 16'h5666;
    defparam add_35_10.INJECT1_0 = "NO";
    defparam add_35_10.INJECT1_1 = "NO";
    CCU2D add_845_16 (.A0(S_0_02[16]), .B0(S_0_03[14]), .C0(GND_net), 
          .D0(GND_net), .A1(S_0_02[17]), .B1(S_0_03[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n19831), .COUT(n19832), .S0(S_1_01_20__N_2205[16]), 
          .S1(S_1_01_20__N_2205[17]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(123[13:48])
    defparam add_845_16.INIT0 = 16'h5666;
    defparam add_845_16.INIT1 = 16'h5666;
    defparam add_845_16.INJECT1_0 = "NO";
    defparam add_845_16.INJECT1_1 = "NO";
    CCU2D add_845_14 (.A0(S_0_02[14]), .B0(S_0_03[12]), .C0(GND_net), 
          .D0(GND_net), .A1(S_0_02[15]), .B1(S_0_03[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n19830), .COUT(n19831), .S0(S_1_01_20__N_2205[14]), 
          .S1(S_1_01_20__N_2205[15]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(123[13:48])
    defparam add_845_14.INIT0 = 16'h5666;
    defparam add_845_14.INIT1 = 16'h5666;
    defparam add_845_14.INJECT1_0 = "NO";
    defparam add_845_14.INJECT1_1 = "NO";
    CCU2D add_35_8 (.A0(S_2_00[14]), .B0(S_2_01[6]), .C0(GND_net), .D0(GND_net), 
          .A1(S_2_00[15]), .B1(S_2_01[7]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19664), .COUT(n19665), .S0(o_p_29__N_2320[14]), .S1(o_p_29__N_2320[15]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(177[13] 178[15])
    defparam add_35_8.INIT0 = 16'h5666;
    defparam add_35_8.INIT1 = 16'h5666;
    defparam add_35_8.INJECT1_0 = "NO";
    defparam add_35_8.INJECT1_1 = "NO";
    CCU2D add_35_6 (.A0(S_2_00[12]), .B0(S_2_01[4]), .C0(GND_net), .D0(GND_net), 
          .A1(S_2_00[13]), .B1(S_2_01[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19663), .COUT(n19664), .S0(o_p_29__N_2320[12]), .S1(o_p_29__N_2320[13]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(177[13] 178[15])
    defparam add_35_6.INIT0 = 16'h5666;
    defparam add_35_6.INIT1 = 16'h5666;
    defparam add_35_6.INJECT1_0 = "NO";
    defparam add_35_6.INJECT1_1 = "NO";
    CCU2D add_845_12 (.A0(S_0_02[12]), .B0(S_0_03[10]), .C0(GND_net), 
          .D0(GND_net), .A1(S_0_02[13]), .B1(S_0_03[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n19829), .COUT(n19830), .S0(S_1_01_20__N_2205[12]), 
          .S1(S_1_01_20__N_2205[13]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(123[13:48])
    defparam add_845_12.INIT0 = 16'h5666;
    defparam add_845_12.INIT1 = 16'h5666;
    defparam add_845_12.INJECT1_0 = "NO";
    defparam add_845_12.INJECT1_1 = "NO";
    CCU2D add_35_4 (.A0(S_2_00[10]), .B0(S_2_01[2]), .C0(GND_net), .D0(GND_net), 
          .A1(S_2_00[11]), .B1(S_2_01[3]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19662), .COUT(n19663), .S0(o_p_29__N_2320[10]), .S1(o_p_29__N_2320[11]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(177[13] 178[15])
    defparam add_35_4.INIT0 = 16'h5666;
    defparam add_35_4.INIT1 = 16'h5666;
    defparam add_35_4.INJECT1_0 = "NO";
    defparam add_35_4.INJECT1_1 = "NO";
    CCU2D add_845_10 (.A0(S_0_02[10]), .B0(S_0_03[8]), .C0(GND_net), .D0(GND_net), 
          .A1(S_0_02[11]), .B1(S_0_03[9]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19828), .COUT(n19829), .S0(S_1_01_20__N_2205[10]), .S1(S_1_01_20__N_2205[11]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(123[13:48])
    defparam add_845_10.INIT0 = 16'h5666;
    defparam add_845_10.INIT1 = 16'h5666;
    defparam add_845_10.INJECT1_0 = "NO";
    defparam add_845_10.INJECT1_1 = "NO";
    CCU2D add_35_2 (.A0(S_2_00[8]), .B0(S_2_01[0]), .C0(GND_net), .D0(GND_net), 
          .A1(S_2_00[9]), .B1(S_2_01[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n19662), .S1(o_p_29__N_2320[9]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(177[13] 178[15])
    defparam add_35_2.INIT0 = 16'h7000;
    defparam add_35_2.INIT1 = 16'h5666;
    defparam add_35_2.INJECT1_0 = "NO";
    defparam add_35_2.INJECT1_1 = "NO";
    CCU2D add_845_8 (.A0(S_0_02[8]), .B0(S_0_03[6]), .C0(GND_net), .D0(GND_net), 
          .A1(S_0_02[9]), .B1(S_0_03[7]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19827), .COUT(n19828), .S0(S_1_01_20__N_2205[8]), .S1(S_1_01_20__N_2205[9]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(123[13:48])
    defparam add_845_8.INIT0 = 16'h5666;
    defparam add_845_8.INIT1 = 16'h5666;
    defparam add_845_8.INJECT1_0 = "NO";
    defparam add_845_8.INJECT1_1 = "NO";
    CCU2D add_845_6 (.A0(S_0_02[6]), .B0(S_0_03[4]), .C0(GND_net), .D0(GND_net), 
          .A1(S_0_02[7]), .B1(S_0_03[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19826), .COUT(n19827), .S0(S_1_01_20__N_2205[6]), .S1(S_1_01_20__N_2205[7]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(123[13:48])
    defparam add_845_6.INIT0 = 16'h5666;
    defparam add_845_6.INIT1 = 16'h5666;
    defparam add_845_6.INJECT1_0 = "NO";
    defparam add_845_6.INJECT1_1 = "NO";
    CCU2D add_845_4 (.A0(S_0_02[4]), .B0(S_0_03[2]), .C0(GND_net), .D0(GND_net), 
          .A1(S_0_02[5]), .B1(S_0_03[3]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19825), .COUT(n19826), .S0(S_1_01_20__N_2205[4]), .S1(S_1_01_20__N_2205[5]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(123[13:48])
    defparam add_845_4.INIT0 = 16'h5666;
    defparam add_845_4.INIT1 = 16'h5666;
    defparam add_845_4.INJECT1_0 = "NO";
    defparam add_845_4.INJECT1_1 = "NO";
    CCU2D add_845_2 (.A0(S_0_02[2]), .B0(S_0_03[0]), .C0(GND_net), .D0(GND_net), 
          .A1(S_0_02[3]), .B1(S_0_03[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n19825), .S1(S_1_01_20__N_2205[3]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(123[13:48])
    defparam add_845_2.INIT0 = 16'h7000;
    defparam add_845_2.INIT1 = 16'h5666;
    defparam add_845_2.INJECT1_0 = "NO";
    defparam add_845_2.INJECT1_1 = "NO";
    CCU2D add_844_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19823), 
          .S0(S_1_02_20__N_2226[20]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(124[13:48])
    defparam add_844_cout.INIT0 = 16'h0000;
    defparam add_844_cout.INIT1 = 16'h0000;
    defparam add_844_cout.INJECT1_0 = "NO";
    defparam add_844_cout.INJECT1_1 = "NO";
    CCU2D add_844_18 (.A0(S_0_05[16]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(S_0_05[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n19822), .COUT(n19823), .S0(S_1_02_20__N_2226[18]), .S1(S_1_02_20__N_2226[19]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(124[13:48])
    defparam add_844_18.INIT0 = 16'hfaaa;
    defparam add_844_18.INIT1 = 16'hfaaa;
    defparam add_844_18.INJECT1_0 = "NO";
    defparam add_844_18.INJECT1_1 = "NO";
    CCU2D add_844_16 (.A0(S_0_04[16]), .B0(S_0_05[14]), .C0(GND_net), 
          .D0(GND_net), .A1(S_0_04[17]), .B1(S_0_05[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n19821), .COUT(n19822), .S0(S_1_02_20__N_2226[16]), 
          .S1(S_1_02_20__N_2226[17]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(124[13:48])
    defparam add_844_16.INIT0 = 16'h5666;
    defparam add_844_16.INIT1 = 16'h5666;
    defparam add_844_16.INJECT1_0 = "NO";
    defparam add_844_16.INJECT1_1 = "NO";
    CCU2D add_844_14 (.A0(S_0_04[14]), .B0(S_0_05[12]), .C0(GND_net), 
          .D0(GND_net), .A1(S_0_04[15]), .B1(S_0_05[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n19820), .COUT(n19821), .S0(S_1_02_20__N_2226[14]), 
          .S1(S_1_02_20__N_2226[15]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(124[13:48])
    defparam add_844_14.INIT0 = 16'h5666;
    defparam add_844_14.INIT1 = 16'h5666;
    defparam add_844_14.INJECT1_0 = "NO";
    defparam add_844_14.INJECT1_1 = "NO";
    CCU2D add_844_12 (.A0(S_0_04[12]), .B0(S_0_05[10]), .C0(GND_net), 
          .D0(GND_net), .A1(S_0_04[13]), .B1(S_0_05[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n19819), .COUT(n19820), .S0(S_1_02_20__N_2226[12]), 
          .S1(S_1_02_20__N_2226[13]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(124[13:48])
    defparam add_844_12.INIT0 = 16'h5666;
    defparam add_844_12.INIT1 = 16'h5666;
    defparam add_844_12.INJECT1_0 = "NO";
    defparam add_844_12.INJECT1_1 = "NO";
    CCU2D add_844_10 (.A0(S_0_04[10]), .B0(S_0_05[8]), .C0(GND_net), .D0(GND_net), 
          .A1(S_0_04[11]), .B1(S_0_05[9]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19818), .COUT(n19819), .S0(S_1_02_20__N_2226[10]), .S1(S_1_02_20__N_2226[11]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(124[13:48])
    defparam add_844_10.INIT0 = 16'h5666;
    defparam add_844_10.INIT1 = 16'h5666;
    defparam add_844_10.INJECT1_0 = "NO";
    defparam add_844_10.INJECT1_1 = "NO";
    CCU2D add_844_8 (.A0(S_0_04[8]), .B0(S_0_05[6]), .C0(GND_net), .D0(GND_net), 
          .A1(S_0_04[9]), .B1(S_0_05[7]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19817), .COUT(n19818), .S0(S_1_02_20__N_2226[8]), .S1(S_1_02_20__N_2226[9]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(124[13:48])
    defparam add_844_8.INIT0 = 16'h5666;
    defparam add_844_8.INIT1 = 16'h5666;
    defparam add_844_8.INJECT1_0 = "NO";
    defparam add_844_8.INJECT1_1 = "NO";
    CCU2D add_844_6 (.A0(S_0_04[6]), .B0(S_0_05[4]), .C0(GND_net), .D0(GND_net), 
          .A1(S_0_04[7]), .B1(S_0_05[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19816), .COUT(n19817), .S0(S_1_02_20__N_2226[6]), .S1(S_1_02_20__N_2226[7]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(124[13:48])
    defparam add_844_6.INIT0 = 16'h5666;
    defparam add_844_6.INIT1 = 16'h5666;
    defparam add_844_6.INJECT1_0 = "NO";
    defparam add_844_6.INJECT1_1 = "NO";
    CCU2D add_844_4 (.A0(S_0_04[4]), .B0(S_0_05[2]), .C0(GND_net), .D0(GND_net), 
          .A1(S_0_04[5]), .B1(S_0_05[3]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19815), .COUT(n19816), .S0(S_1_02_20__N_2226[4]), .S1(S_1_02_20__N_2226[5]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(124[13:48])
    defparam add_844_4.INIT0 = 16'h5666;
    defparam add_844_4.INIT1 = 16'h5666;
    defparam add_844_4.INJECT1_0 = "NO";
    defparam add_844_4.INJECT1_1 = "NO";
    CCU2D add_844_2 (.A0(S_0_04[2]), .B0(S_0_05[0]), .C0(GND_net), .D0(GND_net), 
          .A1(S_0_04[3]), .B1(S_0_05[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n19815), .S1(S_1_02_20__N_2226[3]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(124[13:48])
    defparam add_844_2.INIT0 = 16'h7000;
    defparam add_844_2.INIT1 = 16'h5666;
    defparam add_844_2.INJECT1_0 = "NO";
    defparam add_844_2.INJECT1_1 = "NO";
    CCU2D add_843_22 (.A0(S_1_01[20]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19813), 
          .S0(S_2_00_25__N_2268[24]), .S1(S_2_00_25__N_2268[25]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(152[13:48])
    defparam add_843_22.INIT0 = 16'hfaaa;
    defparam add_843_22.INIT1 = 16'h0000;
    defparam add_843_22.INJECT1_0 = "NO";
    defparam add_843_22.INJECT1_1 = "NO";
    CCU2D add_843_20 (.A0(S_1_01[18]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(S_1_01[19]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n19812), .COUT(n19813), .S0(S_2_00_25__N_2268[22]), .S1(S_2_00_25__N_2268[23]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(152[13:48])
    defparam add_843_20.INIT0 = 16'hfaaa;
    defparam add_843_20.INIT1 = 16'hfaaa;
    defparam add_843_20.INJECT1_0 = "NO";
    defparam add_843_20.INJECT1_1 = "NO";
    CCU2D add_843_18 (.A0(S_1_00[20]), .B0(S_1_01[16]), .C0(GND_net), 
          .D0(GND_net), .A1(S_1_01[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n19811), .COUT(n19812), .S0(S_2_00_25__N_2268[20]), 
          .S1(S_2_00_25__N_2268[21]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(152[13:48])
    defparam add_843_18.INIT0 = 16'h5666;
    defparam add_843_18.INIT1 = 16'hfaaa;
    defparam add_843_18.INJECT1_0 = "NO";
    defparam add_843_18.INJECT1_1 = "NO";
    CCU2D add_843_16 (.A0(S_1_00[18]), .B0(S_1_01[14]), .C0(GND_net), 
          .D0(GND_net), .A1(S_1_00[19]), .B1(S_1_01[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n19810), .COUT(n19811), .S0(S_2_00_25__N_2268[18]), 
          .S1(S_2_00_25__N_2268[19]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(152[13:48])
    defparam add_843_16.INIT0 = 16'h5666;
    defparam add_843_16.INIT1 = 16'h5666;
    defparam add_843_16.INJECT1_0 = "NO";
    defparam add_843_16.INJECT1_1 = "NO";
    CCU2D add_843_14 (.A0(S_1_00[16]), .B0(S_1_01[12]), .C0(GND_net), 
          .D0(GND_net), .A1(S_1_00[17]), .B1(S_1_01[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n19809), .COUT(n19810), .S0(S_2_00_25__N_2268[16]), 
          .S1(S_2_00_25__N_2268[17]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(152[13:48])
    defparam add_843_14.INIT0 = 16'h5666;
    defparam add_843_14.INIT1 = 16'h5666;
    defparam add_843_14.INJECT1_0 = "NO";
    defparam add_843_14.INJECT1_1 = "NO";
    CCU2D add_843_12 (.A0(S_1_00[14]), .B0(S_1_01[10]), .C0(GND_net), 
          .D0(GND_net), .A1(S_1_00[15]), .B1(S_1_01[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n19808), .COUT(n19809), .S0(S_2_00_25__N_2268[14]), 
          .S1(S_2_00_25__N_2268[15]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(152[13:48])
    defparam add_843_12.INIT0 = 16'h5666;
    defparam add_843_12.INIT1 = 16'h5666;
    defparam add_843_12.INJECT1_0 = "NO";
    defparam add_843_12.INJECT1_1 = "NO";
    CCU2D add_843_10 (.A0(S_1_00[12]), .B0(S_1_01[8]), .C0(GND_net), .D0(GND_net), 
          .A1(S_1_00[13]), .B1(S_1_01[9]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19807), .COUT(n19808), .S0(S_2_00_25__N_2268[12]), .S1(S_2_00_25__N_2268[13]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(152[13:48])
    defparam add_843_10.INIT0 = 16'h5666;
    defparam add_843_10.INIT1 = 16'h5666;
    defparam add_843_10.INJECT1_0 = "NO";
    defparam add_843_10.INJECT1_1 = "NO";
    CCU2D add_843_8 (.A0(S_1_00[10]), .B0(S_1_01[6]), .C0(GND_net), .D0(GND_net), 
          .A1(S_1_00[11]), .B1(S_1_01[7]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19806), .COUT(n19807), .S0(S_2_00_25__N_2268[10]), .S1(S_2_00_25__N_2268[11]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(152[13:48])
    defparam add_843_8.INIT0 = 16'h5666;
    defparam add_843_8.INIT1 = 16'h5666;
    defparam add_843_8.INJECT1_0 = "NO";
    defparam add_843_8.INJECT1_1 = "NO";
    CCU2D add_843_6 (.A0(S_1_00[8]), .B0(S_1_01[4]), .C0(GND_net), .D0(GND_net), 
          .A1(S_1_00[9]), .B1(S_1_01[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19805), .COUT(n19806), .S0(S_2_00_25__N_2268[8]), .S1(S_2_00_25__N_2268[9]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(152[13:48])
    defparam add_843_6.INIT0 = 16'h5666;
    defparam add_843_6.INIT1 = 16'h5666;
    defparam add_843_6.INJECT1_0 = "NO";
    defparam add_843_6.INJECT1_1 = "NO";
    CCU2D add_843_4 (.A0(S_1_00[6]), .B0(S_1_01[2]), .C0(GND_net), .D0(GND_net), 
          .A1(S_1_00[7]), .B1(S_1_01[3]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19804), .COUT(n19805), .S0(S_2_00_25__N_2268[6]), .S1(S_2_00_25__N_2268[7]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(152[13:48])
    defparam add_843_4.INIT0 = 16'h5666;
    defparam add_843_4.INIT1 = 16'h5666;
    defparam add_843_4.INJECT1_0 = "NO";
    defparam add_843_4.INJECT1_1 = "NO";
    CCU2D add_843_2 (.A0(S_1_00[4]), .B0(S_1_01[0]), .C0(GND_net), .D0(GND_net), 
          .A1(S_1_00[5]), .B1(S_1_01[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n19804), .S1(S_2_00_25__N_2268[5]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(152[13:48])
    defparam add_843_2.INIT0 = 16'h7000;
    defparam add_843_2.INIT1 = 16'h5666;
    defparam add_843_2.INJECT1_0 = "NO";
    defparam add_843_2.INJECT1_1 = "NO";
    CCU2D add_842_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19763), 
          .S0(S_1_00_20__N_2184[20]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(122[13:48])
    defparam add_842_cout.INIT0 = 16'h0000;
    defparam add_842_cout.INIT1 = 16'h0000;
    defparam add_842_cout.INJECT1_0 = "NO";
    defparam add_842_cout.INJECT1_1 = "NO";
    CCU2D add_842_18 (.A0(S_0_01[16]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(S_0_01[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n19762), .COUT(n19763), .S0(S_1_00_20__N_2184[18]), .S1(S_1_00_20__N_2184[19]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(122[13:48])
    defparam add_842_18.INIT0 = 16'hfaaa;
    defparam add_842_18.INIT1 = 16'hfaaa;
    defparam add_842_18.INJECT1_0 = "NO";
    defparam add_842_18.INJECT1_1 = "NO";
    CCU2D add_842_16 (.A0(S_0_00[16]), .B0(S_0_01[14]), .C0(GND_net), 
          .D0(GND_net), .A1(S_0_00[17]), .B1(S_0_01[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n19761), .COUT(n19762), .S0(S_1_00_20__N_2184[16]), 
          .S1(S_1_00_20__N_2184[17]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(122[13:48])
    defparam add_842_16.INIT0 = 16'h5666;
    defparam add_842_16.INIT1 = 16'h5666;
    defparam add_842_16.INJECT1_0 = "NO";
    defparam add_842_16.INJECT1_1 = "NO";
    CCU2D add_412_18 (.A0(S_1_02[20]), .B0(S_1_03[16]), .C0(GND_net), 
          .D0(GND_net), .A1(S_1_03[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n19607), .S0(S_2_01_25__N_2294[20]), .S1(S_2_01_25__N_2294[21]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(153[13:48])
    defparam add_412_18.INIT0 = 16'h5666;
    defparam add_412_18.INIT1 = 16'hfaaa;
    defparam add_412_18.INJECT1_0 = "NO";
    defparam add_412_18.INJECT1_1 = "NO";
    CCU2D add_412_16 (.A0(S_1_02[18]), .B0(S_1_03[14]), .C0(GND_net), 
          .D0(GND_net), .A1(S_1_02[19]), .B1(S_1_03[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n19606), .COUT(n19607), .S0(S_2_01_25__N_2294[18]), 
          .S1(S_2_01_25__N_2294[19]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(153[13:48])
    defparam add_412_16.INIT0 = 16'h5666;
    defparam add_412_16.INIT1 = 16'h5666;
    defparam add_412_16.INJECT1_0 = "NO";
    defparam add_412_16.INJECT1_1 = "NO";
    CCU2D add_412_14 (.A0(S_1_02[16]), .B0(S_1_03[12]), .C0(GND_net), 
          .D0(GND_net), .A1(S_1_02[17]), .B1(S_1_03[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n19605), .COUT(n19606), .S0(S_2_01_25__N_2294[16]), 
          .S1(S_2_01_25__N_2294[17]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(153[13:48])
    defparam add_412_14.INIT0 = 16'h5666;
    defparam add_412_14.INIT1 = 16'h5666;
    defparam add_412_14.INJECT1_0 = "NO";
    defparam add_412_14.INJECT1_1 = "NO";
    CCU2D add_842_14 (.A0(S_0_00[14]), .B0(S_0_01[12]), .C0(GND_net), 
          .D0(GND_net), .A1(S_0_00[15]), .B1(S_0_01[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n19760), .COUT(n19761), .S0(S_1_00_20__N_2184[14]), 
          .S1(S_1_00_20__N_2184[15]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(122[13:48])
    defparam add_842_14.INIT0 = 16'h5666;
    defparam add_842_14.INIT1 = 16'h5666;
    defparam add_842_14.INJECT1_0 = "NO";
    defparam add_842_14.INJECT1_1 = "NO";
    CCU2D add_842_12 (.A0(S_0_00[12]), .B0(S_0_01[10]), .C0(GND_net), 
          .D0(GND_net), .A1(S_0_00[13]), .B1(S_0_01[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n19759), .COUT(n19760), .S0(S_1_00_20__N_2184[12]), 
          .S1(S_1_00_20__N_2184[13]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(122[13:48])
    defparam add_842_12.INIT0 = 16'h5666;
    defparam add_842_12.INIT1 = 16'h5666;
    defparam add_842_12.INJECT1_0 = "NO";
    defparam add_842_12.INJECT1_1 = "NO";
    CCU2D add_842_10 (.A0(S_0_00[10]), .B0(S_0_01[8]), .C0(GND_net), .D0(GND_net), 
          .A1(S_0_00[11]), .B1(S_0_01[9]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19758), .COUT(n19759), .S0(S_1_00_20__N_2184[10]), .S1(S_1_00_20__N_2184[11]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(122[13:48])
    defparam add_842_10.INIT0 = 16'h5666;
    defparam add_842_10.INIT1 = 16'h5666;
    defparam add_842_10.INJECT1_0 = "NO";
    defparam add_842_10.INJECT1_1 = "NO";
    CCU2D add_842_8 (.A0(S_0_00[8]), .B0(S_0_01[6]), .C0(GND_net), .D0(GND_net), 
          .A1(S_0_00[9]), .B1(S_0_01[7]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19757), .COUT(n19758), .S0(S_1_00_20__N_2184[8]), .S1(S_1_00_20__N_2184[9]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(122[13:48])
    defparam add_842_8.INIT0 = 16'h5666;
    defparam add_842_8.INIT1 = 16'h5666;
    defparam add_842_8.INJECT1_0 = "NO";
    defparam add_842_8.INJECT1_1 = "NO";
    CCU2D add_412_12 (.A0(S_1_02[14]), .B0(S_1_03[10]), .C0(GND_net), 
          .D0(GND_net), .A1(S_1_02[15]), .B1(S_1_03[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n19604), .COUT(n19605), .S0(S_2_01_25__N_2294[14]), 
          .S1(S_2_01_25__N_2294[15]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(153[13:48])
    defparam add_412_12.INIT0 = 16'h5666;
    defparam add_412_12.INIT1 = 16'h5666;
    defparam add_412_12.INJECT1_0 = "NO";
    defparam add_412_12.INJECT1_1 = "NO";
    CCU2D add_842_6 (.A0(S_0_00[6]), .B0(S_0_01[4]), .C0(GND_net), .D0(GND_net), 
          .A1(S_0_00[7]), .B1(S_0_01[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19756), .COUT(n19757), .S0(S_1_00_20__N_2184[6]), .S1(S_1_00_20__N_2184[7]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(122[13:48])
    defparam add_842_6.INIT0 = 16'h5666;
    defparam add_842_6.INIT1 = 16'h5666;
    defparam add_842_6.INJECT1_0 = "NO";
    defparam add_842_6.INJECT1_1 = "NO";
    CCU2D add_412_10 (.A0(S_1_02[12]), .B0(S_1_03[8]), .C0(GND_net), .D0(GND_net), 
          .A1(S_1_02[13]), .B1(S_1_03[9]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19603), .COUT(n19604), .S0(S_2_01_25__N_2294[12]), .S1(S_2_01_25__N_2294[13]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(153[13:48])
    defparam add_412_10.INIT0 = 16'h5666;
    defparam add_412_10.INIT1 = 16'h5666;
    defparam add_412_10.INJECT1_0 = "NO";
    defparam add_412_10.INJECT1_1 = "NO";
    CCU2D add_412_8 (.A0(S_1_02[10]), .B0(S_1_03[6]), .C0(GND_net), .D0(GND_net), 
          .A1(S_1_02[11]), .B1(S_1_03[7]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19602), .COUT(n19603), .S0(S_2_01_25__N_2294[10]), .S1(S_2_01_25__N_2294[11]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(153[13:48])
    defparam add_412_8.INIT0 = 16'h5666;
    defparam add_412_8.INIT1 = 16'h5666;
    defparam add_412_8.INJECT1_0 = "NO";
    defparam add_412_8.INJECT1_1 = "NO";
    CCU2D add_842_4 (.A0(S_0_00[4]), .B0(S_0_01[2]), .C0(GND_net), .D0(GND_net), 
          .A1(S_0_00[5]), .B1(S_0_01[3]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19755), .COUT(n19756), .S0(S_1_00_20__N_2184[4]), .S1(S_1_00_20__N_2184[5]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(122[13:48])
    defparam add_842_4.INIT0 = 16'h5666;
    defparam add_842_4.INIT1 = 16'h5666;
    defparam add_842_4.INJECT1_0 = "NO";
    defparam add_842_4.INJECT1_1 = "NO";
    CCU2D add_412_6 (.A0(S_1_02[8]), .B0(S_1_03[4]), .C0(GND_net), .D0(GND_net), 
          .A1(S_1_02[9]), .B1(S_1_03[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19601), .COUT(n19602), .S0(S_2_01_25__N_2294[8]), .S1(S_2_01_25__N_2294[9]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(153[13:48])
    defparam add_412_6.INIT0 = 16'h5666;
    defparam add_412_6.INIT1 = 16'h5666;
    defparam add_412_6.INJECT1_0 = "NO";
    defparam add_412_6.INJECT1_1 = "NO";
    CCU2D add_842_2 (.A0(S_0_00[2]), .B0(S_0_01[0]), .C0(GND_net), .D0(GND_net), 
          .A1(S_0_00[3]), .B1(S_0_01[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n19755), .S1(S_1_00_20__N_2184[3]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(122[13:48])
    defparam add_842_2.INIT0 = 16'h7000;
    defparam add_842_2.INIT1 = 16'h5666;
    defparam add_842_2.INJECT1_0 = "NO";
    defparam add_842_2.INJECT1_1 = "NO";
    CCU2D add_412_4 (.A0(S_1_02[6]), .B0(S_1_03[2]), .C0(GND_net), .D0(GND_net), 
          .A1(S_1_02[7]), .B1(S_1_03[3]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19600), .COUT(n19601), .S0(S_2_01_25__N_2294[6]), .S1(S_2_01_25__N_2294[7]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(153[13:48])
    defparam add_412_4.INIT0 = 16'h5666;
    defparam add_412_4.INIT1 = 16'h5666;
    defparam add_412_4.INJECT1_0 = "NO";
    defparam add_412_4.INJECT1_1 = "NO";
    CCU2D add_412_2 (.A0(S_1_02[4]), .B0(S_1_03[0]), .C0(GND_net), .D0(GND_net), 
          .A1(S_1_02[5]), .B1(S_1_03[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n19600), .S1(S_2_01_25__N_2294[5]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(153[13:48])
    defparam add_412_2.INIT0 = 16'h7000;
    defparam add_412_2.INIT1 = 16'h5666;
    defparam add_412_2.INJECT1_0 = "NO";
    defparam add_412_2.INJECT1_1 = "NO";
    LUT4 i17610_2_lut (.A(S_2_00[8]), .B(S_2_01[0]), .Z(o_p_29__N_2320[8])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i17610_2_lut.init = 16'h6666;
    LUT4 i17607_2_lut (.A(S_1_02[4]), .B(S_1_03[0]), .Z(S_2_01_25__N_2294[4])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i17607_2_lut.init = 16'h6666;
    LUT4 i17613_2_lut (.A(S_1_00[4]), .B(S_1_01[0]), .Z(S_2_00_25__N_2268[4])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i17613_2_lut.init = 16'h6666;
    LUT4 i17614_2_lut (.A(S_0_04[2]), .B(S_0_05[0]), .Z(S_1_02_20__N_2226[2])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i17614_2_lut.init = 16'h6666;
    LUT4 i17615_2_lut (.A(S_0_02[2]), .B(S_0_03[0]), .Z(S_1_01_20__N_2205[2])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i17615_2_lut.init = 16'h6666;
    LUT4 i17612_2_lut (.A(S_0_00[2]), .B(S_0_01[0]), .Z(S_1_00_20__N_2184[2])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i17612_2_lut.init = 16'h6666;
    FD1S3IX S_3_00__i29 (.D(o_p_29__N_2320[29]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i29.GSR = "DISABLED";
    FD1S3IX S_3_00__i28 (.D(o_p_29__N_2320[28]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i28.GSR = "DISABLED";
    FD1S3IX S_3_00__i27 (.D(o_p_29__N_2320[27]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i27.GSR = "DISABLED";
    FD1S3IX S_3_00__i26 (.D(o_p_29__N_2320[26]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i26.GSR = "DISABLED";
    FD1S3IX S_3_00__i25 (.D(o_p_29__N_2320[25]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i25.GSR = "DISABLED";
    FD1S3IX S_3_00__i24 (.D(o_p_29__N_2320[24]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i24.GSR = "DISABLED";
    FD1S3IX S_3_00__i23 (.D(o_p_29__N_2320[23]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i23.GSR = "DISABLED";
    FD1S3IX S_3_00__i22 (.D(o_p_29__N_2320[22]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i22.GSR = "DISABLED";
    FD1S3IX S_3_00__i21 (.D(o_p_29__N_2320[21]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i21.GSR = "DISABLED";
    FD1S3IX S_3_00__i20 (.D(o_p_29__N_2320[20]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i20.GSR = "DISABLED";
    FD1S3IX S_3_00__i19 (.D(o_p_29__N_2320[19]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i19.GSR = "DISABLED";
    FD1S3IX S_3_00__i18 (.D(o_p_29__N_2320[18]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i18.GSR = "DISABLED";
    FD1S3IX S_3_00__i17 (.D(o_p_29__N_2320[17]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i17.GSR = "DISABLED";
    FD1S3IX S_3_00__i16 (.D(o_p_29__N_2320[16]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i16.GSR = "DISABLED";
    FD1S3IX S_3_00__i15 (.D(o_p_29__N_2320[15]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i15.GSR = "DISABLED";
    FD1S3IX S_3_00__i14 (.D(o_p_29__N_2320[14]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i14.GSR = "DISABLED";
    FD1S3IX S_3_00__i13 (.D(o_p_29__N_2320[13]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i13.GSR = "DISABLED";
    FD1S3IX S_3_00__i12 (.D(o_p_29__N_2320[12]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i12.GSR = "DISABLED";
    FD1S3IX S_3_00__i11 (.D(o_p_29__N_2320[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i11.GSR = "DISABLED";
    FD1S3IX S_3_00__i10 (.D(o_p_29__N_2320[10]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i10.GSR = "DISABLED";
    FD1S3IX S_3_00__i9 (.D(o_p_29__N_2320[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i9.GSR = "DISABLED";
    FD1S3IX S_3_00__i8 (.D(o_p_29__N_2320[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i8.GSR = "DISABLED";
    FD1S3IX S_3_00__i7 (.D(o_p_29__N_2320[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i7.GSR = "DISABLED";
    FD1S3IX S_3_00__i6 (.D(o_p_29__N_2320[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i6.GSR = "DISABLED";
    FD1S3IX S_3_00__i5 (.D(o_p_29__N_2320[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i5.GSR = "DISABLED";
    FD1S3IX S_3_00__i4 (.D(o_p_29__N_2320[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i4.GSR = "DISABLED";
    FD1S3IX S_3_00__i3 (.D(o_p_29__N_2320[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i3.GSR = "DISABLED";
    FD1S3IX S_3_00__i2 (.D(o_p_29__N_2320[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i2.GSR = "DISABLED";
    FD1S3IX S_3_00__i1 (.D(o_p_29__N_2320[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i1.GSR = "DISABLED";
    FD1S3IX S_2_01__i22 (.D(S_2_01_25__N_2294[21]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i22.GSR = "DISABLED";
    FD1S3IX S_2_01__i21 (.D(S_2_01_25__N_2294[20]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i21.GSR = "DISABLED";
    FD1S3IX S_2_01__i20 (.D(S_2_01_25__N_2294[19]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i20.GSR = "DISABLED";
    FD1S3IX S_2_01__i19 (.D(S_2_01_25__N_2294[18]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i19.GSR = "DISABLED";
    FD1S3IX S_2_01__i18 (.D(S_2_01_25__N_2294[17]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i18.GSR = "DISABLED";
    FD1S3IX S_2_01__i17 (.D(S_2_01_25__N_2294[16]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i17.GSR = "DISABLED";
    FD1S3IX S_2_01__i16 (.D(S_2_01_25__N_2294[15]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i16.GSR = "DISABLED";
    FD1S3IX S_2_01__i15 (.D(S_2_01_25__N_2294[14]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i15.GSR = "DISABLED";
    FD1S3IX S_2_01__i14 (.D(S_2_01_25__N_2294[13]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i14.GSR = "DISABLED";
    FD1S3IX S_2_01__i13 (.D(S_2_01_25__N_2294[12]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i13.GSR = "DISABLED";
    FD1S3IX S_2_01__i12 (.D(S_2_01_25__N_2294[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i12.GSR = "DISABLED";
    FD1S3IX S_2_01__i11 (.D(S_2_01_25__N_2294[10]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i11.GSR = "DISABLED";
    FD1S3IX S_2_01__i10 (.D(S_2_01_25__N_2294[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i10.GSR = "DISABLED";
    FD1S3IX S_2_01__i9 (.D(S_2_01_25__N_2294[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i9.GSR = "DISABLED";
    FD1S3IX S_2_01__i8 (.D(S_2_01_25__N_2294[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i8.GSR = "DISABLED";
    FD1S3IX S_2_01__i7 (.D(S_2_01_25__N_2294[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i7.GSR = "DISABLED";
    FD1S3IX S_2_01__i6 (.D(S_2_01_25__N_2294[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i6.GSR = "DISABLED";
    FD1S3IX S_2_01__i5 (.D(S_2_01_25__N_2294[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i5.GSR = "DISABLED";
    FD1S3IX S_2_01__i4 (.D(S_2_01_25__N_2294[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i4.GSR = "DISABLED";
    FD1S3IX S_2_01__i3 (.D(S_2_01_25__N_2294[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i3.GSR = "DISABLED";
    FD1S3IX S_2_01__i2 (.D(S_2_01_25__N_2294[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i2.GSR = "DISABLED";
    FD1S3IX S_2_00__i26 (.D(S_2_00_25__N_2268[25]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i26.GSR = "DISABLED";
    FD1S3IX S_2_00__i25 (.D(S_2_00_25__N_2268[24]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i25.GSR = "DISABLED";
    FD1S3IX S_2_00__i24 (.D(S_2_00_25__N_2268[23]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i24.GSR = "DISABLED";
    FD1S3IX S_2_00__i23 (.D(S_2_00_25__N_2268[22]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i23.GSR = "DISABLED";
    FD1S3IX S_2_00__i22 (.D(S_2_00_25__N_2268[21]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i22.GSR = "DISABLED";
    FD1S3IX S_2_00__i21 (.D(S_2_00_25__N_2268[20]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i21.GSR = "DISABLED";
    FD1S3IX S_2_00__i20 (.D(S_2_00_25__N_2268[19]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i20.GSR = "DISABLED";
    FD1S3IX S_2_00__i19 (.D(S_2_00_25__N_2268[18]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i19.GSR = "DISABLED";
    FD1S3IX S_2_00__i18 (.D(S_2_00_25__N_2268[17]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i18.GSR = "DISABLED";
    FD1S3IX S_2_00__i17 (.D(S_2_00_25__N_2268[16]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i17.GSR = "DISABLED";
    FD1S3IX S_2_00__i16 (.D(S_2_00_25__N_2268[15]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i16.GSR = "DISABLED";
    FD1S3IX S_2_00__i15 (.D(S_2_00_25__N_2268[14]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i15.GSR = "DISABLED";
    FD1S3IX S_2_00__i14 (.D(S_2_00_25__N_2268[13]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i14.GSR = "DISABLED";
    FD1S3IX S_2_00__i13 (.D(S_2_00_25__N_2268[12]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i13.GSR = "DISABLED";
    FD1S3IX S_2_00__i12 (.D(S_2_00_25__N_2268[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i12.GSR = "DISABLED";
    FD1S3IX S_2_00__i11 (.D(S_2_00_25__N_2268[10]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i11.GSR = "DISABLED";
    FD1S3IX S_2_00__i10 (.D(S_2_00_25__N_2268[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i10.GSR = "DISABLED";
    FD1S3IX S_2_00__i9 (.D(S_2_00_25__N_2268[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i9.GSR = "DISABLED";
    FD1S3IX S_2_00__i8 (.D(S_2_00_25__N_2268[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_p_29__N_2320[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i8.GSR = "DISABLED";
    FD1S3IX S_2_00__i7 (.D(S_2_00_25__N_2268[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_p_29__N_2320[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i7.GSR = "DISABLED";
    FD1S3IX S_2_00__i6 (.D(S_2_00_25__N_2268[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_p_29__N_2320[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i6.GSR = "DISABLED";
    FD1S3IX S_2_00__i5 (.D(S_2_00_25__N_2268[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_p_29__N_2320[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i5.GSR = "DISABLED";
    FD1S3IX S_2_00__i4 (.D(S_2_00_25__N_2268[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_p_29__N_2320[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i4.GSR = "DISABLED";
    FD1S3IX S_2_00__i3 (.D(S_2_00_25__N_2268[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_p_29__N_2320[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i3.GSR = "DISABLED";
    FD1S3IX S_2_00__i2 (.D(S_2_00_25__N_2268[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_p_29__N_2320[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i2.GSR = "DISABLED";
    FD1S3IX S_1_03__i18 (.D(S_0_06[17]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_03[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_03__i18.GSR = "DISABLED";
    FD1S3IX S_1_03__i17 (.D(S_0_06[16]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_03[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_03__i17.GSR = "DISABLED";
    FD1S3IX S_1_03__i16 (.D(S_0_06[15]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_03[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_03__i16.GSR = "DISABLED";
    FD1S3IX S_1_03__i15 (.D(S_0_06[14]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_03[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_03__i15.GSR = "DISABLED";
    FD1S3IX S_1_03__i14 (.D(S_0_06[13]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_03[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_03__i14.GSR = "DISABLED";
    FD1S3IX S_1_03__i13 (.D(S_0_06[12]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_03[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_03__i13.GSR = "DISABLED";
    FD1S3IX S_1_03__i12 (.D(S_0_06[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_03[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_03__i12.GSR = "DISABLED";
    FD1S3IX S_1_03__i11 (.D(S_0_06[10]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_03[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_03__i11.GSR = "DISABLED";
    FD1S3IX S_1_03__i10 (.D(S_0_06[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_03[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_03__i10.GSR = "DISABLED";
    FD1S3IX S_1_03__i9 (.D(S_0_06[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_03[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_03__i9.GSR = "DISABLED";
    FD1S3IX S_1_03__i8 (.D(S_0_06[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_03[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_03__i8.GSR = "DISABLED";
    FD1S3IX S_1_03__i7 (.D(S_0_06[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_03[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_03__i7.GSR = "DISABLED";
    FD1S3IX S_1_03__i6 (.D(S_0_06[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_03[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_03__i6.GSR = "DISABLED";
    FD1S3IX S_1_03__i5 (.D(S_0_06[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_03[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_03__i5.GSR = "DISABLED";
    FD1S3IX S_1_03__i4 (.D(S_0_06[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_03[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_03__i4.GSR = "DISABLED";
    FD1S3IX S_1_03__i3 (.D(S_0_06[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_03[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_03__i3.GSR = "DISABLED";
    FD1S3IX S_1_03__i2 (.D(S_0_06[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_03[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_03__i2.GSR = "DISABLED";
    FD1S3IX S_1_02__i21 (.D(S_1_02_20__N_2226[20]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_02[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i21.GSR = "DISABLED";
    FD1S3IX S_1_02__i20 (.D(S_1_02_20__N_2226[19]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_02[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i20.GSR = "DISABLED";
    FD1S3IX S_1_02__i19 (.D(S_1_02_20__N_2226[18]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_02[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i19.GSR = "DISABLED";
    FD1S3IX S_1_02__i18 (.D(S_1_02_20__N_2226[17]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_02[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i18.GSR = "DISABLED";
    FD1S3IX S_1_02__i17 (.D(S_1_02_20__N_2226[16]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_02[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i17.GSR = "DISABLED";
    FD1S3IX S_1_02__i16 (.D(S_1_02_20__N_2226[15]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_02[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i16.GSR = "DISABLED";
    FD1S3IX S_1_02__i15 (.D(S_1_02_20__N_2226[14]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_02[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i15.GSR = "DISABLED";
    FD1S3IX S_1_02__i14 (.D(S_1_02_20__N_2226[13]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_02[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i14.GSR = "DISABLED";
    FD1S3IX S_1_02__i13 (.D(S_1_02_20__N_2226[12]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_02[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i13.GSR = "DISABLED";
    FD1S3IX S_1_02__i12 (.D(S_1_02_20__N_2226[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_02[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i12.GSR = "DISABLED";
    FD1S3IX S_1_02__i11 (.D(S_1_02_20__N_2226[10]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_02[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i11.GSR = "DISABLED";
    FD1S3IX S_1_02__i10 (.D(S_1_02_20__N_2226[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_02[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i10.GSR = "DISABLED";
    FD1S3IX S_1_02__i9 (.D(S_1_02_20__N_2226[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_02[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i9.GSR = "DISABLED";
    FD1S3IX S_1_02__i8 (.D(S_1_02_20__N_2226[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_02[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i8.GSR = "DISABLED";
    FD1S3IX S_1_02__i7 (.D(S_1_02_20__N_2226[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_02[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i7.GSR = "DISABLED";
    FD1S3IX S_1_02__i6 (.D(S_1_02_20__N_2226[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_02[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i6.GSR = "DISABLED";
    FD1S3IX S_1_02__i5 (.D(S_1_02_20__N_2226[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_02[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i5.GSR = "DISABLED";
    FD1S3IX S_1_02__i4 (.D(S_1_02_20__N_2226[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01_25__N_2294[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i4.GSR = "DISABLED";
    FD1S3IX S_1_02__i3 (.D(S_1_02_20__N_2226[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01_25__N_2294[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i3.GSR = "DISABLED";
    FD1S3IX S_1_02__i2 (.D(S_1_02_20__N_2226[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01_25__N_2294[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i2.GSR = "DISABLED";
    FD1S3IX S_1_01__i20 (.D(S_1_01_20__N_2205[20]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i20.GSR = "DISABLED";
    FD1S3IX S_1_01__i19 (.D(S_1_01_20__N_2205[19]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i19.GSR = "DISABLED";
    FD1S3IX S_1_01__i18 (.D(S_1_01_20__N_2205[18]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i18.GSR = "DISABLED";
    FD1S3IX S_1_01__i17 (.D(S_1_01_20__N_2205[17]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i17.GSR = "DISABLED";
    FD1S3IX S_1_01__i16 (.D(S_1_01_20__N_2205[16]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i16.GSR = "DISABLED";
    FD1S3IX S_1_01__i15 (.D(S_1_01_20__N_2205[15]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i15.GSR = "DISABLED";
    FD1S3IX S_1_01__i14 (.D(S_1_01_20__N_2205[14]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i14.GSR = "DISABLED";
    FD1S3IX S_1_01__i13 (.D(S_1_01_20__N_2205[13]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i13.GSR = "DISABLED";
    FD1S3IX S_1_01__i12 (.D(S_1_01_20__N_2205[12]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i12.GSR = "DISABLED";
    FD1S3IX S_1_01__i11 (.D(S_1_01_20__N_2205[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i11.GSR = "DISABLED";
    FD1S3IX S_1_01__i10 (.D(S_1_01_20__N_2205[10]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i10.GSR = "DISABLED";
    FD1S3IX S_1_01__i9 (.D(S_1_01_20__N_2205[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i9.GSR = "DISABLED";
    FD1S3IX S_1_01__i8 (.D(S_1_01_20__N_2205[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i8.GSR = "DISABLED";
    FD1S3IX S_1_01__i7 (.D(S_1_01_20__N_2205[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i7.GSR = "DISABLED";
    FD1S3IX S_1_01__i6 (.D(S_1_01_20__N_2205[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i6.GSR = "DISABLED";
    FD1S3IX S_1_01__i5 (.D(S_1_01_20__N_2205[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i5.GSR = "DISABLED";
    FD1S3IX S_1_01__i4 (.D(S_1_01_20__N_2205[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i4.GSR = "DISABLED";
    FD1S3IX S_1_01__i3 (.D(S_1_01_20__N_2205[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i3.GSR = "DISABLED";
    FD1S3IX S_1_01__i2 (.D(S_1_01_20__N_2205[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i2.GSR = "DISABLED";
    FD1S3IX S_1_01__i1 (.D(S_1_01_20__N_2205[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i1.GSR = "DISABLED";
    FD1S3IX S_1_00__i20 (.D(S_1_00_20__N_2184[20]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_00[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i20.GSR = "DISABLED";
    FD1S3IX S_1_00__i19 (.D(S_1_00_20__N_2184[19]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_00[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i19.GSR = "DISABLED";
    FD1S3IX S_1_00__i18 (.D(S_1_00_20__N_2184[18]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_00[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i18.GSR = "DISABLED";
    FD1S3IX S_1_00__i17 (.D(S_1_00_20__N_2184[17]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_00[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i17.GSR = "DISABLED";
    FD1S3IX S_1_00__i16 (.D(S_1_00_20__N_2184[16]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_00[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i16.GSR = "DISABLED";
    FD1S3IX S_1_00__i15 (.D(S_1_00_20__N_2184[15]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_00[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i15.GSR = "DISABLED";
    FD1S3IX S_1_00__i14 (.D(S_1_00_20__N_2184[14]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_00[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i14.GSR = "DISABLED";
    FD1S3IX S_1_00__i13 (.D(S_1_00_20__N_2184[13]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_00[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i13.GSR = "DISABLED";
    FD1S3IX S_1_00__i12 (.D(S_1_00_20__N_2184[12]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_00[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i12.GSR = "DISABLED";
    FD1S3IX S_1_00__i11 (.D(S_1_00_20__N_2184[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_00[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i11.GSR = "DISABLED";
    FD1S3IX S_1_00__i10 (.D(S_1_00_20__N_2184[10]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_00[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i10.GSR = "DISABLED";
    FD1S3IX S_1_00__i9 (.D(S_1_00_20__N_2184[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_00[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i9.GSR = "DISABLED";
    FD1S3IX S_1_00__i8 (.D(S_1_00_20__N_2184[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_00[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i8.GSR = "DISABLED";
    FD1S3IX S_1_00__i7 (.D(S_1_00_20__N_2184[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_00[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i7.GSR = "DISABLED";
    FD1S3IX S_1_00__i6 (.D(S_1_00_20__N_2184[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_00[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i6.GSR = "DISABLED";
    FD1S3IX S_1_00__i5 (.D(S_1_00_20__N_2184[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_00[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i5.GSR = "DISABLED";
    FD1S3IX S_1_00__i4 (.D(S_1_00_20__N_2184[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_00[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i4.GSR = "DISABLED";
    FD1S3IX S_1_00__i3 (.D(S_1_00_20__N_2184[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00_25__N_2268[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i3.GSR = "DISABLED";
    FD1S3IX S_1_00__i2 (.D(S_1_00_20__N_2184[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00_25__N_2268[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i2.GSR = "DISABLED";
    FD1S3IX S_1_00__i1 (.D(S_1_00_20__N_2184[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00_25__N_2268[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i1.GSR = "DISABLED";
    \bimpy(BW=16)_U6  initialmpy_6_0 (.u_l({u_l}), .\u_s[13] (u_s[13]), 
            .S_0_06({S_0_06}), .dac_clk_p_c(dac_clk_p_c), .n14231(n14231), 
            .n9444(n9444), .\u_s[12] (u_s[12]), .GND_net(GND_net), .i_sw0_c(i_sw0_c)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(90[14:75])
    \bimpy(BW=16)_U7  initialmpy_5_0 (.S_0_05({S_0_05}), .dac_clk_p_c(dac_clk_p_c), 
            .n14231(n14231), .n9446(n9446), .GND_net(GND_net), .u_l({u_l}), 
            .\u_s[11] (u_s[11]), .\u_s[10] (u_s[10]), .i_sw0_c(i_sw0_c)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(87[14:75])
    \bimpy(BW=16)_U8  initialmpy_4_0 (.\S_0_04[0] (S_0_04[0]), .dac_clk_p_c(dac_clk_p_c), 
            .n14231(n14231), .n9448(n9448), .GND_net(GND_net), .u_l({u_l}), 
            .\u_s[9] (u_s[9]), .\u_s[8] (u_s[8]), .\S_0_04[17] (S_0_04[17]), 
            .i_sw0_c(i_sw0_c), .\S_0_04[16] (S_0_04[16]), .\S_0_04[15] (S_0_04[15]), 
            .\S_0_04[14] (S_0_04[14]), .\S_0_04[13] (S_0_04[13]), .\S_0_04[12] (S_0_04[12]), 
            .\S_0_04[11] (S_0_04[11]), .\S_0_04[10] (S_0_04[10]), .\S_0_04[9] (S_0_04[9]), 
            .\S_0_04[8] (S_0_04[8]), .\S_0_04[7] (S_0_04[7]), .\S_0_04[6] (S_0_04[6]), 
            .\S_0_04[5] (S_0_04[5]), .\S_0_04[4] (S_0_04[4]), .\S_0_04[3] (S_0_04[3]), 
            .\S_0_04[2] (S_0_04[2]), .\S_1_02_20__N_2226[1] (S_1_02_20__N_2226[1])) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(84[14:73])
    \bimpy(BW=16)_U9  initialmpy_3_0 (.GND_net(GND_net), .u_l({u_l}), .\u_s[7] (u_s[7]), 
            .S_0_03({S_0_03}), .dac_clk_p_c(dac_clk_p_c), .n14231(n14231), 
            .n9450(n9450), .\u_s[6] (u_s[6]), .i_sw0_c(i_sw0_c)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(81[14:73])
    \bimpy(BW=16)_U10  initialmpy_2_0 (.GND_net(GND_net), .\S_0_02[0] (S_0_02[0]), 
            .dac_clk_p_c(dac_clk_p_c), .n14231(n14231), .n9452(n9452), 
            .u_l({u_l}), .\u_s[5] (u_s[5]), .\u_s[4] (u_s[4]), .\S_0_02[17] (S_0_02[17]), 
            .i_sw0_c(i_sw0_c), .\S_0_02[16] (S_0_02[16]), .\S_0_02[15] (S_0_02[15]), 
            .\S_0_02[14] (S_0_02[14]), .\S_0_02[13] (S_0_02[13]), .\S_0_02[12] (S_0_02[12]), 
            .\S_0_02[11] (S_0_02[11]), .\S_0_02[10] (S_0_02[10]), .\S_0_02[9] (S_0_02[9]), 
            .\S_0_02[8] (S_0_02[8]), .\S_0_02[7] (S_0_02[7]), .\S_0_02[6] (S_0_02[6]), 
            .\S_0_02[5] (S_0_02[5]), .\S_0_02[4] (S_0_02[4]), .\S_0_02[3] (S_0_02[3]), 
            .\S_0_02[2] (S_0_02[2]), .\S_1_01_20__N_2205[1] (S_1_01_20__N_2205[1])) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(78[14:73])
    \bimpy(BW=16)_U11  initialmpy_1_0 (.S_0_01({S_0_01}), .dac_clk_p_c(dac_clk_p_c), 
            .n14231(n14231), .n9454(n9454), .u_l({u_l}), .\u_s[3] (u_s[3]), 
            .\u_s[2] (u_s[2]), .GND_net(GND_net), .i_sw0_c(i_sw0_c)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(75[14:73])
    \bimpy(BW=16)_U12  initialmpy_0_0 (.\S_0_00[0] (S_0_00[0]), .dac_clk_p_c(dac_clk_p_c), 
            .n14231(n14231), .n9456(n9456), .u_l({u_l}), .\u_s[1] (u_s[1]), 
            .\u_s[0] (u_s[0]), .GND_net(GND_net), .\S_0_00[17] (S_0_00[17]), 
            .i_sw0_c(i_sw0_c), .\S_0_00[16] (S_0_00[16]), .\S_0_00[15] (S_0_00[15]), 
            .\S_0_00[14] (S_0_00[14]), .\S_0_00[13] (S_0_00[13]), .\S_0_00[12] (S_0_00[12]), 
            .\S_0_00[11] (S_0_00[11]), .\S_0_00[10] (S_0_00[10]), .\S_0_00[9] (S_0_00[9]), 
            .\S_0_00[8] (S_0_00[8]), .\S_0_00[7] (S_0_00[7]), .\S_0_00[6] (S_0_00[6]), 
            .\S_0_00[5] (S_0_00[5]), .\S_0_00[4] (S_0_00[4]), .\S_0_00[3] (S_0_00[3]), 
            .\S_0_00[2] (S_0_00[2]), .\S_1_00_20__N_2184[1] (S_1_00_20__N_2184[1])) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(72[14:73])
    
endmodule
//
// Verilog Description of module \bimpy(BW=16)_U6 
//

module \bimpy(BW=16)_U6  (u_l, \u_s[13] , S_0_06, dac_clk_p_c, n14231, 
            n9444, \u_s[12] , GND_net, i_sw0_c) /* synthesis syn_module_defined=1 */ ;
    input [15:0]u_l;
    input \u_s[13] ;
    output [17:0]S_0_06;
    input dac_clk_p_c;
    input n14231;
    input n9444;
    input \u_s[12] ;
    input GND_net;
    input i_sw0_c;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[29:38])
    
    wire n29267;
    wire [17:0]o_r_17__N_2438;
    
    wire n19416, n19415;
    wire [14:0]c_15__N_2408;
    wire [14:0]c_15__N_2423;
    
    wire n19414, n19413, n19412, n19411, n19410, n19409, n29266;
    
    LUT4 i12516_2_lut_rep_607 (.A(u_l[0]), .B(\u_s[13] ), .Z(n29267)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(51[18:45])
    defparam i12516_2_lut_rep_607.init = 16'h8888;
    FD1S3IX o_r__i0 (.D(n9444), .CK(dac_clk_p_c), .CD(n14231), .Q(S_0_06[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=90, LSE_RLINE=90 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i0.GSR = "DISABLED";
    LUT4 w_r_16__I_0_i2_2_lut_3_lut_4_lut (.A(u_l[0]), .B(\u_s[13] ), .C(\u_s[12] ), 
         .D(u_l[1]), .Z(o_r_17__N_2438[1])) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(51[18:45])
    defparam w_r_16__I_0_i2_2_lut_3_lut_4_lut.init = 16'h7888;
    CCU2D add_819_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19416), 
          .S0(o_r_17__N_2438[17]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_819_cout.INIT0 = 16'h0000;
    defparam add_819_cout.INIT1 = 16'h0000;
    defparam add_819_cout.INJECT1_0 = "NO";
    defparam add_819_cout.INJECT1_1 = "NO";
    CCU2D add_819_15 (.A0(c_15__N_2408[14]), .B0(c_15__N_2423[14]), .C0(c_15__N_2408[13]), 
          .D0(c_15__N_2423[13]), .A1(u_l[15]), .B1(\u_s[13] ), .C1(c_15__N_2408[14]), 
          .D1(c_15__N_2423[14]), .CIN(n19415), .COUT(n19416), .S0(o_r_17__N_2438[15]), 
          .S1(o_r_17__N_2438[16]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_819_15.INIT0 = 16'h9666;
    defparam add_819_15.INIT1 = 16'h7888;
    defparam add_819_15.INJECT1_0 = "NO";
    defparam add_819_15.INJECT1_1 = "NO";
    CCU2D add_819_13 (.A0(c_15__N_2408[12]), .B0(c_15__N_2423[12]), .C0(c_15__N_2408[11]), 
          .D0(c_15__N_2423[11]), .A1(c_15__N_2408[13]), .B1(c_15__N_2423[13]), 
          .C1(c_15__N_2408[12]), .D1(c_15__N_2423[12]), .CIN(n19414), 
          .COUT(n19415), .S0(o_r_17__N_2438[13]), .S1(o_r_17__N_2438[14]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_819_13.INIT0 = 16'h9666;
    defparam add_819_13.INIT1 = 16'h9666;
    defparam add_819_13.INJECT1_0 = "NO";
    defparam add_819_13.INJECT1_1 = "NO";
    CCU2D add_819_11 (.A0(c_15__N_2408[10]), .B0(c_15__N_2423[10]), .C0(c_15__N_2408[9]), 
          .D0(c_15__N_2423[9]), .A1(c_15__N_2408[11]), .B1(c_15__N_2423[11]), 
          .C1(c_15__N_2408[10]), .D1(c_15__N_2423[10]), .CIN(n19413), 
          .COUT(n19414), .S0(o_r_17__N_2438[11]), .S1(o_r_17__N_2438[12]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_819_11.INIT0 = 16'h9666;
    defparam add_819_11.INIT1 = 16'h9666;
    defparam add_819_11.INJECT1_0 = "NO";
    defparam add_819_11.INJECT1_1 = "NO";
    CCU2D add_819_9 (.A0(c_15__N_2408[8]), .B0(c_15__N_2423[8]), .C0(c_15__N_2408[7]), 
          .D0(c_15__N_2423[7]), .A1(c_15__N_2408[9]), .B1(c_15__N_2423[9]), 
          .C1(c_15__N_2408[8]), .D1(c_15__N_2423[8]), .CIN(n19412), .COUT(n19413), 
          .S0(o_r_17__N_2438[9]), .S1(o_r_17__N_2438[10]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_819_9.INIT0 = 16'h9666;
    defparam add_819_9.INIT1 = 16'h9666;
    defparam add_819_9.INJECT1_0 = "NO";
    defparam add_819_9.INJECT1_1 = "NO";
    CCU2D add_819_7 (.A0(c_15__N_2408[6]), .B0(c_15__N_2423[6]), .C0(c_15__N_2408[5]), 
          .D0(c_15__N_2423[5]), .A1(c_15__N_2408[7]), .B1(c_15__N_2423[7]), 
          .C1(c_15__N_2408[6]), .D1(c_15__N_2423[6]), .CIN(n19411), .COUT(n19412), 
          .S0(o_r_17__N_2438[7]), .S1(o_r_17__N_2438[8]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_819_7.INIT0 = 16'h9666;
    defparam add_819_7.INIT1 = 16'h9666;
    defparam add_819_7.INJECT1_0 = "NO";
    defparam add_819_7.INJECT1_1 = "NO";
    CCU2D add_819_5 (.A0(c_15__N_2408[4]), .B0(c_15__N_2423[4]), .C0(c_15__N_2408[3]), 
          .D0(c_15__N_2423[3]), .A1(c_15__N_2408[5]), .B1(c_15__N_2423[5]), 
          .C1(c_15__N_2408[4]), .D1(c_15__N_2423[4]), .CIN(n19410), .COUT(n19411), 
          .S0(o_r_17__N_2438[5]), .S1(o_r_17__N_2438[6]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_819_5.INIT0 = 16'h9666;
    defparam add_819_5.INIT1 = 16'h9666;
    defparam add_819_5.INJECT1_0 = "NO";
    defparam add_819_5.INJECT1_1 = "NO";
    CCU2D add_819_3 (.A0(c_15__N_2408[2]), .B0(c_15__N_2423[2]), .C0(c_15__N_2408[1]), 
          .D0(c_15__N_2423[1]), .A1(c_15__N_2408[3]), .B1(c_15__N_2423[3]), 
          .C1(c_15__N_2408[2]), .D1(c_15__N_2423[2]), .CIN(n19409), .COUT(n19410), 
          .S0(o_r_17__N_2438[3]), .S1(o_r_17__N_2438[4]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_819_3.INIT0 = 16'h9666;
    defparam add_819_3.INIT1 = 16'h9666;
    defparam add_819_3.INJECT1_0 = "NO";
    defparam add_819_3.INJECT1_1 = "NO";
    LUT4 i13163_2_lut (.A(u_l[14]), .B(\u_s[13] ), .Z(c_15__N_2408[14])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13163_2_lut.init = 16'h8888;
    LUT4 i13149_2_lut (.A(u_l[15]), .B(\u_s[12] ), .Z(c_15__N_2423[14])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13149_2_lut.init = 16'h8888;
    LUT4 i13164_2_lut (.A(u_l[13]), .B(\u_s[13] ), .Z(c_15__N_2408[13])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13164_2_lut.init = 16'h8888;
    LUT4 i13150_2_lut (.A(u_l[14]), .B(\u_s[12] ), .Z(c_15__N_2423[13])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13150_2_lut.init = 16'h8888;
    CCU2D add_819_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(c_15__N_2408[1]), .B1(c_15__N_2423[1]), .C1(n29267), .D1(n29266), 
          .COUT(n19409), .S1(o_r_17__N_2438[2]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_819_1.INIT0 = 16'hF000;
    defparam add_819_1.INIT1 = 16'h9666;
    defparam add_819_1.INJECT1_0 = "NO";
    defparam add_819_1.INJECT1_1 = "NO";
    LUT4 i13165_2_lut (.A(u_l[12]), .B(\u_s[13] ), .Z(c_15__N_2408[12])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13165_2_lut.init = 16'h8888;
    LUT4 i13151_2_lut (.A(u_l[13]), .B(\u_s[12] ), .Z(c_15__N_2423[12])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13151_2_lut.init = 16'h8888;
    LUT4 i13166_2_lut (.A(u_l[11]), .B(\u_s[13] ), .Z(c_15__N_2408[11])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13166_2_lut.init = 16'h8888;
    LUT4 i13152_2_lut (.A(u_l[12]), .B(\u_s[12] ), .Z(c_15__N_2423[11])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13152_2_lut.init = 16'h8888;
    LUT4 i13167_2_lut (.A(u_l[10]), .B(\u_s[13] ), .Z(c_15__N_2408[10])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13167_2_lut.init = 16'h8888;
    LUT4 i13153_2_lut (.A(u_l[11]), .B(\u_s[12] ), .Z(c_15__N_2423[10])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13153_2_lut.init = 16'h8888;
    LUT4 i13168_2_lut (.A(u_l[9]), .B(\u_s[13] ), .Z(c_15__N_2408[9])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13168_2_lut.init = 16'h8888;
    LUT4 i13154_2_lut (.A(u_l[10]), .B(\u_s[12] ), .Z(c_15__N_2423[9])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13154_2_lut.init = 16'h8888;
    LUT4 i13169_2_lut (.A(u_l[8]), .B(\u_s[13] ), .Z(c_15__N_2408[8])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13169_2_lut.init = 16'h8888;
    LUT4 i13155_2_lut (.A(u_l[9]), .B(\u_s[12] ), .Z(c_15__N_2423[8])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13155_2_lut.init = 16'h8888;
    LUT4 i13170_2_lut (.A(u_l[7]), .B(\u_s[13] ), .Z(c_15__N_2408[7])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13170_2_lut.init = 16'h8888;
    LUT4 i13156_2_lut (.A(u_l[8]), .B(\u_s[12] ), .Z(c_15__N_2423[7])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13156_2_lut.init = 16'h8888;
    LUT4 i13171_2_lut (.A(u_l[6]), .B(\u_s[13] ), .Z(c_15__N_2408[6])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13171_2_lut.init = 16'h8888;
    FD1S3IX o_r__i17 (.D(o_r_17__N_2438[17]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_06[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=90, LSE_RLINE=90 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i17.GSR = "DISABLED";
    LUT4 i13157_2_lut (.A(u_l[7]), .B(\u_s[12] ), .Z(c_15__N_2423[6])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13157_2_lut.init = 16'h8888;
    LUT4 i13172_2_lut (.A(u_l[5]), .B(\u_s[13] ), .Z(c_15__N_2408[5])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13172_2_lut.init = 16'h8888;
    LUT4 i13158_2_lut (.A(u_l[6]), .B(\u_s[12] ), .Z(c_15__N_2423[5])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13158_2_lut.init = 16'h8888;
    LUT4 i13174_2_lut (.A(u_l[4]), .B(\u_s[13] ), .Z(c_15__N_2408[4])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13174_2_lut.init = 16'h8888;
    LUT4 i13159_2_lut (.A(u_l[5]), .B(\u_s[12] ), .Z(c_15__N_2423[4])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13159_2_lut.init = 16'h8888;
    LUT4 i13175_2_lut (.A(u_l[3]), .B(\u_s[13] ), .Z(c_15__N_2408[3])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13175_2_lut.init = 16'h8888;
    LUT4 i13160_2_lut (.A(u_l[4]), .B(\u_s[12] ), .Z(c_15__N_2423[3])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13160_2_lut.init = 16'h8888;
    LUT4 i13176_2_lut (.A(u_l[2]), .B(\u_s[13] ), .Z(c_15__N_2408[2])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13176_2_lut.init = 16'h8888;
    LUT4 i13161_2_lut (.A(u_l[3]), .B(\u_s[12] ), .Z(c_15__N_2423[2])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13161_2_lut.init = 16'h8888;
    LUT4 i13177_2_lut (.A(u_l[1]), .B(\u_s[13] ), .Z(c_15__N_2408[1])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13177_2_lut.init = 16'h8888;
    LUT4 i13162_2_lut (.A(u_l[2]), .B(\u_s[12] ), .Z(c_15__N_2423[1])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13162_2_lut.init = 16'h8888;
    FD1S3IX o_r__i16 (.D(o_r_17__N_2438[16]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_06[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=90, LSE_RLINE=90 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i16.GSR = "DISABLED";
    FD1S3IX o_r__i15 (.D(o_r_17__N_2438[15]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_06[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=90, LSE_RLINE=90 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i15.GSR = "DISABLED";
    FD1S3IX o_r__i14 (.D(o_r_17__N_2438[14]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_06[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=90, LSE_RLINE=90 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i14.GSR = "DISABLED";
    FD1S3IX o_r__i13 (.D(o_r_17__N_2438[13]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_06[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=90, LSE_RLINE=90 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i13.GSR = "DISABLED";
    FD1S3IX o_r__i12 (.D(o_r_17__N_2438[12]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_06[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=90, LSE_RLINE=90 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i12.GSR = "DISABLED";
    FD1S3IX o_r__i11 (.D(o_r_17__N_2438[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_06[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=90, LSE_RLINE=90 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i11.GSR = "DISABLED";
    FD1S3IX o_r__i10 (.D(o_r_17__N_2438[10]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_06[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=90, LSE_RLINE=90 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i10.GSR = "DISABLED";
    FD1S3IX o_r__i9 (.D(o_r_17__N_2438[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_06[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=90, LSE_RLINE=90 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i9.GSR = "DISABLED";
    FD1S3IX o_r__i8 (.D(o_r_17__N_2438[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_06[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=90, LSE_RLINE=90 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i8.GSR = "DISABLED";
    FD1S3IX o_r__i7 (.D(o_r_17__N_2438[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_06[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=90, LSE_RLINE=90 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i7.GSR = "DISABLED";
    FD1S3IX o_r__i6 (.D(o_r_17__N_2438[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_06[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=90, LSE_RLINE=90 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i6.GSR = "DISABLED";
    FD1S3IX o_r__i5 (.D(o_r_17__N_2438[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_06[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=90, LSE_RLINE=90 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i5.GSR = "DISABLED";
    FD1S3IX o_r__i4 (.D(o_r_17__N_2438[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_06[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=90, LSE_RLINE=90 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i4.GSR = "DISABLED";
    FD1S3IX o_r__i3 (.D(o_r_17__N_2438[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_06[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=90, LSE_RLINE=90 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i3.GSR = "DISABLED";
    FD1S3IX o_r__i2 (.D(o_r_17__N_2438[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_06[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=90, LSE_RLINE=90 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i2.GSR = "DISABLED";
    FD1S3IX o_r__i1 (.D(o_r_17__N_2438[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_06[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=90, LSE_RLINE=90 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i1.GSR = "DISABLED";
    LUT4 i12517_2_lut_rep_606 (.A(u_l[1]), .B(\u_s[12] ), .Z(n29266)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i12517_2_lut_rep_606.init = 16'h8888;
    
endmodule
//
// Verilog Description of module \bimpy(BW=16)_U7 
//

module \bimpy(BW=16)_U7  (S_0_05, dac_clk_p_c, n14231, n9446, GND_net, 
            u_l, \u_s[11] , \u_s[10] , i_sw0_c) /* synthesis syn_module_defined=1 */ ;
    output [17:0]S_0_05;
    input dac_clk_p_c;
    input n14231;
    input n9446;
    input GND_net;
    input [15:0]u_l;
    input \u_s[11] ;
    input \u_s[10] ;
    input i_sw0_c;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[29:38])
    
    wire n19439;
    wire [17:0]o_r_17__N_2438;
    
    wire n19438;
    wire [14:0]c_15__N_2408;
    wire [14:0]c_15__N_2423;
    
    wire n19437, n19436, n19435, n19434, n19433, n19432, n29291, 
        n29290;
    
    FD1S3IX o_r__i0 (.D(n9446), .CK(dac_clk_p_c), .CD(n14231), .Q(S_0_05[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=87, LSE_RLINE=87 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i0.GSR = "DISABLED";
    CCU2D add_820_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19439), 
          .S0(o_r_17__N_2438[17]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_820_cout.INIT0 = 16'h0000;
    defparam add_820_cout.INIT1 = 16'h0000;
    defparam add_820_cout.INJECT1_0 = "NO";
    defparam add_820_cout.INJECT1_1 = "NO";
    CCU2D add_820_15 (.A0(c_15__N_2408[14]), .B0(c_15__N_2423[14]), .C0(c_15__N_2408[13]), 
          .D0(c_15__N_2423[13]), .A1(u_l[15]), .B1(\u_s[11] ), .C1(c_15__N_2408[14]), 
          .D1(c_15__N_2423[14]), .CIN(n19438), .COUT(n19439), .S0(o_r_17__N_2438[15]), 
          .S1(o_r_17__N_2438[16]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_820_15.INIT0 = 16'h9666;
    defparam add_820_15.INIT1 = 16'h7888;
    defparam add_820_15.INJECT1_0 = "NO";
    defparam add_820_15.INJECT1_1 = "NO";
    CCU2D add_820_13 (.A0(c_15__N_2408[12]), .B0(c_15__N_2423[12]), .C0(c_15__N_2408[11]), 
          .D0(c_15__N_2423[11]), .A1(c_15__N_2408[13]), .B1(c_15__N_2423[13]), 
          .C1(c_15__N_2408[12]), .D1(c_15__N_2423[12]), .CIN(n19437), 
          .COUT(n19438), .S0(o_r_17__N_2438[13]), .S1(o_r_17__N_2438[14]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_820_13.INIT0 = 16'h9666;
    defparam add_820_13.INIT1 = 16'h9666;
    defparam add_820_13.INJECT1_0 = "NO";
    defparam add_820_13.INJECT1_1 = "NO";
    CCU2D add_820_11 (.A0(c_15__N_2408[10]), .B0(c_15__N_2423[10]), .C0(c_15__N_2408[9]), 
          .D0(c_15__N_2423[9]), .A1(c_15__N_2408[11]), .B1(c_15__N_2423[11]), 
          .C1(c_15__N_2408[10]), .D1(c_15__N_2423[10]), .CIN(n19436), 
          .COUT(n19437), .S0(o_r_17__N_2438[11]), .S1(o_r_17__N_2438[12]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_820_11.INIT0 = 16'h9666;
    defparam add_820_11.INIT1 = 16'h9666;
    defparam add_820_11.INJECT1_0 = "NO";
    defparam add_820_11.INJECT1_1 = "NO";
    CCU2D add_820_9 (.A0(c_15__N_2408[8]), .B0(c_15__N_2423[8]), .C0(c_15__N_2408[7]), 
          .D0(c_15__N_2423[7]), .A1(c_15__N_2408[9]), .B1(c_15__N_2423[9]), 
          .C1(c_15__N_2408[8]), .D1(c_15__N_2423[8]), .CIN(n19435), .COUT(n19436), 
          .S0(o_r_17__N_2438[9]), .S1(o_r_17__N_2438[10]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_820_9.INIT0 = 16'h9666;
    defparam add_820_9.INIT1 = 16'h9666;
    defparam add_820_9.INJECT1_0 = "NO";
    defparam add_820_9.INJECT1_1 = "NO";
    CCU2D add_820_7 (.A0(c_15__N_2408[6]), .B0(c_15__N_2423[6]), .C0(c_15__N_2408[5]), 
          .D0(c_15__N_2423[5]), .A1(c_15__N_2408[7]), .B1(c_15__N_2423[7]), 
          .C1(c_15__N_2408[6]), .D1(c_15__N_2423[6]), .CIN(n19434), .COUT(n19435), 
          .S0(o_r_17__N_2438[7]), .S1(o_r_17__N_2438[8]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_820_7.INIT0 = 16'h9666;
    defparam add_820_7.INIT1 = 16'h9666;
    defparam add_820_7.INJECT1_0 = "NO";
    defparam add_820_7.INJECT1_1 = "NO";
    CCU2D add_820_5 (.A0(c_15__N_2408[4]), .B0(c_15__N_2423[4]), .C0(c_15__N_2408[3]), 
          .D0(c_15__N_2423[3]), .A1(c_15__N_2408[5]), .B1(c_15__N_2423[5]), 
          .C1(c_15__N_2408[4]), .D1(c_15__N_2423[4]), .CIN(n19433), .COUT(n19434), 
          .S0(o_r_17__N_2438[5]), .S1(o_r_17__N_2438[6]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_820_5.INIT0 = 16'h9666;
    defparam add_820_5.INIT1 = 16'h9666;
    defparam add_820_5.INJECT1_0 = "NO";
    defparam add_820_5.INJECT1_1 = "NO";
    CCU2D add_820_3 (.A0(c_15__N_2408[2]), .B0(c_15__N_2423[2]), .C0(c_15__N_2408[1]), 
          .D0(c_15__N_2423[1]), .A1(c_15__N_2408[3]), .B1(c_15__N_2423[3]), 
          .C1(c_15__N_2408[2]), .D1(c_15__N_2423[2]), .CIN(n19432), .COUT(n19433), 
          .S0(o_r_17__N_2438[3]), .S1(o_r_17__N_2438[4]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_820_3.INIT0 = 16'h9666;
    defparam add_820_3.INIT1 = 16'h9666;
    defparam add_820_3.INJECT1_0 = "NO";
    defparam add_820_3.INJECT1_1 = "NO";
    CCU2D add_820_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(c_15__N_2408[1]), .B1(c_15__N_2423[1]), .C1(n29291), .D1(n29290), 
          .COUT(n19432), .S1(o_r_17__N_2438[2]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_820_1.INIT0 = 16'hF000;
    defparam add_820_1.INIT1 = 16'h9666;
    defparam add_820_1.INJECT1_0 = "NO";
    defparam add_820_1.INJECT1_1 = "NO";
    LUT4 i13223_2_lut (.A(u_l[14]), .B(\u_s[11] ), .Z(c_15__N_2408[14])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13223_2_lut.init = 16'h8888;
    LUT4 i13209_2_lut (.A(u_l[15]), .B(\u_s[10] ), .Z(c_15__N_2423[14])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13209_2_lut.init = 16'h8888;
    LUT4 i13225_2_lut (.A(u_l[13]), .B(\u_s[11] ), .Z(c_15__N_2408[13])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13225_2_lut.init = 16'h8888;
    LUT4 i13210_2_lut (.A(u_l[14]), .B(\u_s[10] ), .Z(c_15__N_2423[13])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13210_2_lut.init = 16'h8888;
    LUT4 i13226_2_lut (.A(u_l[12]), .B(\u_s[11] ), .Z(c_15__N_2408[12])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13226_2_lut.init = 16'h8888;
    LUT4 i13211_2_lut (.A(u_l[13]), .B(\u_s[10] ), .Z(c_15__N_2423[12])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13211_2_lut.init = 16'h8888;
    LUT4 i13227_2_lut (.A(u_l[11]), .B(\u_s[11] ), .Z(c_15__N_2408[11])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13227_2_lut.init = 16'h8888;
    LUT4 i13212_2_lut (.A(u_l[12]), .B(\u_s[10] ), .Z(c_15__N_2423[11])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13212_2_lut.init = 16'h8888;
    LUT4 i13228_2_lut (.A(u_l[10]), .B(\u_s[11] ), .Z(c_15__N_2408[10])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13228_2_lut.init = 16'h8888;
    LUT4 i13213_2_lut (.A(u_l[11]), .B(\u_s[10] ), .Z(c_15__N_2423[10])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13213_2_lut.init = 16'h8888;
    LUT4 i13229_2_lut (.A(u_l[9]), .B(\u_s[11] ), .Z(c_15__N_2408[9])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13229_2_lut.init = 16'h8888;
    LUT4 i13214_2_lut (.A(u_l[10]), .B(\u_s[10] ), .Z(c_15__N_2423[9])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13214_2_lut.init = 16'h8888;
    LUT4 i13230_2_lut (.A(u_l[8]), .B(\u_s[11] ), .Z(c_15__N_2408[8])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13230_2_lut.init = 16'h8888;
    LUT4 i13215_2_lut (.A(u_l[9]), .B(\u_s[10] ), .Z(c_15__N_2423[8])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13215_2_lut.init = 16'h8888;
    LUT4 i13231_2_lut (.A(u_l[7]), .B(\u_s[11] ), .Z(c_15__N_2408[7])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13231_2_lut.init = 16'h8888;
    LUT4 i13216_2_lut (.A(u_l[8]), .B(\u_s[10] ), .Z(c_15__N_2423[7])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13216_2_lut.init = 16'h8888;
    LUT4 i13232_2_lut (.A(u_l[6]), .B(\u_s[11] ), .Z(c_15__N_2408[6])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13232_2_lut.init = 16'h8888;
    LUT4 i13217_2_lut (.A(u_l[7]), .B(\u_s[10] ), .Z(c_15__N_2423[6])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13217_2_lut.init = 16'h8888;
    LUT4 i13233_2_lut (.A(u_l[5]), .B(\u_s[11] ), .Z(c_15__N_2408[5])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13233_2_lut.init = 16'h8888;
    LUT4 i13218_2_lut (.A(u_l[6]), .B(\u_s[10] ), .Z(c_15__N_2423[5])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13218_2_lut.init = 16'h8888;
    LUT4 i13234_2_lut (.A(u_l[4]), .B(\u_s[11] ), .Z(c_15__N_2408[4])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13234_2_lut.init = 16'h8888;
    LUT4 i13219_2_lut (.A(u_l[5]), .B(\u_s[10] ), .Z(c_15__N_2423[4])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13219_2_lut.init = 16'h8888;
    LUT4 i13235_2_lut (.A(u_l[3]), .B(\u_s[11] ), .Z(c_15__N_2408[3])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13235_2_lut.init = 16'h8888;
    LUT4 i13220_2_lut (.A(u_l[4]), .B(\u_s[10] ), .Z(c_15__N_2423[3])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13220_2_lut.init = 16'h8888;
    LUT4 i13236_2_lut (.A(u_l[2]), .B(\u_s[11] ), .Z(c_15__N_2408[2])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13236_2_lut.init = 16'h8888;
    LUT4 i13221_2_lut (.A(u_l[3]), .B(\u_s[10] ), .Z(c_15__N_2423[2])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13221_2_lut.init = 16'h8888;
    LUT4 i13237_2_lut (.A(u_l[1]), .B(\u_s[11] ), .Z(c_15__N_2408[1])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13237_2_lut.init = 16'h8888;
    LUT4 i13222_2_lut (.A(u_l[2]), .B(\u_s[10] ), .Z(c_15__N_2423[1])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13222_2_lut.init = 16'h8888;
    LUT4 i12515_2_lut_rep_630 (.A(u_l[1]), .B(\u_s[10] ), .Z(n29290)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i12515_2_lut_rep_630.init = 16'h8888;
    LUT4 i12513_2_lut_rep_631 (.A(u_l[0]), .B(\u_s[11] ), .Z(n29291)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(51[18:45])
    defparam i12513_2_lut_rep_631.init = 16'h8888;
    LUT4 w_r_16__I_0_i2_2_lut_3_lut_4_lut (.A(u_l[0]), .B(\u_s[11] ), .C(\u_s[10] ), 
         .D(u_l[1]), .Z(o_r_17__N_2438[1])) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(51[18:45])
    defparam w_r_16__I_0_i2_2_lut_3_lut_4_lut.init = 16'h7888;
    FD1S3IX o_r__i17 (.D(o_r_17__N_2438[17]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_05[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=87, LSE_RLINE=87 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i17.GSR = "DISABLED";
    FD1S3IX o_r__i16 (.D(o_r_17__N_2438[16]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_05[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=87, LSE_RLINE=87 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i16.GSR = "DISABLED";
    FD1S3IX o_r__i15 (.D(o_r_17__N_2438[15]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_05[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=87, LSE_RLINE=87 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i15.GSR = "DISABLED";
    FD1S3IX o_r__i14 (.D(o_r_17__N_2438[14]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_05[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=87, LSE_RLINE=87 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i14.GSR = "DISABLED";
    FD1S3IX o_r__i13 (.D(o_r_17__N_2438[13]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_05[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=87, LSE_RLINE=87 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i13.GSR = "DISABLED";
    FD1S3IX o_r__i12 (.D(o_r_17__N_2438[12]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_05[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=87, LSE_RLINE=87 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i12.GSR = "DISABLED";
    FD1S3IX o_r__i11 (.D(o_r_17__N_2438[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_05[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=87, LSE_RLINE=87 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i11.GSR = "DISABLED";
    FD1S3IX o_r__i10 (.D(o_r_17__N_2438[10]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_05[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=87, LSE_RLINE=87 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i10.GSR = "DISABLED";
    FD1S3IX o_r__i9 (.D(o_r_17__N_2438[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_05[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=87, LSE_RLINE=87 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i9.GSR = "DISABLED";
    FD1S3IX o_r__i8 (.D(o_r_17__N_2438[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_05[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=87, LSE_RLINE=87 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i8.GSR = "DISABLED";
    FD1S3IX o_r__i7 (.D(o_r_17__N_2438[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_05[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=87, LSE_RLINE=87 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i7.GSR = "DISABLED";
    FD1S3IX o_r__i6 (.D(o_r_17__N_2438[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_05[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=87, LSE_RLINE=87 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i6.GSR = "DISABLED";
    FD1S3IX o_r__i5 (.D(o_r_17__N_2438[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_05[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=87, LSE_RLINE=87 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i5.GSR = "DISABLED";
    FD1S3IX o_r__i4 (.D(o_r_17__N_2438[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_05[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=87, LSE_RLINE=87 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i4.GSR = "DISABLED";
    FD1S3IX o_r__i3 (.D(o_r_17__N_2438[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_05[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=87, LSE_RLINE=87 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i3.GSR = "DISABLED";
    FD1S3IX o_r__i2 (.D(o_r_17__N_2438[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_05[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=87, LSE_RLINE=87 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i2.GSR = "DISABLED";
    FD1S3IX o_r__i1 (.D(o_r_17__N_2438[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_05[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=87, LSE_RLINE=87 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i1.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module \bimpy(BW=16)_U8 
//

module \bimpy(BW=16)_U8  (\S_0_04[0] , dac_clk_p_c, n14231, n9448, GND_net, 
            u_l, \u_s[9] , \u_s[8] , \S_0_04[17] , i_sw0_c, \S_0_04[16] , 
            \S_0_04[15] , \S_0_04[14] , \S_0_04[13] , \S_0_04[12] , 
            \S_0_04[11] , \S_0_04[10] , \S_0_04[9] , \S_0_04[8] , \S_0_04[7] , 
            \S_0_04[6] , \S_0_04[5] , \S_0_04[4] , \S_0_04[3] , \S_0_04[2] , 
            \S_1_02_20__N_2226[1] ) /* synthesis syn_module_defined=1 */ ;
    output \S_0_04[0] ;
    input dac_clk_p_c;
    input n14231;
    input n9448;
    input GND_net;
    input [15:0]u_l;
    input \u_s[9] ;
    input \u_s[8] ;
    output \S_0_04[17] ;
    input i_sw0_c;
    output \S_0_04[16] ;
    output \S_0_04[15] ;
    output \S_0_04[14] ;
    output \S_0_04[13] ;
    output \S_0_04[12] ;
    output \S_0_04[11] ;
    output \S_0_04[10] ;
    output \S_0_04[9] ;
    output \S_0_04[8] ;
    output \S_0_04[7] ;
    output \S_0_04[6] ;
    output \S_0_04[5] ;
    output \S_0_04[4] ;
    output \S_0_04[3] ;
    output \S_0_04[2] ;
    output \S_1_02_20__N_2226[1] ;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[29:38])
    
    wire n19447;
    wire [17:0]o_r_17__N_2438;
    
    wire n19446;
    wire [14:0]c_15__N_2408;
    wire [14:0]c_15__N_2423;
    
    wire n19445, n19444, n19443, n19442, n19441, n19440, n29295, 
        n29294;
    
    FD1S3IX o_r__i0 (.D(n9448), .CK(dac_clk_p_c), .CD(n14231), .Q(\S_0_04[0] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=84, LSE_RLINE=84 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i0.GSR = "DISABLED";
    CCU2D add_821_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19447), 
          .S0(o_r_17__N_2438[17]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_821_cout.INIT0 = 16'h0000;
    defparam add_821_cout.INIT1 = 16'h0000;
    defparam add_821_cout.INJECT1_0 = "NO";
    defparam add_821_cout.INJECT1_1 = "NO";
    CCU2D add_821_15 (.A0(c_15__N_2408[14]), .B0(c_15__N_2423[14]), .C0(c_15__N_2408[13]), 
          .D0(c_15__N_2423[13]), .A1(u_l[15]), .B1(\u_s[9] ), .C1(c_15__N_2408[14]), 
          .D1(c_15__N_2423[14]), .CIN(n19446), .COUT(n19447), .S0(o_r_17__N_2438[15]), 
          .S1(o_r_17__N_2438[16]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_821_15.INIT0 = 16'h9666;
    defparam add_821_15.INIT1 = 16'h7888;
    defparam add_821_15.INJECT1_0 = "NO";
    defparam add_821_15.INJECT1_1 = "NO";
    CCU2D add_821_13 (.A0(c_15__N_2408[12]), .B0(c_15__N_2423[12]), .C0(c_15__N_2408[11]), 
          .D0(c_15__N_2423[11]), .A1(c_15__N_2408[13]), .B1(c_15__N_2423[13]), 
          .C1(c_15__N_2408[12]), .D1(c_15__N_2423[12]), .CIN(n19445), 
          .COUT(n19446), .S0(o_r_17__N_2438[13]), .S1(o_r_17__N_2438[14]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_821_13.INIT0 = 16'h9666;
    defparam add_821_13.INIT1 = 16'h9666;
    defparam add_821_13.INJECT1_0 = "NO";
    defparam add_821_13.INJECT1_1 = "NO";
    CCU2D add_821_11 (.A0(c_15__N_2408[10]), .B0(c_15__N_2423[10]), .C0(c_15__N_2408[9]), 
          .D0(c_15__N_2423[9]), .A1(c_15__N_2408[11]), .B1(c_15__N_2423[11]), 
          .C1(c_15__N_2408[10]), .D1(c_15__N_2423[10]), .CIN(n19444), 
          .COUT(n19445), .S0(o_r_17__N_2438[11]), .S1(o_r_17__N_2438[12]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_821_11.INIT0 = 16'h9666;
    defparam add_821_11.INIT1 = 16'h9666;
    defparam add_821_11.INJECT1_0 = "NO";
    defparam add_821_11.INJECT1_1 = "NO";
    CCU2D add_821_9 (.A0(c_15__N_2408[8]), .B0(c_15__N_2423[8]), .C0(c_15__N_2408[7]), 
          .D0(c_15__N_2423[7]), .A1(c_15__N_2408[9]), .B1(c_15__N_2423[9]), 
          .C1(c_15__N_2408[8]), .D1(c_15__N_2423[8]), .CIN(n19443), .COUT(n19444), 
          .S0(o_r_17__N_2438[9]), .S1(o_r_17__N_2438[10]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_821_9.INIT0 = 16'h9666;
    defparam add_821_9.INIT1 = 16'h9666;
    defparam add_821_9.INJECT1_0 = "NO";
    defparam add_821_9.INJECT1_1 = "NO";
    CCU2D add_821_7 (.A0(c_15__N_2408[6]), .B0(c_15__N_2423[6]), .C0(c_15__N_2408[5]), 
          .D0(c_15__N_2423[5]), .A1(c_15__N_2408[7]), .B1(c_15__N_2423[7]), 
          .C1(c_15__N_2408[6]), .D1(c_15__N_2423[6]), .CIN(n19442), .COUT(n19443), 
          .S0(o_r_17__N_2438[7]), .S1(o_r_17__N_2438[8]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_821_7.INIT0 = 16'h9666;
    defparam add_821_7.INIT1 = 16'h9666;
    defparam add_821_7.INJECT1_0 = "NO";
    defparam add_821_7.INJECT1_1 = "NO";
    CCU2D add_821_5 (.A0(c_15__N_2408[4]), .B0(c_15__N_2423[4]), .C0(c_15__N_2408[3]), 
          .D0(c_15__N_2423[3]), .A1(c_15__N_2408[5]), .B1(c_15__N_2423[5]), 
          .C1(c_15__N_2408[4]), .D1(c_15__N_2423[4]), .CIN(n19441), .COUT(n19442), 
          .S0(o_r_17__N_2438[5]), .S1(o_r_17__N_2438[6]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_821_5.INIT0 = 16'h9666;
    defparam add_821_5.INIT1 = 16'h9666;
    defparam add_821_5.INJECT1_0 = "NO";
    defparam add_821_5.INJECT1_1 = "NO";
    CCU2D add_821_3 (.A0(c_15__N_2408[2]), .B0(c_15__N_2423[2]), .C0(c_15__N_2408[1]), 
          .D0(c_15__N_2423[1]), .A1(c_15__N_2408[3]), .B1(c_15__N_2423[3]), 
          .C1(c_15__N_2408[2]), .D1(c_15__N_2423[2]), .CIN(n19440), .COUT(n19441), 
          .S0(o_r_17__N_2438[3]), .S1(o_r_17__N_2438[4]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_821_3.INIT0 = 16'h9666;
    defparam add_821_3.INIT1 = 16'h9666;
    defparam add_821_3.INJECT1_0 = "NO";
    defparam add_821_3.INJECT1_1 = "NO";
    CCU2D add_821_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(c_15__N_2408[1]), .B1(c_15__N_2423[1]), .C1(n29295), .D1(n29294), 
          .COUT(n19440), .S1(o_r_17__N_2438[2]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_821_1.INIT0 = 16'hF000;
    defparam add_821_1.INIT1 = 16'h9666;
    defparam add_821_1.INJECT1_0 = "NO";
    defparam add_821_1.INJECT1_1 = "NO";
    LUT4 i13262_2_lut (.A(u_l[14]), .B(\u_s[9] ), .Z(c_15__N_2408[14])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13262_2_lut.init = 16'h8888;
    LUT4 i13244_2_lut (.A(u_l[15]), .B(\u_s[8] ), .Z(c_15__N_2423[14])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13244_2_lut.init = 16'h8888;
    LUT4 i13263_2_lut (.A(u_l[13]), .B(\u_s[9] ), .Z(c_15__N_2408[13])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13263_2_lut.init = 16'h8888;
    LUT4 i13245_2_lut (.A(u_l[14]), .B(\u_s[8] ), .Z(c_15__N_2423[13])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13245_2_lut.init = 16'h8888;
    LUT4 i13264_2_lut (.A(u_l[12]), .B(\u_s[9] ), .Z(c_15__N_2408[12])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13264_2_lut.init = 16'h8888;
    LUT4 i13247_2_lut (.A(u_l[13]), .B(\u_s[8] ), .Z(c_15__N_2423[12])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13247_2_lut.init = 16'h8888;
    LUT4 i13265_2_lut (.A(u_l[11]), .B(\u_s[9] ), .Z(c_15__N_2408[11])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13265_2_lut.init = 16'h8888;
    LUT4 i13250_2_lut (.A(u_l[12]), .B(\u_s[8] ), .Z(c_15__N_2423[11])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13250_2_lut.init = 16'h8888;
    LUT4 i13266_2_lut (.A(u_l[10]), .B(\u_s[9] ), .Z(c_15__N_2408[10])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13266_2_lut.init = 16'h8888;
    LUT4 i13251_2_lut (.A(u_l[11]), .B(\u_s[8] ), .Z(c_15__N_2423[10])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13251_2_lut.init = 16'h8888;
    LUT4 i13267_2_lut (.A(u_l[9]), .B(\u_s[9] ), .Z(c_15__N_2408[9])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13267_2_lut.init = 16'h8888;
    LUT4 i13252_2_lut (.A(u_l[10]), .B(\u_s[8] ), .Z(c_15__N_2423[9])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13252_2_lut.init = 16'h8888;
    LUT4 i13268_2_lut (.A(u_l[8]), .B(\u_s[9] ), .Z(c_15__N_2408[8])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13268_2_lut.init = 16'h8888;
    LUT4 i13254_2_lut (.A(u_l[9]), .B(\u_s[8] ), .Z(c_15__N_2423[8])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13254_2_lut.init = 16'h8888;
    LUT4 i13269_2_lut (.A(u_l[7]), .B(\u_s[9] ), .Z(c_15__N_2408[7])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13269_2_lut.init = 16'h8888;
    LUT4 i13255_2_lut (.A(u_l[8]), .B(\u_s[8] ), .Z(c_15__N_2423[7])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13255_2_lut.init = 16'h8888;
    LUT4 i13270_2_lut (.A(u_l[6]), .B(\u_s[9] ), .Z(c_15__N_2408[6])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13270_2_lut.init = 16'h8888;
    LUT4 i13256_2_lut (.A(u_l[7]), .B(\u_s[8] ), .Z(c_15__N_2423[6])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13256_2_lut.init = 16'h8888;
    LUT4 i13271_2_lut (.A(u_l[5]), .B(\u_s[9] ), .Z(c_15__N_2408[5])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13271_2_lut.init = 16'h8888;
    LUT4 i13257_2_lut (.A(u_l[6]), .B(\u_s[8] ), .Z(c_15__N_2423[5])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13257_2_lut.init = 16'h8888;
    LUT4 i13272_2_lut (.A(u_l[4]), .B(\u_s[9] ), .Z(c_15__N_2408[4])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13272_2_lut.init = 16'h8888;
    LUT4 i13258_2_lut (.A(u_l[5]), .B(\u_s[8] ), .Z(c_15__N_2423[4])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13258_2_lut.init = 16'h8888;
    LUT4 i13273_2_lut (.A(u_l[3]), .B(\u_s[9] ), .Z(c_15__N_2408[3])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13273_2_lut.init = 16'h8888;
    LUT4 i13259_2_lut (.A(u_l[4]), .B(\u_s[8] ), .Z(c_15__N_2423[3])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13259_2_lut.init = 16'h8888;
    LUT4 i13274_2_lut (.A(u_l[2]), .B(\u_s[9] ), .Z(c_15__N_2408[2])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13274_2_lut.init = 16'h8888;
    LUT4 i13260_2_lut (.A(u_l[3]), .B(\u_s[8] ), .Z(c_15__N_2423[2])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13260_2_lut.init = 16'h8888;
    LUT4 i13275_2_lut (.A(u_l[1]), .B(\u_s[9] ), .Z(c_15__N_2408[1])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13275_2_lut.init = 16'h8888;
    LUT4 i13261_2_lut (.A(u_l[2]), .B(\u_s[8] ), .Z(c_15__N_2423[1])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13261_2_lut.init = 16'h8888;
    LUT4 i12512_2_lut_rep_634 (.A(u_l[1]), .B(\u_s[8] ), .Z(n29294)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i12512_2_lut_rep_634.init = 16'h8888;
    LUT4 i12510_2_lut_rep_635 (.A(u_l[0]), .B(\u_s[9] ), .Z(n29295)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(51[18:45])
    defparam i12510_2_lut_rep_635.init = 16'h8888;
    LUT4 w_r_16__I_0_i2_2_lut_3_lut_4_lut (.A(u_l[0]), .B(\u_s[9] ), .C(\u_s[8] ), 
         .D(u_l[1]), .Z(o_r_17__N_2438[1])) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(51[18:45])
    defparam w_r_16__I_0_i2_2_lut_3_lut_4_lut.init = 16'h7888;
    FD1S3IX o_r__i17 (.D(o_r_17__N_2438[17]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_04[17] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=84, LSE_RLINE=84 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i17.GSR = "DISABLED";
    FD1S3IX o_r__i16 (.D(o_r_17__N_2438[16]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_04[16] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=84, LSE_RLINE=84 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i16.GSR = "DISABLED";
    FD1S3IX o_r__i15 (.D(o_r_17__N_2438[15]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_04[15] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=84, LSE_RLINE=84 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i15.GSR = "DISABLED";
    FD1S3IX o_r__i14 (.D(o_r_17__N_2438[14]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_04[14] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=84, LSE_RLINE=84 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i14.GSR = "DISABLED";
    FD1S3IX o_r__i13 (.D(o_r_17__N_2438[13]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_04[13] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=84, LSE_RLINE=84 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i13.GSR = "DISABLED";
    FD1S3IX o_r__i12 (.D(o_r_17__N_2438[12]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_04[12] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=84, LSE_RLINE=84 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i12.GSR = "DISABLED";
    FD1S3IX o_r__i11 (.D(o_r_17__N_2438[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_04[11] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=84, LSE_RLINE=84 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i11.GSR = "DISABLED";
    FD1S3IX o_r__i10 (.D(o_r_17__N_2438[10]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_04[10] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=84, LSE_RLINE=84 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i10.GSR = "DISABLED";
    FD1S3IX o_r__i9 (.D(o_r_17__N_2438[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_04[9] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=84, LSE_RLINE=84 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i9.GSR = "DISABLED";
    FD1S3IX o_r__i8 (.D(o_r_17__N_2438[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_04[8] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=84, LSE_RLINE=84 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i8.GSR = "DISABLED";
    FD1S3IX o_r__i7 (.D(o_r_17__N_2438[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_04[7] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=84, LSE_RLINE=84 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i7.GSR = "DISABLED";
    FD1S3IX o_r__i6 (.D(o_r_17__N_2438[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_04[6] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=84, LSE_RLINE=84 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i6.GSR = "DISABLED";
    FD1S3IX o_r__i5 (.D(o_r_17__N_2438[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_04[5] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=84, LSE_RLINE=84 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i5.GSR = "DISABLED";
    FD1S3IX o_r__i4 (.D(o_r_17__N_2438[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_04[4] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=84, LSE_RLINE=84 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i4.GSR = "DISABLED";
    FD1S3IX o_r__i3 (.D(o_r_17__N_2438[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_04[3] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=84, LSE_RLINE=84 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i3.GSR = "DISABLED";
    FD1S3IX o_r__i2 (.D(o_r_17__N_2438[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_04[2] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=84, LSE_RLINE=84 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i2.GSR = "DISABLED";
    FD1S3IX o_r__i1 (.D(o_r_17__N_2438[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_1_02_20__N_2226[1] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=84, LSE_RLINE=84 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i1.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module \bimpy(BW=16)_U9 
//

module \bimpy(BW=16)_U9  (GND_net, u_l, \u_s[7] , S_0_03, dac_clk_p_c, 
            n14231, n9450, \u_s[6] , i_sw0_c) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input [15:0]u_l;
    input \u_s[7] ;
    output [17:0]S_0_03;
    input dac_clk_p_c;
    input n14231;
    input n9450;
    input \u_s[6] ;
    input i_sw0_c;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[29:38])
    
    wire n19455;
    wire [17:0]o_r_17__N_2438;
    
    wire n19454;
    wire [14:0]c_15__N_2408;
    wire [14:0]c_15__N_2423;
    
    wire n19453, n19452, n19451, n19450, n19449, n19448, n29306, 
        n29305;
    
    CCU2D add_822_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19455), 
          .S0(o_r_17__N_2438[17]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_822_cout.INIT0 = 16'h0000;
    defparam add_822_cout.INIT1 = 16'h0000;
    defparam add_822_cout.INJECT1_0 = "NO";
    defparam add_822_cout.INJECT1_1 = "NO";
    CCU2D add_822_15 (.A0(c_15__N_2408[14]), .B0(c_15__N_2423[14]), .C0(c_15__N_2408[13]), 
          .D0(c_15__N_2423[13]), .A1(u_l[15]), .B1(\u_s[7] ), .C1(c_15__N_2408[14]), 
          .D1(c_15__N_2423[14]), .CIN(n19454), .COUT(n19455), .S0(o_r_17__N_2438[15]), 
          .S1(o_r_17__N_2438[16]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_822_15.INIT0 = 16'h9666;
    defparam add_822_15.INIT1 = 16'h7888;
    defparam add_822_15.INJECT1_0 = "NO";
    defparam add_822_15.INJECT1_1 = "NO";
    CCU2D add_822_13 (.A0(c_15__N_2408[12]), .B0(c_15__N_2423[12]), .C0(c_15__N_2408[11]), 
          .D0(c_15__N_2423[11]), .A1(c_15__N_2408[13]), .B1(c_15__N_2423[13]), 
          .C1(c_15__N_2408[12]), .D1(c_15__N_2423[12]), .CIN(n19453), 
          .COUT(n19454), .S0(o_r_17__N_2438[13]), .S1(o_r_17__N_2438[14]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_822_13.INIT0 = 16'h9666;
    defparam add_822_13.INIT1 = 16'h9666;
    defparam add_822_13.INJECT1_0 = "NO";
    defparam add_822_13.INJECT1_1 = "NO";
    FD1S3IX o_r__i0 (.D(n9450), .CK(dac_clk_p_c), .CD(n14231), .Q(S_0_03[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=81, LSE_RLINE=81 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i0.GSR = "DISABLED";
    CCU2D add_822_11 (.A0(c_15__N_2408[10]), .B0(c_15__N_2423[10]), .C0(c_15__N_2408[9]), 
          .D0(c_15__N_2423[9]), .A1(c_15__N_2408[11]), .B1(c_15__N_2423[11]), 
          .C1(c_15__N_2408[10]), .D1(c_15__N_2423[10]), .CIN(n19452), 
          .COUT(n19453), .S0(o_r_17__N_2438[11]), .S1(o_r_17__N_2438[12]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_822_11.INIT0 = 16'h9666;
    defparam add_822_11.INIT1 = 16'h9666;
    defparam add_822_11.INJECT1_0 = "NO";
    defparam add_822_11.INJECT1_1 = "NO";
    CCU2D add_822_9 (.A0(c_15__N_2408[8]), .B0(c_15__N_2423[8]), .C0(c_15__N_2408[7]), 
          .D0(c_15__N_2423[7]), .A1(c_15__N_2408[9]), .B1(c_15__N_2423[9]), 
          .C1(c_15__N_2408[8]), .D1(c_15__N_2423[8]), .CIN(n19451), .COUT(n19452), 
          .S0(o_r_17__N_2438[9]), .S1(o_r_17__N_2438[10]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_822_9.INIT0 = 16'h9666;
    defparam add_822_9.INIT1 = 16'h9666;
    defparam add_822_9.INJECT1_0 = "NO";
    defparam add_822_9.INJECT1_1 = "NO";
    CCU2D add_822_7 (.A0(c_15__N_2408[6]), .B0(c_15__N_2423[6]), .C0(c_15__N_2408[5]), 
          .D0(c_15__N_2423[5]), .A1(c_15__N_2408[7]), .B1(c_15__N_2423[7]), 
          .C1(c_15__N_2408[6]), .D1(c_15__N_2423[6]), .CIN(n19450), .COUT(n19451), 
          .S0(o_r_17__N_2438[7]), .S1(o_r_17__N_2438[8]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_822_7.INIT0 = 16'h9666;
    defparam add_822_7.INIT1 = 16'h9666;
    defparam add_822_7.INJECT1_0 = "NO";
    defparam add_822_7.INJECT1_1 = "NO";
    CCU2D add_822_5 (.A0(c_15__N_2408[4]), .B0(c_15__N_2423[4]), .C0(c_15__N_2408[3]), 
          .D0(c_15__N_2423[3]), .A1(c_15__N_2408[5]), .B1(c_15__N_2423[5]), 
          .C1(c_15__N_2408[4]), .D1(c_15__N_2423[4]), .CIN(n19449), .COUT(n19450), 
          .S0(o_r_17__N_2438[5]), .S1(o_r_17__N_2438[6]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_822_5.INIT0 = 16'h9666;
    defparam add_822_5.INIT1 = 16'h9666;
    defparam add_822_5.INJECT1_0 = "NO";
    defparam add_822_5.INJECT1_1 = "NO";
    LUT4 i13292_2_lut (.A(u_l[14]), .B(\u_s[7] ), .Z(c_15__N_2408[14])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13292_2_lut.init = 16'h8888;
    LUT4 i13278_2_lut (.A(u_l[15]), .B(\u_s[6] ), .Z(c_15__N_2423[14])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13278_2_lut.init = 16'h8888;
    LUT4 i13293_2_lut (.A(u_l[13]), .B(\u_s[7] ), .Z(c_15__N_2408[13])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13293_2_lut.init = 16'h8888;
    CCU2D add_822_3 (.A0(c_15__N_2408[2]), .B0(c_15__N_2423[2]), .C0(c_15__N_2408[1]), 
          .D0(c_15__N_2423[1]), .A1(c_15__N_2408[3]), .B1(c_15__N_2423[3]), 
          .C1(c_15__N_2408[2]), .D1(c_15__N_2423[2]), .CIN(n19448), .COUT(n19449), 
          .S0(o_r_17__N_2438[3]), .S1(o_r_17__N_2438[4]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_822_3.INIT0 = 16'h9666;
    defparam add_822_3.INIT1 = 16'h9666;
    defparam add_822_3.INJECT1_0 = "NO";
    defparam add_822_3.INJECT1_1 = "NO";
    LUT4 i13279_2_lut (.A(u_l[14]), .B(\u_s[6] ), .Z(c_15__N_2423[13])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13279_2_lut.init = 16'h8888;
    CCU2D add_822_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(c_15__N_2408[1]), .B1(c_15__N_2423[1]), .C1(n29306), .D1(n29305), 
          .COUT(n19448), .S1(o_r_17__N_2438[2]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_822_1.INIT0 = 16'hF000;
    defparam add_822_1.INIT1 = 16'h9666;
    defparam add_822_1.INJECT1_0 = "NO";
    defparam add_822_1.INJECT1_1 = "NO";
    LUT4 i13294_2_lut (.A(u_l[12]), .B(\u_s[7] ), .Z(c_15__N_2408[12])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13294_2_lut.init = 16'h8888;
    LUT4 i13280_2_lut (.A(u_l[13]), .B(\u_s[6] ), .Z(c_15__N_2423[12])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13280_2_lut.init = 16'h8888;
    LUT4 i13295_2_lut (.A(u_l[11]), .B(\u_s[7] ), .Z(c_15__N_2408[11])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13295_2_lut.init = 16'h8888;
    LUT4 i13281_2_lut (.A(u_l[12]), .B(\u_s[6] ), .Z(c_15__N_2423[11])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13281_2_lut.init = 16'h8888;
    LUT4 i13296_2_lut (.A(u_l[10]), .B(\u_s[7] ), .Z(c_15__N_2408[10])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13296_2_lut.init = 16'h8888;
    LUT4 i13282_2_lut (.A(u_l[11]), .B(\u_s[6] ), .Z(c_15__N_2423[10])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13282_2_lut.init = 16'h8888;
    LUT4 i13297_2_lut (.A(u_l[9]), .B(\u_s[7] ), .Z(c_15__N_2408[9])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13297_2_lut.init = 16'h8888;
    LUT4 i13283_2_lut (.A(u_l[10]), .B(\u_s[6] ), .Z(c_15__N_2423[9])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13283_2_lut.init = 16'h8888;
    LUT4 i13298_2_lut (.A(u_l[8]), .B(\u_s[7] ), .Z(c_15__N_2408[8])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13298_2_lut.init = 16'h8888;
    LUT4 i13284_2_lut (.A(u_l[9]), .B(\u_s[6] ), .Z(c_15__N_2423[8])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13284_2_lut.init = 16'h8888;
    LUT4 i13299_2_lut (.A(u_l[7]), .B(\u_s[7] ), .Z(c_15__N_2408[7])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13299_2_lut.init = 16'h8888;
    LUT4 i13285_2_lut (.A(u_l[8]), .B(\u_s[6] ), .Z(c_15__N_2423[7])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13285_2_lut.init = 16'h8888;
    LUT4 i13300_2_lut (.A(u_l[6]), .B(\u_s[7] ), .Z(c_15__N_2408[6])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13300_2_lut.init = 16'h8888;
    LUT4 i13286_2_lut (.A(u_l[7]), .B(\u_s[6] ), .Z(c_15__N_2423[6])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13286_2_lut.init = 16'h8888;
    LUT4 i13301_2_lut (.A(u_l[5]), .B(\u_s[7] ), .Z(c_15__N_2408[5])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13301_2_lut.init = 16'h8888;
    LUT4 i13287_2_lut (.A(u_l[6]), .B(\u_s[6] ), .Z(c_15__N_2423[5])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13287_2_lut.init = 16'h8888;
    LUT4 i13302_2_lut (.A(u_l[4]), .B(\u_s[7] ), .Z(c_15__N_2408[4])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13302_2_lut.init = 16'h8888;
    LUT4 i13288_2_lut (.A(u_l[5]), .B(\u_s[6] ), .Z(c_15__N_2423[4])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13288_2_lut.init = 16'h8888;
    LUT4 i13303_2_lut (.A(u_l[3]), .B(\u_s[7] ), .Z(c_15__N_2408[3])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13303_2_lut.init = 16'h8888;
    LUT4 i13289_2_lut (.A(u_l[4]), .B(\u_s[6] ), .Z(c_15__N_2423[3])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13289_2_lut.init = 16'h8888;
    LUT4 i13304_2_lut (.A(u_l[2]), .B(\u_s[7] ), .Z(c_15__N_2408[2])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13304_2_lut.init = 16'h8888;
    LUT4 i13290_2_lut (.A(u_l[3]), .B(\u_s[6] ), .Z(c_15__N_2423[2])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13290_2_lut.init = 16'h8888;
    LUT4 i13305_2_lut (.A(u_l[1]), .B(\u_s[7] ), .Z(c_15__N_2408[1])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13305_2_lut.init = 16'h8888;
    LUT4 i13291_2_lut (.A(u_l[2]), .B(\u_s[6] ), .Z(c_15__N_2423[1])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13291_2_lut.init = 16'h8888;
    LUT4 i12509_2_lut_rep_645 (.A(u_l[1]), .B(\u_s[6] ), .Z(n29305)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i12509_2_lut_rep_645.init = 16'h8888;
    LUT4 i12508_2_lut_rep_646 (.A(u_l[0]), .B(\u_s[7] ), .Z(n29306)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(51[18:45])
    defparam i12508_2_lut_rep_646.init = 16'h8888;
    LUT4 w_r_16__I_0_i2_2_lut_3_lut_4_lut (.A(u_l[0]), .B(\u_s[7] ), .C(\u_s[6] ), 
         .D(u_l[1]), .Z(o_r_17__N_2438[1])) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(51[18:45])
    defparam w_r_16__I_0_i2_2_lut_3_lut_4_lut.init = 16'h7888;
    FD1S3IX o_r__i17 (.D(o_r_17__N_2438[17]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_03[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=81, LSE_RLINE=81 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i17.GSR = "DISABLED";
    FD1S3IX o_r__i16 (.D(o_r_17__N_2438[16]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_03[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=81, LSE_RLINE=81 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i16.GSR = "DISABLED";
    FD1S3IX o_r__i15 (.D(o_r_17__N_2438[15]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_03[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=81, LSE_RLINE=81 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i15.GSR = "DISABLED";
    FD1S3IX o_r__i14 (.D(o_r_17__N_2438[14]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_03[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=81, LSE_RLINE=81 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i14.GSR = "DISABLED";
    FD1S3IX o_r__i13 (.D(o_r_17__N_2438[13]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_03[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=81, LSE_RLINE=81 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i13.GSR = "DISABLED";
    FD1S3IX o_r__i12 (.D(o_r_17__N_2438[12]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_03[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=81, LSE_RLINE=81 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i12.GSR = "DISABLED";
    FD1S3IX o_r__i11 (.D(o_r_17__N_2438[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_03[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=81, LSE_RLINE=81 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i11.GSR = "DISABLED";
    FD1S3IX o_r__i10 (.D(o_r_17__N_2438[10]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_03[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=81, LSE_RLINE=81 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i10.GSR = "DISABLED";
    FD1S3IX o_r__i9 (.D(o_r_17__N_2438[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_03[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=81, LSE_RLINE=81 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i9.GSR = "DISABLED";
    FD1S3IX o_r__i8 (.D(o_r_17__N_2438[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_03[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=81, LSE_RLINE=81 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i8.GSR = "DISABLED";
    FD1S3IX o_r__i7 (.D(o_r_17__N_2438[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_03[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=81, LSE_RLINE=81 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i7.GSR = "DISABLED";
    FD1S3IX o_r__i6 (.D(o_r_17__N_2438[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_03[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=81, LSE_RLINE=81 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i6.GSR = "DISABLED";
    FD1S3IX o_r__i5 (.D(o_r_17__N_2438[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_03[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=81, LSE_RLINE=81 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i5.GSR = "DISABLED";
    FD1S3IX o_r__i4 (.D(o_r_17__N_2438[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_03[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=81, LSE_RLINE=81 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i4.GSR = "DISABLED";
    FD1S3IX o_r__i3 (.D(o_r_17__N_2438[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_03[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=81, LSE_RLINE=81 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i3.GSR = "DISABLED";
    FD1S3IX o_r__i2 (.D(o_r_17__N_2438[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_03[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=81, LSE_RLINE=81 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i2.GSR = "DISABLED";
    FD1S3IX o_r__i1 (.D(o_r_17__N_2438[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_03[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=81, LSE_RLINE=81 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i1.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module \bimpy(BW=16)_U10 
//

module \bimpy(BW=16)_U10  (GND_net, \S_0_02[0] , dac_clk_p_c, n14231, 
            n9452, u_l, \u_s[5] , \u_s[4] , \S_0_02[17] , i_sw0_c, 
            \S_0_02[16] , \S_0_02[15] , \S_0_02[14] , \S_0_02[13] , 
            \S_0_02[12] , \S_0_02[11] , \S_0_02[10] , \S_0_02[9] , \S_0_02[8] , 
            \S_0_02[7] , \S_0_02[6] , \S_0_02[5] , \S_0_02[4] , \S_0_02[3] , 
            \S_0_02[2] , \S_1_01_20__N_2205[1] ) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output \S_0_02[0] ;
    input dac_clk_p_c;
    input n14231;
    input n9452;
    input [15:0]u_l;
    input \u_s[5] ;
    input \u_s[4] ;
    output \S_0_02[17] ;
    input i_sw0_c;
    output \S_0_02[16] ;
    output \S_0_02[15] ;
    output \S_0_02[14] ;
    output \S_0_02[13] ;
    output \S_0_02[12] ;
    output \S_0_02[11] ;
    output \S_0_02[10] ;
    output \S_0_02[9] ;
    output \S_0_02[8] ;
    output \S_0_02[7] ;
    output \S_0_02[6] ;
    output \S_0_02[5] ;
    output \S_0_02[4] ;
    output \S_0_02[3] ;
    output \S_0_02[2] ;
    output \S_1_01_20__N_2205[1] ;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[29:38])
    
    wire n19456;
    wire [14:0]c_15__N_2408;
    wire [14:0]c_15__N_2423;
    wire [17:0]o_r_17__N_2438;
    
    wire n19457, n29454, n29453, n19463, n19462, n19461, n19460, 
        n19459, n19458;
    
    CCU2D add_823_3 (.A0(c_15__N_2408[2]), .B0(c_15__N_2423[2]), .C0(c_15__N_2408[1]), 
          .D0(c_15__N_2423[1]), .A1(c_15__N_2408[3]), .B1(c_15__N_2423[3]), 
          .C1(c_15__N_2408[2]), .D1(c_15__N_2423[2]), .CIN(n19456), .COUT(n19457), 
          .S0(o_r_17__N_2438[3]), .S1(o_r_17__N_2438[4]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_823_3.INIT0 = 16'h9666;
    defparam add_823_3.INIT1 = 16'h9666;
    defparam add_823_3.INJECT1_0 = "NO";
    defparam add_823_3.INJECT1_1 = "NO";
    CCU2D add_823_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(c_15__N_2408[1]), .B1(c_15__N_2423[1]), .C1(n29454), .D1(n29453), 
          .COUT(n19456), .S1(o_r_17__N_2438[2]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_823_1.INIT0 = 16'hF000;
    defparam add_823_1.INIT1 = 16'h9666;
    defparam add_823_1.INJECT1_0 = "NO";
    defparam add_823_1.INJECT1_1 = "NO";
    FD1S3IX o_r__i0 (.D(n9452), .CK(dac_clk_p_c), .CD(n14231), .Q(\S_0_02[0] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i0.GSR = "DISABLED";
    LUT4 i13339_2_lut (.A(u_l[2]), .B(\u_s[5] ), .Z(c_15__N_2408[2])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13339_2_lut.init = 16'h8888;
    LUT4 i13325_2_lut (.A(u_l[3]), .B(\u_s[4] ), .Z(c_15__N_2423[2])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13325_2_lut.init = 16'h8888;
    LUT4 i13340_2_lut (.A(u_l[1]), .B(\u_s[5] ), .Z(c_15__N_2408[1])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13340_2_lut.init = 16'h8888;
    LUT4 i13326_2_lut (.A(u_l[2]), .B(\u_s[4] ), .Z(c_15__N_2423[1])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13326_2_lut.init = 16'h8888;
    LUT4 i13338_2_lut (.A(u_l[3]), .B(\u_s[5] ), .Z(c_15__N_2408[3])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13338_2_lut.init = 16'h8888;
    LUT4 i13324_2_lut (.A(u_l[4]), .B(\u_s[4] ), .Z(c_15__N_2423[3])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13324_2_lut.init = 16'h8888;
    FD1S3IX o_r__i17 (.D(o_r_17__N_2438[17]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_02[17] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i17.GSR = "DISABLED";
    FD1S3IX o_r__i16 (.D(o_r_17__N_2438[16]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_02[16] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i16.GSR = "DISABLED";
    FD1S3IX o_r__i15 (.D(o_r_17__N_2438[15]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_02[15] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i15.GSR = "DISABLED";
    FD1S3IX o_r__i14 (.D(o_r_17__N_2438[14]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_02[14] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i14.GSR = "DISABLED";
    FD1S3IX o_r__i13 (.D(o_r_17__N_2438[13]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_02[13] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i13.GSR = "DISABLED";
    FD1S3IX o_r__i12 (.D(o_r_17__N_2438[12]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_02[12] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i12.GSR = "DISABLED";
    FD1S3IX o_r__i11 (.D(o_r_17__N_2438[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_02[11] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i11.GSR = "DISABLED";
    FD1S3IX o_r__i10 (.D(o_r_17__N_2438[10]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_02[10] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i10.GSR = "DISABLED";
    FD1S3IX o_r__i9 (.D(o_r_17__N_2438[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_02[9] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i9.GSR = "DISABLED";
    FD1S3IX o_r__i8 (.D(o_r_17__N_2438[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_02[8] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i8.GSR = "DISABLED";
    FD1S3IX o_r__i7 (.D(o_r_17__N_2438[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_02[7] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i7.GSR = "DISABLED";
    FD1S3IX o_r__i6 (.D(o_r_17__N_2438[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_02[6] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i6.GSR = "DISABLED";
    FD1S3IX o_r__i5 (.D(o_r_17__N_2438[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_02[5] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i5.GSR = "DISABLED";
    FD1S3IX o_r__i4 (.D(o_r_17__N_2438[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_02[4] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i4.GSR = "DISABLED";
    FD1S3IX o_r__i3 (.D(o_r_17__N_2438[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_02[3] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i3.GSR = "DISABLED";
    FD1S3IX o_r__i2 (.D(o_r_17__N_2438[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_02[2] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i2.GSR = "DISABLED";
    FD1S3IX o_r__i1 (.D(o_r_17__N_2438[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_1_01_20__N_2205[1] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i1.GSR = "DISABLED";
    LUT4 i12507_2_lut_rep_793 (.A(u_l[1]), .B(\u_s[4] ), .Z(n29453)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i12507_2_lut_rep_793.init = 16'h8888;
    LUT4 i12506_2_lut_rep_794 (.A(u_l[0]), .B(\u_s[5] ), .Z(n29454)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(51[18:45])
    defparam i12506_2_lut_rep_794.init = 16'h8888;
    LUT4 w_r_16__I_0_i2_2_lut_3_lut_4_lut (.A(u_l[0]), .B(\u_s[5] ), .C(\u_s[4] ), 
         .D(u_l[1]), .Z(o_r_17__N_2438[1])) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(51[18:45])
    defparam w_r_16__I_0_i2_2_lut_3_lut_4_lut.init = 16'h7888;
    LUT4 i13327_2_lut (.A(u_l[14]), .B(\u_s[5] ), .Z(c_15__N_2408[14])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13327_2_lut.init = 16'h8888;
    LUT4 i13313_2_lut (.A(u_l[15]), .B(\u_s[4] ), .Z(c_15__N_2423[14])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13313_2_lut.init = 16'h8888;
    LUT4 i13328_2_lut (.A(u_l[13]), .B(\u_s[5] ), .Z(c_15__N_2408[13])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13328_2_lut.init = 16'h8888;
    LUT4 i13314_2_lut (.A(u_l[14]), .B(\u_s[4] ), .Z(c_15__N_2423[13])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13314_2_lut.init = 16'h8888;
    LUT4 i13329_2_lut (.A(u_l[12]), .B(\u_s[5] ), .Z(c_15__N_2408[12])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13329_2_lut.init = 16'h8888;
    LUT4 i13315_2_lut (.A(u_l[13]), .B(\u_s[4] ), .Z(c_15__N_2423[12])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13315_2_lut.init = 16'h8888;
    LUT4 i13330_2_lut (.A(u_l[11]), .B(\u_s[5] ), .Z(c_15__N_2408[11])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13330_2_lut.init = 16'h8888;
    LUT4 i13316_2_lut (.A(u_l[12]), .B(\u_s[4] ), .Z(c_15__N_2423[11])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13316_2_lut.init = 16'h8888;
    LUT4 i13331_2_lut (.A(u_l[10]), .B(\u_s[5] ), .Z(c_15__N_2408[10])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13331_2_lut.init = 16'h8888;
    LUT4 i13317_2_lut (.A(u_l[11]), .B(\u_s[4] ), .Z(c_15__N_2423[10])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13317_2_lut.init = 16'h8888;
    LUT4 i13332_2_lut (.A(u_l[9]), .B(\u_s[5] ), .Z(c_15__N_2408[9])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13332_2_lut.init = 16'h8888;
    LUT4 i13318_2_lut (.A(u_l[10]), .B(\u_s[4] ), .Z(c_15__N_2423[9])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13318_2_lut.init = 16'h8888;
    LUT4 i13333_2_lut (.A(u_l[8]), .B(\u_s[5] ), .Z(c_15__N_2408[8])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13333_2_lut.init = 16'h8888;
    LUT4 i13319_2_lut (.A(u_l[9]), .B(\u_s[4] ), .Z(c_15__N_2423[8])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13319_2_lut.init = 16'h8888;
    LUT4 i13334_2_lut (.A(u_l[7]), .B(\u_s[5] ), .Z(c_15__N_2408[7])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13334_2_lut.init = 16'h8888;
    LUT4 i13320_2_lut (.A(u_l[8]), .B(\u_s[4] ), .Z(c_15__N_2423[7])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13320_2_lut.init = 16'h8888;
    LUT4 i13335_2_lut (.A(u_l[6]), .B(\u_s[5] ), .Z(c_15__N_2408[6])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13335_2_lut.init = 16'h8888;
    LUT4 i13321_2_lut (.A(u_l[7]), .B(\u_s[4] ), .Z(c_15__N_2423[6])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13321_2_lut.init = 16'h8888;
    LUT4 i13336_2_lut (.A(u_l[5]), .B(\u_s[5] ), .Z(c_15__N_2408[5])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13336_2_lut.init = 16'h8888;
    LUT4 i13322_2_lut (.A(u_l[6]), .B(\u_s[4] ), .Z(c_15__N_2423[5])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13322_2_lut.init = 16'h8888;
    LUT4 i13337_2_lut (.A(u_l[4]), .B(\u_s[5] ), .Z(c_15__N_2408[4])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13337_2_lut.init = 16'h8888;
    LUT4 i13323_2_lut (.A(u_l[5]), .B(\u_s[4] ), .Z(c_15__N_2423[4])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13323_2_lut.init = 16'h8888;
    CCU2D add_823_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19463), 
          .S0(o_r_17__N_2438[17]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_823_cout.INIT0 = 16'h0000;
    defparam add_823_cout.INIT1 = 16'h0000;
    defparam add_823_cout.INJECT1_0 = "NO";
    defparam add_823_cout.INJECT1_1 = "NO";
    CCU2D add_823_15 (.A0(c_15__N_2408[14]), .B0(c_15__N_2423[14]), .C0(c_15__N_2408[13]), 
          .D0(c_15__N_2423[13]), .A1(u_l[15]), .B1(\u_s[5] ), .C1(c_15__N_2408[14]), 
          .D1(c_15__N_2423[14]), .CIN(n19462), .COUT(n19463), .S0(o_r_17__N_2438[15]), 
          .S1(o_r_17__N_2438[16]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_823_15.INIT0 = 16'h9666;
    defparam add_823_15.INIT1 = 16'h7888;
    defparam add_823_15.INJECT1_0 = "NO";
    defparam add_823_15.INJECT1_1 = "NO";
    CCU2D add_823_13 (.A0(c_15__N_2408[12]), .B0(c_15__N_2423[12]), .C0(c_15__N_2408[11]), 
          .D0(c_15__N_2423[11]), .A1(c_15__N_2408[13]), .B1(c_15__N_2423[13]), 
          .C1(c_15__N_2408[12]), .D1(c_15__N_2423[12]), .CIN(n19461), 
          .COUT(n19462), .S0(o_r_17__N_2438[13]), .S1(o_r_17__N_2438[14]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_823_13.INIT0 = 16'h9666;
    defparam add_823_13.INIT1 = 16'h9666;
    defparam add_823_13.INJECT1_0 = "NO";
    defparam add_823_13.INJECT1_1 = "NO";
    CCU2D add_823_11 (.A0(c_15__N_2408[10]), .B0(c_15__N_2423[10]), .C0(c_15__N_2408[9]), 
          .D0(c_15__N_2423[9]), .A1(c_15__N_2408[11]), .B1(c_15__N_2423[11]), 
          .C1(c_15__N_2408[10]), .D1(c_15__N_2423[10]), .CIN(n19460), 
          .COUT(n19461), .S0(o_r_17__N_2438[11]), .S1(o_r_17__N_2438[12]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_823_11.INIT0 = 16'h9666;
    defparam add_823_11.INIT1 = 16'h9666;
    defparam add_823_11.INJECT1_0 = "NO";
    defparam add_823_11.INJECT1_1 = "NO";
    CCU2D add_823_9 (.A0(c_15__N_2408[8]), .B0(c_15__N_2423[8]), .C0(c_15__N_2408[7]), 
          .D0(c_15__N_2423[7]), .A1(c_15__N_2408[9]), .B1(c_15__N_2423[9]), 
          .C1(c_15__N_2408[8]), .D1(c_15__N_2423[8]), .CIN(n19459), .COUT(n19460), 
          .S0(o_r_17__N_2438[9]), .S1(o_r_17__N_2438[10]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_823_9.INIT0 = 16'h9666;
    defparam add_823_9.INIT1 = 16'h9666;
    defparam add_823_9.INJECT1_0 = "NO";
    defparam add_823_9.INJECT1_1 = "NO";
    CCU2D add_823_7 (.A0(c_15__N_2408[6]), .B0(c_15__N_2423[6]), .C0(c_15__N_2408[5]), 
          .D0(c_15__N_2423[5]), .A1(c_15__N_2408[7]), .B1(c_15__N_2423[7]), 
          .C1(c_15__N_2408[6]), .D1(c_15__N_2423[6]), .CIN(n19458), .COUT(n19459), 
          .S0(o_r_17__N_2438[7]), .S1(o_r_17__N_2438[8]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_823_7.INIT0 = 16'h9666;
    defparam add_823_7.INIT1 = 16'h9666;
    defparam add_823_7.INJECT1_0 = "NO";
    defparam add_823_7.INJECT1_1 = "NO";
    CCU2D add_823_5 (.A0(c_15__N_2408[4]), .B0(c_15__N_2423[4]), .C0(c_15__N_2408[3]), 
          .D0(c_15__N_2423[3]), .A1(c_15__N_2408[5]), .B1(c_15__N_2423[5]), 
          .C1(c_15__N_2408[4]), .D1(c_15__N_2423[4]), .CIN(n19457), .COUT(n19458), 
          .S0(o_r_17__N_2438[5]), .S1(o_r_17__N_2438[6]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_823_5.INIT0 = 16'h9666;
    defparam add_823_5.INIT1 = 16'h9666;
    defparam add_823_5.INJECT1_0 = "NO";
    defparam add_823_5.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \bimpy(BW=16)_U11 
//

module \bimpy(BW=16)_U11  (S_0_01, dac_clk_p_c, n14231, n9454, u_l, 
            \u_s[3] , \u_s[2] , GND_net, i_sw0_c) /* synthesis syn_module_defined=1 */ ;
    output [17:0]S_0_01;
    input dac_clk_p_c;
    input n14231;
    input n9454;
    input [15:0]u_l;
    input \u_s[3] ;
    input \u_s[2] ;
    input GND_net;
    input i_sw0_c;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[29:38])
    wire [14:0]c_15__N_2408;
    wire [14:0]c_15__N_2423;
    
    wire n19471;
    wire [17:0]o_r_17__N_2438;
    
    wire n19470, n19469, n19468, n19467, n19466, n19465, n19464, 
        n29248, n29249;
    
    FD1S3IX o_r__i0 (.D(n9454), .CK(dac_clk_p_c), .CD(n14231), .Q(S_0_01[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=75, LSE_RLINE=75 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i0.GSR = "DISABLED";
    LUT4 i13356_2_lut (.A(u_l[14]), .B(\u_s[3] ), .Z(c_15__N_2408[14])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13356_2_lut.init = 16'h8888;
    LUT4 i13342_2_lut (.A(u_l[15]), .B(\u_s[2] ), .Z(c_15__N_2423[14])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13342_2_lut.init = 16'h8888;
    LUT4 i13357_2_lut (.A(u_l[13]), .B(\u_s[3] ), .Z(c_15__N_2408[13])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13357_2_lut.init = 16'h8888;
    LUT4 i13343_2_lut (.A(u_l[14]), .B(\u_s[2] ), .Z(c_15__N_2423[13])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13343_2_lut.init = 16'h8888;
    CCU2D add_824_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19471), 
          .S0(o_r_17__N_2438[17]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_824_cout.INIT0 = 16'h0000;
    defparam add_824_cout.INIT1 = 16'h0000;
    defparam add_824_cout.INJECT1_0 = "NO";
    defparam add_824_cout.INJECT1_1 = "NO";
    CCU2D add_824_15 (.A0(c_15__N_2408[14]), .B0(c_15__N_2423[14]), .C0(c_15__N_2408[13]), 
          .D0(c_15__N_2423[13]), .A1(u_l[15]), .B1(\u_s[3] ), .C1(c_15__N_2408[14]), 
          .D1(c_15__N_2423[14]), .CIN(n19470), .COUT(n19471), .S0(o_r_17__N_2438[15]), 
          .S1(o_r_17__N_2438[16]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_824_15.INIT0 = 16'h9666;
    defparam add_824_15.INIT1 = 16'h7888;
    defparam add_824_15.INJECT1_0 = "NO";
    defparam add_824_15.INJECT1_1 = "NO";
    CCU2D add_824_13 (.A0(c_15__N_2408[12]), .B0(c_15__N_2423[12]), .C0(c_15__N_2408[11]), 
          .D0(c_15__N_2423[11]), .A1(c_15__N_2408[13]), .B1(c_15__N_2423[13]), 
          .C1(c_15__N_2408[12]), .D1(c_15__N_2423[12]), .CIN(n19469), 
          .COUT(n19470), .S0(o_r_17__N_2438[13]), .S1(o_r_17__N_2438[14]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_824_13.INIT0 = 16'h9666;
    defparam add_824_13.INIT1 = 16'h9666;
    defparam add_824_13.INJECT1_0 = "NO";
    defparam add_824_13.INJECT1_1 = "NO";
    CCU2D add_824_11 (.A0(c_15__N_2408[10]), .B0(c_15__N_2423[10]), .C0(c_15__N_2408[9]), 
          .D0(c_15__N_2423[9]), .A1(c_15__N_2408[11]), .B1(c_15__N_2423[11]), 
          .C1(c_15__N_2408[10]), .D1(c_15__N_2423[10]), .CIN(n19468), 
          .COUT(n19469), .S0(o_r_17__N_2438[11]), .S1(o_r_17__N_2438[12]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_824_11.INIT0 = 16'h9666;
    defparam add_824_11.INIT1 = 16'h9666;
    defparam add_824_11.INJECT1_0 = "NO";
    defparam add_824_11.INJECT1_1 = "NO";
    CCU2D add_824_9 (.A0(c_15__N_2408[8]), .B0(c_15__N_2423[8]), .C0(c_15__N_2408[7]), 
          .D0(c_15__N_2423[7]), .A1(c_15__N_2408[9]), .B1(c_15__N_2423[9]), 
          .C1(c_15__N_2408[8]), .D1(c_15__N_2423[8]), .CIN(n19467), .COUT(n19468), 
          .S0(o_r_17__N_2438[9]), .S1(o_r_17__N_2438[10]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_824_9.INIT0 = 16'h9666;
    defparam add_824_9.INIT1 = 16'h9666;
    defparam add_824_9.INJECT1_0 = "NO";
    defparam add_824_9.INJECT1_1 = "NO";
    CCU2D add_824_7 (.A0(c_15__N_2408[6]), .B0(c_15__N_2423[6]), .C0(c_15__N_2408[5]), 
          .D0(c_15__N_2423[5]), .A1(c_15__N_2408[7]), .B1(c_15__N_2423[7]), 
          .C1(c_15__N_2408[6]), .D1(c_15__N_2423[6]), .CIN(n19466), .COUT(n19467), 
          .S0(o_r_17__N_2438[7]), .S1(o_r_17__N_2438[8]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_824_7.INIT0 = 16'h9666;
    defparam add_824_7.INIT1 = 16'h9666;
    defparam add_824_7.INJECT1_0 = "NO";
    defparam add_824_7.INJECT1_1 = "NO";
    CCU2D add_824_5 (.A0(c_15__N_2408[4]), .B0(c_15__N_2423[4]), .C0(c_15__N_2408[3]), 
          .D0(c_15__N_2423[3]), .A1(c_15__N_2408[5]), .B1(c_15__N_2423[5]), 
          .C1(c_15__N_2408[4]), .D1(c_15__N_2423[4]), .CIN(n19465), .COUT(n19466), 
          .S0(o_r_17__N_2438[5]), .S1(o_r_17__N_2438[6]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_824_5.INIT0 = 16'h9666;
    defparam add_824_5.INIT1 = 16'h9666;
    defparam add_824_5.INJECT1_0 = "NO";
    defparam add_824_5.INJECT1_1 = "NO";
    LUT4 i13358_2_lut (.A(u_l[12]), .B(\u_s[3] ), .Z(c_15__N_2408[12])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13358_2_lut.init = 16'h8888;
    LUT4 i13344_2_lut (.A(u_l[13]), .B(\u_s[2] ), .Z(c_15__N_2423[12])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13344_2_lut.init = 16'h8888;
    LUT4 i13359_2_lut (.A(u_l[11]), .B(\u_s[3] ), .Z(c_15__N_2408[11])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13359_2_lut.init = 16'h8888;
    LUT4 i13345_2_lut (.A(u_l[12]), .B(\u_s[2] ), .Z(c_15__N_2423[11])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13345_2_lut.init = 16'h8888;
    LUT4 i13360_2_lut (.A(u_l[10]), .B(\u_s[3] ), .Z(c_15__N_2408[10])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13360_2_lut.init = 16'h8888;
    LUT4 i13346_2_lut (.A(u_l[11]), .B(\u_s[2] ), .Z(c_15__N_2423[10])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13346_2_lut.init = 16'h8888;
    LUT4 i13361_2_lut (.A(u_l[9]), .B(\u_s[3] ), .Z(c_15__N_2408[9])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13361_2_lut.init = 16'h8888;
    LUT4 i13347_2_lut (.A(u_l[10]), .B(\u_s[2] ), .Z(c_15__N_2423[9])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13347_2_lut.init = 16'h8888;
    LUT4 i13362_2_lut (.A(u_l[8]), .B(\u_s[3] ), .Z(c_15__N_2408[8])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13362_2_lut.init = 16'h8888;
    LUT4 i13348_2_lut (.A(u_l[9]), .B(\u_s[2] ), .Z(c_15__N_2423[8])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13348_2_lut.init = 16'h8888;
    LUT4 i13363_2_lut (.A(u_l[7]), .B(\u_s[3] ), .Z(c_15__N_2408[7])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13363_2_lut.init = 16'h8888;
    LUT4 i13349_2_lut (.A(u_l[8]), .B(\u_s[2] ), .Z(c_15__N_2423[7])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13349_2_lut.init = 16'h8888;
    LUT4 i13364_2_lut (.A(u_l[6]), .B(\u_s[3] ), .Z(c_15__N_2408[6])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13364_2_lut.init = 16'h8888;
    LUT4 i13350_2_lut (.A(u_l[7]), .B(\u_s[2] ), .Z(c_15__N_2423[6])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13350_2_lut.init = 16'h8888;
    LUT4 i13365_2_lut (.A(u_l[5]), .B(\u_s[3] ), .Z(c_15__N_2408[5])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13365_2_lut.init = 16'h8888;
    LUT4 i13351_2_lut (.A(u_l[6]), .B(\u_s[2] ), .Z(c_15__N_2423[5])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13351_2_lut.init = 16'h8888;
    LUT4 i13366_2_lut (.A(u_l[4]), .B(\u_s[3] ), .Z(c_15__N_2408[4])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13366_2_lut.init = 16'h8888;
    LUT4 i13352_2_lut (.A(u_l[5]), .B(\u_s[2] ), .Z(c_15__N_2423[4])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13352_2_lut.init = 16'h8888;
    CCU2D add_824_3 (.A0(c_15__N_2408[2]), .B0(c_15__N_2423[2]), .C0(c_15__N_2408[1]), 
          .D0(c_15__N_2423[1]), .A1(c_15__N_2408[3]), .B1(c_15__N_2423[3]), 
          .C1(c_15__N_2408[2]), .D1(c_15__N_2423[2]), .CIN(n19464), .COUT(n19465), 
          .S0(o_r_17__N_2438[3]), .S1(o_r_17__N_2438[4]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_824_3.INIT0 = 16'h9666;
    defparam add_824_3.INIT1 = 16'h9666;
    defparam add_824_3.INJECT1_0 = "NO";
    defparam add_824_3.INJECT1_1 = "NO";
    FD1S3IX o_r__i17 (.D(o_r_17__N_2438[17]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_01[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=75, LSE_RLINE=75 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i17.GSR = "DISABLED";
    LUT4 i13367_2_lut (.A(u_l[3]), .B(\u_s[3] ), .Z(c_15__N_2408[3])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13367_2_lut.init = 16'h8888;
    LUT4 i13353_2_lut (.A(u_l[4]), .B(\u_s[2] ), .Z(c_15__N_2423[3])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13353_2_lut.init = 16'h8888;
    FD1S3IX o_r__i16 (.D(o_r_17__N_2438[16]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_01[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=75, LSE_RLINE=75 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i16.GSR = "DISABLED";
    FD1S3IX o_r__i15 (.D(o_r_17__N_2438[15]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_01[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=75, LSE_RLINE=75 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i15.GSR = "DISABLED";
    FD1S3IX o_r__i14 (.D(o_r_17__N_2438[14]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_01[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=75, LSE_RLINE=75 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i14.GSR = "DISABLED";
    FD1S3IX o_r__i13 (.D(o_r_17__N_2438[13]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_01[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=75, LSE_RLINE=75 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i13.GSR = "DISABLED";
    FD1S3IX o_r__i12 (.D(o_r_17__N_2438[12]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_01[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=75, LSE_RLINE=75 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i12.GSR = "DISABLED";
    FD1S3IX o_r__i11 (.D(o_r_17__N_2438[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_01[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=75, LSE_RLINE=75 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i11.GSR = "DISABLED";
    FD1S3IX o_r__i10 (.D(o_r_17__N_2438[10]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_01[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=75, LSE_RLINE=75 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i10.GSR = "DISABLED";
    FD1S3IX o_r__i9 (.D(o_r_17__N_2438[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_01[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=75, LSE_RLINE=75 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i9.GSR = "DISABLED";
    FD1S3IX o_r__i8 (.D(o_r_17__N_2438[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_01[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=75, LSE_RLINE=75 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i8.GSR = "DISABLED";
    FD1S3IX o_r__i7 (.D(o_r_17__N_2438[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_01[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=75, LSE_RLINE=75 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i7.GSR = "DISABLED";
    FD1S3IX o_r__i6 (.D(o_r_17__N_2438[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_01[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=75, LSE_RLINE=75 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i6.GSR = "DISABLED";
    FD1S3IX o_r__i5 (.D(o_r_17__N_2438[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_01[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=75, LSE_RLINE=75 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i5.GSR = "DISABLED";
    FD1S3IX o_r__i4 (.D(o_r_17__N_2438[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_01[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=75, LSE_RLINE=75 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i4.GSR = "DISABLED";
    FD1S3IX o_r__i3 (.D(o_r_17__N_2438[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_01[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=75, LSE_RLINE=75 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i3.GSR = "DISABLED";
    FD1S3IX o_r__i2 (.D(o_r_17__N_2438[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_01[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=75, LSE_RLINE=75 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i2.GSR = "DISABLED";
    FD1S3IX o_r__i1 (.D(o_r_17__N_2438[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_01[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=75, LSE_RLINE=75 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i1.GSR = "DISABLED";
    LUT4 i13368_2_lut (.A(u_l[2]), .B(\u_s[3] ), .Z(c_15__N_2408[2])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13368_2_lut.init = 16'h8888;
    LUT4 i13354_2_lut (.A(u_l[3]), .B(\u_s[2] ), .Z(c_15__N_2423[2])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13354_2_lut.init = 16'h8888;
    LUT4 i13369_2_lut (.A(u_l[1]), .B(\u_s[3] ), .Z(c_15__N_2408[1])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13369_2_lut.init = 16'h8888;
    LUT4 i13355_2_lut (.A(u_l[2]), .B(\u_s[2] ), .Z(c_15__N_2423[1])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13355_2_lut.init = 16'h8888;
    LUT4 i12505_2_lut_rep_588 (.A(u_l[1]), .B(\u_s[2] ), .Z(n29248)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i12505_2_lut_rep_588.init = 16'h8888;
    LUT4 i12504_2_lut_rep_589 (.A(u_l[0]), .B(\u_s[3] ), .Z(n29249)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(51[18:45])
    defparam i12504_2_lut_rep_589.init = 16'h8888;
    LUT4 w_r_16__I_0_i2_2_lut_3_lut_4_lut (.A(u_l[0]), .B(\u_s[3] ), .C(\u_s[2] ), 
         .D(u_l[1]), .Z(o_r_17__N_2438[1])) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(51[18:45])
    defparam w_r_16__I_0_i2_2_lut_3_lut_4_lut.init = 16'h7888;
    CCU2D add_824_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(c_15__N_2408[1]), .B1(c_15__N_2423[1]), .C1(n29249), .D1(n29248), 
          .COUT(n19464), .S1(o_r_17__N_2438[2]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_824_1.INIT0 = 16'hF000;
    defparam add_824_1.INIT1 = 16'h9666;
    defparam add_824_1.INJECT1_0 = "NO";
    defparam add_824_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \bimpy(BW=16)_U12 
//

module \bimpy(BW=16)_U12  (\S_0_00[0] , dac_clk_p_c, n14231, n9456, 
            u_l, \u_s[1] , \u_s[0] , GND_net, \S_0_00[17] , i_sw0_c, 
            \S_0_00[16] , \S_0_00[15] , \S_0_00[14] , \S_0_00[13] , 
            \S_0_00[12] , \S_0_00[11] , \S_0_00[10] , \S_0_00[9] , \S_0_00[8] , 
            \S_0_00[7] , \S_0_00[6] , \S_0_00[5] , \S_0_00[4] , \S_0_00[3] , 
            \S_0_00[2] , \S_1_00_20__N_2184[1] ) /* synthesis syn_module_defined=1 */ ;
    output \S_0_00[0] ;
    input dac_clk_p_c;
    input n14231;
    input n9456;
    input [15:0]u_l;
    input \u_s[1] ;
    input \u_s[0] ;
    input GND_net;
    output \S_0_00[17] ;
    input i_sw0_c;
    output \S_0_00[16] ;
    output \S_0_00[15] ;
    output \S_0_00[14] ;
    output \S_0_00[13] ;
    output \S_0_00[12] ;
    output \S_0_00[11] ;
    output \S_0_00[10] ;
    output \S_0_00[9] ;
    output \S_0_00[8] ;
    output \S_0_00[7] ;
    output \S_0_00[6] ;
    output \S_0_00[5] ;
    output \S_0_00[4] ;
    output \S_0_00[3] ;
    output \S_0_00[2] ;
    output \S_1_00_20__N_2184[1] ;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[29:38])
    wire [14:0]c_15__N_2408;
    wire [14:0]c_15__N_2423;
    
    wire n19479;
    wire [17:0]o_r_17__N_2438;
    
    wire n19478, n19477, n19476, n19475, n19474, n19473, n19472, 
        n29263, n29262;
    
    FD1S3IX o_r__i0 (.D(n9456), .CK(dac_clk_p_c), .CD(n14231), .Q(\S_0_00[0] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i0.GSR = "DISABLED";
    LUT4 i13390_2_lut (.A(u_l[12]), .B(\u_s[1] ), .Z(c_15__N_2408[12])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13390_2_lut.init = 16'h8888;
    LUT4 i13375_2_lut (.A(u_l[13]), .B(\u_s[0] ), .Z(c_15__N_2423[12])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13375_2_lut.init = 16'h8888;
    LUT4 i13391_2_lut (.A(u_l[11]), .B(\u_s[1] ), .Z(c_15__N_2408[11])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13391_2_lut.init = 16'h8888;
    LUT4 i13376_2_lut (.A(u_l[12]), .B(\u_s[0] ), .Z(c_15__N_2423[11])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13376_2_lut.init = 16'h8888;
    LUT4 i13392_2_lut (.A(u_l[10]), .B(\u_s[1] ), .Z(c_15__N_2408[10])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13392_2_lut.init = 16'h8888;
    LUT4 i13377_2_lut (.A(u_l[11]), .B(\u_s[0] ), .Z(c_15__N_2423[10])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13377_2_lut.init = 16'h8888;
    LUT4 i13393_2_lut (.A(u_l[9]), .B(\u_s[1] ), .Z(c_15__N_2408[9])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13393_2_lut.init = 16'h8888;
    LUT4 i13378_2_lut (.A(u_l[10]), .B(\u_s[0] ), .Z(c_15__N_2423[9])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13378_2_lut.init = 16'h8888;
    LUT4 i13394_2_lut (.A(u_l[8]), .B(\u_s[1] ), .Z(c_15__N_2408[8])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13394_2_lut.init = 16'h8888;
    LUT4 i13379_2_lut (.A(u_l[9]), .B(\u_s[0] ), .Z(c_15__N_2423[8])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13379_2_lut.init = 16'h8888;
    LUT4 i13395_2_lut (.A(u_l[7]), .B(\u_s[1] ), .Z(c_15__N_2408[7])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13395_2_lut.init = 16'h8888;
    LUT4 i13380_2_lut (.A(u_l[8]), .B(\u_s[0] ), .Z(c_15__N_2423[7])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13380_2_lut.init = 16'h8888;
    LUT4 i13396_2_lut (.A(u_l[6]), .B(\u_s[1] ), .Z(c_15__N_2408[6])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13396_2_lut.init = 16'h8888;
    LUT4 i13381_2_lut (.A(u_l[7]), .B(\u_s[0] ), .Z(c_15__N_2423[6])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13381_2_lut.init = 16'h8888;
    LUT4 i13397_2_lut (.A(u_l[5]), .B(\u_s[1] ), .Z(c_15__N_2408[5])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13397_2_lut.init = 16'h8888;
    LUT4 i13382_2_lut (.A(u_l[6]), .B(\u_s[0] ), .Z(c_15__N_2423[5])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13382_2_lut.init = 16'h8888;
    LUT4 i13398_2_lut (.A(u_l[4]), .B(\u_s[1] ), .Z(c_15__N_2408[4])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13398_2_lut.init = 16'h8888;
    LUT4 i13383_2_lut (.A(u_l[5]), .B(\u_s[0] ), .Z(c_15__N_2423[4])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13383_2_lut.init = 16'h8888;
    LUT4 i13399_2_lut (.A(u_l[3]), .B(\u_s[1] ), .Z(c_15__N_2408[3])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13399_2_lut.init = 16'h8888;
    LUT4 i13384_2_lut (.A(u_l[4]), .B(\u_s[0] ), .Z(c_15__N_2423[3])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13384_2_lut.init = 16'h8888;
    LUT4 i13400_2_lut (.A(u_l[2]), .B(\u_s[1] ), .Z(c_15__N_2408[2])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13400_2_lut.init = 16'h8888;
    LUT4 i13386_2_lut (.A(u_l[3]), .B(\u_s[0] ), .Z(c_15__N_2423[2])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13386_2_lut.init = 16'h8888;
    LUT4 i13401_2_lut (.A(u_l[1]), .B(\u_s[1] ), .Z(c_15__N_2408[1])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13401_2_lut.init = 16'h8888;
    LUT4 i13387_2_lut (.A(u_l[2]), .B(\u_s[0] ), .Z(c_15__N_2423[1])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13387_2_lut.init = 16'h8888;
    CCU2D add_825_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19479), 
          .S0(o_r_17__N_2438[17]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_825_cout.INIT0 = 16'h0000;
    defparam add_825_cout.INIT1 = 16'h0000;
    defparam add_825_cout.INJECT1_0 = "NO";
    defparam add_825_cout.INJECT1_1 = "NO";
    CCU2D add_825_15 (.A0(c_15__N_2408[14]), .B0(c_15__N_2423[14]), .C0(c_15__N_2408[13]), 
          .D0(c_15__N_2423[13]), .A1(u_l[15]), .B1(\u_s[1] ), .C1(c_15__N_2408[14]), 
          .D1(c_15__N_2423[14]), .CIN(n19478), .COUT(n19479), .S0(o_r_17__N_2438[15]), 
          .S1(o_r_17__N_2438[16]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_825_15.INIT0 = 16'h9666;
    defparam add_825_15.INIT1 = 16'h7888;
    defparam add_825_15.INJECT1_0 = "NO";
    defparam add_825_15.INJECT1_1 = "NO";
    CCU2D add_825_13 (.A0(c_15__N_2408[12]), .B0(c_15__N_2423[12]), .C0(c_15__N_2408[11]), 
          .D0(c_15__N_2423[11]), .A1(c_15__N_2408[13]), .B1(c_15__N_2423[13]), 
          .C1(c_15__N_2408[12]), .D1(c_15__N_2423[12]), .CIN(n19477), 
          .COUT(n19478), .S0(o_r_17__N_2438[13]), .S1(o_r_17__N_2438[14]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_825_13.INIT0 = 16'h9666;
    defparam add_825_13.INIT1 = 16'h9666;
    defparam add_825_13.INJECT1_0 = "NO";
    defparam add_825_13.INJECT1_1 = "NO";
    CCU2D add_825_11 (.A0(c_15__N_2408[10]), .B0(c_15__N_2423[10]), .C0(c_15__N_2408[9]), 
          .D0(c_15__N_2423[9]), .A1(c_15__N_2408[11]), .B1(c_15__N_2423[11]), 
          .C1(c_15__N_2408[10]), .D1(c_15__N_2423[10]), .CIN(n19476), 
          .COUT(n19477), .S0(o_r_17__N_2438[11]), .S1(o_r_17__N_2438[12]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_825_11.INIT0 = 16'h9666;
    defparam add_825_11.INIT1 = 16'h9666;
    defparam add_825_11.INJECT1_0 = "NO";
    defparam add_825_11.INJECT1_1 = "NO";
    CCU2D add_825_9 (.A0(c_15__N_2408[8]), .B0(c_15__N_2423[8]), .C0(c_15__N_2408[7]), 
          .D0(c_15__N_2423[7]), .A1(c_15__N_2408[9]), .B1(c_15__N_2423[9]), 
          .C1(c_15__N_2408[8]), .D1(c_15__N_2423[8]), .CIN(n19475), .COUT(n19476), 
          .S0(o_r_17__N_2438[9]), .S1(o_r_17__N_2438[10]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_825_9.INIT0 = 16'h9666;
    defparam add_825_9.INIT1 = 16'h9666;
    defparam add_825_9.INJECT1_0 = "NO";
    defparam add_825_9.INJECT1_1 = "NO";
    CCU2D add_825_7 (.A0(c_15__N_2408[6]), .B0(c_15__N_2423[6]), .C0(c_15__N_2408[5]), 
          .D0(c_15__N_2423[5]), .A1(c_15__N_2408[7]), .B1(c_15__N_2423[7]), 
          .C1(c_15__N_2408[6]), .D1(c_15__N_2423[6]), .CIN(n19474), .COUT(n19475), 
          .S0(o_r_17__N_2438[7]), .S1(o_r_17__N_2438[8]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_825_7.INIT0 = 16'h9666;
    defparam add_825_7.INIT1 = 16'h9666;
    defparam add_825_7.INJECT1_0 = "NO";
    defparam add_825_7.INJECT1_1 = "NO";
    CCU2D add_825_5 (.A0(c_15__N_2408[4]), .B0(c_15__N_2423[4]), .C0(c_15__N_2408[3]), 
          .D0(c_15__N_2423[3]), .A1(c_15__N_2408[5]), .B1(c_15__N_2423[5]), 
          .C1(c_15__N_2408[4]), .D1(c_15__N_2423[4]), .CIN(n19473), .COUT(n19474), 
          .S0(o_r_17__N_2438[5]), .S1(o_r_17__N_2438[6]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_825_5.INIT0 = 16'h9666;
    defparam add_825_5.INIT1 = 16'h9666;
    defparam add_825_5.INJECT1_0 = "NO";
    defparam add_825_5.INJECT1_1 = "NO";
    CCU2D add_825_3 (.A0(c_15__N_2408[2]), .B0(c_15__N_2423[2]), .C0(c_15__N_2408[1]), 
          .D0(c_15__N_2423[1]), .A1(c_15__N_2408[3]), .B1(c_15__N_2423[3]), 
          .C1(c_15__N_2408[2]), .D1(c_15__N_2423[2]), .CIN(n19472), .COUT(n19473), 
          .S0(o_r_17__N_2438[3]), .S1(o_r_17__N_2438[4]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_825_3.INIT0 = 16'h9666;
    defparam add_825_3.INIT1 = 16'h9666;
    defparam add_825_3.INJECT1_0 = "NO";
    defparam add_825_3.INJECT1_1 = "NO";
    CCU2D add_825_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(c_15__N_2408[1]), .B1(c_15__N_2423[1]), .C1(n29263), .D1(n29262), 
          .COUT(n19472), .S1(o_r_17__N_2438[2]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_825_1.INIT0 = 16'hF000;
    defparam add_825_1.INIT1 = 16'h9666;
    defparam add_825_1.INJECT1_0 = "NO";
    defparam add_825_1.INJECT1_1 = "NO";
    LUT4 i13388_2_lut (.A(u_l[14]), .B(\u_s[1] ), .Z(c_15__N_2408[14])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13388_2_lut.init = 16'h8888;
    LUT4 i13373_2_lut (.A(u_l[15]), .B(\u_s[0] ), .Z(c_15__N_2423[14])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13373_2_lut.init = 16'h8888;
    LUT4 i13389_2_lut (.A(u_l[13]), .B(\u_s[1] ), .Z(c_15__N_2408[13])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13389_2_lut.init = 16'h8888;
    LUT4 i13374_2_lut (.A(u_l[14]), .B(\u_s[0] ), .Z(c_15__N_2423[13])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13374_2_lut.init = 16'h8888;
    FD1S3IX o_r__i17 (.D(o_r_17__N_2438[17]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_00[17] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i17.GSR = "DISABLED";
    FD1S3IX o_r__i16 (.D(o_r_17__N_2438[16]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_00[16] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i16.GSR = "DISABLED";
    FD1S3IX o_r__i15 (.D(o_r_17__N_2438[15]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_00[15] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i15.GSR = "DISABLED";
    FD1S3IX o_r__i14 (.D(o_r_17__N_2438[14]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_00[14] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i14.GSR = "DISABLED";
    FD1S3IX o_r__i13 (.D(o_r_17__N_2438[13]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_00[13] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i13.GSR = "DISABLED";
    FD1S3IX o_r__i12 (.D(o_r_17__N_2438[12]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_00[12] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i12.GSR = "DISABLED";
    FD1S3IX o_r__i11 (.D(o_r_17__N_2438[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_00[11] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i11.GSR = "DISABLED";
    FD1S3IX o_r__i10 (.D(o_r_17__N_2438[10]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_00[10] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i10.GSR = "DISABLED";
    FD1S3IX o_r__i9 (.D(o_r_17__N_2438[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_00[9] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i9.GSR = "DISABLED";
    FD1S3IX o_r__i8 (.D(o_r_17__N_2438[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_00[8] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i8.GSR = "DISABLED";
    FD1S3IX o_r__i7 (.D(o_r_17__N_2438[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_00[7] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i7.GSR = "DISABLED";
    FD1S3IX o_r__i6 (.D(o_r_17__N_2438[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_00[6] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i6.GSR = "DISABLED";
    FD1S3IX o_r__i5 (.D(o_r_17__N_2438[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_00[5] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i5.GSR = "DISABLED";
    FD1S3IX o_r__i4 (.D(o_r_17__N_2438[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_00[4] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i4.GSR = "DISABLED";
    FD1S3IX o_r__i3 (.D(o_r_17__N_2438[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_00[3] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i3.GSR = "DISABLED";
    FD1S3IX o_r__i2 (.D(o_r_17__N_2438[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_00[2] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i2.GSR = "DISABLED";
    FD1S3IX o_r__i1 (.D(o_r_17__N_2438[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_1_00_20__N_2184[1] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i1.GSR = "DISABLED";
    LUT4 i12503_2_lut_rep_602 (.A(u_l[1]), .B(\u_s[0] ), .Z(n29262)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i12503_2_lut_rep_602.init = 16'h8888;
    LUT4 i12502_2_lut_rep_603 (.A(u_l[0]), .B(\u_s[1] ), .Z(n29263)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(51[18:45])
    defparam i12502_2_lut_rep_603.init = 16'h8888;
    LUT4 w_r_16__I_0_i2_2_lut_3_lut_4_lut (.A(u_l[0]), .B(\u_s[1] ), .C(\u_s[0] ), 
         .D(u_l[1]), .Z(o_r_17__N_2438[1])) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(51[18:45])
    defparam w_r_16__I_0_i2_2_lut_3_lut_4_lut.init = 16'h7888;
    
endmodule
//
// Verilog Description of module dds
//

module dds (dac_clk_p_c, i_sw0_c, \addr_space[1][0] , \addr_space[1][30] , 
            \addr_space[1][29] , \addr_space[1][28] , \addr_space[1][27] , 
            \addr_space[1][26] , \addr_space[1][25] , \addr_space[1][24] , 
            \addr_space[1][23] , \addr_space[1][22] , \addr_space[1][21] , 
            \addr_space[1][20] , \addr_space[1][19] , \addr_space[1][18] , 
            \addr_space[1][17] , \addr_space[1][16] , \addr_space[1][15] , 
            \addr_space[1][14] , \addr_space[1][13] , \addr_space[1][12] , 
            \addr_space[1][11] , \addr_space[1][10] , \addr_space[1][9] , 
            \addr_space[1][8] , \addr_space[1][7] , \addr_space[1][6] , 
            \addr_space[1][5] , \addr_space[1][4] , \addr_space[1][3] , 
            \addr_space[1][2] , \addr_space[1][1] , dac_clk_p_c_enable_630, 
            modulation_output, \quarter_wave_sample_register_i[15] , GND_net) /* synthesis syn_module_defined=1 */ ;
    input dac_clk_p_c;
    input i_sw0_c;
    input \addr_space[1][0] ;
    input \addr_space[1][30] ;
    input \addr_space[1][29] ;
    input \addr_space[1][28] ;
    input \addr_space[1][27] ;
    input \addr_space[1][26] ;
    input \addr_space[1][25] ;
    input \addr_space[1][24] ;
    input \addr_space[1][23] ;
    input \addr_space[1][22] ;
    input \addr_space[1][21] ;
    input \addr_space[1][20] ;
    input \addr_space[1][19] ;
    input \addr_space[1][18] ;
    input \addr_space[1][17] ;
    input \addr_space[1][16] ;
    input \addr_space[1][15] ;
    input \addr_space[1][14] ;
    input \addr_space[1][13] ;
    input \addr_space[1][12] ;
    input \addr_space[1][11] ;
    input \addr_space[1][10] ;
    input \addr_space[1][9] ;
    input \addr_space[1][8] ;
    input \addr_space[1][7] ;
    input \addr_space[1][6] ;
    input \addr_space[1][5] ;
    input \addr_space[1][4] ;
    input \addr_space[1][3] ;
    input \addr_space[1][2] ;
    input \addr_space[1][1] ;
    input dac_clk_p_c_enable_630;
    output [15:0]modulation_output;
    input \quarter_wave_sample_register_i[15] ;
    input GND_net;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[29:38])
    wire [15:0]modulation_output_c /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(86[39:56])
    wire [30:0]increment;   // d:/documents/git_local/fm_modulator/rtl/dds.v(14[31:40])
    wire [11:0]o_phase;   // d:/documents/git_local/fm_modulator/rtl/dds.v(18[26:33])
    
    FD1S3DX increment_i0 (.D(\addr_space[1][0] ), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[0])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=96, LSE_RLINE=96 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i0.GSR = "DISABLED";
    FD1S3DX increment_i30 (.D(\addr_space[1][30] ), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[30])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=96, LSE_RLINE=96 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i30.GSR = "DISABLED";
    FD1S3DX increment_i29 (.D(\addr_space[1][29] ), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[29])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=96, LSE_RLINE=96 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i29.GSR = "DISABLED";
    FD1S3DX increment_i28 (.D(\addr_space[1][28] ), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[28])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=96, LSE_RLINE=96 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i28.GSR = "DISABLED";
    FD1S3DX increment_i27 (.D(\addr_space[1][27] ), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[27])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=96, LSE_RLINE=96 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i27.GSR = "DISABLED";
    FD1S3DX increment_i26 (.D(\addr_space[1][26] ), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[26])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=96, LSE_RLINE=96 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i26.GSR = "DISABLED";
    FD1S3DX increment_i25 (.D(\addr_space[1][25] ), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[25])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=96, LSE_RLINE=96 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i25.GSR = "DISABLED";
    FD1S3DX increment_i24 (.D(\addr_space[1][24] ), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[24])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=96, LSE_RLINE=96 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i24.GSR = "DISABLED";
    FD1S3DX increment_i23 (.D(\addr_space[1][23] ), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[23])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=96, LSE_RLINE=96 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i23.GSR = "DISABLED";
    FD1S3DX increment_i22 (.D(\addr_space[1][22] ), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[22])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=96, LSE_RLINE=96 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i22.GSR = "DISABLED";
    FD1S3DX increment_i21 (.D(\addr_space[1][21] ), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[21])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=96, LSE_RLINE=96 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i21.GSR = "DISABLED";
    FD1S3DX increment_i20 (.D(\addr_space[1][20] ), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[20])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=96, LSE_RLINE=96 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i20.GSR = "DISABLED";
    FD1S3DX increment_i19 (.D(\addr_space[1][19] ), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[19])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=96, LSE_RLINE=96 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i19.GSR = "DISABLED";
    FD1S3DX increment_i18 (.D(\addr_space[1][18] ), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[18])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=96, LSE_RLINE=96 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i18.GSR = "DISABLED";
    FD1S3DX increment_i17 (.D(\addr_space[1][17] ), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[17])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=96, LSE_RLINE=96 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i17.GSR = "DISABLED";
    FD1S3DX increment_i16 (.D(\addr_space[1][16] ), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[16])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=96, LSE_RLINE=96 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i16.GSR = "DISABLED";
    FD1S3DX increment_i15 (.D(\addr_space[1][15] ), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[15])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=96, LSE_RLINE=96 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i15.GSR = "DISABLED";
    FD1S3DX increment_i14 (.D(\addr_space[1][14] ), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[14])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=96, LSE_RLINE=96 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i14.GSR = "DISABLED";
    FD1S3DX increment_i13 (.D(\addr_space[1][13] ), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[13])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=96, LSE_RLINE=96 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i13.GSR = "DISABLED";
    FD1S3DX increment_i12 (.D(\addr_space[1][12] ), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[12])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=96, LSE_RLINE=96 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i12.GSR = "DISABLED";
    FD1S3DX increment_i11 (.D(\addr_space[1][11] ), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[11])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=96, LSE_RLINE=96 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i11.GSR = "DISABLED";
    FD1S3DX increment_i10 (.D(\addr_space[1][10] ), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[10])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=96, LSE_RLINE=96 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i10.GSR = "DISABLED";
    FD1S3DX increment_i9 (.D(\addr_space[1][9] ), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[9])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=96, LSE_RLINE=96 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i9.GSR = "DISABLED";
    FD1S3DX increment_i8 (.D(\addr_space[1][8] ), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[8])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=96, LSE_RLINE=96 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i8.GSR = "DISABLED";
    FD1S3DX increment_i7 (.D(\addr_space[1][7] ), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[7])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=96, LSE_RLINE=96 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i7.GSR = "DISABLED";
    FD1S3DX increment_i6 (.D(\addr_space[1][6] ), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[6])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=96, LSE_RLINE=96 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i6.GSR = "DISABLED";
    FD1S3DX increment_i5 (.D(\addr_space[1][5] ), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[5])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=96, LSE_RLINE=96 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i5.GSR = "DISABLED";
    FD1S3DX increment_i4 (.D(\addr_space[1][4] ), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[4])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=96, LSE_RLINE=96 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i4.GSR = "DISABLED";
    FD1S3DX increment_i3 (.D(\addr_space[1][3] ), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[3])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=96, LSE_RLINE=96 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i3.GSR = "DISABLED";
    FD1S3DX increment_i2 (.D(\addr_space[1][2] ), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[2])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=96, LSE_RLINE=96 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i2.GSR = "DISABLED";
    FD1S3DX increment_i1 (.D(\addr_space[1][1] ), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[1])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=96, LSE_RLINE=96 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i1.GSR = "DISABLED";
    quarter_wave_sine_lookup qtr_inst (.dac_clk_p_c(dac_clk_p_c), .dac_clk_p_c_enable_630(dac_clk_p_c_enable_630), 
            .o_phase({o_phase}), .i_sw0_c(i_sw0_c), .modulation_output({modulation_output}), 
            .\quarter_wave_sample_register_i[15] (\quarter_wave_sample_register_i[15] ), 
            .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(21[70:134])
    \nco(OW=12)  nco_inst (.increment({increment}), .GND_net(GND_net), .o_phase({o_phase}), 
            .dac_clk_p_c(dac_clk_p_c), .i_sw0_c(i_sw0_c)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(20[49:100])
    
endmodule
//
// Verilog Description of module quarter_wave_sine_lookup
//

module quarter_wave_sine_lookup (dac_clk_p_c, dac_clk_p_c_enable_630, o_phase, 
            i_sw0_c, modulation_output, \quarter_wave_sample_register_i[15] , 
            GND_net) /* synthesis syn_module_defined=1 */ ;
    input dac_clk_p_c;
    input dac_clk_p_c_enable_630;
    input [11:0]o_phase;
    input i_sw0_c;
    output [15:0]modulation_output;
    input \quarter_wave_sample_register_i[15] ;
    input GND_net;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[29:38])
    wire [15:0]modulation_output_c /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(86[39:56])
    wire [15:0]\o_val_pipeline_i[0]  /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(15[24:40])
    wire [9:0]index_i;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(31[17:24])
    
    wire n844, n24561, n24562, n24577, n24563, n24564, n24578, 
        n24929, n24930, n24937, n24565, n24566, n24579, n26586, 
        n29221, n26587, n24567, n24568, n24580, n24935, n24936, 
        n24940, n24569, n24570, n24581, n24573, n24574, n24583, 
        n23575, n23576, n23577, n23578, n23579, n23580, n23581, 
        n23582, n23583, n23584, n23585, n23586, n24592, n24593, 
        n24608, n24594, n24595, n24609, n24596, n24597, n24610, 
        n23590, n23591, n23592, n24600, n24601, n24612, n24602, 
        n24603, n24613, n29225, n26584, n26585, n23596, n23597, 
        n23598, n24604, n24605, n24614, n24606, n24607, n24615, 
        n747, n762, n25351, n23599, n23600, n23601, n23602, n23603, 
        n23604, n26565, n26562, n26566, n13518, n25354, n397, 
        n475, n23833, n318, n381, n23275;
    wire [11:0]phase_i;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(11[17:24])
    wire [1:0]phase_negation_i;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(23[12:28])
    wire [9:0]index_i_9__N_1748;
    wire [15:0]quarter_wave_sample_register_i;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(22[24:54])
    wire [14:0]quarter_wave_sample_register_i_15__N_1768;
    
    wire n26564, n475_adj_3470, n25111, n25112, n25123, n25113, 
        n25114, n25124, n25115, n25116, n25125, n23820, n23823, 
        n25148, n13449, n23826, n25149, n29242, n26561, n23456, 
        n13562, n13563, n24301, n13461, n23832, n23835, n25151, 
        n574, n23838, n25152, n23841, n764, n25153, n797, n828, 
        n24635, n24623, n24624, n24639, n24625, n24626, n24640, 
        n25177, n25178, n25181, n26559, n26557, n26560, n25179, 
        n25180, n25182, n26558, n285, n526, n541, n25344, n24627, 
        n24628, n24641, n24629, n24630, n24642, n23572, n620, 
        n635, n636, n24631, n24632, n24643, n24637, n24638, n24646, 
        n251, n443, n23831, n26556, n26555, n781, n29415, n29414, 
        n29325, n189, n875, n29229, n29412, n61, n30605, n29568, 
        n812, n27643, n28719, n24656, n24657, n24671, n397_adj_3471, 
        n23482, n24658, n24659, n24672, n716, n24660, n24661, 
        n24673, n24662, n24663, n24674, n24664, n24665, n24675, 
        n25345, n25360, n25346, n25347, n25361, n25348, n25349, 
        n25362, n25350, n25363, n23443, n29218, n526_adj_3472, n542, 
        n635_adj_3473, n23837, n25352, n25353, n25364, n25355, n25365, 
        n475_adj_3474, n23483, n859, n23444, n23567, n27403, n27405, 
        n25356, n25357, n25366, n25358, n25359, n25367, n316, 
        n94, n23562, n24686, n26553, n26550, n26554, n32037, n29413, 
        n270, n762_adj_3475, n23565, n23568, n24687, n762_adj_3476, 
        n379, n23571, n317, n24689, n28298, n13485, n349, n23574, 
        n24690, n890, n13515, n428, n252, n46, n716_adj_3477, 
        n604, n781_adj_3478, n443_adj_3479, n24691, n24692, n29150, 
        n29141, n24694, n860, n892, n23595, n700, n24695, n32050, 
        n7, n15, n24697, n23513, n924, n23607, n24699, n684, 
        n987, n23610, n24700, n124, n24907, n29061, n109, n24909, 
        n460, n890_adj_3480, n29233, n29337, n23852, n29152, n29056, 
        n701, n29257, n475_adj_3481, n32027, n23459, n29256, n653, 
        n32032, n684_adj_3482, n23854, n24908, n29215, n19993, n29239, 
        n19992, n412, n29156, n445, n32040, n924_adj_3483, n956, 
        n699, n24759, n24760, n24763, n16698, n23830, n684_adj_3484, 
        n24761, n24762, n24764, n723, n23563, n32041, n142, n157, 
        n32042, n23477, n24766, n24767, n24770, n32043, n301, 
        n24768, n24769, n24771, n32044, n32045, n985, n986, n29343, 
        n971, n29207, n939, n26552, n26551, n29588, n23561, n32059, 
        n32030, n923, n29525, n23573, n29151, n29082, n29524, 
        n29234, n251_adj_3485, n844_adj_3486, n860_adj_3487, n29362, 
        n444, n46_adj_3488, n23819, n747_adj_3489, n124_adj_3490, 
        n32046, n29222, n404, n23465, n173, n364, n23485, n32048, 
        n29261, n605, n29528, n23525, n32049, n396, n23531, n29084, 
        n29027, n716_adj_3491, n731, n732, n23530, n23532, n23528, 
        n23524, n23526, n653_adj_3492, n669, n142_adj_3493, n604_adj_3494, 
        n605_adj_3495, n29527, n173_adj_3496, n189_adj_3497, n29490, 
        n29491, n29492, n508, n32058, n23552, n23553, n29531, 
        n23548, n23549, n23550, n23506, n23569, n29169, n25186, 
        n796, n23519, n29076, n29075, n25155, n29530, n23518, 
        n23520, n26549, n29344, n23516, n29339, n676, n23515, 
        n23517, n476, n26477, n26478, n32051, n254, n29252, n29363, 
        n16890, n653_adj_3498, n32052, n397_adj_3499, n954, n413, 
        n29247, n22136, n27645, n29349, n29255, n908, n668, n316_adj_3500, 
        n317_adj_3501, n270_adj_3502, n286, n30481, n30482, n29182, 
        n32038, n30484, n29582, n29583, n29584, n26439, n29046, 
        n78, n467, n23593, n142_adj_3503, n15533, n158, n26548, 
        n30596, n30597, n30598, n30599, n29103, n30600, n30601, 
        n30602, n30603, n30604, n348, n29033, n23507, n23508, 
        n286_adj_3504, n29231, n716_adj_3505, n23533, n29485, n23535, 
        n29037, n27771, n29562, n444_adj_3506, n26481, n31735, n25183, 
        n27775, n908_adj_3507, n924_adj_3508, n23503, n541_adj_3509, 
        n890_adj_3510, n891, n23501, n669_adj_3511, n891_adj_3512, 
        n13497, n23594, n23521, n23522, n23523, n32053, n460_adj_3513, 
        n476_adj_3514, n844_adj_3515, n859_adj_3516, n860_adj_3517, 
        n491, n16936, n890_adj_3518, n891_adj_3519, n29228, n23489, 
        n27818, n23488, n812_adj_3520, n15423, n828_adj_3521, n700_adj_3522, 
        n23490, n29043, n797_adj_3523, n23486, n23487, n21724, n1018, 
        n882, n890_adj_3524, n29359, n891_adj_3525, n653_adj_3526, 
        n668_adj_3527, n669_adj_3528, n29556, n27819, n27824, n23484, 
        n23479, n413_adj_3529, n29085, n574_adj_3530, n29230, n542_adj_3531, 
        n93, n15523, n286_adj_3532, n460_adj_3533, n700_adj_3534, 
        n12501, n252_adj_3535, n23473, n28720, n25106, n23471, n23470, 
        n23468, n747_adj_3536, n763, n29092, n158_adj_3537, n23464, 
        n29345, n23462, n638, n23307, n27928, n16816, n28122, 
        n29030, n23461, n23463, n15_adj_3538, n30, n31, n29350, 
        n62, n29097, n31_adj_3539, n23458, n23460, n620_adj_3540, 
        n30_adj_3541, n31_adj_3542, n30485, n23453, n23452, n382, 
        n509, n27930, n23301, n27931, n32062, n13509, n13510, 
        n27951, n26482, n27953, n27954, n23818, n23450, n30_adj_3543, 
        n125, n332, n23449, n23821, n23822, n731_adj_3544, n732_adj_3545, 
        n28302, n30_adj_3546, n28509, n24305, n13453, n542_adj_3547, 
        n573, n27453, n23864, n23865, n16886, n21719, n24542, 
        n541_adj_3548, n29340, n141, n23435, n29240, n23434, n29214, 
        n23432, n23834, n23836, n557, n572, n23839, n23840, n29162, 
        n23842, n23843, n23844, n412_adj_3549, n29341, n23431, n23845, 
        n23846, n23847, n23848, n23849, n23850, n173_adj_3550, n732_adj_3551, 
        n23276, n732_adj_3552, n24668, n28941, n24677, n28182, n13454, 
        n25154, n23851, n23853, n684_adj_3553, n700_adj_3554, n29546, 
        n23855, n23856, n29545, n511, n16658, n1021, n317_adj_3555, 
        n413_adj_3556, n93_adj_3557, n28507, n731_adj_3558, n412_adj_3559, 
        n23857, n23858, n23859, n26606, n637, n28920, n24667, 
        n24676, n23860, n23861, n23862, n10789, n16938, n25150, 
        n25157, n25156, n25158, n25159, n25161, n26609, n25130, 
        n25109, n25122, n25108, n25121, n1002, n29098, n16734, 
        n252_adj_3560, n29555, n25104, n25119, n25038, n668_adj_3561, 
        n24619, n24939, n24942, n24938, n24941, n24548, n24549, 
        n24555, n24546, n24547, n24554, n638_adj_3562, n766, n22122, 
        n23066, n29554, n62_adj_3563, n25370, n25371, n25373, n25368, 
        n25369, n25372, n25160, n125_adj_3564, n31732, n252_adj_3565, 
        n31730, n31733, n28184, n24588, n24582, n24587, n24590, 
        n29035, n22166, n28127, n23277, n23065, n29060, n29055, 
        n189_adj_3566, n1022, n221, n24914, n93_adj_3567, n24915, 
        n29219, n23474, n29417, n124_adj_3568, n28506, n24680, n24681, 
        n24683, n24678, n24679, n24682, n285_adj_3569, n13559, n13560, 
        n24132, n13456, n29226, n23608, n24649, n24650, n24652, 
        n24647, n24648, n24651, n24585, n24586, n24589, n557_adj_3570, 
        n573_adj_3571, n573_adj_3572, n23278, n24711, n24712, n24714, 
        n24709, n24710, n24713, n491_adj_3573, n860_adj_3574, n443_adj_3575, 
        n32064, n23514, n1002_adj_3576, n506, n860_adj_3577, n29561, 
        n29560, n28519, n28522, n27772, n27773, n24906, n24910, 
        n23504, n23505, n26779, n26780, n32063, n24911, n908_adj_3578, 
        n653_adj_3579, n29532, n26781, n26784, n29487, n29488, n29489, 
        n124_adj_3580, n25054, n23476, n23500, n23502, n25053, n25052, 
        n684_adj_3581, n700_adj_3582, n669_adj_3583, n25051, n29237, 
        n25047, n506_adj_3584, n29189, n29526, n108, n25046, n986_adj_3585, 
        n25045, n25044, n29212, n25040, n25039, n286_adj_3586, n25037, 
        n23480, n94_adj_3587, n157_adj_3588, n24917, n15_adj_3589, 
        n954_adj_3590, n635_adj_3591, n16239, n636_adj_3592, n29567, 
        n188, n24918, n620_adj_3593, n348_adj_3594, n349_adj_3595, 
        n28758, n491_adj_3596, n26870, n26867, n26871, n28759, n26869, 
        n26868, n875_adj_3597, n379_adj_3598, n891_adj_3599, n859_adj_3600, 
        n860_adj_3601, n29083, n26866, n26865, n23609, n24913, n29566, 
        n908_adj_3602, n635_adj_3603, n23545, n23546, n23547, n23478, 
        n157_adj_3604, n29208, n636_adj_3605, n19995, n19996, n19997, 
        n28940, n28938, n507, n589, n476_adj_3606, n572_adj_3607, 
        n28939, n28937, n28936, n397_adj_3608, n413_adj_3609, n349_adj_3610, 
        n20007, n20008, n20009, n109_adj_3611, n125_adj_3612, n94_adj_3613, 
        n28919, n28916, n28918, n28917, n700_adj_3614, n32065, n26853, 
        n26851, n26854, n29044, n28915, n23540, n732_adj_3615, n221_adj_3616, 
        n142_adj_3617, n158_adj_3618, n506_adj_3619, n333, n348_adj_3620, 
        n24923, n26849, n15481, n924_adj_3621, n26852, n24924, n397_adj_3622, 
        n24925, n24926, n23433, n475_adj_3623, n24927, n23436, n253, 
        n12561, n24928, n190, n26850, n812_adj_3624, n26607, n29223, 
        n24130, n23605, n13452, n24912, n22204, n24553, n828_adj_3625, 
        n16238, n491_adj_3626, n507_adj_3627, n23466, n23469, n23472, 
        n23475, n573_adj_3628, n605_adj_3629, n491_adj_3630, n24571, 
        n29236, n23481, n24572, n333_adj_3631, n348_adj_3632, n364_adj_3633, 
        n397_adj_3634, n24916, n797_adj_3635, n931, n24931, n27507, 
        n24934, n29051, n572_adj_3636, n573_adj_3637, n19745;
    wire [15:0]o_val_pipeline_i_0__15__N_1799;
    
    wire n19744, n23542, n19743, n25041, n221_adj_3638, n252_adj_3639, 
        n25042, n19742, n19741, n19740, n25048, n19739, n891_adj_3640, 
        n19738, n25049, n25055, n25056, n763_adj_3641, n22568, n668_adj_3642, 
        n26785, n62_adj_3643, n892_adj_3644, n747_adj_3645, n716_adj_3646, 
        n32061, n93_adj_3647, n828_adj_3648, n32060, n28521, n28520, 
        n526_adj_3649, n684_adj_3650, n699_adj_3651, n23606, n28510, 
        n28508, n23467, n491_adj_3652, n23554, n23543, n23570, n23555, 
        n23556, n23544, n24943, n25374, n31734, n31731, n25127, 
        n25128, n25131, n15399, n491_adj_3653, n94_adj_3654, n24707, 
        n24708, n24701, n24702, n24705, n24706, n28301, n24558, 
        n24556, n24557, n24559, n25120, n23539, n23541, n27451, 
        n24644, n24633, n24634, n62_adj_3655, n28303, n24645, n221_adj_3656, 
        n24696, n24698, n24703, n24704, n875_adj_3657, n796_adj_3658, 
        n25043, n25050, n25057, n26608, n24550, n24551, n24552, 
        n25129, n30487, n27648, n28183, n28181, n27407, n24636, 
        n763_adj_3659, n24685, n28180, n29105, n28126, n348_adj_3660, 
        n23440, n23441, n23442, n29529, n23445, n23451, n62_adj_3661, 
        n27955, n27952, n23454, n27932, n27929, n27506, n25132;
    wire [15:0]n672;
    
    wire n29271, n19994, n23566, n444_adj_3662, n254_adj_3663, n285_adj_3664, 
        n23564, n23529, n13501, n1017, n22324, n30486, n30483, 
        n27647, n27644, n27646, n349_adj_3665, n23512, n507_adj_3666, 
        n27452, n93_adj_3667, n23527, n763_adj_3668, n205, n27406, 
        n27404, n348_adj_3669;
    
    LUT4 i13434_2_lut_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), .C(index_i[1]), 
         .D(index_i[0]), .Z(n844)) /* synthesis lut_function=(A ((C (D)+!C !(D))+!B)+!A (B+(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i13434_2_lut_3_lut_4_lut.init = 16'hf66f;
    L6MUX21 i22076 (.D0(n24561), .D1(n24562), .SD(index_i[6]), .Z(n24577));
    L6MUX21 i22077 (.D0(n24563), .D1(n24564), .SD(index_i[6]), .Z(n24578));
    L6MUX21 i22436 (.D0(n24929), .D1(n24930), .SD(index_i[6]), .Z(n24937));
    L6MUX21 i22078 (.D0(n24565), .D1(n24566), .SD(index_i[6]), .Z(n24579));
    PFUMX i24953 (.BLUT(n26586), .ALUT(n29221), .C0(index_i[5]), .Z(n26587));
    L6MUX21 i22079 (.D0(n24567), .D1(n24568), .SD(index_i[6]), .Z(n24580));
    L6MUX21 i22439 (.D0(n24935), .D1(n24936), .SD(index_i[6]), .Z(n24940));
    L6MUX21 i22080 (.D0(n24569), .D1(n24570), .SD(index_i[6]), .Z(n24581));
    L6MUX21 i22082 (.D0(n24573), .D1(n24574), .SD(index_i[6]), .Z(n24583));
    PFUMX i21095 (.BLUT(n23575), .ALUT(n23576), .C0(index_i[4]), .Z(n23577));
    PFUMX i21098 (.BLUT(n23578), .ALUT(n23579), .C0(index_i[4]), .Z(n23580));
    PFUMX i21101 (.BLUT(n23581), .ALUT(n23582), .C0(index_i[4]), .Z(n23583));
    PFUMX i21104 (.BLUT(n23584), .ALUT(n23585), .C0(index_i[4]), .Z(n23586));
    L6MUX21 i22107 (.D0(n24592), .D1(n24593), .SD(index_i[6]), .Z(n24608));
    L6MUX21 i22108 (.D0(n24594), .D1(n24595), .SD(index_i[6]), .Z(n24609));
    L6MUX21 i22109 (.D0(n24596), .D1(n24597), .SD(index_i[6]), .Z(n24610));
    PFUMX i21110 (.BLUT(n23590), .ALUT(n23591), .C0(index_i[4]), .Z(n23592));
    PFUMX i22111 (.BLUT(n24600), .ALUT(n24601), .C0(index_i[6]), .Z(n24612));
    L6MUX21 i22112 (.D0(n24602), .D1(n24603), .SD(index_i[6]), .Z(n24613));
    PFUMX i24951 (.BLUT(n29225), .ALUT(n26584), .C0(index_i[2]), .Z(n26585));
    PFUMX i21116 (.BLUT(n23596), .ALUT(n23597), .C0(index_i[4]), .Z(n23598));
    L6MUX21 i22113 (.D0(n24604), .D1(n24605), .SD(index_i[6]), .Z(n24614));
    PFUMX i22114 (.BLUT(n24606), .ALUT(n24607), .C0(index_i[6]), .Z(n24615));
    PFUMX i22850 (.BLUT(n747), .ALUT(n762), .C0(index_i[4]), .Z(n25351));
    PFUMX i21119 (.BLUT(n23599), .ALUT(n23600), .C0(index_i[4]), .Z(n23601));
    PFUMX i21122 (.BLUT(n23602), .ALUT(n23603), .C0(index_i[4]), .Z(n23604));
    L6MUX21 i24945 (.D0(n26565), .D1(n26562), .SD(index_i[5]), .Z(n26566));
    PFUMX i22853 (.BLUT(n844), .ALUT(n13518), .C0(index_i[4]), .Z(n25354));
    LUT4 i21351_3_lut (.A(n397), .B(n475), .C(index_i[4]), .Z(n23833)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21351_3_lut.init = 16'hcaca;
    PFUMX i20793 (.BLUT(n318), .ALUT(n381), .C0(index_i[6]), .Z(n23275));
    FD1P3AX phase_i_i0_i0 (.D(o_phase[0]), .SP(dac_clk_p_c_enable_630), 
            .CK(dac_clk_p_c), .Q(phase_i[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam phase_i_i0_i0.GSR = "DISABLED";
    FD1S3DX phase_negation_i_i0 (.D(phase_i[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(phase_negation_i[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam phase_negation_i_i0.GSR = "DISABLED";
    FD1S3DX index_i_i0 (.D(index_i_9__N_1748[0]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(index_i[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam index_i_i0.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i1 (.D(\o_val_pipeline_i[0] [0]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(modulation_output[0])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i1.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i0 (.D(quarter_wave_sample_register_i_15__N_1768[0]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_i[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_i_i0.GSR = "DISABLED";
    PFUMX i24943 (.BLUT(n26564), .ALUT(n475_adj_3470), .C0(index_i[4]), 
          .Z(n26565));
    L6MUX21 i22622 (.D0(n25111), .D1(n25112), .SD(index_i[6]), .Z(n25123));
    L6MUX21 i22623 (.D0(n25113), .D1(n25114), .SD(index_i[6]), .Z(n25124));
    L6MUX21 i22624 (.D0(n25115), .D1(n25116), .SD(index_i[6]), .Z(n25125));
    L6MUX21 i22647 (.D0(n23820), .D1(n23823), .SD(index_i[6]), .Z(n25148));
    PFUMX i22648 (.BLUT(n13449), .ALUT(n23826), .C0(index_i[6]), .Z(n25149));
    LUT4 mux_208_Mux_6_i378_3_lut_4_lut_3_lut_rep_582 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29242)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_6_i378_3_lut_4_lut_3_lut_rep_582.init = 16'h4949;
    PFUMX i24940 (.BLUT(n26561), .ALUT(n23456), .C0(index_i[4]), .Z(n26562));
    PFUMX i11165 (.BLUT(n13562), .ALUT(n13563), .C0(n24301), .Z(n13461));
    L6MUX21 i22650 (.D0(n23832), .D1(n23835), .SD(index_i[6]), .Z(n25151));
    L6MUX21 i22651 (.D0(n574), .D1(n23838), .SD(index_i[6]), .Z(n25152));
    L6MUX21 i22652 (.D0(n23841), .D1(n764), .SD(index_i[6]), .Z(n25153));
    PFUMX i22134 (.BLUT(n797), .ALUT(n828), .C0(index_i[5]), .Z(n24635));
    L6MUX21 i22138 (.D0(n24623), .D1(n24624), .SD(index_i[6]), .Z(n24639));
    L6MUX21 i22139 (.D0(n24625), .D1(n24626), .SD(index_i[6]), .Z(n24640));
    PFUMX i22680 (.BLUT(n25177), .ALUT(n25178), .C0(index_i[6]), .Z(n25181));
    L6MUX21 i24938 (.D0(n26559), .D1(n26557), .SD(index_i[5]), .Z(n26560));
    PFUMX i22681 (.BLUT(n25179), .ALUT(n25180), .C0(index_i[6]), .Z(n25182));
    PFUMX i24936 (.BLUT(n26558), .ALUT(n285), .C0(index_i[4]), .Z(n26559));
    PFUMX i22843 (.BLUT(n526), .ALUT(n541), .C0(index_i[4]), .Z(n25344));
    L6MUX21 i22140 (.D0(n24627), .D1(n24628), .SD(index_i[6]), .Z(n24641));
    L6MUX21 i22141 (.D0(n24629), .D1(n24630), .SD(index_i[6]), .Z(n24642));
    LUT4 i21090_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n23572)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (D))+!A !(B (C (D))+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21090_3_lut_3_lut_4_lut.init = 16'h4933;
    PFUMX mux_208_Mux_1_i636 (.BLUT(n620), .ALUT(n635), .C0(index_i[4]), 
          .Z(n636)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    L6MUX21 i22142 (.D0(n24631), .D1(n24632), .SD(index_i[6]), .Z(n24643));
    L6MUX21 i22145 (.D0(n24637), .D1(n24638), .SD(index_i[6]), .Z(n24646));
    LUT4 i21114_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n23596)) /* synthesis lut_function=(A (B (C)+!B (C (D)+!C !(D)))+!A !(B (C+!(D))+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21114_3_lut_4_lut_4_lut.init = 16'ha593;
    LUT4 i21349_3_lut (.A(n251), .B(n443), .C(index_i[4]), .Z(n23831)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21349_3_lut.init = 16'hcaca;
    PFUMX i24934 (.BLUT(n26556), .ALUT(n26555), .C0(index_i[4]), .Z(n26557));
    LUT4 mux_208_Mux_6_i781_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n781)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+(D)))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_6_i781_3_lut_4_lut_4_lut_4_lut.init = 16'h9993;
    LUT4 mux_208_Mux_4_i93_3_lut_4_lut_4_lut_3_lut_rep_755_4_lut (.A(index_i[0]), 
         .B(index_i[3]), .C(index_i[1]), .D(index_i[2]), .Z(n29415)) /* synthesis lut_function=(!(A (B+(C (D)))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_4_i93_3_lut_4_lut_4_lut_3_lut_rep_755_4_lut.init = 16'h4666;
    LUT4 mux_208_Mux_4_i236_3_lut_4_lut_3_lut_rep_754_4_lut (.A(index_i[0]), 
         .B(index_i[3]), .C(index_i[1]), .D(index_i[2]), .Z(n29414)) /* synthesis lut_function=(A (B)+!A !(B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_4_i236_3_lut_4_lut_3_lut_rep_754_4_lut.init = 16'h999d;
    LUT4 i11197_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[4]), .D(n29325), .Z(n189)) /* synthesis lut_function=(A (B (C (D)))+!A !(B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11197_3_lut_4_lut_4_lut_4_lut.init = 16'h9555;
    LUT4 i11210_3_lut_4_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[1]), .Z(n875)) /* synthesis lut_function=(A (B (C))+!A !(B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11210_3_lut_4_lut_3_lut_4_lut.init = 16'h95d5;
    LUT4 mux_208_Mux_4_i61_3_lut (.A(n29229), .B(n29412), .C(index_i[3]), 
         .Z(n61)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_4_i61_3_lut.init = 16'hcaca;
    LUT4 i24136_3_lut (.A(n30605), .B(n29568), .C(index_i[5]), .Z(n24606)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24136_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_4_i812_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[4]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n812)) /* synthesis lut_function=(A (B (C+(D)))+!A !(B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_4_i812_3_lut_3_lut_4_lut.init = 16'h9995;
    LUT4 n293_bdd_3_lut_26924_3_lut_4_lut (.A(index_i[0]), .B(index_i[3]), 
         .C(index_i[1]), .D(index_i[2]), .Z(n27643)) /* synthesis lut_function=(!(A (B+(C (D)+!C !(D)))+!A !(B+!((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n293_bdd_3_lut_26924_3_lut_4_lut.init = 16'h4674;
    LUT4 n162_bdd_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[2]), .C(index_i[1]), 
         .D(index_i[3]), .Z(n28719)) /* synthesis lut_function=(!(A (B)+!A !(B (C+(D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n162_bdd_4_lut_4_lut_4_lut.init = 16'h6763;
    L6MUX21 i22170 (.D0(n24656), .D1(n24657), .SD(index_i[6]), .Z(n24671));
    LUT4 mux_208_Mux_3_i397_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n397_adj_3471)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !(B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_3_i397_3_lut_4_lut_4_lut.init = 16'ha95a;
    LUT4 mux_208_Mux_0_i747_3_lut_4_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[1]), .Z(n747)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C+(D)))+!A !(B ((D)+!C)+!B (C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_0_i747_3_lut_4_lut_3_lut_4_lut.init = 16'h5596;
    LUT4 i21000_3_lut_4_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[3]), 
         .C(index_i[1]), .D(index_i[2]), .Z(n23482)) /* synthesis lut_function=(!(A (B)+!A !(B (C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21000_3_lut_4_lut_3_lut_4_lut.init = 16'h6662;
    L6MUX21 i22171 (.D0(n24658), .D1(n24659), .SD(index_i[6]), .Z(n24672));
    LUT4 mux_208_Mux_1_i716_3_lut_3_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[1]), .D(index_i[3]), .Z(n716)) /* synthesis lut_function=(!(A (B (D)+!B !(C))+!A !(B (C (D))+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_1_i716_3_lut_3_lut_4_lut_4_lut.init = 16'h70a9;
    L6MUX21 i22172 (.D0(n24660), .D1(n24661), .SD(index_i[6]), .Z(n24673));
    L6MUX21 i22173 (.D0(n24662), .D1(n24663), .SD(index_i[6]), .Z(n24674));
    L6MUX21 i22174 (.D0(n24664), .D1(n24665), .SD(index_i[6]), .Z(n24675));
    L6MUX21 i22859 (.D0(n25344), .D1(n25345), .SD(index_i[5]), .Z(n25360));
    L6MUX21 i22860 (.D0(n25346), .D1(n25347), .SD(index_i[5]), .Z(n25361));
    L6MUX21 i22861 (.D0(n25348), .D1(n25349), .SD(index_i[5]), .Z(n25362));
    L6MUX21 i22862 (.D0(n25350), .D1(n25351), .SD(index_i[5]), .Z(n25363));
    LUT4 i20961_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[1]), .Z(n23443)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+!(D)))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20961_3_lut_4_lut_4_lut_4_lut.init = 16'h9399;
    LUT4 mux_208_Mux_8_i542_3_lut_4_lut (.A(n29218), .B(index_i[3]), .C(index_i[4]), 
         .D(n526_adj_3472), .Z(n542)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_8_i542_3_lut_4_lut.init = 16'h6f60;
    LUT4 i21355_3_lut_4_lut (.A(n29218), .B(index_i[3]), .C(index_i[4]), 
         .D(n635_adj_3473), .Z(n23837)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21355_3_lut_4_lut.init = 16'hf606;
    L6MUX21 i22863 (.D0(n25352), .D1(n25353), .SD(index_i[5]), .Z(n25364));
    L6MUX21 i22864 (.D0(n25354), .D1(n25355), .SD(index_i[5]), .Z(n25365));
    LUT4 mux_208_Mux_5_i475_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[1]), .Z(n475_adj_3474)) /* synthesis lut_function=(A (B ((D)+!C))+!A (B (C)+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_5_i475_3_lut_4_lut_4_lut.init = 16'hd949;
    LUT4 i21001_3_lut_4_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[1]), .Z(n23483)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C))+!A (B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21001_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'h29a9;
    LUT4 mux_208_Mux_3_i859_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n859)) /* synthesis lut_function=(!(A (B (D)+!B !(D))+!A (B (C+(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_3_i859_3_lut_3_lut_4_lut.init = 16'h339c;
    LUT4 i20962_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n23444)) /* synthesis lut_function=(A (C)+!A !(B (C)+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20962_3_lut_4_lut_4_lut.init = 16'hb4b5;
    LUT4 i21085_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n23567)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B (C+(D))+!B (C)))) */ ;
    defparam i21085_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h7c78;
    LUT4 n78_bdd_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n27403)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A !((C)+!B))) */ ;
    defparam n78_bdd_3_lut_4_lut_4_lut_4_lut.init = 16'h7173;
    LUT4 n285_bdd_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n27405)) /* synthesis lut_function=(A (B (C)+!B ((D)+!C))+!A (B+!(C))) */ ;
    defparam n285_bdd_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'he7c7;
    L6MUX21 i22865 (.D0(n25356), .D1(n25357), .SD(index_i[5]), .Z(n25366));
    L6MUX21 i22866 (.D0(n25358), .D1(n25359), .SD(index_i[5]), .Z(n25367));
    LUT4 mux_208_Mux_9_i316_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), 
         .B(index_i[2]), .C(index_i[3]), .D(index_i[0]), .Z(n316)) /* synthesis lut_function=(!(A (B (C)+!B !(C+(D)))+!A !(B+(C)))) */ ;
    defparam mux_208_Mux_9_i316_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h7e7c;
    PFUMX i22185 (.BLUT(n94), .ALUT(n23562), .C0(index_i[5]), .Z(n24686));
    L6MUX21 i24931 (.D0(n26553), .D1(n26550), .SD(index_i[5]), .Z(n26554));
    LUT4 mux_208_Mux_4_i270_3_lut (.A(n32037), .B(n29413), .C(index_i[3]), 
         .Z(n270)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_4_i270_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_7_i762_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), 
         .B(index_i[2]), .C(index_i[3]), .D(index_i[0]), .Z(n762_adj_3475)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B ((D)+!C)+!B !(C)))) */ ;
    defparam mux_208_Mux_7_i762_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h3878;
    L6MUX21 i22186 (.D0(n23565), .D1(n23568), .SD(index_i[5]), .Z(n24687));
    LUT4 mux_208_Mux_8_i443_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n443)) /* synthesis lut_function=(A (B (C+!(D))+!B !((D)+!C))+!A !(B (D)+!B ((D)+!C))) */ ;
    defparam mux_208_Mux_8_i443_3_lut_4_lut_4_lut.init = 16'h80fc;
    LUT4 i11203_3_lut_3_lut_4_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n762_adj_3476)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11203_3_lut_3_lut_4_lut_3_lut_4_lut.init = 16'h1999;
    LUT4 mux_208_Mux_0_i379_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n379)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !((D)+!C))+!A !(B ((D)+!C)+!B (D))) */ ;
    defparam mux_208_Mux_0_i379_3_lut_4_lut_4_lut.init = 16'h8079;
    PFUMX i22188 (.BLUT(n23571), .ALUT(n317), .C0(index_i[5]), .Z(n24689));
    LUT4 n589_bdd_3_lut_26394_4_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[4]), .D(index_i[1]), .Z(n28298)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n589_bdd_3_lut_26394_4_lut_4_lut_4_lut.init = 16'h8387;
    LUT4 i11189_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n13485)) /* synthesis lut_function=(!(A (B (C)+!B ((D)+!C))+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11189_3_lut_4_lut_4_lut.init = 16'h4969;
    PFUMX i22189 (.BLUT(n349), .ALUT(n23574), .C0(index_i[5]), .Z(n24690));
    LUT4 mux_208_Mux_2_i890_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n890)) /* synthesis lut_function=(A (B (C)+!B !(C+!(D)))+!A !(B (C+(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_2_i890_3_lut_4_lut_4_lut.init = 16'h9394;
    LUT4 i11219_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n13515)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))+!A !(B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11219_3_lut_4_lut_4_lut.init = 16'hb5b3;
    LUT4 mux_208_Mux_0_i428_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[2]), 
         .B(index_i[1]), .C(index_i[0]), .D(index_i[3]), .Z(n428)) /* synthesis lut_function=(A (B (C+!(D))+!B !((D)+!C))+!A (B (D)+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_0_i428_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hd5a9;
    LUT4 mux_208_Mux_5_i252_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[4]), .Z(n252)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+(D)))+!A (B (C (D))+!B !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_5_i252_3_lut_4_lut.init = 16'hc993;
    LUT4 mux_208_Mux_0_i46_3_lut_4_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n46)) /* synthesis lut_function=(A (B)+!A ((C+(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_0_i46_3_lut_4_lut_4_lut_4_lut.init = 16'hddd9;
    LUT4 mux_208_Mux_8_i716_3_lut_4_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n716_adj_3477)) /* synthesis lut_function=(!(A (B)+!A !(B+(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_8_i716_3_lut_4_lut_4_lut_4_lut.init = 16'h7776;
    LUT4 mux_208_Mux_0_i604_3_lut_4_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[1]), .D(index_i[3]), .Z(n604)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A !(B (D)+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_0_i604_3_lut_4_lut_4_lut_4_lut.init = 16'h5439;
    LUT4 mux_208_Mux_0_i781_4_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n781_adj_3478)) /* synthesis lut_function=(!(A (B+!((D)+!C))+!A !(B (C)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_0_i781_4_lut_4_lut_4_lut.init = 16'h6252;
    LUT4 i21109_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[2]), .C(index_i[3]), 
         .D(index_i[1]), .Z(n23591)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+!(D)))+!A !(B+!(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21109_3_lut_4_lut_4_lut.init = 16'h6c67;
    LUT4 i11222_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n13518)) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B ((D)+!C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11222_3_lut_4_lut_4_lut.init = 16'hcdad;
    LUT4 mux_208_Mux_0_i443_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n443_adj_3479)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(D))+!A (B (D)+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_0_i443_3_lut_4_lut_4_lut_4_lut.init = 16'h32d5;
    L6MUX21 i22190 (.D0(n23577), .D1(n23580), .SD(index_i[5]), .Z(n24691));
    L6MUX21 i22191 (.D0(n23583), .D1(n23586), .SD(index_i[5]), .Z(n24692));
    LUT4 i22679_3_lut_4_lut_4_lut (.A(n29150), .B(index_i[4]), .C(index_i[5]), 
         .D(n29141), .Z(n25180)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C)+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i22679_3_lut_4_lut_4_lut.init = 16'h0434;
    L6MUX21 i22193 (.D0(n23592), .D1(n636), .SD(index_i[5]), .Z(n24694));
    LUT4 mux_208_Mux_8_i892_3_lut_4_lut (.A(n29150), .B(index_i[4]), .C(index_i[5]), 
         .D(n860), .Z(n892)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_8_i892_3_lut_4_lut.init = 16'h4f40;
    PFUMX i22194 (.BLUT(n23595), .ALUT(n700), .C0(index_i[5]), .Z(n24695));
    LUT4 mux_208_Mux_4_i15_3_lut (.A(n32050), .B(n7), .C(index_i[3]), 
         .Z(n15)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_4_i15_3_lut.init = 16'hcaca;
    L6MUX21 i22196 (.D0(n23598), .D1(n23601), .SD(index_i[5]), .Z(n24697));
    LUT4 i21031_3_lut_4_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[1]), 
         .C(index_i[0]), .D(index_i[3]), .Z(n23513)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C+!(D)))+!A !(((D)+!C)+!B)) */ ;
    defparam i21031_3_lut_4_lut_4_lut_4_lut.init = 16'ha86a;
    PFUMX i22198 (.BLUT(n924), .ALUT(n23607), .C0(index_i[5]), .Z(n24699));
    LUT4 mux_208_Mux_1_i684_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n684)) /* synthesis lut_function=(A (B ((D)+!C)+!B !((D)+!C))+!A !(B (C+(D))+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_1_i684_3_lut_4_lut_4_lut.init = 16'h992d;
    PFUMX i22199 (.BLUT(n987), .ALUT(n23610), .C0(index_i[5]), .Z(n24700));
    LUT4 mux_208_Mux_8_i124_3_lut_3_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n124)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (B (C+!(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_8_i124_3_lut_3_lut_4_lut_4_lut.init = 16'h07a1;
    LUT4 i22406_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n24907)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i22406_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hf81f;
    LUT4 mux_208_Mux_8_i61_3_lut_rep_401_4_lut_4_lut_4_lut (.A(index_i[1]), 
         .B(index_i[0]), .C(index_i[2]), .D(index_i[3]), .Z(n29061)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A (B (C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_8_i61_3_lut_rep_401_4_lut_4_lut_4_lut.init = 16'he0f8;
    LUT4 mux_208_Mux_8_i109_3_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n109)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (B (C+!(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_8_i109_3_lut_4_lut_4_lut.init = 16'hf85e;
    LUT4 i22408_3_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[0]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n24909)) /* synthesis lut_function=(A (B (C+!(D))+!B !((D)+!C))+!A !(B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i22408_3_lut_4_lut_4_lut.init = 16'h81f8;
    LUT4 mux_208_Mux_8_i251_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), 
         .B(index_i[0]), .C(index_i[2]), .D(index_i[3]), .Z(n251)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_8_i251_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h07e0;
    LUT4 mux_208_Mux_0_i460_3_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n460)) /* synthesis lut_function=(A (B+(C))+!A (C (D)+!C !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_0_i460_3_lut_4_lut_4_lut.init = 16'hf8ad;
    LUT4 mux_208_Mux_0_i890_3_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n890_adj_3480)) /* synthesis lut_function=(!(A (B (D)+!B !(C))+!A !(B (C (D)+!C !(D))+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_0_i890_3_lut_4_lut_4_lut.init = 16'h70ac;
    LUT4 i21115_3_lut (.A(n29229), .B(n29233), .C(index_i[3]), .Z(n23597)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21115_3_lut.init = 16'hcaca;
    LUT4 i21370_3_lut_4_lut_4_lut_4_lut (.A(n29337), .B(index_i[2]), .C(index_i[3]), 
         .D(index_i[4]), .Z(n23852)) /* synthesis lut_function=(A (B)+!A (B (C (D))+!B !(C (D)))) */ ;
    defparam i21370_3_lut_4_lut_4_lut_4_lut.init = 16'hc999;
    LUT4 mux_208_Mux_10_i701_4_lut_4_lut (.A(n29152), .B(index_i[4]), .C(index_i[5]), 
         .D(n29056), .Z(n701)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B (C (D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_10_i701_4_lut_4_lut.init = 16'h3efe;
    LUT4 mux_208_Mux_7_i475_3_lut_4_lut (.A(n29337), .B(index_i[2]), .C(index_i[3]), 
         .D(n29257), .Z(n475_adj_3481)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+(D)))) */ ;
    defparam mux_208_Mux_7_i475_3_lut_4_lut.init = 16'h9f90;
    LUT4 i20977_3_lut_4_lut (.A(n29337), .B(index_i[2]), .C(index_i[3]), 
         .D(n32027), .Z(n23459)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;
    defparam i20977_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_208_Mux_7_i653_3_lut_4_lut (.A(n29337), .B(index_i[2]), .C(index_i[3]), 
         .D(n29256), .Z(n653)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam mux_208_Mux_7_i653_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_208_Mux_2_i684_3_lut_4_lut (.A(n29337), .B(index_i[2]), .C(index_i[3]), 
         .D(n32032), .Z(n684_adj_3482)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;
    defparam mux_208_Mux_2_i684_3_lut_4_lut.init = 16'h6f60;
    LUT4 i21372_4_lut_4_lut_4_lut (.A(n29337), .B(index_i[2]), .C(index_i[4]), 
         .D(index_i[3]), .Z(n23854)) /* synthesis lut_function=(A (B)+!A !(B (C+(D))+!B !(C+(D)))) */ ;
    defparam i21372_4_lut_4_lut_4_lut.init = 16'h999c;
    LUT4 i22407_3_lut_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n24908)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C+!(D))+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i22407_3_lut_3_lut_4_lut_4_lut.init = 16'h1f81;
    LUT4 i17679_3_lut (.A(n29215), .B(n29242), .C(index_i[3]), .Z(n19993)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17679_3_lut.init = 16'hcaca;
    LUT4 i21120_3_lut_4_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n23602)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(D))+!A !(B (D)+!B ((D)+!C)))) */ ;
    defparam i21120_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'h7f01;
    LUT4 i17678_3_lut (.A(n29242), .B(n29239), .C(index_i[3]), .Z(n19992)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17678_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_0_i412_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .D(index_i[3]), .Z(n412)) /* synthesis lut_function=(A (B (D)+!B (C+(D)))+!A !(B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;
    defparam mux_208_Mux_0_i412_3_lut_4_lut_4_lut_4_lut.init = 16'hab70;
    LUT4 mux_208_Mux_11_i445_3_lut_4_lut_4_lut_4_lut (.A(index_i[3]), .B(index_i[4]), 
         .C(index_i[5]), .D(n29156), .Z(n445)) /* synthesis lut_function=(!(A (B (C))+!A !(B+(C+(D))))) */ ;
    defparam mux_208_Mux_11_i445_3_lut_4_lut_4_lut_4_lut.init = 16'h7f7e;
    LUT4 mux_208_Mux_3_i676_3_lut_4_lut_3_lut_rep_839 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n32040)) /* synthesis lut_function=(A (B (C))+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_3_i676_3_lut_4_lut_3_lut_rep_839.init = 16'h9494;
    LUT4 mux_208_Mux_7_i956_3_lut_3_lut_4_lut (.A(n29152), .B(index_i[4]), 
         .C(n924_adj_3483), .D(index_i[5]), .Z(n956)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_7_i956_3_lut_3_lut_4_lut.init = 16'h11f0;
    LUT4 mux_208_Mux_7_i699_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n699)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (D))) */ ;
    defparam mux_208_Mux_7_i699_3_lut_4_lut_4_lut_4_lut.init = 16'hf70e;
    PFUMX i22262 (.BLUT(n24759), .ALUT(n24760), .C0(index_i[5]), .Z(n24763));
    LUT4 i21348_3_lut (.A(n397), .B(n16698), .C(index_i[4]), .Z(n23830)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;
    defparam i21348_3_lut.init = 16'h3a3a;
    LUT4 mux_208_Mux_3_i684_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[4]), .Z(n684_adj_3484)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A !(B ((D)+!C)+!B (C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_3_i684_3_lut_3_lut_4_lut.init = 16'h5594;
    PFUMX i22263 (.BLUT(n24761), .ALUT(n24762), .C0(index_i[5]), .Z(n24764));
    LUT4 i21081_3_lut (.A(n723), .B(n29233), .C(index_i[3]), .Z(n23563)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21081_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_6_i29_3_lut_4_lut_3_lut_rep_840 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n32041)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_6_i29_3_lut_4_lut_3_lut_rep_840.init = 16'h6969;
    LUT4 mux_208_Mux_0_i142_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n142)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C))+!A !(B (C (D)+!C !(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_0_i142_3_lut_4_lut_4_lut.init = 16'ha569;
    LUT4 n26585_bdd_3_lut (.A(n26585), .B(n157), .C(index_i[4]), .Z(n26586)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n26585_bdd_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_6_i60_3_lut_4_lut_3_lut_rep_841 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n32042)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_6_i60_3_lut_4_lut_3_lut_rep_841.init = 16'hd6d6;
    LUT4 i20995_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n23477)) /* synthesis lut_function=(A (B (C)+!B !(C (D)+!C !(D)))+!A (B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20995_3_lut_4_lut_4_lut.init = 16'hd6a5;
    PFUMX i22269 (.BLUT(n24766), .ALUT(n24767), .C0(index_i[5]), .Z(n24770));
    LUT4 mux_208_Mux_6_i262_3_lut_4_lut_3_lut_rep_842 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n32043)) /* synthesis lut_function=(A ((C)+!B)+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_6_i262_3_lut_4_lut_3_lut_rep_842.init = 16'hb6b6;
    LUT4 mux_208_Mux_1_i301_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n301)) /* synthesis lut_function=(A (B (C+(D))+!B !(D))+!A !(B (C+(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_1_i301_3_lut_4_lut_4_lut.init = 16'h99b6;
    PFUMX i22270 (.BLUT(n24768), .ALUT(n24769), .C0(index_i[5]), .Z(n24771));
    LUT4 mux_208_Mux_6_i467_3_lut_3_lut_3_lut_rep_843 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n32044)) /* synthesis lut_function=(!(A (B)+!A (B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_6_i467_3_lut_3_lut_3_lut_rep_843.init = 16'h3636;
    LUT4 mux_208_Mux_0_i986_3_lut (.A(n32045), .B(n985), .C(index_i[3]), 
         .Z(n986)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_0_i986_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_0_i971_3_lut (.A(n32044), .B(n29343), .C(index_i[3]), 
         .Z(n971)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_0_i971_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_0_i939_4_lut (.A(n7), .B(n29207), .C(index_i[3]), 
         .D(index_i[2]), .Z(n939)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_0_i939_4_lut.init = 16'hfaca;
    PFUMX i24929 (.BLUT(n26552), .ALUT(n26551), .C0(index_i[4]), .Z(n26553));
    LUT4 i24013_3_lut (.A(n29588), .B(n23561), .C(index_i[4]), .Z(n23562)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24013_3_lut.init = 16'hcaca;
    LUT4 i21342_3_lut_else_4_lut (.A(index_i[4]), .B(index_i[0]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n32059)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A !(C (D)+!C !(D)))) */ ;
    defparam i21342_3_lut_else_4_lut.init = 16'h5a85;
    LUT4 mux_208_Mux_0_i923_3_lut (.A(n32030), .B(n29257), .C(index_i[3]), 
         .Z(n923)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_0_i923_3_lut.init = 16'hcaca;
    LUT4 i26830_then_4_lut (.A(index_i[2]), .B(index_i[1]), .C(index_i[4]), 
         .D(index_i[3]), .Z(n29525)) /* synthesis lut_function=(A (B (C+(D))+!B !(C))+!A !(B (C+(D))+!B !(C+!(D)))) */ ;
    defparam i26830_then_4_lut.init = 16'h9a97;
    LUT4 i21091_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n23573)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(D))+!A (B (D)+!B ((D)+!C))) */ ;
    defparam i21091_3_lut_4_lut_4_lut.init = 16'hd52b;
    LUT4 i22677_3_lut_4_lut_4_lut (.A(n29151), .B(index_i[4]), .C(index_i[5]), 
         .D(n29082), .Z(n25178)) /* synthesis lut_function=(A ((C+!(D))+!B)+!A (B (C+!(D))+!B !(C))) */ ;
    defparam i22677_3_lut_4_lut_4_lut.init = 16'he3ef;
    LUT4 mux_208_Mux_6_i157_3_lut_4_lut (.A(n29207), .B(index_i[2]), .C(index_i[3]), 
         .D(n29413), .Z(n157)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_6_i157_3_lut_4_lut.init = 16'hf606;
    LUT4 i26830_else_4_lut (.A(index_i[2]), .B(index_i[1]), .C(index_i[4]), 
         .D(index_i[3]), .Z(n29524)) /* synthesis lut_function=(!(A (B (C)+!B (C+(D)))+!A !(B (C (D)+!C !(D))+!B (C+!(D))))) */ ;
    defparam i26830_else_4_lut.init = 16'h581f;
    LUT4 mux_208_Mux_6_i251_3_lut_4_lut (.A(n29207), .B(index_i[2]), .C(index_i[3]), 
         .D(n29234), .Z(n251_adj_3485)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_6_i251_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_208_Mux_6_i860_3_lut_3_lut (.A(n29061), .B(index_i[4]), .C(n844_adj_3486), 
         .Z(n860_adj_3487)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam mux_208_Mux_6_i860_3_lut_3_lut.init = 16'h7474;
    LUT4 i11183_3_lut_4_lut (.A(n29207), .B(index_i[2]), .C(n29362), .D(n29234), 
         .Z(n444)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11183_3_lut_4_lut.init = 16'h6f60;
    LUT4 i21337_3_lut_3_lut (.A(n29061), .B(index_i[4]), .C(n46_adj_3488), 
         .Z(n23819)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam i21337_3_lut_3_lut.init = 16'h7474;
    LUT4 mux_208_Mux_4_i747_3_lut_4_lut (.A(n29207), .B(index_i[2]), .C(index_i[3]), 
         .D(n32043), .Z(n747_adj_3489)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_4_i747_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_208_Mux_6_i475_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n475_adj_3470)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A !(B (C+(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_6_i475_3_lut_4_lut_4_lut.init = 16'h9936;
    LUT4 mux_208_Mux_6_i483_3_lut_3_lut_rep_844 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n32045)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_6_i483_3_lut_3_lut_rep_844.init = 16'h6c6c;
    LUT4 mux_208_Mux_0_i124_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n124_adj_3490)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A !(B (D)+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_0_i124_3_lut_4_lut_4_lut.init = 16'h6c99;
    LUT4 mux_208_Mux_5_i363_3_lut_4_lut_3_lut_rep_845 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n32046)) /* synthesis lut_function=(A (B+!(C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_5_i363_3_lut_4_lut_3_lut_rep_845.init = 16'hdbdb;
    LUT4 i20983_3_lut_4_lut (.A(n29222), .B(index_i[1]), .C(index_i[3]), 
         .D(n404), .Z(n23465)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20983_3_lut_4_lut.init = 16'hdfd0;
    LUT4 mux_208_Mux_0_i173_3_lut_4_lut (.A(n29222), .B(index_i[1]), .C(index_i[3]), 
         .D(n29239), .Z(n173)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_0_i173_3_lut_4_lut.init = 16'hdfd0;
    LUT4 mux_208_Mux_1_i620_3_lut_4_lut (.A(n29222), .B(index_i[1]), .C(index_i[3]), 
         .D(n32037), .Z(n620)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_1_i620_3_lut_4_lut.init = 16'hdfd0;
    LUT4 mux_208_Mux_0_i364_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n364)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A ((C+!(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_0_i364_3_lut_3_lut_4_lut.init = 16'hdb55;
    LUT4 mux_208_Mux_6_i844_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n844_adj_3486)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (B (C)+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_6_i844_3_lut_4_lut_4_lut.init = 16'hc1e0;
    LUT4 i21003_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n23485)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A !(B (C+!(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21003_3_lut_4_lut_4_lut.init = 16'ha52b;
    LUT4 i12920_3_lut_3_lut_rep_847 (.A(index_i[2]), .B(index_i[0]), .C(index_i[1]), 
         .Z(n32048)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12920_3_lut_3_lut_rep_847.init = 16'hd0d0;
    LUT4 i11171_3_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[0]), .C(index_i[1]), 
         .D(n29261), .Z(n605)) /* synthesis lut_function=(A (B (C)+!B !(C+!(D)))+!A (B (C)+!B !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11171_3_lut_4_lut_4_lut.init = 16'hc3d0;
    LUT4 mux_208_Mux_5_i781_3_lut_4_lut_4_lut_then_4_lut (.A(index_i[3]), 
         .B(index_i[0]), .C(index_i[4]), .D(index_i[2]), .Z(n29528)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_5_i781_3_lut_4_lut_4_lut_then_4_lut.init = 16'hece0;
    LUT4 i21043_3_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[0]), .C(index_i[1]), 
         .D(index_i[3]), .Z(n23525)) /* synthesis lut_function=(A (B (C)+!B !(C+!(D)))+!A (B (C)+!B !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21043_3_lut_4_lut_4_lut.init = 16'hc3d0;
    LUT4 mux_208_Mux_4_i340_3_lut_rep_848 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n32049)) /* synthesis lut_function=(A (B+!(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_4_i340_3_lut_rep_848.init = 16'hdada;
    LUT4 i21049_3_lut (.A(n396), .B(n29233), .C(index_i[3]), .Z(n23531)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21049_3_lut.init = 16'hcaca;
    LUT4 n589_bdd_4_lut (.A(n29084), .B(index_i[4]), .C(n28298), .D(index_i[5]), 
         .Z(n29027)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (B (C (D))+!B (C+!(D)))) */ ;
    defparam n589_bdd_4_lut.init = 16'hf099;
    LUT4 i23503_3_lut (.A(n716_adj_3491), .B(n731), .C(index_i[4]), .Z(n732)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23503_3_lut.init = 16'hcaca;
    LUT4 i23560_3_lut (.A(n23530), .B(n23531), .C(index_i[4]), .Z(n23532)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23560_3_lut.init = 16'hcaca;
    LUT4 i21046_3_lut (.A(n32040), .B(n32043), .C(index_i[3]), .Z(n23528)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21046_3_lut.init = 16'hcaca;
    LUT4 i23568_3_lut (.A(n23524), .B(n23525), .C(index_i[4]), .Z(n23526)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23568_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_2_i669_3_lut (.A(n653_adj_3492), .B(n475_adj_3470), 
         .C(index_i[4]), .Z(n669)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_2_i669_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_2_i605_3_lut (.A(n142_adj_3493), .B(n604_adj_3494), 
         .C(index_i[4]), .Z(n605_adj_3495)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_2_i605_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_5_i781_3_lut_4_lut_4_lut_else_4_lut (.A(index_i[3]), 
         .B(index_i[0]), .C(index_i[4]), .Z(n29527)) /* synthesis lut_function=(!(A (C)+!A (B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_5_i781_3_lut_4_lut_4_lut_else_4_lut.init = 16'h1f1f;
    LUT4 mux_208_Mux_2_i189_3_lut_3_lut_4_lut (.A(index_i[1]), .B(n29325), 
         .C(n173_adj_3496), .D(index_i[4]), .Z(n189_adj_3497)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(C+(D)))) */ ;
    defparam mux_208_Mux_2_i189_3_lut_3_lut_4_lut.init = 16'h77f0;
    PFUMX i27078 (.BLUT(n29490), .ALUT(n29491), .C0(index_i[0]), .Z(n29492));
    LUT4 i12768_2_lut_3_lut_4_lut (.A(index_i[1]), .B(n29325), .C(index_i[5]), 
         .D(index_i[4]), .Z(n508)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;
    defparam i12768_2_lut_3_lut_4_lut.init = 16'hf080;
    LUT4 i23510_3_lut (.A(n32058), .B(n23552), .C(index_i[4]), .Z(n23553)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23510_3_lut.init = 16'hcaca;
    LUT4 i25127_then_3_lut (.A(index_i[0]), .B(index_i[4]), .C(index_i[3]), 
         .Z(n29531)) /* synthesis lut_function=(A (B)+!A (B (C)+!B !(C))) */ ;
    defparam i25127_then_3_lut.init = 16'hc9c9;
    LUT4 i23512_3_lut (.A(n23548), .B(n23549), .C(index_i[4]), .Z(n23550)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23512_3_lut.init = 16'hcaca;
    LUT4 i21024_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n23506)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21024_3_lut_4_lut_4_lut.init = 16'hda5a;
    LUT4 mux_208_Mux_5_i505_3_lut_3_lut_rep_849 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n32050)) /* synthesis lut_function=(A (B+(C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_5_i505_3_lut_3_lut_rep_849.init = 16'hadad;
    LUT4 i21087_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n23569)) /* synthesis lut_function=(!(A (B (C (D))+!B (C (D)+!C !(D)))+!A !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21087_3_lut_4_lut_4_lut.init = 16'h5aad;
    LUT4 i22685_4_lut_4_lut (.A(n29082), .B(n29169), .C(index_i[5]), .D(index_i[4]), 
         .Z(n25186)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C+(D))+!B !(C (D)+!C !(D)))) */ ;
    defparam i22685_4_lut_4_lut.init = 16'hcf50;
    LUT4 mux_208_Mux_0_i796_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n796)) /* synthesis lut_function=(A (B (C+(D))+!B (C (D)))+!A !(B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_0_i796_3_lut_4_lut_4_lut.init = 16'hadc0;
    LUT4 i21037_3_lut (.A(n32046), .B(n29413), .C(index_i[3]), .Z(n23519)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21037_3_lut.init = 16'hcaca;
    LUT4 i22654_3_lut_4_lut (.A(n29076), .B(n29075), .C(index_i[5]), .D(index_i[6]), 
         .Z(n25155)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (B+((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i22654_3_lut_4_lut.init = 16'hffc5;
    LUT4 i25127_else_3_lut (.A(index_i[2]), .B(index_i[0]), .C(index_i[4]), 
         .D(index_i[3]), .Z(n29530)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)+!C !(D)))+!A (B (C+!(D))+!B !(C)))) */ ;
    defparam i25127_else_3_lut.init = 16'h1e38;
    LUT4 i21036_3_lut (.A(n32044), .B(n29242), .C(index_i[3]), .Z(n23518)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21036_3_lut.init = 16'hcaca;
    LUT4 i23581_3_lut (.A(n23518), .B(n23519), .C(index_i[4]), .Z(n23520)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23581_3_lut.init = 16'hcaca;
    LUT4 n53_bdd_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n26549)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n53_bdd_3_lut_4_lut_4_lut.init = 16'ha5ad;
    LUT4 i21034_3_lut (.A(n32048), .B(n29344), .C(index_i[3]), .Z(n23516)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21034_3_lut.init = 16'hcaca;
    LUT4 i21033_3_lut (.A(n29339), .B(n676), .C(index_i[3]), .Z(n23515)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21033_3_lut.init = 16'hcaca;
    LUT4 i23584_3_lut (.A(n23515), .B(n23516), .C(index_i[4]), .Z(n23517)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23584_3_lut.init = 16'hcaca;
    LUT4 n476_bdd_3_lut_25126 (.A(n476), .B(n26477), .C(index_i[5]), .Z(n26478)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n476_bdd_3_lut_25126.init = 16'hcaca;
    LUT4 mux_208_Mux_5_i308_3_lut_4_lut_3_lut_rep_850 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n32051)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_5_i308_3_lut_4_lut_3_lut_rep_850.init = 16'h4d4d;
    LUT4 i12729_2_lut_3_lut_4_lut (.A(n29156), .B(n29261), .C(index_i[6]), 
         .D(index_i[5]), .Z(n254)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i12729_2_lut_3_lut_4_lut.init = 16'hfef0;
    LUT4 mux_208_Mux_8_i763_3_lut_4_lut (.A(n29252), .B(n29363), .C(index_i[4]), 
         .D(n29151), .Z(n16890)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam mux_208_Mux_8_i763_3_lut_4_lut.init = 16'hfe0e;
    LUT4 mux_208_Mux_3_i653_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n653_adj_3498)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A !(B (D)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_3_i653_3_lut_4_lut_4_lut.init = 16'h4d99;
    LUT4 mux_208_Mux_4_i356_3_lut_rep_851 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n32052)) /* synthesis lut_function=(A (C)+!A !((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_4_i356_3_lut_rep_851.init = 16'ha4a4;
    LUT4 mux_208_Mux_2_i413_3_lut (.A(n397_adj_3499), .B(n954), .C(index_i[4]), 
         .Z(n413)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_2_i413_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_4_lut (.A(n29337), .B(n29325), .C(index_i[4]), .D(n29247), 
         .Z(n22136)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;
    defparam i1_3_lut_4_lut.init = 16'hfff8;
    LUT4 n53_bdd_3_lut_25892 (.A(n29343), .B(n32048), .C(index_i[3]), 
         .Z(n27645)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n53_bdd_3_lut_25892.init = 16'hcaca;
    LUT4 mux_208_Mux_0_i908_3_lut_4_lut_4_lut (.A(n29349), .B(n29255), .C(index_i[3]), 
         .D(index_i[0]), .Z(n908)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B ((D)+!C)+!B (C (D))))) */ ;
    defparam mux_208_Mux_0_i908_3_lut_4_lut_4_lut.init = 16'h5c0c;
    LUT4 i21067_3_lut (.A(n404), .B(n32051), .C(index_i[3]), .Z(n23549)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21067_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_2_i317_3_lut (.A(n668), .B(n316_adj_3500), .C(index_i[4]), 
         .Z(n317_adj_3501)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_2_i317_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_2_i286_3_lut (.A(n270_adj_3502), .B(n653_adj_3498), 
         .C(index_i[4]), .Z(n286)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_2_i286_3_lut.init = 16'hcaca;
    LUT4 index_i_2__bdd_4_lut_27866 (.A(index_i[2]), .B(index_i[0]), .C(index_i[4]), 
         .D(index_i[1]), .Z(n30481)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((C (D))+!B))) */ ;
    defparam index_i_2__bdd_4_lut_27866.init = 16'h0cec;
    LUT4 index_i_2__bdd_3_lut_27865 (.A(index_i[2]), .B(index_i[0]), .C(index_i[4]), 
         .Z(n30482)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B (C)+!B !(C)))) */ ;
    defparam index_i_2__bdd_3_lut_27865.init = 16'h6969;
    LUT4 n29253_bdd_3_lut_28201 (.A(n29182), .B(n32038), .C(index_i[4]), 
         .Z(n30484)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n29253_bdd_3_lut_28201.init = 16'hcaca;
    PFUMX i27139 (.BLUT(n29582), .ALUT(n29583), .C0(index_i[1]), .Z(n29584));
    LUT4 n172_bdd_3_lut_4_lut (.A(n29337), .B(index_i[2]), .C(index_i[3]), 
         .D(n29256), .Z(n26439)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n172_bdd_3_lut_4_lut.init = 16'hf707;
    LUT4 i24749_2_lut_rep_386_3_lut_4_lut (.A(n29337), .B(index_i[2]), .C(index_i[5]), 
         .D(n29261), .Z(n29046)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i24749_2_lut_rep_386_3_lut_4_lut.init = 16'h0f7f;
    LUT4 mux_208_Mux_8_i78_3_lut_4_lut (.A(n29337), .B(index_i[2]), .C(index_i[3]), 
         .D(n29256), .Z(n78)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_8_i78_3_lut_4_lut.init = 16'h8f80;
    LUT4 i21111_3_lut_3_lut_4_lut (.A(n29337), .B(index_i[2]), .C(n467), 
         .D(index_i[3]), .Z(n23593)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21111_3_lut_3_lut_4_lut.init = 16'hf077;
    LUT4 i23533_3_lut (.A(n142_adj_3503), .B(n15533), .C(index_i[4]), 
         .Z(n158)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23533_3_lut.init = 16'hcaca;
    PFUMX i24926 (.BLUT(n26549), .ALUT(n26548), .C0(index_i[4]), .Z(n26550));
    LUT4 mux_208_Mux_3_i828_3_lut_3_lut_4_lut_4_lut_4_lut (.A(n29337), .B(index_i[2]), 
         .C(index_i[4]), .D(index_i[3]), .Z(n828)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C (D)+!C !(D)))+!A !(B (C+!(D))+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_3_i828_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h70c7;
    LUT4 index_i_6__bdd_1_lut (.A(index_i[5]), .Z(n30596)) /* synthesis lut_function=(!(A)) */ ;
    defparam index_i_6__bdd_1_lut.init = 16'h5555;
    LUT4 index_i_6__bdd_4_lut_27901 (.A(index_i[6]), .B(index_i[5]), .C(index_i[1]), 
         .D(index_i[0]), .Z(n30597)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C))+!A (B (C)+!B !(C)))) */ ;
    defparam index_i_6__bdd_4_lut_27901.init = 16'h3cbc;
    LUT4 index_i_5__bdd_3_lut_28313 (.A(index_i[5]), .B(n30598), .C(index_i[3]), 
         .Z(n30599)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam index_i_5__bdd_3_lut_28313.init = 16'hcaca;
    LUT4 n29337_bdd_3_lut_28553 (.A(n29103), .B(index_i[6]), .C(index_i[5]), 
         .Z(n30600)) /* synthesis lut_function=(!(A (B)+!A (C))) */ ;
    defparam n29337_bdd_3_lut_28553.init = 16'h2727;
    LUT4 n29337_bdd_4_lut (.A(n29337), .B(index_i[6]), .C(index_i[2]), 
         .D(index_i[5]), .Z(n30601)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A !(B (C+(D))+!B (D)))) */ ;
    defparam n29337_bdd_4_lut.init = 16'h5fe0;
    LUT4 n30602_bdd_3_lut (.A(n30602), .B(n30599), .C(index_i[4]), .Z(n30603)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n30602_bdd_3_lut.init = 16'hcaca;
    LUT4 index_i_1__bdd_4_lut_28579 (.A(index_i[1]), .B(index_i[3]), .C(index_i[0]), 
         .D(index_i[2]), .Z(n30604)) /* synthesis lut_function=(A (B (C+(D))+!B (C (D)))+!A !(B (C)+!B !(C+(D)))) */ ;
    defparam index_i_1__bdd_4_lut_28579.init = 16'hbd94;
    LUT4 n30604_bdd_3_lut (.A(n30604), .B(index_i[1]), .C(index_i[4]), 
         .Z(n30605)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n30604_bdd_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_4_i348_3_lut (.A(n32049), .B(n29239), .C(index_i[3]), 
         .Z(n348)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_4_i348_3_lut.init = 16'hcaca;
    LUT4 i14492_2_lut_rep_373_3_lut_4_lut (.A(n29082), .B(index_i[4]), .C(index_i[6]), 
         .D(index_i[5]), .Z(n29033)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i14492_2_lut_rep_373_3_lut_4_lut.init = 16'hf080;
    LUT4 i21025_3_lut (.A(n32043), .B(n396), .C(index_i[3]), .Z(n23507)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21025_3_lut.init = 16'hcaca;
    LUT4 i23660_3_lut (.A(n23506), .B(n23507), .C(index_i[4]), .Z(n23508)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23660_3_lut.init = 16'hcaca;
    LUT4 i17714_4_lut (.A(index_i[0]), .B(index_i[4]), .C(index_i[1]), 
         .D(n29363), .Z(n286_adj_3504)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i17714_4_lut.init = 16'hccc8;
    LUT4 mux_208_Mux_0_i716_3_lut (.A(n29231), .B(n29412), .C(index_i[3]), 
         .Z(n716_adj_3505)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_0_i716_3_lut.init = 16'hcaca;
    LUT4 i23558_3_lut (.A(n23533), .B(n29485), .C(index_i[4]), .Z(n23535)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23558_3_lut.init = 16'hcaca;
    LUT4 n23278_bdd_3_lut_26842 (.A(n29037), .B(n701), .C(index_i[6]), 
         .Z(n27771)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n23278_bdd_3_lut_26842.init = 16'hacac;
    LUT4 i7128_2_lut (.A(phase_i[0]), .B(phase_i[10]), .Z(index_i_9__N_1748[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(60[14] 63[8])
    defparam i7128_2_lut.init = 16'h6666;
    LUT4 n26480_bdd_3_lut (.A(n29562), .B(n444_adj_3506), .C(index_i[5]), 
         .Z(n26481)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n26480_bdd_3_lut.init = 16'hcaca;
    LUT4 n27774_bdd_3_lut (.A(n31735), .B(n25183), .C(index_i[8]), .Z(n27775)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n27774_bdd_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_3_i924_3_lut (.A(n908_adj_3507), .B(index_i[0]), .C(index_i[4]), 
         .Z(n924_adj_3508)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_3_i924_3_lut.init = 16'hcaca;
    LUT4 i21021_3_lut (.A(n7), .B(n29229), .C(index_i[3]), .Z(n23503)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21021_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_3_i891_3_lut (.A(n541_adj_3509), .B(n890_adj_3510), 
         .C(index_i[4]), .Z(n891)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_3_i891_3_lut.init = 16'hcaca;
    LUT4 i21019_3_lut (.A(n723), .B(n396), .C(index_i[3]), .Z(n23501)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21019_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_3_i669_3_lut (.A(n653_adj_3498), .B(n668), .C(index_i[4]), 
         .Z(n669_adj_3511)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_3_i669_3_lut.init = 16'hcaca;
    PFUMX mux_208_Mux_2_i891 (.BLUT(n875), .ALUT(n890), .C0(index_i[4]), 
          .Z(n891_adj_3512)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 i11201_4_lut (.A(n29349), .B(n29182), .C(index_i[3]), .D(index_i[4]), 
         .Z(n13497)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B ((D)+!C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11201_4_lut.init = 16'h3afa;
    LUT4 i21112_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n23594)) /* synthesis lut_function=(!(A ((D)+!C)+!A !(B ((D)+!C)+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21112_3_lut_3_lut_4_lut.init = 16'h55a4;
    LUT4 i23570_3_lut (.A(n23521), .B(n23522), .C(index_i[4]), .Z(n23523)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23570_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_5_i483_rep_852 (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .Z(n32053)) /* synthesis lut_function=(!(A (C)+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_5_i483_rep_852.init = 16'h4a4a;
    LUT4 mux_208_Mux_3_i476_3_lut (.A(n460_adj_3513), .B(n285), .C(index_i[4]), 
         .Z(n476_adj_3514)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_3_i476_3_lut.init = 16'hcaca;
    PFUMX mux_208_Mux_2_i860 (.BLUT(n844_adj_3515), .ALUT(n859_adj_3516), 
          .C0(index_i[4]), .Z(n860_adj_3517)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 mux_208_Mux_5_i491_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n491)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A !(B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_5_i491_3_lut_4_lut_4_lut.init = 16'ha54a;
    LUT4 i14500_2_lut_3_lut_4_lut (.A(n29084), .B(index_i[4]), .C(index_i[6]), 
         .D(index_i[5]), .Z(n16936)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i14500_2_lut_3_lut_4_lut.init = 16'hfef0;
    LUT4 mux_208_Mux_6_i891_3_lut (.A(n78), .B(n890_adj_3518), .C(index_i[4]), 
         .Z(n891_adj_3519)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_6_i891_3_lut.init = 16'hcaca;
    LUT4 i21007_3_lut (.A(n29239), .B(n29228), .C(index_i[3]), .Z(n23489)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21007_3_lut.init = 16'hcaca;
    LUT4 n254_bdd_4_lut_26807 (.A(index_i[5]), .B(index_i[3]), .C(index_i[6]), 
         .D(index_i[4]), .Z(n27818)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;
    defparam n254_bdd_4_lut_26807.init = 16'hf8f0;
    LUT4 i21006_3_lut (.A(n32052), .B(n396), .C(index_i[3]), .Z(n23488)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21006_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_6_i828_4_lut (.A(n812_adj_3520), .B(n15423), .C(index_i[4]), 
         .D(index_i[2]), .Z(n828_adj_3521)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_6_i828_4_lut.init = 16'hfaca;
    LUT4 mux_208_Mux_2_i700_3_lut_4_lut (.A(index_i[1]), .B(n29363), .C(index_i[4]), 
         .D(n684_adj_3482), .Z(n700_adj_3522)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_2_i700_3_lut_4_lut.init = 16'hefe0;
    LUT4 i23672_3_lut (.A(n23488), .B(n23489), .C(index_i[4]), .Z(n23490)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23672_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_6_i797_3_lut (.A(n781), .B(n29043), .C(index_i[4]), 
         .Z(n797_adj_3523)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_6_i797_3_lut.init = 16'hcaca;
    LUT4 i21004_3_lut (.A(n32042), .B(n29413), .C(index_i[3]), .Z(n23486)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21004_3_lut.init = 16'hcaca;
    LUT4 i23676_3_lut (.A(n23485), .B(n23486), .C(index_i[4]), .Z(n23487)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23676_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_3_i1018_3_lut_4_lut (.A(index_i[1]), .B(n29363), .C(index_i[4]), 
         .D(n21724), .Z(n1018)) /* synthesis lut_function=(A (C+!(D))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_3_i1018_3_lut_4_lut.init = 16'he0ef;
    PFUMX mux_208_Mux_1_i891 (.BLUT(n882), .ALUT(n890_adj_3524), .C0(n29359), 
          .Z(n891_adj_3525)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 mux_208_Mux_6_i669_3_lut (.A(n653_adj_3526), .B(n668_adj_3527), 
         .C(index_i[4]), .Z(n669_adj_3528)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_6_i669_3_lut.init = 16'hcaca;
    LUT4 n27823_bdd_3_lut (.A(n29556), .B(n27819), .C(index_i[7]), .Z(n27824)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n27823_bdd_3_lut.init = 16'hcaca;
    LUT4 i23680_3_lut (.A(n23482), .B(n23483), .C(index_i[4]), .Z(n23484)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23680_3_lut.init = 16'hcaca;
    LUT4 i20997_3_lut (.A(n29228), .B(n32046), .C(index_i[3]), .Z(n23479)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20997_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_3_i413_3_lut (.A(n397_adj_3471), .B(n29414), .C(index_i[4]), 
         .Z(n413_adj_3529)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_3_i413_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_10_i574_4_lut_4_lut (.A(n29084), .B(index_i[4]), .C(index_i[5]), 
         .D(n29085), .Z(n574_adj_3530)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B !(C+(D))))) */ ;
    defparam mux_208_Mux_10_i574_4_lut_4_lut.init = 16'h1f1c;
    LUT4 mux_208_Mux_6_i542_3_lut (.A(n29230), .B(n541_adj_3509), .C(index_i[4]), 
         .Z(n542_adj_3531)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_6_i542_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_3_i286_4_lut (.A(n93), .B(index_i[2]), .C(index_i[4]), 
         .D(n15523), .Z(n286_adj_3532)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_3_i286_4_lut.init = 16'h3aca;
    LUT4 mux_208_Mux_5_i700_3_lut (.A(n460_adj_3533), .B(n32041), .C(index_i[4]), 
         .Z(n700_adj_3534)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_5_i700_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_6_i252_4_lut (.A(index_i[2]), .B(n251_adj_3485), .C(index_i[4]), 
         .D(n12501), .Z(n252_adj_3535)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_6_i252_4_lut.init = 16'hc5ca;
    LUT4 i20991_3_lut (.A(n396), .B(n32046), .C(index_i[3]), .Z(n23473)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20991_3_lut.init = 16'hcaca;
    LUT4 i24108_3_lut (.A(n28720), .B(n252_adj_3535), .C(index_i[5]), 
         .Z(n25106)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24108_3_lut.init = 16'hcaca;
    LUT4 i20989_3_lut (.A(n29242), .B(n32043), .C(index_i[3]), .Z(n23471)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20989_3_lut.init = 16'hcaca;
    LUT4 i20988_3_lut (.A(n29233), .B(n32044), .C(index_i[3]), .Z(n23470)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20988_3_lut.init = 16'hcaca;
    LUT4 i20986_3_lut (.A(n32051), .B(n32044), .C(index_i[3]), .Z(n23468)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20986_3_lut.init = 16'hcaca;
    PFUMX mux_208_Mux_3_i763 (.BLUT(n747_adj_3536), .ALUT(n762_adj_3476), 
          .C0(index_i[4]), .Z(n763)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 mux_208_Mux_3_i158_3_lut (.A(n142_adj_3493), .B(n29092), .C(index_i[4]), 
         .Z(n158_adj_3537)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_3_i158_3_lut.init = 16'hcaca;
    LUT4 i20982_3_lut (.A(n29228), .B(n32044), .C(index_i[3]), .Z(n23464)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20982_3_lut.init = 16'hcaca;
    LUT4 i20980_3_lut (.A(n29345), .B(n32048), .C(index_i[3]), .Z(n23462)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20980_3_lut.init = 16'hcaca;
    LUT4 n638_bdd_3_lut_26751 (.A(n638), .B(n23307), .C(index_i[7]), .Z(n27928)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n638_bdd_3_lut_26751.init = 16'hcaca;
    LUT4 index_i_7__bdd_4_lut_28237 (.A(index_i[7]), .B(n16816), .C(n28122), 
         .D(index_i[5]), .Z(n29030)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(B (C+(D))+!B !((D)+!C)))) */ ;
    defparam index_i_7__bdd_4_lut_28237.init = 16'h66f0;
    LUT4 i23599_3_lut (.A(n23461), .B(n23462), .C(index_i[4]), .Z(n23463)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23599_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_5_i31_3_lut (.A(n15_adj_3538), .B(n30), .C(index_i[4]), 
         .Z(n31)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_5_i31_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_4_i62_4_lut (.A(n29350), .B(n61), .C(index_i[4]), 
         .D(index_i[3]), .Z(n62)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_4_i62_4_lut.init = 16'hc5ca;
    LUT4 mux_208_Mux_4_i31_4_lut (.A(n15), .B(n29097), .C(index_i[4]), 
         .D(index_i[3]), .Z(n31_adj_3539)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_4_i31_4_lut.init = 16'h3aca;
    LUT4 i23576_3_lut (.A(n23458), .B(n23459), .C(index_i[4]), .Z(n23460)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23576_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_7_i620_3_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n620_adj_3540)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_7_i620_3_lut_4_lut_4_lut.init = 16'h85a5;
    LUT4 mux_208_Mux_3_i31_3_lut (.A(n781), .B(n30_adj_3541), .C(index_i[4]), 
         .Z(n31_adj_3542)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_3_i31_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_7_i490_3_lut_rep_826 (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[2]), .Z(n32027)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_7_i490_3_lut_rep_826.init = 16'h5858;
    LUT4 i20974_3_lut (.A(n404), .B(n29233), .C(index_i[3]), .Z(n23456)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20974_3_lut.init = 16'hcaca;
    LUT4 n29253_bdd_2_lut_4_lut (.A(index_i[1]), .B(index_i[0]), .C(index_i[2]), 
         .D(index_i[4]), .Z(n30485)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n29253_bdd_2_lut_4_lut.init = 16'h5800;
    LUT4 i20971_3_lut (.A(n404), .B(n29215), .C(index_i[3]), .Z(n23453)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20971_3_lut.init = 16'hcaca;
    LUT4 i20970_3_lut (.A(n29239), .B(n396), .C(index_i[3]), .Z(n23452)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20970_3_lut.init = 16'hcaca;
    LUT4 n23301_bdd_3_lut_26118 (.A(n382), .B(n509), .C(index_i[7]), .Z(n27930)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n23301_bdd_3_lut_26118.init = 16'hcaca;
    LUT4 n23301_bdd_3_lut (.A(n23301), .B(n30603), .C(index_i[7]), .Z(n27931)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n23301_bdd_3_lut.init = 16'hcaca;
    LUT4 index_i_0__bdd_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n32062)) /* synthesis lut_function=(A (B (D)+!B !((D)+!C))+!A !(B (C+!(D))+!B (D))) */ ;
    defparam index_i_0__bdd_4_lut.init = 16'h8c31;
    LUT4 i11214_3_lut (.A(n13509), .B(n32037), .C(index_i[3]), .Z(n13510)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11214_3_lut.init = 16'hcaca;
    LUT4 n24619_bdd_3_lut (.A(n24612), .B(n24613), .C(index_i[7]), .Z(n27951)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n24619_bdd_3_lut.init = 16'hcaca;
    LUT4 n24608_bdd_3_lut_26138 (.A(n24610), .B(n26482), .C(index_i[7]), 
         .Z(n27953)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n24608_bdd_3_lut_26138.init = 16'hcaca;
    LUT4 n24608_bdd_3_lut (.A(n24608), .B(n24609), .C(index_i[7]), .Z(n27954)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n24608_bdd_3_lut.init = 16'hcaca;
    PFUMX i21338 (.BLUT(n23818), .ALUT(n23819), .C0(index_i[5]), .Z(n23820));
    LUT4 i20968_3_lut (.A(n29239), .B(n29215), .C(index_i[3]), .Z(n23450)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20968_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_3_i125_3_lut (.A(n46_adj_3488), .B(n30_adj_3543), .C(index_i[4]), 
         .Z(n125)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_3_i125_3_lut.init = 16'hcaca;
    LUT4 i20967_3_lut (.A(n396), .B(n332), .C(index_i[3]), .Z(n23449)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20967_3_lut.init = 16'hcaca;
    PFUMX i21341 (.BLUT(n23821), .ALUT(n23822), .C0(index_i[5]), .Z(n23823));
    PFUMX mux_208_Mux_5_i732 (.BLUT(n13485), .ALUT(n731_adj_3544), .C0(index_i[4]), 
          .Z(n732_adj_3545)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 n589_bdd_3_lut_4_lut_4_lut (.A(n29218), .B(index_i[3]), .C(index_i[4]), 
         .D(n29182), .Z(n28302)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C))+!A !(B (C+(D))+!B (C))) */ ;
    defparam n589_bdd_3_lut_4_lut_4_lut.init = 16'h838f;
    LUT4 i22260_3_lut_3_lut_4_lut_4_lut (.A(n29218), .B(index_i[3]), .C(index_i[4]), 
         .D(n29156), .Z(n24761)) /* synthesis lut_function=(!(A (B (C)+!B ((D)+!C))+!A (B+((D)+!C)))) */ ;
    defparam i22260_3_lut_3_lut_4_lut_4_lut.init = 16'h0838;
    LUT4 n62_bdd_3_lut_4_lut (.A(n29218), .B(index_i[3]), .C(index_i[4]), 
         .D(n30_adj_3546), .Z(n28509)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;
    defparam n62_bdd_3_lut_4_lut.init = 16'hf808;
    LUT4 i21804_2_lut (.A(index_i[3]), .B(index_i[5]), .Z(n24305)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21804_2_lut.init = 16'h8888;
    LUT4 i11157_3_lut_4_lut_4_lut (.A(n29218), .B(index_i[3]), .C(index_i[5]), 
         .D(n29103), .Z(n13453)) /* synthesis lut_function=(A (B+(C (D)))+!A (B (C)+!B (C (D)))) */ ;
    defparam i11157_3_lut_4_lut_4_lut.init = 16'hf8c8;
    PFUMX i21350 (.BLUT(n23830), .ALUT(n23831), .C0(index_i[5]), .Z(n23832));
    LUT4 i24142_3_lut (.A(n542_adj_3547), .B(n573), .C(index_i[5]), .Z(n24600)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24142_3_lut.init = 16'hcaca;
    LUT4 i24165_3_lut (.A(n27453), .B(n23864), .C(index_i[5]), .Z(n23865)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24165_3_lut.init = 16'hcaca;
    LUT4 i19377_4_lut (.A(n29362), .B(n16886), .C(index_i[6]), .D(index_i[5]), 
         .Z(n21719)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D))))) */ ;
    defparam i19377_4_lut.init = 16'h3a35;
    LUT4 i24398_3_lut (.A(n21719), .B(n22136), .C(index_i[7]), .Z(n24542)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24398_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_7_i235_3_lut_rep_829 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n32030)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_7_i235_3_lut_rep_829.init = 16'he3e3;
    LUT4 mux_208_Mux_7_i541_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n541_adj_3548)) /* synthesis lut_function=(A (B (C)+!B ((D)+!C))+!A (B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_7_i541_3_lut_4_lut_4_lut.init = 16'he3c3;
    LUT4 i20953_3_lut (.A(n29340), .B(n141), .C(index_i[3]), .Z(n23435)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20953_3_lut.init = 16'hcaca;
    LUT4 i20952_3_lut (.A(n29240), .B(n32030), .C(index_i[3]), .Z(n23434)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20952_3_lut.init = 16'hcaca;
    LUT4 i20950_3_lut (.A(n29340), .B(n29214), .C(index_i[3]), .Z(n23432)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20950_3_lut.init = 16'hcaca;
    PFUMX i21353 (.BLUT(n23833), .ALUT(n23834), .C0(index_i[5]), .Z(n23835));
    PFUMX i21356 (.BLUT(n23836), .ALUT(n23837), .C0(index_i[5]), .Z(n23838));
    PFUMX i22844 (.BLUT(n557), .ALUT(n572), .C0(index_i[4]), .Z(n25345));
    PFUMX i21359 (.BLUT(n23839), .ALUT(n23840), .C0(index_i[5]), .Z(n23841));
    LUT4 index_i_4__bdd_4_lut_27395 (.A(index_i[4]), .B(n29162), .C(index_i[7]), 
         .D(n29152), .Z(n28122)) /* synthesis lut_function=(A ((C)+!B)+!A ((D)+!C)) */ ;
    defparam index_i_4__bdd_4_lut_27395.init = 16'hf7a7;
    LUT4 i12725_3_lut_4_lut (.A(n29033), .B(index_i[7]), .C(index_i[8]), 
         .D(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_1768[14])) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (D))) */ ;
    defparam i12725_3_lut_4_lut.init = 16'hffe0;
    PFUMX i21362 (.BLUT(n23842), .ALUT(n23843), .C0(index_i[5]), .Z(n23844));
    LUT4 mux_208_Mux_7_i412_3_lut (.A(n32030), .B(n32027), .C(index_i[3]), 
         .Z(n412_adj_3549)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_7_i412_3_lut.init = 16'hcaca;
    LUT4 i20949_3_lut (.A(n29341), .B(n141), .C(index_i[3]), .Z(n23431)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20949_3_lut.init = 16'hcaca;
    PFUMX i21365 (.BLUT(n23845), .ALUT(n23846), .C0(index_i[5]), .Z(n23847));
    PFUMX i21368 (.BLUT(n23848), .ALUT(n23849), .C0(index_i[5]), .Z(n23850));
    LUT4 mux_208_Mux_7_i173_3_lut (.A(n29240), .B(n29214), .C(index_i[3]), 
         .Z(n173_adj_3550)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_7_i173_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_6_i732_3_lut_4_lut (.A(n29339), .B(index_i[3]), .C(index_i[4]), 
         .D(n412_adj_3549), .Z(n732_adj_3551)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_6_i732_3_lut_4_lut.init = 16'hf909;
    PFUMX i20794 (.BLUT(n445), .ALUT(n508), .C0(index_i[6]), .Z(n23276));
    LUT4 mux_208_Mux_1_i732_3_lut (.A(n716), .B(n491), .C(index_i[4]), 
         .Z(n732_adj_3552)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_1_i732_3_lut.init = 16'hcaca;
    LUT4 i24370_3_lut (.A(n24668), .B(n28941), .C(index_i[6]), .Z(n24677)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24370_3_lut.init = 16'hcaca;
    LUT4 n26439_bdd_3_lut (.A(n26439), .B(n954), .C(index_i[4]), .Z(n28182)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n26439_bdd_3_lut.init = 16'hcaca;
    LUT4 i24306_3_lut (.A(n13454), .B(n892), .C(index_i[6]), .Z(n25154)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24306_3_lut.init = 16'hcaca;
    PFUMX i21371 (.BLUT(n23851), .ALUT(n23852), .C0(index_i[5]), .Z(n23853));
    LUT4 mux_208_Mux_6_i700_3_lut_4_lut (.A(n29339), .B(index_i[3]), .C(index_i[4]), 
         .D(n684_adj_3553), .Z(n700_adj_3554)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_6_i700_3_lut_4_lut.init = 16'h9f90;
    LUT4 mux_208_Mux_9_i62_3_lut_3_lut_4_lut_then_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[1]), .D(index_i[4]), .Z(n29546)) /* synthesis lut_function=(!(A (B+(C+!(D)))+!A !(B (D)+!B ((D)+!C)))) */ ;
    defparam mux_208_Mux_9_i62_3_lut_3_lut_4_lut_then_4_lut.init = 16'h5701;
    PFUMX i21374 (.BLUT(n23854), .ALUT(n23855), .C0(index_i[5]), .Z(n23856));
    LUT4 mux_208_Mux_9_i62_3_lut_3_lut_4_lut_else_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[1]), .D(index_i[4]), .Z(n29545)) /* synthesis lut_function=(A+(B (C+!(D))+!B !(D))) */ ;
    defparam mux_208_Mux_9_i62_3_lut_3_lut_4_lut_else_4_lut.init = 16'heaff;
    LUT4 mux_208_Mux_13_i511_4_lut_4_lut (.A(n29033), .B(index_i[7]), .C(index_i[8]), 
         .D(n254), .Z(n511)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (B (C+!(D))+!B !(C)))) */ ;
    defparam mux_208_Mux_13_i511_4_lut_4_lut.init = 16'h1c10;
    LUT4 i12806_4_lut (.A(n16658), .B(index_i[7]), .C(n16886), .D(index_i[6]), 
         .Z(n1021)) /* synthesis lut_function=(A (B+(C (D)))+!A (B+(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12806_4_lut.init = 16'hfcdd;
    LUT4 mux_208_Mux_10_i317_3_lut_3_lut_4_lut (.A(n29103), .B(index_i[3]), 
         .C(n29141), .D(index_i[4]), .Z(n317_adj_3555)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;
    defparam mux_208_Mux_10_i317_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 i22267_3_lut_4_lut (.A(n29156), .B(index_i[3]), .C(index_i[4]), 
         .D(n29150), .Z(n24768)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i22267_3_lut_4_lut.init = 16'hfe0e;
    LUT4 mux_208_Mux_10_i413_3_lut_3_lut_4_lut (.A(n29156), .B(index_i[3]), 
         .C(n29141), .D(index_i[4]), .Z(n413_adj_3556)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_10_i413_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 i21358_3_lut_3_lut_4_lut (.A(n29103), .B(index_i[3]), .C(n93_adj_3557), 
         .D(index_i[4]), .Z(n23840)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;
    defparam i21358_3_lut_3_lut_4_lut.init = 16'h11f0;
    LUT4 n124_bdd_3_lut_4_lut (.A(n29103), .B(index_i[3]), .C(index_i[4]), 
         .D(n93_adj_3557), .Z(n28507)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam n124_bdd_3_lut_4_lut.init = 16'hfe0e;
    LUT4 i22259_3_lut_3_lut_4_lut (.A(n29103), .B(index_i[3]), .C(n316), 
         .D(index_i[4]), .Z(n24760)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;
    defparam i22259_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 mux_208_Mux_0_i731_3_lut_4_lut (.A(n29252), .B(index_i[2]), .C(index_i[3]), 
         .D(n29340), .Z(n731_adj_3558)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_0_i731_3_lut_4_lut.init = 16'h4f40;
    LUT4 i22265_3_lut_3_lut_4_lut (.A(n29156), .B(index_i[3]), .C(n412_adj_3559), 
         .D(index_i[4]), .Z(n24766)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i22265_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 i21118_3_lut_4_lut (.A(n29252), .B(index_i[2]), .C(index_i[3]), 
         .D(n32045), .Z(n23600)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21118_3_lut_4_lut.init = 16'hf404;
    PFUMX i21377 (.BLUT(n23857), .ALUT(n23858), .C0(index_i[5]), .Z(n23859));
    LUT4 i14432_1_lut_2_lut_3_lut_4_lut (.A(n29156), .B(index_i[3]), .C(index_i[5]), 
         .D(index_i[4]), .Z(n381)) /* synthesis lut_function=(!(A (C+(D))+!A (B (C+(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i14432_1_lut_2_lut_3_lut_4_lut.init = 16'h010f;
    LUT4 n699_bdd_4_lut_24964_4_lut (.A(n29103), .B(index_i[3]), .C(index_i[2]), 
         .D(index_i[6]), .Z(n26606)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C+(D)))+!A (B ((D)+!C)+!B !((D)+!C))) */ ;
    defparam n699_bdd_4_lut_24964_4_lut.init = 16'hee3c;
    LUT4 mux_208_Mux_10_i637_3_lut_4_lut_4_lut (.A(n29169), .B(index_i[4]), 
         .C(index_i[5]), .D(n29084), .Z(n637)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B !(C+(D))))) */ ;
    defparam mux_208_Mux_10_i637_3_lut_4_lut_4_lut.init = 16'h1f1c;
    LUT4 i22175_3_lut (.A(n28920), .B(n24667), .C(index_i[6]), .Z(n24676)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22175_3_lut.init = 16'hcaca;
    PFUMX i21380 (.BLUT(n23860), .ALUT(n23861), .C0(index_i[5]), .Z(n23862));
    LUT4 i14502_3_lut_4_lut (.A(n29103), .B(index_i[3]), .C(n10789), .D(index_i[6]), 
         .Z(n16938)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (D))) */ ;
    defparam i14502_3_lut_4_lut.init = 16'hffe0;
    LUT4 i22656_3_lut (.A(n25150), .B(n25151), .C(index_i[7]), .Z(n25157)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22656_3_lut.init = 16'hcaca;
    LUT4 i22655_3_lut (.A(n25148), .B(n25149), .C(index_i[7]), .Z(n25156)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22655_3_lut.init = 16'hcaca;
    LUT4 i22660_3_lut (.A(n25158), .B(n25159), .C(index_i[8]), .Z(n25161)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22660_3_lut.init = 16'hcaca;
    LUT4 i22629_3_lut (.A(n25125), .B(n26609), .C(index_i[7]), .Z(n25130)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22629_3_lut.init = 16'hcaca;
    LUT4 i22621_3_lut (.A(n25109), .B(n26566), .C(index_i[6]), .Z(n25122)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22621_3_lut.init = 16'hcaca;
    LUT4 i22620_3_lut (.A(n26560), .B(n25108), .C(index_i[6]), .Z(n25121)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22620_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_0_i1002_3_lut_3_lut_4_lut (.A(n29252), .B(index_i[2]), 
         .C(n467), .D(index_i[3]), .Z(n1002)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_0_i1002_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 mux_208_Mux_6_i890_3_lut_3_lut_4_lut (.A(n29252), .B(index_i[2]), 
         .C(n29343), .D(index_i[3]), .Z(n890_adj_3518)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_6_i890_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 mux_208_Mux_3_i252_3_lut_4_lut (.A(n29098), .B(index_i[3]), .C(index_i[4]), 
         .D(n16734), .Z(n252_adj_3560)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;
    defparam mux_208_Mux_3_i252_3_lut_4_lut.init = 16'h08f8;
    LUT4 index_i_8__bdd_3_lut_26125_then_4_lut (.A(index_i[4]), .B(index_i[6]), 
         .C(index_i[5]), .D(n29082), .Z(n29555)) /* synthesis lut_function=(!(A (B (C+(D)))+!A (B (C)))) */ ;
    defparam index_i_8__bdd_3_lut_26125_then_4_lut.init = 16'h373f;
    LUT4 mux_208_Mux_3_i93_3_lut_4_lut (.A(n29252), .B(index_i[2]), .C(index_i[3]), 
         .D(n29256), .Z(n93)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_3_i93_3_lut_4_lut.init = 16'hefe0;
    LUT4 i22618_3_lut (.A(n26554), .B(n25104), .C(index_i[6]), .Z(n25119)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22618_3_lut.init = 16'hcaca;
    LUT4 i22537_3_lut_3_lut (.A(n29339), .B(index_i[3]), .C(n32048), .Z(n25038)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam i22537_3_lut_3_lut.init = 16'h7474;
    LUT4 mux_208_Mux_4_i668_3_lut_3_lut (.A(n29339), .B(index_i[3]), .C(n32048), 
         .Z(n668_adj_3561)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;
    defparam mux_208_Mux_4_i668_3_lut_3_lut.init = 16'hd1d1;
    LUT4 i22118_3_lut (.A(n24614), .B(n24615), .C(index_i[7]), .Z(n24619)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22118_3_lut.init = 16'hcaca;
    LUT4 i24006_3_lut (.A(n23572), .B(n23573), .C(index_i[4]), .Z(n23574)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24006_3_lut.init = 16'hcaca;
    LUT4 i22441_3_lut (.A(n24939), .B(n24940), .C(index_i[7]), .Z(n24942)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22441_3_lut.init = 16'hcaca;
    LUT4 i22440_3_lut (.A(n24937), .B(n24938), .C(index_i[7]), .Z(n24941)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22440_3_lut.init = 16'hcaca;
    LUT4 i22054_3_lut (.A(n24548), .B(n24549), .C(index_i[7]), .Z(n24555)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22054_3_lut.init = 16'hcaca;
    LUT4 i22053_3_lut (.A(n24546), .B(n24547), .C(index_i[7]), .Z(n24554)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22053_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_11_i766_3_lut (.A(n638_adj_3562), .B(n16938), .C(index_i[7]), 
         .Z(n766)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_11_i766_3_lut.init = 16'h3a3a;
    LUT4 i24444_3_lut (.A(n766), .B(n22122), .C(index_i[8]), .Z(n23066)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24444_3_lut.init = 16'hcaca;
    LUT4 index_i_8__bdd_3_lut_26125_else_4_lut (.A(n29162), .B(index_i[4]), 
         .C(index_i[6]), .D(index_i[5]), .Z(n29554)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;
    defparam index_i_8__bdd_3_lut_26125_else_4_lut.init = 16'hf080;
    LUT4 mux_208_Mux_8_i860_3_lut_4_lut (.A(n29098), .B(index_i[3]), .C(index_i[4]), 
         .D(n29151), .Z(n860)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;
    defparam mux_208_Mux_8_i860_3_lut_4_lut.init = 16'h08f8;
    LUT4 mux_208_Mux_10_i62_3_lut_3_lut_4_lut (.A(n29098), .B(index_i[3]), 
         .C(n29151), .D(index_i[4]), .Z(n62_adj_3563)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C+!(D))) */ ;
    defparam mux_208_Mux_10_i62_3_lut_3_lut_4_lut.init = 16'hf077;
    LUT4 i22872_3_lut (.A(n25370), .B(n25371), .C(index_i[7]), .Z(n25373)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22872_3_lut.init = 16'hcaca;
    LUT4 i22871_3_lut (.A(n25368), .B(n25369), .C(index_i[7]), .Z(n25372)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22871_3_lut.init = 16'hcaca;
    LUT4 i24429_3_lut (.A(n25156), .B(n25157), .C(index_i[8]), .Z(n25160)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24429_3_lut.init = 16'hcaca;
    LUT4 n62_bdd_3_lut (.A(n62_adj_3563), .B(n125_adj_3564), .C(index_i[6]), 
         .Z(n31732)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n62_bdd_3_lut.init = 16'hcaca;
    LUT4 n25186_bdd_4_lut (.A(n252_adj_3565), .B(n29152), .C(index_i[4]), 
         .D(index_i[5]), .Z(n31730)) /* synthesis lut_function=(A (B (D)+!B ((D)+!C))+!A !(B+(C+(D)))) */ ;
    defparam n25186_bdd_4_lut.init = 16'haa03;
    LUT4 n62_bdd_4_lut (.A(n29363), .B(n29162), .C(index_i[6]), .D(index_i[4]), 
         .Z(n31733)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C+(D)))+!A (B ((D)+!C)+!B !(C)))) */ ;
    defparam n62_bdd_4_lut.init = 16'h3af0;
    LUT4 i22087_3_lut (.A(n24583), .B(n28184), .C(index_i[7]), .Z(n24588)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22087_3_lut.init = 16'hcaca;
    LUT4 i22086_3_lut (.A(n24581), .B(n24582), .C(index_i[7]), .Z(n24587)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22086_3_lut.init = 16'hcaca;
    LUT4 i24470_3_lut (.A(n24587), .B(n24588), .C(index_i[8]), .Z(n24590)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24470_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut (.A(index_i[7]), .B(n29035), .C(index_i[6]), .D(index_i[8]), 
         .Z(n22166)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_4_lut.init = 16'hfffe;
    LUT4 i14498_2_lut_rep_375_3_lut_4_lut (.A(n29098), .B(index_i[3]), .C(index_i[5]), 
         .D(index_i[4]), .Z(n29035)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;
    defparam i14498_2_lut_rep_375_3_lut_4_lut.init = 16'hf080;
    LUT4 i20583_3_lut (.A(n28127), .B(n23277), .C(index_i[8]), .Z(n23065)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20583_3_lut.init = 16'hcaca;
    LUT4 index_i_6__bdd_3_lut_25413_rep_395_4_lut (.A(n29098), .B(index_i[3]), 
         .C(index_i[4]), .D(n29060), .Z(n29055)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam index_i_6__bdd_3_lut_25413_rep_395_4_lut.init = 16'h8f80;
    LUT4 mux_208_Mux_3_i189_3_lut_3_lut_4_lut (.A(n29098), .B(index_i[3]), 
         .C(index_i[4]), .D(n29141), .Z(n189_adj_3566)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;
    defparam mux_208_Mux_3_i189_3_lut_3_lut_4_lut.init = 16'h08f8;
    LUT4 i12754_4_lut (.A(n16936), .B(index_i[8]), .C(n16938), .D(index_i[7]), 
         .Z(n1022)) /* synthesis lut_function=(A (B+(C (D)))+!A (B+(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12754_4_lut.init = 16'hfcdd;
    LUT4 mux_208_Mux_3_i221_3_lut_4_lut (.A(n29182), .B(index_i[3]), .C(index_i[4]), 
         .D(n29152), .Z(n221)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;
    defparam mux_208_Mux_3_i221_3_lut_4_lut.init = 16'h08f8;
    LUT4 i22413_3_lut_4_lut (.A(n29182), .B(index_i[3]), .C(index_i[4]), 
         .D(n46), .Z(n24914)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam i22413_3_lut_4_lut.init = 16'h8f80;
    LUT4 i22414_3_lut_3_lut_4_lut (.A(n29182), .B(index_i[3]), .C(n93_adj_3567), 
         .D(index_i[4]), .Z(n24915)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C+!(D))) */ ;
    defparam i22414_3_lut_3_lut_4_lut.init = 16'hf077;
    LUT4 i21079_3_lut_4_lut (.A(n29219), .B(index_i[2]), .C(index_i[3]), 
         .D(n29242), .Z(n23561)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21079_3_lut_4_lut.init = 16'hf606;
    LUT4 i20992_3_lut_4_lut (.A(n29219), .B(index_i[2]), .C(index_i[3]), 
         .D(n32043), .Z(n23474)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20992_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_208_Mux_3_i460_3_lut_4_lut (.A(n29219), .B(index_i[2]), .C(index_i[3]), 
         .D(n29229), .Z(n460_adj_3513)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_3_i460_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_208_Mux_6_i285_3_lut_4_lut (.A(n29219), .B(index_i[2]), .C(index_i[3]), 
         .D(n32041), .Z(n285)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_6_i285_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_208_Mux_1_i700_3_lut_4_lut (.A(n29417), .B(index_i[3]), .C(index_i[4]), 
         .D(n684), .Z(n700)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_1_i700_3_lut_4_lut.init = 16'hefe0;
    LUT4 n124_bdd_3_lut_26575_4_lut (.A(n29349), .B(index_i[3]), .C(index_i[4]), 
         .D(n124_adj_3568), .Z(n28506)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n124_bdd_3_lut_26575_4_lut.init = 16'hf101;
    LUT4 mux_208_Mux_4_i573_3_lut_4_lut_4_lut_4_lut (.A(n29349), .B(index_i[3]), 
         .C(n29156), .D(index_i[4]), .Z(n573)) /* synthesis lut_function=(!(A (B (D)+!B ((D)+!C))+!A (B (D)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_4_i573_3_lut_4_lut_4_lut_4_lut.init = 16'h11fc;
    LUT4 mux_208_Mux_10_i252_3_lut_4_lut_4_lut (.A(n29182), .B(index_i[3]), 
         .C(index_i[4]), .D(n29156), .Z(n252_adj_3565)) /* synthesis lut_function=(!(A (B (C)+!B !(C+(D)))+!A !(B+(C+(D))))) */ ;
    defparam mux_208_Mux_10_i252_3_lut_4_lut_4_lut.init = 16'h7f7c;
    LUT4 i22182_3_lut (.A(n24680), .B(n24681), .C(index_i[8]), .Z(n24683)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22182_3_lut.init = 16'hcaca;
    LUT4 i22181_3_lut (.A(n24678), .B(n24679), .C(index_i[8]), .Z(n24682)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22181_3_lut.init = 16'hcaca;
    LUT4 i22258_3_lut_4_lut (.A(n29349), .B(index_i[3]), .C(index_i[4]), 
         .D(n285_adj_3569), .Z(n24759)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i22258_3_lut_4_lut.init = 16'hfe0e;
    LUT4 mux_208_Mux_10_i125_3_lut_4_lut_4_lut (.A(n29349), .B(index_i[3]), 
         .C(index_i[4]), .D(n29182), .Z(n125_adj_3564)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B (C (D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_10_i125_3_lut_4_lut_4_lut.init = 16'h3efe;
    PFUMX i11160 (.BLUT(n13559), .ALUT(n13560), .C0(n24132), .Z(n13456));
    LUT4 i21126_3_lut (.A(n29413), .B(n29226), .C(index_i[3]), .Z(n23608)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21126_3_lut.init = 16'hcaca;
    LUT4 i22151_3_lut (.A(n24649), .B(n24650), .C(index_i[8]), .Z(n24652)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22151_3_lut.init = 16'hcaca;
    LUT4 i22150_3_lut (.A(n24647), .B(n24648), .C(index_i[8]), .Z(n24651)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22150_3_lut.init = 16'hcaca;
    LUT4 i22088_3_lut (.A(n24585), .B(n24586), .C(index_i[8]), .Z(n24589)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22088_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_2_i573_3_lut_3_lut_4_lut (.A(n29349), .B(index_i[3]), 
         .C(n557_adj_3570), .D(index_i[4]), .Z(n573_adj_3571)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_2_i573_3_lut_3_lut_4_lut.init = 16'h11f0;
    LUT4 mux_208_Mux_3_i573_3_lut_3_lut_4_lut (.A(n29349), .B(index_i[3]), 
         .C(n397), .D(index_i[4]), .Z(n573_adj_3572)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_3_i573_3_lut_3_lut_4_lut.init = 16'h11f0;
    LUT4 i24481_3_lut (.A(n574_adj_3530), .B(n637), .C(index_i[6]), .Z(n23278)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24481_3_lut.init = 16'hcaca;
    LUT4 i22213_3_lut (.A(n24711), .B(n24712), .C(index_i[8]), .Z(n24714)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22213_3_lut.init = 16'hcaca;
    LUT4 i22212_3_lut (.A(n24709), .B(n24710), .C(index_i[8]), .Z(n24713)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22212_3_lut.init = 16'hcaca;
    LUT4 n476_bdd_3_lut_24865_4_lut (.A(index_i[2]), .B(n29252), .C(index_i[4]), 
         .D(n491_adj_3573), .Z(n26477)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+(D)))) */ ;
    defparam n476_bdd_3_lut_24865_4_lut.init = 16'h9f90;
    LUT4 i21042_3_lut_3_lut_4_lut (.A(index_i[2]), .B(n29252), .C(n29214), 
         .D(index_i[3]), .Z(n23524)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (B (C (D))+!B (C+!(D)))) */ ;
    defparam i21042_3_lut_3_lut_4_lut.init = 16'hf099;
    LUT4 mux_208_Mux_3_i860_3_lut_4_lut (.A(index_i[2]), .B(n29252), .C(index_i[4]), 
         .D(n859), .Z(n860_adj_3574)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam mux_208_Mux_3_i860_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_208_Mux_7_i443_3_lut_4_lut (.A(index_i[2]), .B(n29252), .C(index_i[3]), 
         .D(n32030), .Z(n443_adj_3575)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;
    defparam mux_208_Mux_7_i443_3_lut_4_lut.init = 16'h6f60;
    LUT4 i20976_3_lut_3_lut_4_lut (.A(index_i[2]), .B(n29252), .C(n32030), 
         .D(index_i[3]), .Z(n23458)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (B (C (D))+!B (C+!(D)))) */ ;
    defparam i20976_3_lut_3_lut_4_lut.init = 16'hf099;
    LUT4 i11235_3_lut_then_4_lut (.A(index_i[4]), .B(index_i[0]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n32064)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11235_3_lut_then_4_lut.init = 16'hd4a5;
    LUT4 index_i_0__bdd_4_lut_28945 (.A(index_i[0]), .B(index_i[3]), .C(index_i[1]), 
         .D(index_i[2]), .Z(n32058)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C (D)))+!A !(B (C+!(D))+!B !(C+(D))))) */ ;
    defparam index_i_0__bdd_4_lut_28945.init = 16'h4ae7;
    LUT4 i21121_3_lut_4_lut (.A(n29337), .B(index_i[2]), .C(index_i[3]), 
         .D(n29233), .Z(n23603)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21121_3_lut_4_lut.init = 16'hdfd0;
    LUT4 i22106_4_lut (.A(n23514), .B(n1002_adj_3576), .C(index_i[5]), 
         .D(index_i[4]), .Z(n24607)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;
    defparam i22106_4_lut.init = 16'hfaca;
    LUT4 mux_208_Mux_4_i860_3_lut (.A(n506), .B(n26552), .C(index_i[4]), 
         .Z(n860_adj_3577)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_4_i860_3_lut.init = 16'hcaca;
    LUT4 i24866_then_4_lut (.A(index_i[0]), .B(index_i[4]), .C(index_i[1]), 
         .D(index_i[3]), .Z(n29561)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam i24866_then_4_lut.init = 16'h3c69;
    LUT4 i24866_else_4_lut (.A(index_i[0]), .B(index_i[4]), .C(index_i[1]), 
         .D(index_i[3]), .Z(n29560)) /* synthesis lut_function=(!(A (B (C)+!B !(C (D)+!C !(D)))+!A (B ((D)+!C)+!B !((D)+!C)))) */ ;
    defparam i24866_else_4_lut.init = 16'h394b;
    LUT4 n699_bdd_4_lut (.A(n29056), .B(index_i[6]), .C(n29151), .D(index_i[5]), 
         .Z(n28519)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C+!(D))+!B (D))) */ ;
    defparam n699_bdd_4_lut.init = 16'hd1cc;
    LUT4 n28522_bdd_3_lut (.A(n28522), .B(n28519), .C(index_i[4]), .Z(n23307)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n28522_bdd_3_lut.init = 16'hcaca;
    LUT4 n27772_bdd_3_lut_3_lut (.A(n1021), .B(index_i[8]), .C(n27772), 
         .Z(n27773)) /* synthesis lut_function=(A (B+(C))+!A !(B+!(C))) */ ;
    defparam n27772_bdd_3_lut_3_lut.init = 16'hb8b8;
    PFUMX i22409 (.BLUT(n24906), .ALUT(n24907), .C0(index_i[4]), .Z(n24910));
    LUT4 i23662_3_lut (.A(n23503), .B(n23504), .C(index_i[4]), .Z(n23505)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23662_3_lut.init = 16'hcaca;
    LUT4 n26779_bdd_3_lut (.A(n26779), .B(n476), .C(index_i[5]), .Z(n26780)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n26779_bdd_3_lut.init = 16'hcaca;
    LUT4 i11235_3_lut_else_4_lut (.A(index_i[4]), .B(index_i[0]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n32063)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A !(B (C (D)+!C !(D))+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11235_3_lut_else_4_lut.init = 16'h5a95;
    LUT4 i13040_3_lut_rep_831 (.A(index_i[2]), .B(index_i[1]), .C(index_i[0]), 
         .Z(n32032)) /* synthesis lut_function=(!(A (B)+!A (B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i13040_3_lut_rep_831.init = 16'h2323;
    PFUMX i22410 (.BLUT(n24908), .ALUT(n24909), .C0(index_i[4]), .Z(n24911));
    LUT4 mux_208_Mux_2_i908_3_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[1]), 
         .C(index_i[0]), .D(index_i[3]), .Z(n908_adj_3578)) /* synthesis lut_function=(!(A (B)+!A !(B (D)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_2_i908_3_lut_4_lut_4_lut.init = 16'h6623;
    LUT4 mux_208_Mux_0_i653_3_lut (.A(n29214), .B(n29413), .C(index_i[3]), 
         .Z(n653_adj_3579)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_0_i653_3_lut.init = 16'hcaca;
    LUT4 i21108_3_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[1]), .C(index_i[0]), 
         .D(index_i[3]), .Z(n23590)) /* synthesis lut_function=(!(A (B (D)+!B !(D))+!A (B+(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21108_3_lut_4_lut_4_lut.init = 16'h2388;
    LUT4 n26783_bdd_3_lut (.A(n29532), .B(n26781), .C(index_i[5]), .Z(n26784)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n26783_bdd_3_lut.init = 16'hcaca;
    PFUMX i27076 (.BLUT(n29487), .ALUT(n29488), .C0(index_i[0]), .Z(n29489));
    LUT4 mux_208_Mux_5_i124_3_lut (.A(n29214), .B(n29345), .C(index_i[3]), 
         .Z(n124_adj_3580)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_5_i124_3_lut.init = 16'hcaca;
    LUT4 i22553_3_lut (.A(n141), .B(n32027), .C(index_i[3]), .Z(n25054)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22553_3_lut.init = 16'hcaca;
    LUT4 i20994_3_lut_4_lut (.A(index_i[0]), .B(n29349), .C(index_i[3]), 
         .D(n29229), .Z(n23476)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A ((D)+!C)) */ ;
    defparam i20994_3_lut_4_lut.init = 16'hfd0d;
    LUT4 i23664_3_lut (.A(n23500), .B(n23501), .C(index_i[4]), .Z(n23502)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23664_3_lut.init = 16'hcaca;
    LUT4 i22552_3_lut (.A(n676), .B(n29340), .C(index_i[3]), .Z(n25053)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22552_3_lut.init = 16'hcaca;
    LUT4 i22551_3_lut (.A(n32032), .B(n29339), .C(index_i[3]), .Z(n25052)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22551_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_4_i700_3_lut (.A(n684_adj_3581), .B(index_i[1]), .C(index_i[4]), 
         .Z(n700_adj_3582)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_4_i700_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_4_i669_3_lut (.A(n781), .B(n668_adj_3561), .C(index_i[4]), 
         .Z(n669_adj_3583)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_4_i669_3_lut.init = 16'hcaca;
    LUT4 i22550_3_lut (.A(n32027), .B(n29257), .C(index_i[3]), .Z(n25051)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22550_3_lut.init = 16'hcaca;
    LUT4 i22546_3_lut (.A(n29237), .B(n29257), .C(index_i[3]), .Z(n25047)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22546_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_4_i542_3_lut (.A(n30_adj_3543), .B(n506_adj_3584), 
         .C(index_i[4]), .Z(n542_adj_3547)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_4_i542_3_lut.init = 16'hcaca;
    LUT4 i22100_4_lut (.A(n29189), .B(n29526), .C(index_i[5]), .D(index_i[4]), 
         .Z(n24601)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam i22100_4_lut.init = 16'hc5ca;
    LUT4 i22545_3_lut (.A(n32032), .B(n108), .C(index_i[3]), .Z(n25046)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22545_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_1_i986_3_lut (.A(n29340), .B(n32038), .C(index_i[3]), 
         .Z(n986_adj_3585)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_1_i986_3_lut.init = 16'hcaca;
    LUT4 i22544_3_lut (.A(n676), .B(n29339), .C(index_i[3]), .Z(n25045)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22544_3_lut.init = 16'hcaca;
    LUT4 i22543_3_lut (.A(n29214), .B(n29240), .C(index_i[3]), .Z(n25044)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22543_3_lut.init = 16'hcaca;
    LUT4 i12876_2_lut_rep_552 (.A(index_i[0]), .B(index_i[1]), .Z(n29212)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12876_2_lut_rep_552.init = 16'h4444;
    LUT4 i22539_3_lut (.A(n29257), .B(n29341), .C(index_i[3]), .Z(n25040)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22539_3_lut.init = 16'hcaca;
    LUT4 i22538_3_lut (.A(n467), .B(n29237), .C(index_i[3]), .Z(n25039)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22538_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_4_i286_3_lut (.A(n270), .B(n15), .C(index_i[4]), 
         .Z(n286_adj_3586)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_4_i286_3_lut.init = 16'hcaca;
    LUT4 i22536_3_lut (.A(n29341), .B(n29214), .C(index_i[3]), .Z(n25037)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22536_3_lut.init = 16'hcaca;
    LUT4 i20998_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n23480)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A (B (C (D)+!C !(D))+!B (D))) */ ;
    defparam i20998_3_lut_4_lut.init = 16'hd926;
    LUT4 mux_208_Mux_4_i94_3_lut (.A(n61), .B(n29415), .C(index_i[4]), 
         .Z(n94_adj_3587)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_4_i94_3_lut.init = 16'hcaca;
    PFUMX i22416 (.BLUT(n142), .ALUT(n157_adj_3588), .C0(index_i[4]), 
          .Z(n24917));
    LUT4 mux_208_Mux_8_i15_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n15_adj_3589)) /* synthesis lut_function=(A (B (C)+!B !(C (D)+!C !(D)))+!A !(B ((D)+!C)+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_8_i15_3_lut_4_lut_4_lut.init = 16'h83e0;
    LUT4 mux_208_Mux_0_i954_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n954_adj_3590)) /* synthesis lut_function=(A (D)+!A !(B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_0_i954_3_lut_4_lut_4_lut.init = 16'haf40;
    LUT4 mux_208_Mux_6_i636_4_lut_4_lut (.A(index_i[1]), .B(index_i[4]), 
         .C(n635_adj_3591), .D(n16239), .Z(n636_adj_3592)) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_6_i636_4_lut_4_lut.init = 16'hf3d1;
    LUT4 i23658_3_lut_then_4_lut (.A(index_i[2]), .B(n29337), .C(index_i[3]), 
         .D(n29339), .Z(n29567)) /* synthesis lut_function=(A (C+(D))+!A !(B (C+!(D))+!B !(C+(D)))) */ ;
    defparam i23658_3_lut_then_4_lut.init = 16'hbfb0;
    PFUMX i22417 (.BLUT(n173), .ALUT(n188), .C0(index_i[4]), .Z(n24918));
    LUT4 mux_208_Mux_0_i620_3_lut (.A(n29340), .B(n32037), .C(index_i[3]), 
         .Z(n620_adj_3593)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_0_i620_3_lut.init = 16'hcaca;
    LUT4 n476_bdd_3_lut_25942_3_lut (.A(index_i[1]), .B(index_i[4]), .C(n124_adj_3580), 
         .Z(n26779)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n476_bdd_3_lut_25942_3_lut.init = 16'hd1d1;
    LUT4 mux_208_Mux_3_i349_3_lut_3_lut (.A(index_i[1]), .B(index_i[4]), 
         .C(n348_adj_3594), .Z(n349_adj_3595)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_3_i349_3_lut_3_lut.init = 16'hd1d1;
    LUT4 i12998_2_lut_rep_547_2_lut (.A(index_i[1]), .B(index_i[0]), .Z(n29207)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12998_2_lut_rep_547_2_lut.init = 16'h4444;
    LUT4 i21357_3_lut_4_lut (.A(n29156), .B(n29103), .C(index_i[3]), .D(index_i[4]), 
         .Z(n23839)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C (D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21357_3_lut_4_lut.init = 16'hf03a;
    LUT4 n396_bdd_3_lut_26821 (.A(n29339), .B(n467), .C(index_i[3]), .Z(n28758)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B+(C)))) */ ;
    defparam n396_bdd_3_lut_26821.init = 16'h5c5c;
    LUT4 mux_208_Mux_6_i411_3_lut_4_lut_4_lut_3_lut_rep_555 (.A(index_i[1]), 
         .B(index_i[2]), .C(index_i[0]), .Z(n29215)) /* synthesis lut_function=(!(A (B+(C))+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_6_i411_3_lut_4_lut_4_lut_3_lut_rep_555.init = 16'h4242;
    LUT4 mux_208_Mux_0_i491_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .D(index_i[3]), .Z(n491_adj_3596)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !(B (C)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_0_i491_3_lut_4_lut.init = 16'h42f0;
    LUT4 i14253_2_lut_rep_558 (.A(index_i[1]), .B(index_i[2]), .Z(n29218)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14253_2_lut_rep_558.init = 16'heeee;
    LUT4 mux_208_Mux_9_i93_3_lut_3_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .Z(n93_adj_3557)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B !(C))) */ ;
    defparam mux_208_Mux_9_i93_3_lut_3_lut_3_lut.init = 16'hc1c1;
    L6MUX21 i25205 (.D0(n26870), .D1(n26867), .SD(index_i[5]), .Z(n26871));
    LUT4 i12918_2_lut_rep_437_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[0]), 
         .Z(n29097)) /* synthesis lut_function=(A (C)+!A ((C)+!B)) */ ;
    defparam i12918_2_lut_rep_437_3_lut.init = 16'hf1f1;
    LUT4 n396_bdd_3_lut_26921 (.A(n32048), .B(n32032), .C(index_i[3]), 
         .Z(n28759)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n396_bdd_3_lut_26921.init = 16'hcaca;
    PFUMX i25203 (.BLUT(n26869), .ALUT(n26868), .C0(index_i[4]), .Z(n26870));
    LUT4 i21100_3_lut (.A(n32050), .B(n29234), .C(index_i[3]), .Z(n23582)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21100_3_lut.init = 16'hcaca;
    LUT4 i14441_2_lut_rep_509_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[3]), 
         .Z(n29169)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i14441_2_lut_rep_509_3_lut.init = 16'he0e0;
    LUT4 mux_208_Mux_5_i891_3_lut (.A(n875_adj_3597), .B(n379_adj_3598), 
         .C(index_i[4]), .Z(n891_adj_3599)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_5_i891_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_5_i860_3_lut (.A(n15_adj_3538), .B(n859_adj_3600), 
         .C(index_i[4]), .Z(n860_adj_3601)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_5_i860_3_lut.init = 16'hcaca;
    LUT4 i14443_2_lut_rep_423_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[4]), .D(index_i[3]), .Z(n29083)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i14443_2_lut_rep_423_3_lut_4_lut.init = 16'hfef0;
    PFUMX i25200 (.BLUT(n26866), .ALUT(n26865), .C0(index_i[4]), .Z(n26867));
    LUT4 i21127_3_lut_3_lut_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[3]), 
         .Z(n23609)) /* synthesis lut_function=(A (C)+!A (B+!(C))) */ ;
    defparam i21127_3_lut_3_lut_3_lut.init = 16'he5e5;
    LUT4 i12996_2_lut_rep_559 (.A(index_i[0]), .B(index_i[1]), .Z(n29219)) /* synthesis lut_function=((B)+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12996_2_lut_rep_559.init = 16'hdddd;
    LUT4 i22412_3_lut (.A(n541_adj_3548), .B(n32062), .C(index_i[4]), 
         .Z(n24913)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22412_3_lut.init = 16'hcaca;
    LUT4 i23658_3_lut_else_4_lut (.A(n29255), .B(n676), .C(index_i[3]), 
         .Z(n29566)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23658_3_lut_else_4_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_1_i908_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n908_adj_3602)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+(D)))+!A (B (C+(D))+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_1_i908_3_lut_4_lut_4_lut_4_lut.init = 16'h332d;
    LUT4 mux_208_Mux_0_i635_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n635_adj_3603)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_0_i635_3_lut_4_lut_4_lut.init = 16'hfd0a;
    LUT4 i21093_3_lut (.A(n29229), .B(n32046), .C(index_i[3]), .Z(n23575)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21093_3_lut.init = 16'hcaca;
    LUT4 i23520_3_lut (.A(n23545), .B(n23546), .C(index_i[4]), .Z(n23547)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23520_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_0_i157_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n157_adj_3588)) /* synthesis lut_function=(A (B (C+!(D))+!B !(D))+!A (B (D)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_0_i157_3_lut_4_lut.init = 16'hd4aa;
    LUT4 i23713_3_lut (.A(n23476), .B(n23477), .C(index_i[4]), .Z(n23478)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23713_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_5_i636_4_lut (.A(n157_adj_3604), .B(n29208), .C(index_i[4]), 
         .D(index_i[3]), .Z(n636_adj_3605)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_5_i636_4_lut.init = 16'h3aca;
    LUT4 i5339_2_lut_rep_561 (.A(index_i[0]), .B(index_i[2]), .Z(n29221)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i5339_2_lut_rep_561.init = 16'h6666;
    LUT4 i23716_3_lut (.A(n19995), .B(n19996), .C(index_i[4]), .Z(n19997)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23716_3_lut.init = 16'hcaca;
    L6MUX21 i26995 (.D0(n28940), .D1(n28938), .SD(index_i[5]), .Z(n28941));
    LUT4 mux_208_Mux_5_i507_3_lut (.A(n491), .B(n506), .C(index_i[4]), 
         .Z(n507)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_5_i507_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_0_i589_3_lut (.A(n29257), .B(n7), .C(index_i[3]), 
         .Z(n589)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_0_i589_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_5_i476_3_lut (.A(n460_adj_3533), .B(n475_adj_3474), 
         .C(index_i[4]), .Z(n476_adj_3606)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_5_i476_3_lut.init = 16'hcaca;
    LUT4 i23994_3_lut (.A(n23608), .B(n23609), .C(index_i[4]), .Z(n23610)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23994_3_lut.init = 16'hcaca;
    PFUMX i26993 (.BLUT(n572_adj_3607), .ALUT(n28939), .C0(index_i[4]), 
          .Z(n28940));
    PFUMX i26990 (.BLUT(n28937), .ALUT(n28936), .C0(index_i[4]), .Z(n28938));
    LUT4 mux_208_Mux_5_i413_3_lut (.A(n397_adj_3608), .B(n251_adj_3485), 
         .C(index_i[4]), .Z(n413_adj_3609)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_5_i413_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_4_i349_3_lut_4_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[4]), .D(n348), .Z(n349_adj_3610)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_4_i349_3_lut_4_lut.init = 16'hf606;
    LUT4 i17682_3_lut_3_lut (.A(index_i[0]), .B(index_i[2]), .C(index_i[3]), 
         .Z(n19996)) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i17682_3_lut_3_lut.init = 16'h6a6a;
    LUT4 i13079_2_lut_rep_562 (.A(index_i[2]), .B(index_i[0]), .Z(n29222)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i13079_2_lut_rep_562.init = 16'heeee;
    LUT4 i1_2_lut_rep_438_3_lut (.A(index_i[2]), .B(index_i[0]), .C(index_i[1]), 
         .Z(n29098)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_2_lut_rep_438_3_lut.init = 16'hfefe;
    LUT4 mux_208_Mux_2_i173_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[2]), 
         .B(index_i[0]), .C(index_i[3]), .D(index_i[1]), .Z(n173_adj_3496)) /* synthesis lut_function=(!(A (C)+!A (B (C+!(D))+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_2_i173_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h0f1a;
    LUT4 i17695_3_lut (.A(n20007), .B(n20008), .C(index_i[4]), .Z(n20009)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17695_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_5_i954_3_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[1]), .Z(n954)) /* synthesis lut_function=(!(A (C)+!A (B+((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_5_i954_3_lut_4_lut_4_lut.init = 16'h0a1a;
    LUT4 i14435_2_lut_rep_424_3_lut_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[1]), .Z(n29084)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i14435_2_lut_rep_424_3_lut_4_lut.init = 16'hf0e0;
    LUT4 mux_208_Mux_5_i125_3_lut (.A(n109_adj_3611), .B(n124_adj_3580), 
         .C(index_i[4]), .Z(n125_adj_3612)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_5_i125_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_9_i285_3_lut_3_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[1]), .Z(n285_adj_3569)) /* synthesis lut_function=(A (C)+!A !(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_9_i285_3_lut_3_lut_4_lut_4_lut.init = 16'ha0a1;
    LUT4 mux_208_Mux_5_i94_3_lut (.A(n653_adj_3526), .B(n635_adj_3591), 
         .C(index_i[4]), .Z(n94_adj_3613)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_5_i94_3_lut.init = 16'hcaca;
    L6MUX21 i26974 (.D0(n28919), .D1(n28916), .SD(index_i[5]), .Z(n28920));
    PFUMX i26972 (.BLUT(n28918), .ALUT(n28917), .C0(index_i[4]), .Z(n28919));
    LUT4 index_i_1__bdd_4_lut_27143 (.A(index_i[1]), .B(index_i[3]), .C(index_i[0]), 
         .D(index_i[2]), .Z(n29485)) /* synthesis lut_function=(!(A (B (D)+!B (C))+!A (B (C+!(D))+!B !(C+!(D))))) */ ;
    defparam index_i_1__bdd_4_lut_27143.init = 16'h169b;
    LUT4 mux_208_Mux_3_i700_3_lut_4_lut (.A(index_i[4]), .B(index_i[3]), 
         .C(n684_adj_3484), .D(n32053), .Z(n700_adj_3614)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_3_i700_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i28946 (.BLUT(n32063), .ALUT(n32064), .C0(index_i[1]), .Z(n32065));
    L6MUX21 i25190 (.D0(n26853), .D1(n26851), .SD(index_i[4]), .Z(n26854));
    PFUMX i26969 (.BLUT(n29044), .ALUT(n28915), .C0(index_i[4]), .Z(n28916));
    LUT4 i21058_3_lut_4_lut_4_lut (.A(index_i[2]), .B(n141), .C(index_i[3]), 
         .D(n29337), .Z(n23540)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21058_3_lut_4_lut_4_lut.init = 16'hc5c0;
    LUT4 mux_208_Mux_8_i732_3_lut (.A(index_i[3]), .B(n16890), .C(index_i[5]), 
         .Z(n732_adj_3615)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_8_i732_3_lut.init = 16'h3a3a;
    PFUMX i22063 (.BLUT(n221_adj_3616), .ALUT(n252), .C0(index_i[5]), 
          .Z(n24564));
    LUT4 n300_bdd_3_lut_26971_4_lut_4_lut (.A(index_i[2]), .B(n676), .C(index_i[3]), 
         .D(n29337), .Z(n28917)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B ((D)+!C)+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n300_bdd_3_lut_26971_4_lut_4_lut.init = 16'h5c0c;
    LUT4 mux_208_Mux_4_i158_3_lut (.A(n142_adj_3617), .B(n157_adj_3604), 
         .C(index_i[4]), .Z(n158_adj_3618)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_4_i158_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_7_i506_3_lut_4_lut_4_lut (.A(index_i[2]), .B(n29340), 
         .C(index_i[3]), .D(n29337), .Z(n506_adj_3619)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B ((D)+!C)+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_7_i506_3_lut_4_lut_4_lut.init = 16'h5c0c;
    PFUMX i22422 (.BLUT(n333), .ALUT(n348_adj_3620), .C0(index_i[4]), 
          .Z(n24923));
    LUT4 n518_bdd_3_lut_25185 (.A(n32044), .B(n32041), .C(index_i[3]), 
         .Z(n26849)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n518_bdd_3_lut_25185.init = 16'hcaca;
    LUT4 mux_208_Mux_4_i491_3_lut_4_lut_4_lut (.A(index_i[2]), .B(n29340), 
         .C(index_i[3]), .D(n29252), .Z(n491_adj_3573)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_4_i491_3_lut_4_lut_4_lut.init = 16'hfc5c;
    LUT4 mux_208_Mux_5_i924_4_lut_3_lut (.A(index_i[2]), .B(n15481), .C(index_i[4]), 
         .Z(n924_adj_3621)) /* synthesis lut_function=(!(A (B+(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_5_i924_4_lut_3_lut.init = 16'h5656;
    PFUMX i25188 (.BLUT(n29085), .ALUT(n26852), .C0(index_i[5]), .Z(n26853));
    PFUMX i22423 (.BLUT(n364), .ALUT(n379), .C0(index_i[4]), .Z(n24924));
    PFUMX i22424 (.BLUT(n397_adj_3622), .ALUT(n412), .C0(index_i[4]), 
          .Z(n24925));
    PFUMX i22425 (.BLUT(n428), .ALUT(n443_adj_3479), .C0(index_i[4]), 
          .Z(n24926));
    LUT4 i23749_3_lut (.A(n23431), .B(n23432), .C(index_i[4]), .Z(n23433)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i23749_3_lut.init = 16'hcaca;
    LUT4 i13082_3_lut_3_lut (.A(index_i[2]), .B(index_i[0]), .C(index_i[1]), 
         .Z(n467)) /* synthesis lut_function=(A (C)+!A (B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i13082_3_lut_3_lut.init = 16'hf4f4;
    PFUMX i22426 (.BLUT(n460), .ALUT(n475_adj_3623), .C0(index_i[4]), 
          .Z(n24927));
    L6MUX21 mux_208_Mux_7_i253 (.D0(n13456), .D1(n23436), .SD(index_i[5]), 
            .Z(n253)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    PFUMX i22427 (.BLUT(n491_adj_3596), .ALUT(n12561), .C0(index_i[4]), 
          .Z(n24928));
    PFUMX mux_208_Mux_7_i190 (.BLUT(n23433), .ALUT(n173_adj_3550), .C0(index_i[5]), 
          .Z(n190)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    PFUMX i25186 (.BLUT(n26850), .ALUT(n26849), .C0(index_i[5]), .Z(n26851));
    LUT4 mux_208_Mux_0_i397_3_lut (.A(n29257), .B(n32043), .C(index_i[3]), 
         .Z(n397_adj_3622)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_0_i397_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_0_i812_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n812_adj_3624)) /* synthesis lut_function=(A (B (C+(D))+!B !(C))+!A (B (D)+!B !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_0_i812_3_lut_4_lut_4_lut_4_lut.init = 16'hcf92;
    LUT4 n699_bdd_4_lut_26313_4_lut (.A(n29156), .B(index_i[3]), .C(n29349), 
         .D(index_i[6]), .Z(n26607)) /* synthesis lut_function=(!(A (B+(C (D)+!C !(D)))+!A (B (D)+!B (C (D)+!C !(D))))) */ ;
    defparam n699_bdd_4_lut_26313_4_lut.init = 16'h0374;
    LUT4 i12997_2_lut_rep_563 (.A(index_i[0]), .B(index_i[1]), .Z(n29223)) /* synthesis lut_function=(A+!(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12997_2_lut_rep_563.init = 16'hbbbb;
    PFUMX i22093 (.BLUT(n158_adj_3618), .ALUT(n189), .C0(index_i[5]), 
          .Z(n24594));
    LUT4 mux_208_Mux_2_i955_then_4_lut (.A(index_i[4]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n29488)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B (C+!(D))+!B !(C (D)))) */ ;
    defparam mux_208_Mux_2_i955_then_4_lut.init = 16'he95d;
    PFUMX mux_208_Mux_8_i764 (.BLUT(n716_adj_3477), .ALUT(n732_adj_3615), 
          .C0(n24130), .Z(n764)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 mux_208_Mux_4_i723_3_lut_4_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n723)) /* synthesis lut_function=(A ((C)+!B)+!A !(B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_4_i723_3_lut_4_lut_4_lut_3_lut.init = 16'hb2b2;
    LUT4 i21123_3_lut (.A(n467), .B(n7), .C(index_i[3]), .Z(n23605)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21123_3_lut.init = 16'hcaca;
    PFUMX mux_208_Mux_8_i574 (.BLUT(n542), .ALUT(n13452), .C0(index_i[5]), 
          .Z(n574)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 n300_bdd_3_lut_26992 (.A(n32049), .B(n32044), .C(index_i[3]), 
         .Z(n28918)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n300_bdd_3_lut_26992.init = 16'hcaca;
    PFUMX i27129 (.BLUT(n29566), .ALUT(n29567), .C0(index_i[4]), .Z(n29568));
    LUT4 i21070_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n23552)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D))+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21070_3_lut_4_lut.init = 16'hccdb;
    LUT4 i5217_2_lut_rep_565 (.A(index_i[0]), .B(index_i[1]), .Z(n29225)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i5217_2_lut_rep_565.init = 16'h6666;
    PFUMX i22845 (.BLUT(n589), .ALUT(n604), .C0(index_i[4]), .Z(n25346));
    LUT4 n442_bdd_3_lut_26998 (.A(n29228), .B(n32048), .C(index_i[3]), 
         .Z(n28937)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n442_bdd_3_lut_26998.init = 16'hcaca;
    L6MUX21 i22411 (.D0(n24910), .D1(n24911), .SD(index_i[5]), .Z(n24912));
    LUT4 i11261_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n13560)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B ((D)+!C)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11261_3_lut_4_lut_4_lut.init = 16'h6c3c;
    LUT4 mux_208_Mux_2_i955_else_4_lut (.A(index_i[4]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n29487)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+(D)))+!A !(B (C+!(D))+!B !(C+!(D))))) */ ;
    defparam mux_208_Mux_2_i955_else_4_lut.init = 16'h49c6;
    PFUMX i22052 (.BLUT(n956), .ALUT(n22204), .C0(index_i[6]), .Z(n24553));
    LUT4 mux_208_Mux_5_i828_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[4]), .D(n29363), .Z(n828_adj_3625)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_5_i828_4_lut_4_lut.init = 16'hc66c;
    LUT4 mux_208_Mux_5_i356_3_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n396)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_5_i356_3_lut_4_lut_3_lut.init = 16'h6d6d;
    PFUMX i22061 (.BLUT(n94_adj_3613), .ALUT(n125_adj_3612), .C0(index_i[5]), 
          .Z(n24562));
    PFUMX i22062 (.BLUT(n20009), .ALUT(n16238), .C0(index_i[5]), .Z(n24563));
    LUT4 n300_bdd_3_lut (.A(n32049), .B(n7), .C(index_i[3]), .Z(n28939)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n300_bdd_3_lut.init = 16'hacac;
    LUT4 mux_208_Mux_3_i507_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[4]), .D(n491_adj_3626), .Z(n507_adj_3627)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_3_i507_3_lut_4_lut.init = 16'h6f60;
    LUT4 i11263_3_lut_4_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[4]), .Z(n13562)) /* synthesis lut_function=(!(A (B)+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11263_3_lut_4_lut_4_lut_3_lut.init = 16'h6262;
    LUT4 i22261_3_lut_4_lut_4_lut (.A(n29156), .B(index_i[3]), .C(n29098), 
         .D(index_i[4]), .Z(n24762)) /* synthesis lut_function=(A (B (C (D))+!B !((D)+!C))+!A (B (C+!(D))+!B !((D)+!C))) */ ;
    defparam i22261_3_lut_4_lut_4_lut.init = 16'hc074;
    LUT4 mux_208_Mux_7_i156_3_lut_3_lut_rep_554_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29214)) /* synthesis lut_function=(!(A (B)+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_7_i156_3_lut_3_lut_rep_554_3_lut.init = 16'h6363;
    LUT4 mux_208_Mux_1_i882_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n882)) /* synthesis lut_function=(A ((C)+!B)+!A !((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_1_i882_3_lut_3_lut.init = 16'ha6a6;
    L6MUX21 i22064 (.D0(n23466), .D1(n23469), .SD(index_i[5]), .Z(n24565));
    LUT4 mux_208_Mux_7_i108_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n108)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_7_i108_3_lut_3_lut.init = 16'hc6c6;
    LUT4 i11181_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(n29325), .D(index_i[4]), .Z(n221_adj_3616)) /* synthesis lut_function=(!(A (B)+!A (B (C+(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11181_3_lut_4_lut_4_lut_4_lut.init = 16'h3336;
    L6MUX21 i22065 (.D0(n23472), .D1(n23475), .SD(index_i[5]), .Z(n24566));
    LUT4 mux_208_Mux_5_i459_3_lut_4_lut_3_lut_rep_566 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29226)) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_5_i459_3_lut_4_lut_3_lut_rep_566.init = 16'h6b6b;
    PFUMX i22066 (.BLUT(n413_adj_3609), .ALUT(n444), .C0(index_i[5]), 
          .Z(n24567));
    LUT4 mux_208_Mux_5_i773_rep_568 (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .Z(n29228)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_5_i773_rep_568.init = 16'h6464;
    LUT4 mux_208_Mux_5_i652_3_lut_3_lut_rep_569 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29229)) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_5_i652_3_lut_3_lut_rep_569.init = 16'h6a6a;
    LUT4 mux_208_Mux_3_i963_3_lut_4_lut_4_lut_3_lut_rep_571 (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[2]), .Z(n29231)) /* synthesis lut_function=(!(A (B)+!A ((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_3_i963_3_lut_4_lut_4_lut_3_lut_rep_571.init = 16'h2626;
    PFUMX i22067 (.BLUT(n476_adj_3606), .ALUT(n507), .C0(index_i[5]), 
          .Z(n24568));
    LUT4 i21051_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n23533)) /* synthesis lut_function=(!(A (B)+!A (B (C+(D))+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21051_3_lut_3_lut_4_lut.init = 16'h3326;
    PFUMX i22068 (.BLUT(n19997), .ALUT(n573_adj_3628), .C0(index_i[5]), 
          .Z(n24569));
    LUT4 n23537_bdd_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(n29363), 
         .D(index_i[4]), .Z(n26781)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+(D)))+!A (B (D)+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n23537_bdd_3_lut_3_lut_4_lut.init = 16'h336c;
    PFUMX i22069 (.BLUT(n605_adj_3629), .ALUT(n636_adj_3605), .C0(index_i[5]), 
          .Z(n24570));
    LUT4 mux_208_Mux_2_i491_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n491_adj_3630)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A !(B (C)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_2_i491_3_lut_4_lut_4_lut.init = 16'h6a5a;
    PFUMX i22070 (.BLUT(n23478), .ALUT(n700_adj_3534), .C0(index_i[5]), 
          .Z(n24571));
    LUT4 i21018_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n23500)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21018_3_lut_4_lut.init = 16'h64cc;
    LUT4 n22_bdd_3_lut_25172_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n26552)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C))+!A !(B (C+!(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n22_bdd_3_lut_25172_4_lut_4_lut.init = 16'h5ad6;
    LUT4 mux_208_Mux_5_i460_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n460_adj_3533)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A !(B (C)+!B !(C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_5_i460_3_lut_4_lut_4_lut.init = 16'h6b5a;
    LUT4 n396_bdd_3_lut_25426 (.A(n29339), .B(n29236), .C(index_i[3]), 
         .Z(n26869)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n396_bdd_3_lut_25426.init = 16'hcaca;
    LUT4 mux_208_Mux_5_i277_3_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n404)) /* synthesis lut_function=(A (B+!(C))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_5_i277_3_lut_4_lut_3_lut.init = 16'h9b9b;
    L6MUX21 i22071 (.D0(n732_adj_3545), .D1(n23481), .SD(index_i[5]), 
            .Z(n24572));
    PFUMX i22428 (.BLUT(n24913), .ALUT(n24914), .C0(index_i[5]), .Z(n24929));
    LUT4 mux_208_Mux_7_i333_3_lut (.A(n29339), .B(n29214), .C(index_i[3]), 
         .Z(n333_adj_3631)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_7_i333_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_7_i348_3_lut (.A(n29340), .B(n29257), .C(index_i[3]), 
         .Z(n348_adj_3632)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_7_i348_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_7_i364_3_lut (.A(n29339), .B(n29340), .C(index_i[3]), 
         .Z(n364_adj_3633)) /* synthesis lut_function=(A (B (C))+!A (B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_7_i364_3_lut.init = 16'hc5c5;
    LUT4 mux_208_Mux_7_i379_3_lut (.A(n29257), .B(n29339), .C(index_i[3]), 
         .Z(n379_adj_3598)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_7_i379_3_lut.init = 16'h3a3a;
    LUT4 mux_208_Mux_7_i397_3_lut (.A(n29340), .B(n29339), .C(index_i[3]), 
         .Z(n397_adj_3634)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_7_i397_3_lut.init = 16'hcaca;
    PFUMX i22429 (.BLUT(n24915), .ALUT(n24916), .C0(index_i[5]), .Z(n24930));
    PFUMX i22072 (.BLUT(n797_adj_3635), .ALUT(n828_adj_3625), .C0(index_i[5]), 
          .Z(n24573));
    LUT4 mux_208_Mux_0_i188_3_lut (.A(n29341), .B(n931), .C(index_i[3]), 
         .Z(n188)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_0_i188_3_lut.init = 16'hcaca;
    PFUMX i22073 (.BLUT(n860_adj_3601), .ALUT(n891_adj_3599), .C0(index_i[5]), 
          .Z(n24574));
    PFUMX i26822 (.BLUT(n28759), .ALUT(n28758), .C0(index_i[4]), .Z(n476));
    L6MUX21 i22430 (.D0(n24917), .D1(n24918), .SD(index_i[5]), .Z(n24931));
    LUT4 mux_208_Mux_1_i987_3_lut_4_lut (.A(n32027), .B(index_i[3]), .C(index_i[4]), 
         .D(n986_adj_3585), .Z(n987)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_1_i987_3_lut_4_lut.init = 16'hf202;
    LUT4 n155_bdd_3_lut_26757_4_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .Z(n26584)) /* synthesis lut_function=(A (B)+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n155_bdd_3_lut_26757_4_lut_3_lut.init = 16'hd9d9;
    LUT4 i23709_3_lut (.A(n27507), .B(n124_adj_3490), .C(index_i[4]), 
         .Z(n24916)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23709_3_lut.init = 16'hcaca;
    L6MUX21 i22433 (.D0(n24923), .D1(n24924), .SD(index_i[5]), .Z(n24934));
    L6MUX21 i22434 (.D0(n24925), .D1(n24926), .SD(index_i[5]), .Z(n24935));
    L6MUX21 i22435 (.D0(n24927), .D1(n24928), .SD(index_i[5]), .Z(n24936));
    LUT4 i24599_2_lut (.A(index_i[3]), .B(index_i[2]), .Z(n24132)) /* synthesis lut_function=(A+!(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i24599_2_lut.init = 16'hbbbb;
    PFUMX i26786 (.BLUT(n28719), .ALUT(n29221), .C0(index_i[4]), .Z(n28720));
    LUT4 mux_208_Mux_11_i638_4_lut_4_lut (.A(n29051), .B(index_i[5]), .C(index_i[6]), 
         .D(n29083), .Z(n638_adj_3562)) /* synthesis lut_function=(A (B (C (D))+!B !(C))+!A (B ((D)+!C)+!B !(C))) */ ;
    defparam mux_208_Mux_11_i638_4_lut_4_lut.init = 16'hc707;
    PFUMX i22846 (.BLUT(n620_adj_3593), .ALUT(n635_adj_3603), .C0(index_i[4]), 
          .Z(n25347));
    LUT4 i21099_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n23581)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !(B (C+!(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21099_3_lut_4_lut_4_lut.init = 16'ha5a9;
    LUT4 mux_208_Mux_6_i573_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[4]), .D(n572_adj_3636), .Z(n573_adj_3637)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_6_i573_3_lut_4_lut.init = 16'hf909;
    LUT4 mux_208_Mux_5_i109_3_lut_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .Z(n109_adj_3611)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_5_i109_3_lut_3_lut_3_lut.init = 16'h3939;
    CCU2D unary_minus_10_add_3_17 (.A0(\quarter_wave_sample_register_i[15] ), 
          .B0(GND_net), .C0(GND_net), .D0(GND_net), .A1(GND_net), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n19745), .S0(o_val_pipeline_i_0__15__N_1799[15]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam unary_minus_10_add_3_17.INIT0 = 16'hf555;
    defparam unary_minus_10_add_3_17.INIT1 = 16'h0000;
    defparam unary_minus_10_add_3_17.INJECT1_0 = "NO";
    defparam unary_minus_10_add_3_17.INJECT1_1 = "NO";
    PFUMX i22092 (.BLUT(n94_adj_3587), .ALUT(n23484), .C0(index_i[5]), 
          .Z(n24593));
    CCU2D unary_minus_10_add_3_15 (.A0(quarter_wave_sample_register_i[13]), 
          .B0(GND_net), .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[14]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19744), .COUT(n19745), 
          .S0(o_val_pipeline_i_0__15__N_1799[13]), .S1(o_val_pipeline_i_0__15__N_1799[14]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam unary_minus_10_add_3_15.INIT0 = 16'hf555;
    defparam unary_minus_10_add_3_15.INIT1 = 16'hf555;
    defparam unary_minus_10_add_3_15.INJECT1_0 = "NO";
    defparam unary_minus_10_add_3_15.INJECT1_1 = "NO";
    LUT4 i21060_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n23542)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C))+!A !(B ((D)+!C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21060_3_lut_4_lut_4_lut.init = 16'h925a;
    CCU2D unary_minus_10_add_3_13 (.A0(quarter_wave_sample_register_i[11]), 
          .B0(GND_net), .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[12]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19743), .COUT(n19744), 
          .S0(o_val_pipeline_i_0__15__N_1799[11]), .S1(o_val_pipeline_i_0__15__N_1799[12]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam unary_minus_10_add_3_13.INIT0 = 16'hf555;
    defparam unary_minus_10_add_3_13.INIT1 = 16'hf555;
    defparam unary_minus_10_add_3_13.INJECT1_0 = "NO";
    defparam unary_minus_10_add_3_13.INJECT1_1 = "NO";
    PFUMX i22540 (.BLUT(n25037), .ALUT(n25038), .C0(index_i[4]), .Z(n25041));
    PFUMX i22094 (.BLUT(n221_adj_3638), .ALUT(n252_adj_3639), .C0(index_i[5]), 
          .Z(n24595));
    PFUMX i22095 (.BLUT(n286_adj_3586), .ALUT(n23487), .C0(index_i[5]), 
          .Z(n24596));
    PFUMX i22541 (.BLUT(n25039), .ALUT(n25040), .C0(index_i[4]), .Z(n25042));
    CCU2D unary_minus_10_add_3_11 (.A0(quarter_wave_sample_register_i[9]), 
          .B0(GND_net), .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[10]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19742), .COUT(n19743), 
          .S0(o_val_pipeline_i_0__15__N_1799[9]), .S1(o_val_pipeline_i_0__15__N_1799[10]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam unary_minus_10_add_3_11.INIT0 = 16'hf555;
    defparam unary_minus_10_add_3_11.INIT1 = 16'hf555;
    defparam unary_minus_10_add_3_11.INJECT1_0 = "NO";
    defparam unary_minus_10_add_3_11.INJECT1_1 = "NO";
    CCU2D unary_minus_10_add_3_9 (.A0(quarter_wave_sample_register_i[7]), 
          .B0(GND_net), .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[8]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19741), .COUT(n19742), 
          .S0(o_val_pipeline_i_0__15__N_1799[7]), .S1(o_val_pipeline_i_0__15__N_1799[8]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam unary_minus_10_add_3_9.INIT0 = 16'hf555;
    defparam unary_minus_10_add_3_9.INIT1 = 16'hf555;
    defparam unary_minus_10_add_3_9.INJECT1_0 = "NO";
    defparam unary_minus_10_add_3_9.INJECT1_1 = "NO";
    PFUMX i22096 (.BLUT(n349_adj_3610), .ALUT(n23490), .C0(index_i[5]), 
          .Z(n24597));
    CCU2D unary_minus_10_add_3_7 (.A0(quarter_wave_sample_register_i[5]), 
          .B0(GND_net), .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[6]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19740), .COUT(n19741), 
          .S0(o_val_pipeline_i_0__15__N_1799[5]), .S1(o_val_pipeline_i_0__15__N_1799[6]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam unary_minus_10_add_3_7.INIT0 = 16'hf555;
    defparam unary_minus_10_add_3_7.INIT1 = 16'hf555;
    defparam unary_minus_10_add_3_7.INJECT1_0 = "NO";
    defparam unary_minus_10_add_3_7.INJECT1_1 = "NO";
    PFUMX i22547 (.BLUT(n25044), .ALUT(n25045), .C0(index_i[4]), .Z(n25048));
    CCU2D unary_minus_10_add_3_5 (.A0(quarter_wave_sample_register_i[3]), 
          .B0(GND_net), .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[4]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19739), .COUT(n19740), 
          .S0(o_val_pipeline_i_0__15__N_1799[3]), .S1(o_val_pipeline_i_0__15__N_1799[4]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam unary_minus_10_add_3_5.INIT0 = 16'hf555;
    defparam unary_minus_10_add_3_5.INIT1 = 16'hf555;
    defparam unary_minus_10_add_3_5.INJECT1_0 = "NO";
    defparam unary_minus_10_add_3_5.INJECT1_1 = "NO";
    LUT4 mux_208_Mux_7_i891_3_lut_4_lut_4_lut (.A(n29182), .B(index_i[3]), 
         .C(n29103), .D(index_i[4]), .Z(n891_adj_3640)) /* synthesis lut_function=(A (B (C+!(D))+!B !((D)+!C))+!A (B (C+!(D))+!B (C+(D)))) */ ;
    defparam mux_208_Mux_7_i891_3_lut_4_lut_4_lut.init = 16'hd1fc;
    CCU2D unary_minus_10_add_3_3 (.A0(quarter_wave_sample_register_i[1]), 
          .B0(GND_net), .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[2]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19738), .COUT(n19739), 
          .S0(o_val_pipeline_i_0__15__N_1799[1]), .S1(o_val_pipeline_i_0__15__N_1799[2]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam unary_minus_10_add_3_3.INIT0 = 16'hf555;
    defparam unary_minus_10_add_3_3.INIT1 = 16'hf555;
    defparam unary_minus_10_add_3_3.INJECT1_0 = "NO";
    defparam unary_minus_10_add_3_3.INJECT1_1 = "NO";
    PFUMX i22548 (.BLUT(n25046), .ALUT(n25047), .C0(index_i[4]), .Z(n25049));
    CCU2D unary_minus_10_add_3_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(quarter_wave_sample_register_i[0]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .COUT(n19738), .S1(o_val_pipeline_i_0__15__N_1799[0]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam unary_minus_10_add_3_1.INIT0 = 16'hF000;
    defparam unary_minus_10_add_3_1.INIT1 = 16'h0aaa;
    defparam unary_minus_10_add_3_1.INJECT1_0 = "NO";
    defparam unary_minus_10_add_3_1.INJECT1_1 = "NO";
    PFUMX i22101 (.BLUT(n669_adj_3583), .ALUT(n700_adj_3582), .C0(index_i[5]), 
          .Z(n24602));
    PFUMX i22554 (.BLUT(n25051), .ALUT(n25052), .C0(index_i[4]), .Z(n25055));
    PFUMX i22555 (.BLUT(n25053), .ALUT(n25054), .C0(index_i[4]), .Z(n25056));
    PFUMX i22102 (.BLUT(n23502), .ALUT(n763_adj_3641), .C0(index_i[5]), 
          .Z(n24603));
    LUT4 i24600_2_lut (.A(index_i[5]), .B(index_i[4]), .Z(n24130)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i24600_2_lut.init = 16'heeee;
    LUT4 i1_3_lut (.A(index_i[0]), .B(index_i[4]), .C(index_i[2]), .Z(n22568)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_3_lut.init = 16'hfefe;
    PFUMX i22847 (.BLUT(n653_adj_3579), .ALUT(n668_adj_3642), .C0(index_i[4]), 
          .Z(n25348));
    PFUMX i25129 (.BLUT(n26784), .ALUT(n26780), .C0(index_i[6]), .Z(n26785));
    LUT4 mux_208_Mux_6_i505_3_lut_rep_573 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29233)) /* synthesis lut_function=(A (B)+!A (B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_6_i505_3_lut_rep_573.init = 16'hc9c9;
    LUT4 mux_208_Mux_7_i892_3_lut (.A(n62_adj_3643), .B(n891_adj_3640), 
         .C(index_i[5]), .Z(n892_adj_3644)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_7_i892_3_lut.init = 16'hcaca;
    LUT4 i21379_3_lut (.A(n747_adj_3645), .B(n762_adj_3475), .C(index_i[4]), 
         .Z(n23861)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21379_3_lut.init = 16'hcaca;
    LUT4 i21378_3_lut (.A(n716_adj_3646), .B(n16698), .C(index_i[4]), 
         .Z(n23860)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21378_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_6_i653_3_lut (.A(n29344), .B(n676), .C(index_i[3]), 
         .Z(n653_adj_3526)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_6_i653_3_lut.init = 16'hcaca;
    LUT4 i24100_3_lut (.A(n32061), .B(n29492), .C(index_i[5]), .Z(n23826)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24100_3_lut.init = 16'hcaca;
    LUT4 i21376_3_lut (.A(n93_adj_3647), .B(n699), .C(index_i[4]), .Z(n23858)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21376_3_lut.init = 16'hcaca;
    LUT4 i21375_3_lut (.A(n653), .B(n29061), .C(index_i[4]), .Z(n23857)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21375_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_6_i250_3_lut_4_lut_3_lut_rep_574 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29234)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_6_i250_3_lut_4_lut_3_lut_rep_574.init = 16'h9696;
    LUT4 mux_208_Mux_4_i684_3_lut (.A(n676), .B(n108), .C(index_i[3]), 
         .Z(n684_adj_3581)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_4_i684_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_5_i397_3_lut (.A(n29242), .B(n332), .C(index_i[3]), 
         .Z(n397_adj_3608)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_5_i397_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_5_i506_3_lut (.A(n29413), .B(n32050), .C(index_i[3]), 
         .Z(n506)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_5_i506_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_5_i761_3_lut_4_lut_3_lut_rep_576 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29236)) /* synthesis lut_function=(A (B)+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_5_i761_3_lut_4_lut_3_lut_rep_576.init = 16'hd9d9;
    PFUMX i22103 (.BLUT(n23505), .ALUT(n828_adj_3648), .C0(index_i[5]), 
          .Z(n24604));
    LUT4 mux_208_Mux_7_i116_3_lut_3_lut_3_lut_rep_577 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29237)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_7_i116_3_lut_3_lut_3_lut_rep_577.init = 16'h3939;
    LUT4 mux_208_Mux_6_i363_3_lut_4_lut_4_lut_3_lut_rep_579 (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[2]), .Z(n29239)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_6_i363_3_lut_4_lut_4_lut_3_lut_rep_579.init = 16'h9292;
    PFUMX i27125 (.BLUT(n29560), .ALUT(n29561), .C0(index_i[2]), .Z(n29562));
    LUT4 mux_208_Mux_5_i15_3_lut (.A(n29240), .B(n32032), .C(index_i[3]), 
         .Z(n15_adj_3538)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_5_i15_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_5_i859_3_lut (.A(n141), .B(n29240), .C(index_i[3]), 
         .Z(n859_adj_3600)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_5_i859_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_5_i875_3_lut (.A(n29214), .B(n29340), .C(index_i[3]), 
         .Z(n875_adj_3597)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_5_i875_3_lut.init = 16'hcaca;
    LUT4 i21342_3_lut_then_4_lut (.A(index_i[4]), .B(index_i[0]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n32060)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A !(B (C)+!B !((D)+!C))) */ ;
    defparam i21342_3_lut_then_4_lut.init = 16'h95a5;
    PFUMX i26589 (.BLUT(n28521), .ALUT(n28520), .C0(index_i[5]), .Z(n28522));
    LUT4 i21369_3_lut (.A(n526_adj_3649), .B(n541_adj_3548), .C(index_i[4]), 
         .Z(n23851)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21369_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_7_i77_3_lut_3_lut_rep_580 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29240)) /* synthesis lut_function=(A (B)+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_7_i77_3_lut_3_lut_rep_580.init = 16'h9c9c;
    LUT4 i21343_3_lut_then_4_lut (.A(index_i[4]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n29491)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)+!C !(D)))+!A !(B (C+!(D))+!B (C (D)+!C !(D))))) */ ;
    defparam i21343_3_lut_then_4_lut.init = 16'h5a65;
    LUT4 i21343_3_lut_else_4_lut (.A(index_i[4]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n29490)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A !(B (C+!(D))+!B ((D)+!C)))) */ ;
    defparam i21343_3_lut_else_4_lut.init = 16'h59e5;
    PFUMX i22848 (.BLUT(n684_adj_3650), .ALUT(n699_adj_3651), .C0(index_i[4]), 
          .Z(n25349));
    PFUMX i22104 (.BLUT(n860_adj_3577), .ALUT(n23508), .C0(index_i[5]), 
          .Z(n24605));
    LUT4 i21366_3_lut (.A(n397_adj_3634), .B(n475_adj_3481), .C(index_i[4]), 
         .Z(n23848)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21366_3_lut.init = 16'hcaca;
    LUT4 i23996_3_lut (.A(n23605), .B(n23606), .C(index_i[4]), .Z(n23607)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23996_3_lut.init = 16'hcaca;
    LUT4 i21364_3_lut (.A(n348_adj_3632), .B(n443_adj_3575), .C(index_i[4]), 
         .Z(n23846)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21364_3_lut.init = 16'hcaca;
    L6MUX21 i26580 (.D0(n28510), .D1(n28508), .SD(index_i[6]), .Z(n23301));
    PFUMX i26578 (.BLUT(n28509), .ALUT(n62_adj_3643), .C0(index_i[5]), 
          .Z(n28510));
    LUT4 i21363_3_lut (.A(n397_adj_3634), .B(n412_adj_3549), .C(index_i[4]), 
         .Z(n23845)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21363_3_lut.init = 16'hcaca;
    LUT4 i21361_3_lut (.A(n364_adj_3633), .B(n379_adj_3598), .C(index_i[4]), 
         .Z(n23843)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21361_3_lut.init = 16'hcaca;
    PFUMX i26576 (.BLUT(n28507), .ALUT(n28506), .C0(index_i[5]), .Z(n28508));
    LUT4 i21360_3_lut (.A(n333_adj_3631), .B(n348_adj_3632), .C(index_i[4]), 
         .Z(n23842)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21360_3_lut.init = 16'hcaca;
    LUT4 i20985_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n23467)) /* synthesis lut_function=(A (B (C (D))+!B !(C (D)))+!A !(B (D)+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20985_3_lut_4_lut_4_lut.init = 16'h9366;
    LUT4 mux_208_Mux_2_i604_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n604_adj_3494)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)+!C !(D)))+!A (B (D)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_2_i604_3_lut_4_lut_4_lut_4_lut.init = 16'h39cf;
    LUT4 i21352_3_lut (.A(n491_adj_3652), .B(n506_adj_3584), .C(index_i[4]), 
         .Z(n23834)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21352_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_5_i731_3_lut (.A(n32046), .B(n32043), .C(index_i[3]), 
         .Z(n731_adj_3544)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_5_i731_3_lut.init = 16'hcaca;
    LUT4 i21339_3_lut (.A(n78), .B(n93_adj_3647), .C(index_i[4]), .Z(n23821)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21339_3_lut.init = 16'hcaca;
    LUT4 i21336_3_lut (.A(n15_adj_3589), .B(n30_adj_3543), .C(index_i[4]), 
         .Z(n23818)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21336_3_lut.init = 16'hcaca;
    LUT4 i21072_3_lut (.A(n404), .B(n32052), .C(index_i[3]), .Z(n23554)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21072_3_lut.init = 16'hcaca;
    LUT4 i21061_3_lut (.A(n32051), .B(n29345), .C(index_i[3]), .Z(n23543)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21061_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_6_i572_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n572_adj_3636)) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_6_i572_3_lut_4_lut.init = 16'hccd9;
    LUT4 i21088_3_lut_4_lut (.A(index_i[0]), .B(n29218), .C(index_i[3]), 
         .D(n32042), .Z(n23570)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21088_3_lut_4_lut.init = 16'hfb0b;
    LUT4 n676_bdd_3_lut_25788_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n26866)) /* synthesis lut_function=(A (B (C+(D)))+!A (B ((D)+!C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n676_bdd_3_lut_25788_4_lut.init = 16'hcc94;
    LUT4 mux_208_Mux_2_i653_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n653_adj_3492)) /* synthesis lut_function=(A (B (C+!(D))+!B !(D))+!A !(B (C+!(D))+!B !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_2_i653_3_lut_4_lut.init = 16'h94aa;
    LUT4 i23508_3_lut (.A(n23554), .B(n23555), .C(index_i[4]), .Z(n23556)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23508_3_lut.init = 16'hcaca;
    LUT4 i23522_3_lut (.A(n23542), .B(n23543), .C(index_i[4]), .Z(n23544)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23522_3_lut.init = 16'hcaca;
    LUT4 n396_bdd_3_lut_25202_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n26868)) /* synthesis lut_function=(A (B (C+(D))+!B ((D)+!C))+!A !(B (C+(D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n396_bdd_3_lut_25202_4_lut.init = 16'haa96;
    LUT4 i21124_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n23606)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C+(D)))+!A (B (C)+!B !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21124_3_lut_4_lut_4_lut.init = 16'hc95a;
    PFUMX i22214 (.BLUT(n24713), .ALUT(n24714), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_1768[1]));
    PFUMX i22090 (.BLUT(n24589), .ALUT(n24590), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_1768[5]));
    PFUMX i22152 (.BLUT(n24651), .ALUT(n24652), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_1768[3]));
    PFUMX i22183 (.BLUT(n24682), .ALUT(n24683), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_1768[2]));
    PFUMX i27121 (.BLUT(n29554), .ALUT(n29555), .C0(index_i[8]), .Z(n29556));
    LUT4 i21063_3_lut_3_lut_4_lut (.A(n29222), .B(index_i[1]), .C(index_i[3]), 
         .D(n29103), .Z(n23545)) /* synthesis lut_function=(!(A (C (D))+!A (B (C (D))+!B ((D)+!C)))) */ ;
    defparam i21063_3_lut_3_lut_4_lut.init = 16'h0efe;
    L6MUX21 i14977388_i1 (.D0(n24943), .D1(n25374), .SD(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_1768[0]));
    PFUMX i20585 (.BLUT(n23065), .ALUT(n23066), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_1768[11]));
    L6MUX21 i28733 (.D0(n31734), .D1(n31731), .SD(index_i[7]), .Z(n31735));
    PFUMX mux_208_Mux_13_i1023 (.BLUT(n511), .ALUT(n22166), .C0(index_i[9]), 
          .Z(quarter_wave_sample_register_i_15__N_1768[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    PFUMX i28731 (.BLUT(n31733), .ALUT(n31732), .C0(index_i[5]), .Z(n31734));
    LUT4 i21354_4_lut_4_lut_3_lut_4_lut (.A(n29222), .B(index_i[1]), .C(index_i[4]), 
         .D(index_i[3]), .Z(n23836)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B !((D)+!C)))) */ ;
    defparam i21354_4_lut_4_lut_3_lut_4_lut.init = 16'h11ef;
    PFUMX i28729 (.BLUT(n25186), .ALUT(n31730), .C0(index_i[6]), .Z(n31731));
    L6MUX21 i22630 (.D0(n25127), .D1(n25128), .SD(index_i[8]), .Z(n25131));
    PFUMX i22661 (.BLUT(n25160), .ALUT(n25161), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_1768[8]));
    LUT4 i23858_3_lut (.A(n620_adj_3540), .B(n15399), .C(index_i[4]), 
         .Z(n23855)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23858_3_lut.init = 16'hcaca;
    LUT4 i23863_3_lut (.A(n491_adj_3653), .B(n506_adj_3619), .C(index_i[4]), 
         .Z(n23849)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23863_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_3_i747_3_lut (.A(n29228), .B(n404), .C(index_i[3]), 
         .Z(n747_adj_3536)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_3_i747_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_3_i94_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[4]), .D(n93), .Z(n94_adj_3654)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_3_i94_3_lut_4_lut.init = 16'hf606;
    PFUMX i22873 (.BLUT(n25372), .ALUT(n25373), .C0(index_i[8]), .Z(n25374));
    LUT4 i11156_4_lut_4_lut (.A(n29222), .B(index_i[1]), .C(index_i[3]), 
         .D(n22568), .Z(n13452)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A (B (C)+!B ((D)+!C)))) */ ;
    defparam i11156_4_lut_4_lut.init = 16'h0e3e;
    LUT4 mux_208_Mux_9_i124_3_lut_3_lut_4_lut (.A(n29222), .B(index_i[1]), 
         .C(index_i[3]), .D(n29182), .Z(n124_adj_3568)) /* synthesis lut_function=(!(A (C (D))+!A (B (C (D))+!B ((D)+!C)))) */ ;
    defparam mux_208_Mux_9_i124_3_lut_3_lut_4_lut.init = 16'h0efe;
    L6MUX21 i22211 (.D0(n24707), .D1(n24708), .SD(index_i[7]), .Z(n24712));
    LUT4 i23879_3_lut (.A(n109), .B(n124), .C(index_i[4]), .Z(n23822)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23879_3_lut.init = 16'hcaca;
    LUT4 i22208_3_lut (.A(n24701), .B(n24702), .C(index_i[7]), .Z(n24709)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22208_3_lut.init = 16'hcaca;
    LUT4 i22201_3_lut (.A(n24687), .B(n26854), .C(index_i[6]), .Z(n24702)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22201_3_lut.init = 16'hcaca;
    LUT4 i22210_3_lut (.A(n24705), .B(n24706), .C(index_i[7]), .Z(n24711)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22210_3_lut.init = 16'hcaca;
    LUT4 i12995_2_lut_rep_665 (.A(index_i[2]), .B(index_i[3]), .Z(n29325)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12995_2_lut_rep_665.init = 16'h8888;
    LUT4 i22204_3_lut (.A(n26871), .B(n24694), .C(index_i[6]), .Z(n24705)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22204_3_lut.init = 16'hcaca;
    LUT4 n589_bdd_3_lut_26395_3_lut_4_lut (.A(n29222), .B(index_i[1]), .C(index_i[4]), 
         .D(index_i[3]), .Z(n28301)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B ((D)+!C))) */ ;
    defparam n589_bdd_3_lut_26395_3_lut_4_lut.init = 16'hf10f;
    LUT4 i22268_3_lut_3_lut_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[4]), .D(index_i[1]), .Z(n24769)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i22268_3_lut_3_lut_3_lut_4_lut.init = 16'h878f;
    LUT4 i21800_1_lut_2_lut (.A(index_i[2]), .B(index_i[3]), .Z(n24301)) /* synthesis lut_function=(!(A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21800_1_lut_2_lut.init = 16'h7777;
    LUT4 i17693_3_lut_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), .C(index_i[1]), 
         .D(index_i[0]), .Z(n20007)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i17693_3_lut_3_lut_4_lut.init = 16'hf078;
    LUT4 i13041_2_lut_rep_481_3_lut (.A(index_i[2]), .B(index_i[3]), .C(index_i[1]), 
         .Z(n29141)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i13041_2_lut_rep_481_3_lut.init = 16'h8080;
    LUT4 i14459_2_lut_rep_416_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[4]), .D(n29337), .Z(n29076)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i14459_2_lut_rep_416_3_lut_4_lut.init = 16'hf8f0;
    LUT4 i9147_3_lut_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), .C(index_i[1]), 
         .D(index_i[0]), .Z(n157_adj_3604)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(D))+!A !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9147_3_lut_3_lut_4_lut.init = 16'h7780;
    PFUMX i22057 (.BLUT(n24554), .ALUT(n24555), .C0(index_i[8]), .Z(n24558));
    L6MUX21 i22058 (.D0(n24556), .D1(n24557), .SD(index_i[8]), .Z(n24559));
    PFUMX i22442 (.BLUT(n24941), .ALUT(n24942), .C0(index_i[8]), .Z(n24943));
    LUT4 i1_2_lut_rep_492_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), .C(index_i[0]), 
         .D(index_i[1]), .Z(n29152)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_2_lut_rep_492_3_lut_4_lut.init = 16'h8000;
    LUT4 mux_208_Mux_8_i475_3_lut_3_lut_4_lut (.A(n29222), .B(index_i[1]), 
         .C(index_i[3]), .D(n29182), .Z(n475)) /* synthesis lut_function=(A (C+!(D))+!A (B (C+!(D))+!B !(C+(D)))) */ ;
    defparam mux_208_Mux_8_i475_3_lut_3_lut_4_lut.init = 16'he0ef;
    PFUMX i22626 (.BLUT(n25119), .ALUT(n25120), .C0(index_i[7]), .Z(n25127));
    PFUMX i22627 (.BLUT(n25121), .ALUT(n25122), .C0(index_i[7]), .Z(n25128));
    LUT4 i17694_3_lut_3_lut_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n20008)) /* synthesis lut_function=(!(A (B (C)+!B !(C (D)+!C !(D)))+!A !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i17694_3_lut_3_lut_3_lut_4_lut.init = 16'h780f;
    LUT4 i11169_3_lut_3_lut_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n541_adj_3509)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11169_3_lut_3_lut_3_lut_4_lut.init = 16'h870f;
    LUT4 i23529_3_lut (.A(n23539), .B(n23540), .C(index_i[4]), .Z(n23541)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23529_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_7_i924_3_lut_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[4]), .D(n29337), .Z(n924_adj_3483)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_7_i924_3_lut_3_lut_4_lut.init = 16'h878f;
    LUT4 n20197_bdd_4_lut_then_4_lut (.A(index_i[3]), .B(index_i[4]), .C(index_i[0]), 
         .D(index_i[2]), .Z(n29583)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B+(C (D)+!C !(D)))) */ ;
    defparam n20197_bdd_4_lut_then_4_lut.init = 16'hf44f;
    LUT4 n45_bdd_2_lut_3_lut_4_lut_4_lut (.A(index_i[3]), .B(index_i[1]), 
         .C(index_i[0]), .D(index_i[2]), .Z(n27451)) /* synthesis lut_function=(!(A+!(B+(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n45_bdd_2_lut_3_lut_4_lut_4_lut.init = 16'h5554;
    LUT4 i10306_4_lut_4_lut (.A(index_i[3]), .B(index_i[0]), .C(index_i[1]), 
         .D(index_i[2]), .Z(n12561)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (D)+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i10306_4_lut_4_lut.init = 16'h0bf4;
    LUT4 i22148_3_lut (.A(n24643), .B(n24644), .C(index_i[7]), .Z(n24649)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22148_3_lut.init = 16'hcaca;
    LUT4 i22143_3_lut (.A(n24633), .B(n24634), .C(index_i[6]), .Z(n24644)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22143_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_0_i572_3_lut_4_lut (.A(n29222), .B(index_i[1]), .C(index_i[3]), 
         .D(n32044), .Z(n572)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam mux_208_Mux_0_i572_3_lut_4_lut.init = 16'hefe0;
    LUT4 mux_208_Mux_3_i62_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[4]), .D(n812_adj_3520), .Z(n62_adj_3655)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_3_i62_3_lut_4_lut.init = 16'h6f60;
    L6MUX21 i26398 (.D0(n28303), .D1(n29027), .SD(index_i[6]), .Z(n638));
    PFUMX i26396 (.BLUT(n28302), .ALUT(n28301), .C0(index_i[5]), .Z(n28303));
    LUT4 i22177_3_lut (.A(n26785), .B(n24671), .C(index_i[7]), .Z(n24678)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22177_3_lut.init = 16'hcaca;
    L6MUX21 i22149 (.D0(n24645), .D1(n24646), .SD(index_i[7]), .Z(n24650));
    LUT4 i22266_3_lut_4_lut_3_lut (.A(index_i[3]), .B(index_i[4]), .C(n29182), 
         .Z(n24767)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i22266_3_lut_4_lut_3_lut.init = 16'h6464;
    LUT4 mux_208_Mux_3_i251_3_lut_4_lut (.A(n29222), .B(index_i[1]), .C(index_i[3]), 
         .D(n29156), .Z(n16734)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam mux_208_Mux_3_i251_3_lut_4_lut.init = 16'hfe0e;
    L6MUX21 i22178 (.D0(n24672), .D1(n24673), .SD(index_i[7]), .Z(n24679));
    LUT4 mux_208_Mux_2_i221_4_lut_4_lut (.A(index_i[3]), .B(index_i[4]), 
         .C(n29103), .D(n29085), .Z(n221_adj_3656)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (B+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_2_i221_4_lut_4_lut.init = 16'hf7c4;
    L6MUX21 i22179 (.D0(n24674), .D1(n24675), .SD(index_i[7]), .Z(n24680));
    PFUMX i22180 (.BLUT(n24676), .ALUT(n24677), .C0(index_i[7]), .Z(n24681));
    L6MUX21 i22205 (.D0(n24695), .D1(n24696), .SD(index_i[6]), .Z(n24706));
    L6MUX21 i22206 (.D0(n24697), .D1(n24698), .SD(index_i[6]), .Z(n24707));
    L6MUX21 i22209 (.D0(n24703), .D1(n24704), .SD(index_i[7]), .Z(n24710));
    LUT4 i13014_2_lut_3_lut_3_lut (.A(index_i[3]), .B(index_i[0]), .C(index_i[1]), 
         .Z(n15423)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i13014_2_lut_3_lut_3_lut.init = 16'h4040;
    LUT4 i13403_2_lut_4_lut_4_lut_4_lut (.A(index_i[3]), .B(index_i[2]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n668_adj_3642)) /* synthesis lut_function=(!(A+!(B (C)+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i13403_2_lut_4_lut_4_lut_4_lut.init = 16'h5041;
    LUT4 i21096_3_lut_3_lut_4_lut (.A(n29222), .B(index_i[1]), .C(n29103), 
         .D(index_i[3]), .Z(n23578)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;
    defparam i21096_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 i13447_4_lut_4_lut (.A(index_i[3]), .B(index_i[2]), .C(index_i[0]), 
         .D(index_i[1]), .Z(n875_adj_3657)) /* synthesis lut_function=((B (C)+!B (D))+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i13447_4_lut_4_lut.init = 16'hf7d5;
    LUT4 i21382_4_lut_3_lut (.A(index_i[3]), .B(index_i[4]), .C(n29103), 
         .Z(n23864)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21382_4_lut_3_lut.init = 16'h6565;
    LUT4 i11264_3_lut_4_lut_4_lut_4_lut (.A(index_i[3]), .B(index_i[2]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n13563)) /* synthesis lut_function=(!(A ((D)+!C)+!A !(B (C+!(D))+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11264_3_lut_4_lut_4_lut_4_lut.init = 16'h51e5;
    LUT4 i11158_3_lut_3_lut (.A(index_i[3]), .B(index_i[4]), .C(n13453), 
         .Z(n13454)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11158_3_lut_3_lut.init = 16'h7474;
    LUT4 i8558_2_lut (.A(index_i[4]), .B(index_i[5]), .Z(n10789)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i8558_2_lut.init = 16'h8888;
    LUT4 mux_208_Mux_3_i796_3_lut_3_lut (.A(index_i[4]), .B(n412_adj_3549), 
         .C(index_i[2]), .Z(n796_adj_3658)) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam mux_208_Mux_3_i796_3_lut_3_lut.init = 16'he4e4;
    LUT4 i22167_4_lut_4_lut (.A(index_i[4]), .B(index_i[5]), .C(n29489), 
         .D(n908_adj_3578), .Z(n24668)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam i22167_4_lut_4_lut.init = 16'hd1c0;
    LUT4 i11153_4_lut_4_lut (.A(index_i[4]), .B(n24305), .C(n32065), .D(n29256), 
         .Z(n13449)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam i11153_4_lut_4_lut.init = 16'hf4b0;
    LUT4 i14496_2_lut_rep_391_3_lut_4_lut (.A(n29222), .B(index_i[1]), .C(index_i[4]), 
         .D(index_i[3]), .Z(n29051)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i14496_2_lut_rep_391_3_lut_4_lut.init = 16'hfef0;
    LUT4 i1_2_lut_rep_587 (.A(index_i[5]), .B(index_i[6]), .Z(n29247)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_2_lut_rep_587.init = 16'heeee;
    LUT4 i1_3_lut_4_lut_adj_192 (.A(index_i[5]), .B(index_i[6]), .C(index_i[7]), 
         .D(n29362), .Z(n22122)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_3_lut_4_lut_adj_192.init = 16'hfffe;
    LUT4 i22081_3_lut (.A(n24571), .B(n24572), .C(index_i[6]), .Z(n24582)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22081_3_lut.init = 16'hcaca;
    L6MUX21 i22542 (.D0(n25041), .D1(n25042), .SD(index_i[5]), .Z(n25043));
    L6MUX21 i22549 (.D0(n25048), .D1(n25049), .SD(index_i[5]), .Z(n25050));
    L6MUX21 i20795 (.D0(n23275), .D1(n23276), .SD(index_i[7]), .Z(n23277));
    L6MUX21 i22556 (.D0(n25055), .D1(n25056), .SD(index_i[5]), .Z(n25057));
    LUT4 mux_208_Mux_6_i452_3_lut_3_lut_3_lut_rep_837 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n32038)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_6_i452_3_lut_3_lut_3_lut_rep_837.init = 16'h9393;
    PFUMX i27115 (.BLUT(n29545), .ALUT(n29546), .C0(index_i[3]), .Z(n62_adj_3643));
    LUT4 n26608_bdd_3_lut_4_lut (.A(n29055), .B(index_i[6]), .C(index_i[5]), 
         .D(n26608), .Z(n26609)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam n26608_bdd_3_lut_4_lut.init = 16'hefe0;
    LUT4 n20197_bdd_4_lut_else_4_lut (.A(index_i[3]), .B(index_i[4]), .C(index_i[0]), 
         .D(index_i[2]), .Z(n29582)) /* synthesis lut_function=(!(A (B (D)+!B ((D)+!C))+!A !(B+!((D)+!C)))) */ ;
    defparam n20197_bdd_4_lut_else_4_lut.init = 16'h44fc;
    L6MUX21 i22055 (.D0(n24550), .D1(n24551), .SD(index_i[7]), .Z(n24556));
    L6MUX21 i22056 (.D0(n24552), .D1(n24553), .SD(index_i[7]), .Z(n24557));
    L6MUX21 i22084 (.D0(n24577), .D1(n24578), .SD(index_i[7]), .Z(n24585));
    L6MUX21 i22085 (.D0(n24579), .D1(n24580), .SD(index_i[7]), .Z(n24586));
    L6MUX21 i22628 (.D0(n25123), .D1(n25124), .SD(index_i[7]), .Z(n25129));
    L6MUX21 i22657 (.D0(n25152), .D1(n25153), .SD(index_i[7]), .Z(n25158));
    PFUMX i22658 (.BLUT(n25154), .ALUT(n25155), .C0(index_i[7]), .Z(n25159));
    LUT4 i22046_3_lut (.A(n190), .B(n253), .C(index_i[6]), .Z(n24547)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22046_3_lut.init = 16'hcaca;
    LUT4 i22047_3_lut (.A(n25057), .B(n23844), .C(index_i[6]), .Z(n24548)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22047_3_lut.init = 16'hcaca;
    LUT4 i22437_3_lut (.A(n24931), .B(n30487), .C(index_i[6]), .Z(n24938)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22437_3_lut.init = 16'hcaca;
    LUT4 i22438_3_lut (.A(n27648), .B(n24934), .C(index_i[6]), .Z(n24939)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22438_3_lut.init = 16'hcaca;
    L6MUX21 i26318 (.D0(n28183), .D1(n28181), .SD(index_i[6]), .Z(n28184));
    LUT4 i22649_3_lut (.A(n27407), .B(n24912), .C(index_i[6]), .Z(n25150)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22649_3_lut.init = 16'hcaca;
    PFUMX i26316 (.BLUT(n924_adj_3621), .ALUT(n28182), .C0(index_i[5]), 
          .Z(n28183));
    LUT4 n22_bdd_3_lut_24928 (.A(n32053), .B(n32041), .C(index_i[3]), 
         .Z(n26551)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n22_bdd_3_lut_24928.init = 16'hcaca;
    L6MUX21 i22682 (.D0(n25181), .D1(n25182), .SD(index_i[7]), .Z(n25183));
    L6MUX21 i22144 (.D0(n24635), .D1(n24636), .SD(index_i[6]), .Z(n24645));
    L6MUX21 i22146 (.D0(n24639), .D1(n24640), .SD(index_i[7]), .Z(n24647));
    L6MUX21 i22147 (.D0(n24641), .D1(n24642), .SD(index_i[7]), .Z(n24648));
    L6MUX21 i22867 (.D0(n25360), .D1(n25361), .SD(index_i[6]), .Z(n25368));
    L6MUX21 i22868 (.D0(n25362), .D1(n25363), .SD(index_i[6]), .Z(n25369));
    L6MUX21 i22869 (.D0(n25364), .D1(n25365), .SD(index_i[6]), .Z(n25370));
    L6MUX21 i22870 (.D0(n25366), .D1(n25367), .SD(index_i[6]), .Z(n25371));
    PFUMX i22195 (.BLUT(n732_adj_3552), .ALUT(n763_adj_3659), .C0(index_i[5]), 
          .Z(n24696));
    L6MUX21 i22197 (.D0(n23604), .D1(n891_adj_3525), .SD(index_i[5]), 
            .Z(n24698));
    L6MUX21 i22200 (.D0(n24685), .D1(n24686), .SD(index_i[6]), .Z(n24701));
    L6MUX21 i22202 (.D0(n24689), .D1(n24690), .SD(index_i[6]), .Z(n24703));
    L6MUX21 i22203 (.D0(n24691), .D1(n24692), .SD(index_i[6]), .Z(n24704));
    L6MUX21 i22207 (.D0(n24699), .D1(n24700), .SD(index_i[6]), .Z(n24708));
    L6MUX21 i22264 (.D0(n24763), .D1(n24764), .SD(index_i[6]), .Z(n382));
    L6MUX21 i22271 (.D0(n24770), .D1(n24771), .SD(index_i[6]), .Z(n509));
    LUT4 n308_bdd_3_lut (.A(n32051), .B(n32038), .C(index_i[3]), .Z(n26564)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n308_bdd_3_lut.init = 16'hacac;
    PFUMX i26314 (.BLUT(n28180), .ALUT(n29105), .C0(index_i[5]), .Z(n28181));
    LUT4 i1_2_lut_rep_592 (.A(index_i[1]), .B(index_i[0]), .Z(n29252)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_2_lut_rep_592.init = 16'h8888;
    L6MUX21 i26269 (.D0(n28126), .D1(n29030), .SD(index_i[6]), .Z(n28127));
    PFUMX i26267 (.BLUT(n29035), .ALUT(n29046), .C0(index_i[7]), .Z(n28126));
    LUT4 mux_208_Mux_1_i348_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n348_adj_3660)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_1_i348_3_lut_4_lut_4_lut_4_lut.init = 16'h58f0;
    LUT4 i12879_3_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .Z(n12501)) /* synthesis lut_function=(!((B (C))+!A)) */ ;
    defparam i12879_3_lut.init = 16'h2a2a;
    LUT4 i13114_3_lut (.A(index_i[3]), .B(index_i[1]), .C(index_i[0]), 
         .Z(n15523)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i13114_3_lut.init = 16'hc8c8;
    LUT4 mux_208_Mux_3_i348_3_lut (.A(n32038), .B(n29233), .C(index_i[3]), 
         .Z(n348_adj_3594)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_3_i348_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_6_i668_3_lut (.A(n108), .B(n29341), .C(index_i[3]), 
         .Z(n668_adj_3527)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_6_i668_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_6_i684_3_lut (.A(n29214), .B(n32048), .C(index_i[3]), 
         .Z(n684_adj_3553)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_6_i684_3_lut.init = 16'hcaca;
    PFUMX i20954 (.BLUT(n23434), .ALUT(n23435), .C0(index_i[4]), .Z(n23436));
    LUT4 mux_208_Mux_3_i908_3_lut (.A(n29226), .B(n29412), .C(index_i[3]), 
         .Z(n908_adj_3507)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_3_i908_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_4_i828_3_lut_4_lut (.A(index_i[4]), .B(index_i[3]), 
         .C(n812), .D(n32053), .Z(n828_adj_3648)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_4_i828_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i20960 (.BLUT(n23440), .ALUT(n23441), .C0(index_i[4]), .Z(n23442));
    LUT4 mux_208_Mux_5_i797_3_lut_4_lut (.A(index_i[4]), .B(index_i[3]), 
         .C(n29529), .D(n29228), .Z(n797_adj_3635)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_5_i797_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i11260_3_lut_4_lut_3_lut (.A(index_i[1]), .B(index_i[0]), .C(index_i[4]), 
         .Z(n13559)) /* synthesis lut_function=(A (B)+!A !(B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11260_3_lut_4_lut_3_lut.init = 16'h9898;
    LUT4 mux_208_Mux_1_i763_3_lut_4_lut (.A(index_i[4]), .B(index_i[3]), 
         .C(n29584), .D(n29228), .Z(n763_adj_3659)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_1_i763_3_lut_4_lut.init = 16'hf1e0;
    L6MUX21 i22045 (.D0(n25043), .D1(n25050), .SD(index_i[6]), .Z(n24546));
    L6MUX21 i22048 (.D0(n23847), .D1(n23850), .SD(index_i[6]), .Z(n24549));
    L6MUX21 i22049 (.D0(n23853), .D1(n23856), .SD(index_i[6]), .Z(n24550));
    L6MUX21 i22050 (.D0(n23859), .D1(n23862), .SD(index_i[6]), .Z(n24551));
    PFUMX i22051 (.BLUT(n23865), .ALUT(n892_adj_3644), .C0(index_i[6]), 
          .Z(n24552));
    LUT4 i14388_2_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[0]), .C(n29362), 
         .D(index_i[2]), .Z(n16816)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i14388_2_lut_3_lut_4_lut.init = 16'hf080;
    LUT4 mux_208_Mux_7_i491_3_lut_4_lut_4_lut_4_lut_4_lut (.A(index_i[1]), 
         .B(index_i[0]), .C(index_i[2]), .D(index_i[3]), .Z(n491_adj_3653)) /* synthesis lut_function=(!(A (B (C+!(D))+!B ((D)+!C))+!A !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_7_i491_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'h5870;
    PFUMX i20963 (.BLUT(n23443), .ALUT(n23444), .C0(index_i[4]), .Z(n23445));
    LUT4 mux_208_Mux_7_i747_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), 
         .B(index_i[0]), .C(index_i[3]), .D(index_i[2]), .Z(n747_adj_3645)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))+!A (C (D)+!C !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_7_i747_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hf0a7;
    LUT4 i12990_3_lut_3_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n15399)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (D))+!A (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12990_3_lut_3_lut_3_lut_4_lut.init = 16'h00f7;
    LUT4 mux_208_Mux_2_i270_3_lut (.A(n29240), .B(n29237), .C(index_i[3]), 
         .Z(n270_adj_3502)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_2_i270_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_2_i316_3_lut (.A(n32040), .B(n29229), .C(index_i[3]), 
         .Z(n316_adj_3500)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_2_i316_3_lut.init = 16'hcaca;
    PFUMX i22123 (.BLUT(n94_adj_3654), .ALUT(n125), .C0(index_i[5]), .Z(n24624));
    PFUMX i20969 (.BLUT(n23449), .ALUT(n23450), .C0(index_i[4]), .Z(n23451));
    PFUMX i22184 (.BLUT(n13510), .ALUT(n62_adj_3661), .C0(index_i[5]), 
          .Z(n24685));
    L6MUX21 i26141 (.D0(n27955), .D1(n27952), .SD(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_1768[4]));
    LUT4 index_i_6__bdd_3_lut_26692_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(n29325), .D(index_i[6]), .Z(n28521)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam index_i_6__bdd_3_lut_26692_4_lut.init = 16'hf07f;
    PFUMX i26139 (.BLUT(n27954), .ALUT(n27953), .C0(index_i[8]), .Z(n27955));
    PFUMX i20972 (.BLUT(n23452), .ALUT(n23453), .C0(index_i[4]), .Z(n23454));
    PFUMX i26136 (.BLUT(n27951), .ALUT(n24619), .C0(index_i[8]), .Z(n27952));
    L6MUX21 i26121 (.D0(n27932), .D1(n27929), .SD(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_1768[9]));
    PFUMX i26119 (.BLUT(n27931), .ALUT(n27930), .C0(index_i[8]), .Z(n27932));
    LUT4 n518_bdd_3_lut_4_lut_4_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n26850)) /* synthesis lut_function=(A (B (C)+!B !(D))+!A !(D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n518_bdd_3_lut_4_lut_4_lut_3_lut_4_lut.init = 16'h80f7;
    PFUMX i22122 (.BLUT(n31_adj_3542), .ALUT(n62_adj_3655), .C0(index_i[5]), 
          .Z(n24623));
    PFUMX i26116 (.BLUT(n27928), .ALUT(n24542), .C0(index_i[8]), .Z(n27929));
    PFUMX i22091 (.BLUT(n31_adj_3539), .ALUT(n62), .C0(index_i[5]), .Z(n24592));
    PFUMX i22060 (.BLUT(n31), .ALUT(n23463), .C0(index_i[5]), .Z(n24561));
    LUT4 mux_208_Mux_6_i812_3_lut_4_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n812_adj_3520)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(D))+!A !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_6_i812_3_lut_4_lut_3_lut_4_lut.init = 16'h7780;
    LUT4 mux_208_Mux_2_i397_3_lut (.A(n32048), .B(n32030), .C(index_i[3]), 
         .Z(n397_adj_3499)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_2_i397_3_lut.init = 16'hcaca;
    LUT4 i12871_2_lut_rep_677 (.A(index_i[0]), .B(index_i[1]), .Z(n29337)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12871_2_lut_rep_677.init = 16'heeee;
    PFUMX i20984 (.BLUT(n23464), .ALUT(n23465), .C0(index_i[4]), .Z(n23466));
    LUT4 i14437_2_lut_rep_425_3_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n29085)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i14437_2_lut_rep_425_3_lut_4_lut.init = 16'hf080;
    LUT4 i12719_2_lut_rep_422_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n29082)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12719_2_lut_rep_422_3_lut_4_lut.init = 16'hfef0;
    LUT4 mux_208_Mux_7_i572_3_lut_rep_383_3_lut_3_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n29043)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_7_i572_3_lut_rep_383_3_lut_3_lut_4_lut.init = 16'hfe01;
    LUT4 i12718_2_lut_rep_496_3_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .Z(n29156)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12718_2_lut_rep_496_3_lut.init = 16'he0e0;
    LUT4 i14232_1_lut_rep_384_2_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n29044)) /* synthesis lut_function=(!(A (C+(D))+!A (B (C+(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i14232_1_lut_rep_384_2_lut_3_lut_4_lut.init = 16'h010f;
    PFUMX i22124 (.BLUT(n158_adj_3537), .ALUT(n189_adj_3566), .C0(index_i[5]), 
          .Z(n24625));
    LUT4 n179_bdd_3_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .Z(n27506)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n179_bdd_3_lut_4_lut_3_lut.init = 16'h6161;
    LUT4 i13124_3_lut_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n15533)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i13124_3_lut_3_lut_3_lut_4_lut.init = 16'h10ff;
    LUT4 mux_208_Mux_2_i931_3_lut_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n931)) /* synthesis lut_function=(!(A (B (C))+!A (B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_2_i931_3_lut_3_lut_3_lut.init = 16'h3e3e;
    LUT4 mux_208_Mux_0_i333_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n333)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_0_i333_3_lut_3_lut_4_lut.init = 16'hf10e;
    LUT4 mux_208_Mux_3_i30_3_lut_3_lut_4_lut_3_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n30_adj_3541)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_3_i30_3_lut_3_lut_4_lut_3_lut_4_lut.init = 16'hfe11;
    LUT4 i21103_3_lut_4_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n23585)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)+!C !(D)))+!A (B (C+!(D))+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21103_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'h0e30;
    LUT4 i22059_3_lut (.A(n24558), .B(n24559), .C(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_1768[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22059_3_lut.init = 16'hcaca;
    LUT4 i21057_3_lut_3_lut_4_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n23539)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21057_3_lut_3_lut_4_lut_3_lut_4_lut.init = 16'h11ef;
    LUT4 mux_208_Mux_8_i397_3_lut_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n397)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_8_i397_3_lut_3_lut_3_lut_4_lut.init = 16'hf10f;
    LUT4 i22632_3_lut (.A(n25131), .B(n25132), .C(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_1768[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22632_3_lut.init = 16'hcaca;
    LUT4 i22631_3_lut (.A(n25129), .B(n25130), .C(index_i[8]), .Z(n25132)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22631_3_lut.init = 16'hcaca;
    LUT4 i13018_2_lut_rep_491_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n29151)) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i13018_2_lut_rep_491_3_lut_4_lut.init = 16'he000;
    LUT4 mux_208_Mux_2_i142_3_lut_4_lut_4_lut_4_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n142_adj_3503)) /* synthesis lut_function=(!(A (B (D)+!B (C (D)+!C !(D)))+!A (B (D)+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_2_i142_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'h03ec;
    LUT4 mux_208_Mux_7_i141_3_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n141)) /* synthesis lut_function=(A ((C)+!B)+!A (B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_7_i141_3_lut_4_lut_3_lut.init = 16'he7e7;
    LUT4 n348_bdd_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n28915)) /* synthesis lut_function=(A (B (C)+!B (C+(D)))+!A (B (C)+!B !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n348_bdd_3_lut_4_lut_4_lut_4_lut.init = 16'he3f0;
    PFUMX i20987 (.BLUT(n23467), .ALUT(n23468), .C0(index_i[4]), .Z(n23469));
    LUT4 mux_208_Mux_3_i157_3_lut_3_lut_rep_432_3_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n29092)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_3_i157_3_lut_3_lut_rep_432_3_lut_4_lut.init = 16'h1ff0;
    L6MUX21 i22603 (.D0(n23442), .D1(n23445), .SD(index_i[5]), .Z(n25104));
    LUT4 mux_162_i16_3_lut (.A(\quarter_wave_sample_register_i[15] ), .B(o_val_pipeline_i_0__15__N_1799[15]), 
         .C(phase_negation_i[1]), .Z(n672[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam mux_162_i16_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_8_i46_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n46_adj_3488)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (D)+!B !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_8_i46_3_lut_4_lut_4_lut.init = 16'hcf10;
    PFUMX i22125 (.BLUT(n221), .ALUT(n252_adj_3560), .C0(index_i[5]), 
          .Z(n24626));
    LUT4 mux_162_i15_3_lut (.A(quarter_wave_sample_register_i[14]), .B(o_val_pipeline_i_0__15__N_1799[14]), 
         .C(phase_negation_i[1]), .Z(n672[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam mux_162_i15_3_lut.init = 16'hcaca;
    PFUMX i20990 (.BLUT(n23470), .ALUT(n23471), .C0(index_i[4]), .Z(n23472));
    LUT4 mux_162_i14_3_lut (.A(quarter_wave_sample_register_i[13]), .B(o_val_pipeline_i_0__15__N_1799[13]), 
         .C(phase_negation_i[1]), .Z(n672[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam mux_162_i14_3_lut.init = 16'hcaca;
    PFUMX i20993 (.BLUT(n23473), .ALUT(n23474), .C0(index_i[4]), .Z(n23475));
    LUT4 mux_162_i13_3_lut (.A(quarter_wave_sample_register_i[12]), .B(o_val_pipeline_i_0__15__N_1799[12]), 
         .C(phase_negation_i[1]), .Z(n672[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam mux_162_i13_3_lut.init = 16'hcaca;
    LUT4 mux_162_i12_3_lut (.A(quarter_wave_sample_register_i[11]), .B(o_val_pipeline_i_0__15__N_1799[11]), 
         .C(phase_negation_i[1]), .Z(n672[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam mux_162_i12_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_8_i506_3_lut_4_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n506_adj_3584)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_8_i506_3_lut_4_lut_3_lut_4_lut.init = 16'h0ef0;
    LUT4 mux_208_Mux_2_i716_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n716_adj_3491)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)+!C !(D)))+!A (B (D)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_2_i716_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h31cf;
    LUT4 i13067_2_lut_rep_611 (.A(index_i[2]), .B(index_i[0]), .Z(n29271)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i13067_2_lut_rep_611.init = 16'h8888;
    LUT4 i24386_3_lut (.A(n26587), .B(n25106), .C(index_i[6]), .Z(n25120)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24386_3_lut.init = 16'hcaca;
    LUT4 mux_162_i11_3_lut (.A(quarter_wave_sample_register_i[10]), .B(o_val_pipeline_i_0__15__N_1799[10]), 
         .C(phase_negation_i[1]), .Z(n672[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam mux_162_i11_3_lut.init = 16'hcaca;
    LUT4 mux_162_i10_3_lut (.A(quarter_wave_sample_register_i[9]), .B(o_val_pipeline_i_0__15__N_1799[9]), 
         .C(phase_negation_i[1]), .Z(n672[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam mux_162_i10_3_lut.init = 16'hcaca;
    L6MUX21 i22607 (.D0(n23451), .D1(n19994), .SD(index_i[5]), .Z(n25108));
    LUT4 mux_162_i9_3_lut (.A(quarter_wave_sample_register_i[8]), .B(o_val_pipeline_i_0__15__N_1799[8]), 
         .C(phase_negation_i[1]), .Z(n672[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam mux_162_i9_3_lut.init = 16'hcaca;
    LUT4 mux_162_i8_3_lut (.A(quarter_wave_sample_register_i[7]), .B(o_val_pipeline_i_0__15__N_1799[7]), 
         .C(phase_negation_i[1]), .Z(n672[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam mux_162_i8_3_lut.init = 16'hcaca;
    L6MUX21 i22608 (.D0(n23454), .D1(n13461), .SD(index_i[5]), .Z(n25109));
    LUT4 index_i_1__bdd_4_lut_27788 (.A(index_i[1]), .B(index_i[0]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n29588)) /* synthesis lut_function=(!(A (B (D)+!B (C+!(D)))+!A !(B (C (D)+!C !(D))+!B !((D)+!C)))) */ ;
    defparam index_i_1__bdd_4_lut_27788.init = 16'h429c;
    PFUMX i22126 (.BLUT(n286_adj_3532), .ALUT(n23517), .C0(index_i[5]), 
          .Z(n24627));
    LUT4 mux_162_i7_3_lut (.A(quarter_wave_sample_register_i[6]), .B(o_val_pipeline_i_0__15__N_1799[6]), 
         .C(phase_negation_i[1]), .Z(n672[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam mux_162_i7_3_lut.init = 16'hcaca;
    LUT4 mux_162_i6_3_lut (.A(quarter_wave_sample_register_i[5]), .B(o_val_pipeline_i_0__15__N_1799[5]), 
         .C(phase_negation_i[1]), .Z(n672[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam mux_162_i6_3_lut.init = 16'hcaca;
    LUT4 mux_162_i5_3_lut (.A(quarter_wave_sample_register_i[4]), .B(o_val_pipeline_i_0__15__N_1799[4]), 
         .C(phase_negation_i[1]), .Z(n672[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam mux_162_i5_3_lut.init = 16'hcaca;
    LUT4 mux_162_i4_3_lut (.A(quarter_wave_sample_register_i[3]), .B(o_val_pipeline_i_0__15__N_1799[3]), 
         .C(phase_negation_i[1]), .Z(n672[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam mux_162_i4_3_lut.init = 16'hcaca;
    PFUMX i22610 (.BLUT(n542_adj_3531), .ALUT(n573_adj_3637), .C0(index_i[5]), 
          .Z(n25111));
    LUT4 mux_162_i3_3_lut (.A(quarter_wave_sample_register_i[2]), .B(o_val_pipeline_i_0__15__N_1799[2]), 
         .C(phase_negation_i[1]), .Z(n672[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam mux_162_i3_3_lut.init = 16'hcaca;
    LUT4 mux_162_i2_3_lut (.A(quarter_wave_sample_register_i[1]), .B(o_val_pipeline_i_0__15__N_1799[1]), 
         .C(phase_negation_i[1]), .Z(n672[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam mux_162_i2_3_lut.init = 16'hcaca;
    LUT4 mux_162_i1_3_lut (.A(quarter_wave_sample_register_i[0]), .B(o_val_pipeline_i_0__15__N_1799[0]), 
         .C(phase_negation_i[1]), .Z(n672[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam mux_162_i1_3_lut.init = 16'hcaca;
    LUT4 i7131_2_lut (.A(phase_i[9]), .B(phase_i[10]), .Z(index_i_9__N_1748[9])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(60[14] 63[8])
    defparam i7131_2_lut.init = 16'h6666;
    LUT4 i7132_2_lut (.A(phase_i[8]), .B(phase_i[10]), .Z(index_i_9__N_1748[8])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(60[14] 63[8])
    defparam i7132_2_lut.init = 16'h6666;
    LUT4 i7133_2_lut (.A(phase_i[7]), .B(phase_i[10]), .Z(index_i_9__N_1748[7])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(60[14] 63[8])
    defparam i7133_2_lut.init = 16'h6666;
    LUT4 i7134_2_lut (.A(phase_i[6]), .B(phase_i[10]), .Z(index_i_9__N_1748[6])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(60[14] 63[8])
    defparam i7134_2_lut.init = 16'h6666;
    LUT4 i7135_2_lut (.A(phase_i[5]), .B(phase_i[10]), .Z(index_i_9__N_1748[5])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(60[14] 63[8])
    defparam i7135_2_lut.init = 16'h6666;
    LUT4 i7136_2_lut (.A(phase_i[4]), .B(phase_i[10]), .Z(index_i_9__N_1748[4])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(60[14] 63[8])
    defparam i7136_2_lut.init = 16'h6666;
    LUT4 i7137_2_lut (.A(phase_i[3]), .B(phase_i[10]), .Z(index_i_9__N_1748[3])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(60[14] 63[8])
    defparam i7137_2_lut.init = 16'h6666;
    PFUMX i22127 (.BLUT(n349_adj_3595), .ALUT(n23520), .C0(index_i[5]), 
          .Z(n24628));
    LUT4 i7138_2_lut (.A(phase_i[2]), .B(phase_i[10]), .Z(index_i_9__N_1748[2])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(60[14] 63[8])
    defparam i7138_2_lut.init = 16'h6666;
    LUT4 i13180_2_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n635)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A (B (C+!(D))+!B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i13180_2_lut_4_lut_4_lut.init = 16'hf1fc;
    LUT4 i21094_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n23576)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B ((D)+!C)+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21094_3_lut_4_lut_4_lut.init = 16'hfc1c;
    LUT4 i22405_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n24906)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A !(C (D)+!C !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i22405_3_lut_4_lut_4_lut_4_lut.init = 16'h85f0;
    LUT4 i7139_2_lut (.A(phase_i[1]), .B(phase_i[10]), .Z(index_i_9__N_1748[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(60[14] 63[8])
    defparam i7139_2_lut.init = 16'h6666;
    LUT4 i21084_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n23566)) /* synthesis lut_function=(A (B (D)+!B ((D)+!C))+!A (B (D)+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21084_3_lut_4_lut_4_lut_4_lut.init = 16'hfe13;
    PFUMX i22128 (.BLUT(n413_adj_3529), .ALUT(n444_adj_3662), .C0(index_i[5]), 
          .Z(n24629));
    PFUMX i20999 (.BLUT(n23479), .ALUT(n23480), .C0(index_i[4]), .Z(n23481));
    PFUMX i22611 (.BLUT(n605), .ALUT(n636_adj_3592), .C0(index_i[5]), 
          .Z(n25112));
    PFUMX i28943 (.BLUT(n32059), .ALUT(n32060), .C0(index_i[1]), .Z(n32061));
    LUT4 mux_208_Mux_7_i92_3_lut_rep_679 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29339)) /* synthesis lut_function=(A (B+!(C))+!A !((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_7_i92_3_lut_rep_679.init = 16'h8e8e;
    LUT4 mux_208_Mux_7_i300_3_lut_rep_680 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29340)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_7_i300_3_lut_rep_680.init = 16'h1c1c;
    PFUMX i26025 (.BLUT(n27824), .ALUT(n1022), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_1768[12]));
    LUT4 mux_208_Mux_7_i134_3_lut_4_lut_3_lut_rep_681 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29341)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_7_i134_3_lut_4_lut_3_lut_rep_681.init = 16'h1818;
    PFUMX i22849 (.BLUT(n716_adj_3505), .ALUT(n731_adj_3558), .C0(index_i[4]), 
          .Z(n25350));
    LUT4 mux_208_Mux_7_i691_3_lut_rep_683 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29343)) /* synthesis lut_function=(!(A (B (C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_7_i691_3_lut_rep_683.init = 16'h7e7e;
    LUT4 mux_208_Mux_6_i645_3_lut_3_lut_4_lut_3_lut_rep_684 (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[2]), .Z(n29344)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_6_i645_3_lut_3_lut_4_lut_3_lut_rep_684.init = 16'h1919;
    PFUMX i22612 (.BLUT(n669_adj_3528), .ALUT(n700_adj_3554), .C0(index_i[5]), 
          .Z(n25113));
    PFUMX i24868 (.BLUT(n26481), .ALUT(n26478), .C0(index_i[6]), .Z(n26482));
    PFUMX i22613 (.BLUT(n732_adj_3551), .ALUT(n23460), .C0(index_i[5]), 
          .Z(n25114));
    PFUMX i22614 (.BLUT(n797_adj_3523), .ALUT(n828_adj_3521), .C0(index_i[5]), 
          .Z(n25115));
    LUT4 mux_208_Mux_5_i53_3_lut_4_lut_3_lut_rep_685 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29345)) /* synthesis lut_function=(A ((C)+!B)+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_5_i53_3_lut_4_lut_3_lut_rep_685.init = 16'he6e6;
    PFUMX i22615 (.BLUT(n860_adj_3487), .ALUT(n891_adj_3519), .C0(index_i[5]), 
          .Z(n25116));
    LUT4 mux_208_Mux_0_i557_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n557)) /* synthesis lut_function=(A ((D)+!C)+!A !((D)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_0_i557_3_lut_4_lut.init = 16'haa4e;
    LUT4 mux_208_Mux_6_i635_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n635_adj_3591)) /* synthesis lut_function=(A (B (C+(D))+!B !(D))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_6_i635_3_lut_4_lut.init = 16'hcce6;
    LUT4 i20979_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n23461)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(D))+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20979_3_lut_3_lut_4_lut.init = 16'h3319;
    PFUMX i26021 (.BLUT(n254_adj_3663), .ALUT(n27818), .C0(index_i[8]), 
          .Z(n27819));
    LUT4 mux_208_Mux_8_i30_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n30_adj_3543)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A !(B ((D)+!C)+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_8_i30_3_lut_3_lut_4_lut.init = 16'h7e0f;
    LUT4 mux_208_Mux_8_i285_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n285_adj_3664)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C (D)+!C !(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_8_i285_3_lut_3_lut_4_lut.init = 16'h0fc1;
    PFUMX i22129 (.BLUT(n476_adj_3514), .ALUT(n507_adj_3627), .C0(index_i[5]), 
          .Z(n24630));
    LUT4 mux_208_Mux_2_i557_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n557_adj_3570)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C+!(D))+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_2_i557_3_lut_3_lut_4_lut.init = 16'h0f18;
    LUT4 i21082_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n23564)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A (B (D)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21082_3_lut_4_lut.init = 16'h18cc;
    LUT4 i21040_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n23522)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21040_3_lut_3_lut_4_lut.init = 16'h0f1c;
    LUT4 i21117_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n23599)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C (D)))+!A (B (C+(D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21117_4_lut_4_lut_4_lut.init = 16'h301c;
    PFUMX i22130 (.BLUT(n23523), .ALUT(n573_adj_3572), .C0(index_i[5]), 
          .Z(n24631));
    LUT4 mux_208_Mux_0_i699_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n699_adj_3651)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (D))+!A (B (C+!(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_0_i699_3_lut_3_lut_4_lut.init = 16'h1c33;
    LUT4 i21039_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n23521)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)))+!A !(B (C+!(D))+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21039_3_lut_3_lut_4_lut.init = 16'h71cc;
    LUT4 mux_208_Mux_7_i716_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n716_adj_3646)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C+!(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_7_i716_3_lut_3_lut_4_lut.init = 16'h0f81;
    LUT4 mux_208_Mux_8_i635_3_lut_4_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n635_adj_3473)) /* synthesis lut_function=(!(A (B (C (D))+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_8_i635_3_lut_4_lut_3_lut_4_lut.init = 16'h0ff8;
    PFUMX i22131 (.BLUT(n13497), .ALUT(n23526), .C0(index_i[5]), .Z(n24632));
    LUT4 i21102_3_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[0]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n23584)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21102_3_lut_4_lut_4_lut.init = 16'h5a8a;
    LUT4 i14255_2_lut_rep_689 (.A(index_i[1]), .B(index_i[2]), .Z(n29349)) /* synthesis lut_function=(A (B)) */ ;
    defparam i14255_2_lut_rep_689.init = 16'h8888;
    PFUMX i22132 (.BLUT(n669_adj_3511), .ALUT(n700_adj_3614), .C0(index_i[5]), 
          .Z(n24633));
    LUT4 mux_208_Mux_9_i30_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .D(index_i[3]), .Z(n30_adj_3546)) /* synthesis lut_function=(A (B (C (D))+!B !(D))+!A !(B+(D))) */ ;
    defparam mux_208_Mux_9_i30_3_lut_4_lut_4_lut_4_lut.init = 16'h8033;
    L6MUX21 i22133 (.D0(n23529), .D1(n763), .SD(index_i[5]), .Z(n24634));
    LUT4 i12916_2_lut_rep_443_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[0]), 
         .Z(n29103)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i12916_2_lut_rep_443_3_lut.init = 16'h8080;
    LUT4 n699_bdd_4_lut_26588_4_lut_4_lut (.A(index_i[0]), .B(n29349), .C(index_i[4]), 
         .D(index_i[3]), .Z(n28180)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (D))+!A (B (C (D)+!C !(D))+!B (D)))) */ ;
    defparam n699_bdd_4_lut_26588_4_lut_4_lut.init = 16'h0c73;
    PFUMX i22135 (.BLUT(n860_adj_3574), .ALUT(n891), .C0(index_i[5]), 
          .Z(n24636));
    LUT4 i11205_2_lut_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[3]), 
         .Z(n13501)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i11205_2_lut_3_lut.init = 16'h8080;
    LUT4 mux_208_Mux_9_i412_3_lut_3_lut_4_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .Z(n412_adj_3559)) /* synthesis lut_function=(!(A (B (C))+!A !(B+(C)))) */ ;
    defparam mux_208_Mux_9_i412_3_lut_3_lut_4_lut_3_lut.init = 16'h7e7e;
    LUT4 mux_208_Mux_3_i142_3_lut_3_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .Z(n142_adj_3493)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B+!(C)))) */ ;
    defparam mux_208_Mux_3_i142_3_lut_3_lut_3_lut.init = 16'h3838;
    PFUMX i25989 (.BLUT(n27775), .ALUT(n27773), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_1768[10]));
    LUT4 i14439_2_lut_rep_396_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n29056)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;
    defparam i14439_2_lut_rep_396_3_lut_4_lut.init = 16'hf8f0;
    LUT4 i17681_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n19995)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C (D)+!C !(D)))+!A !(B (D)+!B (C (D)+!C !(D)))) */ ;
    defparam i17681_3_lut_4_lut_4_lut_4_lut.init = 16'h83fc;
    LUT4 mux_208_Mux_8_i491_3_lut_4_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .D(index_i[3]), .Z(n491_adj_3652)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(D))+!A !(D))) */ ;
    defparam mux_208_Mux_8_i491_3_lut_4_lut_3_lut_4_lut.init = 16'h7780;
    LUT4 i12788_2_lut_rep_529_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[3]), 
         .Z(n29189)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam i12788_2_lut_rep_529_3_lut.init = 16'hf8f8;
    PFUMX i22136 (.BLUT(n924_adj_3508), .ALUT(n23532), .C0(index_i[5]), 
          .Z(n24637));
    LUT4 i13827_2_lut_rep_548_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[0]), 
         .Z(n29208)) /* synthesis lut_function=(A (B+!(C))+!A !(C)) */ ;
    defparam i13827_2_lut_rep_548_3_lut.init = 16'h8f8f;
    LUT4 i12764_3_lut_4_lut (.A(index_i[0]), .B(n29349), .C(n29261), .D(index_i[5]), 
         .Z(n318)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (C (D))) */ ;
    defparam i12764_3_lut_4_lut.init = 16'hf800;
    LUT4 i21022_3_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[3]), 
         .D(index_i[0]), .Z(n23504)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D))) */ ;
    defparam i21022_3_lut_3_lut_4_lut.init = 16'hf80f;
    LUT4 i21064_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .D(index_i[3]), .Z(n23546)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(D))+!A (B+!(D)))) */ ;
    defparam i21064_3_lut_4_lut_4_lut_4_lut.init = 16'h3380;
    LUT4 mux_208_Mux_8_i412_3_lut_4_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .Z(n16698)) /* synthesis lut_function=(A (B+!(C))+!A !((C)+!B)) */ ;
    defparam mux_208_Mux_8_i412_3_lut_4_lut_3_lut.init = 16'h8e8e;
    LUT4 i12914_2_lut_rep_690 (.A(index_i[1]), .B(index_i[2]), .C(index_i[0]), 
         .Z(n29350)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i12914_2_lut_rep_690.init = 16'h7070;
    LUT4 mux_208_Mux_0_i1017_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .D(index_i[3]), .Z(n1017)) /* synthesis lut_function=(A (B (D)+!B !((D)+!C))+!A (C+(D))) */ ;
    defparam mux_208_Mux_0_i1017_4_lut_4_lut_4_lut.init = 16'hdd70;
    PFUMX i22137 (.BLUT(n23535), .ALUT(n1018), .C0(index_i[5]), .Z(n24638));
    LUT4 index_i_6__bdd_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[6]), .D(n29363), .Z(n28520)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam index_i_6__bdd_4_lut_4_lut_4_lut.init = 16'h0f7a;
    PFUMX i25987 (.BLUT(n23278), .ALUT(n27771), .C0(index_i[7]), .Z(n27772));
    LUT4 i24597_2_lut_rep_699 (.A(index_i[4]), .B(index_i[3]), .Z(n29359)) /* synthesis lut_function=((B)+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i24597_2_lut_rep_699.init = 16'hdddd;
    LUT4 mux_208_Mux_3_i797_3_lut_4_lut (.A(index_i[4]), .B(index_i[3]), 
         .C(n796_adj_3658), .D(n29256), .Z(n797)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_3_i797_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i27894 (.BLUT(n30601), .ALUT(n30600), .C0(index_i[3]), .Z(n30602));
    PFUMX i27892 (.BLUT(n30597), .ALUT(n30596), .C0(index_i[2]), .Z(n30598));
    PFUMX i22155 (.BLUT(n158), .ALUT(n189_adj_3497), .C0(index_i[5]), 
          .Z(n24656));
    LUT4 i14233_2_lut_rep_702 (.A(index_i[3]), .B(index_i[4]), .Z(n29362)) /* synthesis lut_function=(A (B)) */ ;
    defparam i14233_2_lut_rep_702.init = 16'h8888;
    LUT4 i14239_2_lut_3_lut (.A(index_i[3]), .B(index_i[4]), .C(index_i[5]), 
         .Z(n16658)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam i14239_2_lut_3_lut.init = 16'hf8f8;
    LUT4 i22678_3_lut_3_lut_4_lut (.A(index_i[3]), .B(index_i[4]), .C(n413_adj_3556), 
         .D(index_i[5]), .Z(n25179)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(C+(D)))) */ ;
    defparam i22678_3_lut_3_lut_4_lut.init = 16'h77f0;
    PFUMX i22156 (.BLUT(n221_adj_3656), .ALUT(n23541), .C0(index_i[5]), 
          .Z(n24657));
    LUT4 i1_2_lut_3_lut (.A(index_i[3]), .B(index_i[4]), .C(index_i[5]), 
         .Z(n22324)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h8080;
    LUT4 i11199_3_lut_3_lut_3_lut_4_lut (.A(index_i[3]), .B(index_i[4]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n444_adj_3506)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C))+!A (C))) */ ;
    defparam i11199_3_lut_3_lut_3_lut_4_lut.init = 16'h0f87;
    LUT4 i1_2_lut_rep_703 (.A(index_i[3]), .B(index_i[2]), .Z(n29363)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_2_lut_rep_703.init = 16'heeee;
    LUT4 i11167_3_lut_3_lut_rep_570_4_lut (.A(index_i[3]), .B(index_i[2]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n29230)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11167_3_lut_3_lut_rep_570_4_lut.init = 16'h1ef0;
    LUT4 i11208_3_lut_4_lut_3_lut_4_lut (.A(index_i[3]), .B(index_i[2]), 
         .C(index_i[0]), .D(index_i[1]), .Z(n844_adj_3515)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11208_3_lut_4_lut_3_lut_4_lut.init = 16'hf00e;
    LUT4 i24725_2_lut_rep_490_3_lut_4_lut (.A(index_i[3]), .B(index_i[2]), 
         .C(index_i[0]), .D(index_i[1]), .Z(n29150)) /* synthesis lut_function=(!(A+(B+(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i24725_2_lut_rep_490_3_lut_4_lut.init = 16'h0111;
    LUT4 n526_bdd_3_lut_25828_3_lut_3_lut_4_lut (.A(index_i[3]), .B(index_i[2]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n26852)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n526_bdd_3_lut_25828_3_lut_3_lut_4_lut.init = 16'h0fe1;
    LUT4 i12988_2_lut_rep_502_3_lut (.A(index_i[3]), .B(index_i[2]), .C(index_i[1]), 
         .Z(n29162)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12988_2_lut_rep_502_3_lut.init = 16'hfefe;
    LUT4 mux_208_Mux_8_i653_3_lut_rep_400_4_lut (.A(index_i[0]), .B(n29349), 
         .C(index_i[3]), .D(n29156), .Z(n29060)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(C+(D)))) */ ;
    defparam mux_208_Mux_8_i653_3_lut_rep_400_4_lut.init = 16'h7f70;
    L6MUX21 i27819 (.D0(n30486), .D1(n30483), .SD(index_i[5]), .Z(n30487));
    PFUMX i27817 (.BLUT(n30485), .ALUT(n30484), .C0(index_i[3]), .Z(n30486));
    PFUMX i27815 (.BLUT(n30482), .ALUT(n30481), .C0(index_i[3]), .Z(n30483));
    PFUMX i22157 (.BLUT(n286), .ALUT(n317_adj_3501), .C0(index_i[5]), 
          .Z(n24658));
    LUT4 i13072_3_lut (.A(index_i[3]), .B(index_i[1]), .C(index_i[0]), 
         .Z(n15481)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i13072_3_lut.init = 16'hecec;
    PFUMX i27105 (.BLUT(n29530), .ALUT(n29531), .C0(index_i[1]), .Z(n29532));
    L6MUX21 i25895 (.D0(n27647), .D1(n27644), .SD(index_i[5]), .Z(n27648));
    PFUMX i25893 (.BLUT(n27646), .ALUT(n27645), .C0(index_i[4]), .Z(n27647));
    PFUMX i25890 (.BLUT(n27643), .ALUT(n908_adj_3602), .C0(index_i[4]), 
          .Z(n27644));
    LUT4 mux_208_Mux_3_i668_3_lut_4_lut (.A(n29212), .B(index_i[2]), .C(index_i[3]), 
         .D(n29239), .Z(n668)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_3_i668_3_lut_4_lut.init = 16'h6f60;
    LUT4 n53_bdd_3_lut_24925_4_lut (.A(n29212), .B(index_i[2]), .C(n32042), 
         .D(index_i[3]), .Z(n26548)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n53_bdd_3_lut_24925_4_lut.init = 16'hf066;
    LUT4 n676_bdd_2_lut_25787_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n26865)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n676_bdd_2_lut_25787_4_lut_4_lut_4_lut.init = 16'h0058;
    PFUMX i22158 (.BLUT(n349_adj_3665), .ALUT(n23544), .C0(index_i[5]), 
          .Z(n24659));
    PFUMX i22159 (.BLUT(n413), .ALUT(n23547), .C0(index_i[5]), .Z(n24660));
    PFUMX i21032 (.BLUT(n23512), .ALUT(n23513), .C0(index_i[4]), .Z(n23514));
    LUT4 mux_208_Mux_4_i763_3_lut_4_lut (.A(n29212), .B(index_i[2]), .C(index_i[4]), 
         .D(n747_adj_3489), .Z(n763_adj_3641)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_4_i763_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_208_Mux_2_i731_3_lut_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n731)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(B (C)+!B !(C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_2_i731_3_lut_3_lut_4_lut.init = 16'h69f0;
    LUT4 mux_208_Mux_8_i526_3_lut_3_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n526_adj_3472)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_8_i526_3_lut_3_lut_3_lut_4_lut.init = 16'h0f70;
    LUT4 mux_208_Mux_1_i924_3_lut (.A(n908_adj_3602), .B(n412_adj_3559), 
         .C(index_i[4]), .Z(n924)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_1_i924_3_lut.init = 16'hcaca;
    PFUMX i22160 (.BLUT(n23550), .ALUT(n507_adj_3666), .C0(index_i[5]), 
          .Z(n24661));
    LUT4 i23999_3_lut (.A(n23593), .B(n23594), .C(index_i[4]), .Z(n23595)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23999_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_rep_445_4_lut (.A(index_i[1]), .B(index_i[0]), .C(index_i[2]), 
         .D(n29261), .Z(n29105)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_3_lut_rep_445_4_lut.init = 16'hfff8;
    PFUMX i22161 (.BLUT(n23553), .ALUT(n573_adj_3571), .C0(index_i[5]), 
          .Z(n24662));
    LUT4 mux_208_Mux_12_i254_4_lut (.A(n29046), .B(n22324), .C(index_i[6]), 
         .D(n29182), .Z(n254_adj_3663)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_12_i254_4_lut.init = 16'hca0a;
    FD1S3BX quarter_wave_sample_register_i_i14 (.D(quarter_wave_sample_register_i_15__N_1768[14]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_i[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_i_i14.GSR = "DISABLED";
    PFUMX i27103 (.BLUT(n29527), .ALUT(n29528), .C0(index_i[1]), .Z(n29529));
    LUT4 mux_208_Mux_3_i1002_3_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n21724)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (D))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_3_i1002_3_lut_3_lut_4_lut.init = 16'hf708;
    LUT4 mux_208_Mux_1_i349_3_lut (.A(n506_adj_3584), .B(n348_adj_3660), 
         .C(index_i[4]), .Z(n349)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_1_i349_3_lut.init = 16'hcaca;
    LUT4 i24008_3_lut (.A(n23569), .B(n23570), .C(index_i[4]), .Z(n23571)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24008_3_lut.init = 16'hcaca;
    FD1S3BX quarter_wave_sample_register_i_i13 (.D(quarter_wave_sample_register_i_15__N_1768[13]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_i[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_i_i13.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i12 (.D(quarter_wave_sample_register_i_15__N_1768[12]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_i[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_i_i12.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i11 (.D(quarter_wave_sample_register_i_15__N_1768[11]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_i[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_i_i11.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i10 (.D(quarter_wave_sample_register_i_15__N_1768[10]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_i[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_i_i10.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i9 (.D(quarter_wave_sample_register_i_15__N_1768[9]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_i[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_i_i9.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i8 (.D(quarter_wave_sample_register_i_15__N_1768[8]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_i[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_i_i8.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i7 (.D(quarter_wave_sample_register_i_15__N_1768[7]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_i[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_i_i7.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i6 (.D(quarter_wave_sample_register_i_15__N_1768[6]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_i[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_i_i6.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i5 (.D(quarter_wave_sample_register_i_15__N_1768[5]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_i[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_i_i5.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i4 (.D(quarter_wave_sample_register_i_15__N_1768[4]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_i[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_i_i4.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i3 (.D(quarter_wave_sample_register_i_15__N_1768[3]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_i[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_i_i3.GSR = "DISABLED";
    PFUMX i22162 (.BLUT(n605_adj_3495), .ALUT(n23556), .C0(index_i[5]), 
          .Z(n24663));
    FD1S3BX quarter_wave_sample_register_i_i2 (.D(quarter_wave_sample_register_i_15__N_1768[2]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_i[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_i_i2.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i1 (.D(quarter_wave_sample_register_i_15__N_1768[1]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_i[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_i_i1.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i32 (.D(n672[15]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_i[0] [15])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i32.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i31 (.D(n672[14]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_i[0] [14])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i31.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i30 (.D(n672[13]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_i[0] [13])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i30.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i29 (.D(n672[12]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_i[0] [12])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i29.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i28 (.D(n672[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_i[0] [11])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i28.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i27 (.D(n672[10]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_i[0] [10])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i27.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i26 (.D(n672[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_i[0] [9])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i26.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i25 (.D(n672[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_i[0] [8])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i25.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i24 (.D(n672[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_i[0] [7])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i24.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i23 (.D(n672[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_i[0] [6])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i23.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i22 (.D(n672[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_i[0] [5])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i22.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i21 (.D(n672[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_i[0] [4])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i21.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i20 (.D(n672[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_i[0] [3])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i20.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i19 (.D(n672[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_i[0] [2])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i19.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i18 (.D(n672[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_i[0] [1])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i18.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i17 (.D(n672[0]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_i[0] [0])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i17.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i16 (.D(\o_val_pipeline_i[0] [15]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(modulation_output[15])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i16.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i15 (.D(\o_val_pipeline_i[0] [14]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(modulation_output[14])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i15.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i14 (.D(\o_val_pipeline_i[0] [13]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(modulation_output[13])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i14.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i13 (.D(\o_val_pipeline_i[0] [12]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(modulation_output[12])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i13.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i12 (.D(\o_val_pipeline_i[0] [11]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(modulation_output[11])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i12.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i11 (.D(\o_val_pipeline_i[0] [10]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(modulation_output[10])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i11.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i10 (.D(\o_val_pipeline_i[0] [9]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(modulation_output[9])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i10.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i9 (.D(\o_val_pipeline_i[0] [8]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(modulation_output[8])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i9.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i8 (.D(\o_val_pipeline_i[0] [7]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(modulation_output[7])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i8.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i7 (.D(\o_val_pipeline_i[0] [6]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(modulation_output[6])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i7.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i6 (.D(\o_val_pipeline_i[0] [5]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(modulation_output[5])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i6.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i5 (.D(\o_val_pipeline_i[0] [4]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(modulation_output[4])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i5.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i4 (.D(\o_val_pipeline_i[0] [3]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(modulation_output[3])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i4.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i3 (.D(\o_val_pipeline_i[0] [2]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(modulation_output[2])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i3.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i2 (.D(\o_val_pipeline_i[0] [1]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(modulation_output[1])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i2.GSR = "DISABLED";
    FD1S3DX index_i_i9 (.D(index_i_9__N_1748[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(index_i[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam index_i_i9.GSR = "DISABLED";
    FD1S3DX index_i_i8 (.D(index_i_9__N_1748[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(index_i[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam index_i_i8.GSR = "DISABLED";
    LUT4 n45_bdd_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n27452)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n45_bdd_3_lut_4_lut_4_lut_4_lut.init = 16'h0f58;
    FD1S3DX index_i_i7 (.D(index_i_9__N_1748[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(index_i[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam index_i_i7.GSR = "DISABLED";
    FD1S3DX index_i_i6 (.D(index_i_9__N_1748[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(index_i[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam index_i_i6.GSR = "DISABLED";
    FD1S3DX index_i_i5 (.D(index_i_9__N_1748[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(index_i[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam index_i_i5.GSR = "DISABLED";
    FD1S3DX index_i_i4 (.D(index_i_9__N_1748[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(index_i[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam index_i_i4.GSR = "DISABLED";
    LUT4 mux_208_Mux_7_i526_3_lut_4_lut_4_lut_3_lut_4_lut (.A(index_i[1]), 
         .B(index_i[0]), .C(index_i[3]), .D(index_i[2]), .Z(n526_adj_3649)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(D))+!A !(D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_7_i526_3_lut_4_lut_4_lut_3_lut_4_lut.init = 16'h887f;
    FD1S3DX index_i_i3 (.D(index_i_9__N_1748[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(index_i[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam index_i_i3.GSR = "DISABLED";
    FD1S3DX index_i_i2 (.D(index_i_9__N_1748[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(index_i[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam index_i_i2.GSR = "DISABLED";
    FD1S3DX index_i_i1 (.D(index_i_9__N_1748[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(index_i[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam index_i_i1.GSR = "DISABLED";
    FD1S3DX phase_negation_i_i1 (.D(phase_negation_i[0]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(phase_negation_i[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam phase_negation_i_i1.GSR = "DISABLED";
    PFUMX i22163 (.BLUT(n669), .ALUT(n700_adj_3522), .C0(index_i[5]), 
          .Z(n24664));
    LUT4 mux_208_Mux_4_i1002_3_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n1002_adj_3576)) /* synthesis lut_function=(A (B (C (D))+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_4_i1002_3_lut_3_lut_4_lut.init = 16'hf007;
    LUT4 mux_208_Mux_1_i94_3_lut (.A(index_i[0]), .B(n93_adj_3667), .C(index_i[4]), 
         .Z(n94)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_1_i94_3_lut.init = 16'hcaca;
    LUT4 n269_bdd_3_lut_24933 (.A(n32052), .B(index_i[3]), .C(n29234), 
         .Z(n26555)) /* synthesis lut_function=(A (B+(C))+!A !(B+!(C))) */ ;
    defparam n269_bdd_3_lut_24933.init = 16'hb8b8;
    LUT4 i21097_3_lut_4_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n23579)) /* synthesis lut_function=(!(A (B (C)+!B (C+(D)))+!A !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21097_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'h585f;
    PFUMX i25756 (.BLUT(n27506), .ALUT(n32048), .C0(index_i[3]), .Z(n27507));
    FD1P3AX phase_i_i0_i11 (.D(o_phase[11]), .SP(dac_clk_p_c_enable_630), 
            .CK(dac_clk_p_c), .Q(phase_i[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam phase_i_i0_i11.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i10 (.D(o_phase[10]), .SP(dac_clk_p_c_enable_630), 
            .CK(dac_clk_p_c), .Q(phase_i[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam phase_i_i0_i10.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i9 (.D(o_phase[9]), .SP(dac_clk_p_c_enable_630), 
            .CK(dac_clk_p_c), .Q(phase_i[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam phase_i_i0_i9.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i8 (.D(o_phase[8]), .SP(dac_clk_p_c_enable_630), 
            .CK(dac_clk_p_c), .Q(phase_i[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam phase_i_i0_i8.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i7 (.D(o_phase[7]), .SP(dac_clk_p_c_enable_630), 
            .CK(dac_clk_p_c), .Q(phase_i[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam phase_i_i0_i7.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i6 (.D(o_phase[6]), .SP(dac_clk_p_c_enable_630), 
            .CK(dac_clk_p_c), .Q(phase_i[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam phase_i_i0_i6.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i5 (.D(o_phase[5]), .SP(dac_clk_p_c_enable_630), 
            .CK(dac_clk_p_c), .Q(phase_i[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam phase_i_i0_i5.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i4 (.D(o_phase[4]), .SP(dac_clk_p_c_enable_630), 
            .CK(dac_clk_p_c), .Q(phase_i[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam phase_i_i0_i4.GSR = "DISABLED";
    PFUMX i21047 (.BLUT(n23527), .ALUT(n23528), .C0(index_i[4]), .Z(n23529));
    FD1P3AX phase_i_i0_i3 (.D(o_phase[3]), .SP(dac_clk_p_c_enable_630), 
            .CK(dac_clk_p_c), .Q(phase_i[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam phase_i_i0_i3.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i2 (.D(o_phase[2]), .SP(dac_clk_p_c_enable_630), 
            .CK(dac_clk_p_c), .Q(phase_i[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam phase_i_i0_i2.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i1 (.D(o_phase[1]), .SP(dac_clk_p_c_enable_630), 
            .CK(dac_clk_p_c), .Q(phase_i[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam phase_i_i0_i1.GSR = "DISABLED";
    PFUMX i22164 (.BLUT(n732), .ALUT(n763_adj_3668), .C0(index_i[5]), 
          .Z(n24665));
    LUT4 i14454_3_lut_4_lut (.A(n29325), .B(index_i[4]), .C(index_i[5]), 
         .D(n29337), .Z(n16886)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i14454_3_lut_4_lut.init = 16'hf8f0;
    LUT4 i12763_2_lut_rep_522_3_lut (.A(index_i[1]), .B(index_i[0]), .C(index_i[2]), 
         .Z(n29182)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12763_2_lut_rep_522_3_lut.init = 16'hf8f8;
    LUT4 i12801_2_lut_rep_415_3_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[4]), .D(n29325), .Z(n29075)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12801_2_lut_rep_415_3_lut_4_lut.init = 16'hf8f0;
    LUT4 mux_208_Mux_0_i475_3_lut_4_lut (.A(n29271), .B(index_i[1]), .C(index_i[3]), 
         .D(n29182), .Z(n475_adj_3623)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_0_i475_3_lut_4_lut.init = 16'h4f40;
    PFUMX i25703 (.BLUT(n27452), .ALUT(n27451), .C0(index_i[4]), .Z(n27453));
    LUT4 mux_208_Mux_2_i836_3_lut_4_lut_3_lut_rep_595 (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[2]), .Z(n29255)) /* synthesis lut_function=(A (B)+!A !(B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_2_i836_3_lut_4_lut_3_lut_rep_595.init = 16'h9898;
    PFUMX i27101 (.BLUT(n29524), .ALUT(n29525), .C0(index_i[0]), .Z(n29526));
    LUT4 mux_208_Mux_3_i491_3_lut_4_lut (.A(n29271), .B(index_i[1]), .C(index_i[3]), 
         .D(n32038), .Z(n491_adj_3626)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_3_i491_3_lut_4_lut.init = 16'h4f40;
    LUT4 mux_208_Mux_8_i172_3_lut_3_lut_rep_596 (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[2]), .Z(n29256)) /* synthesis lut_function=(!(A (B (C))+!A !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_8_i172_3_lut_3_lut_rep_596.init = 16'h7a7a;
    LUT4 mux_208_Mux_7_i347_3_lut_3_lut_3_lut_rep_597 (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[2]), .Z(n29257)) /* synthesis lut_function=(A ((C)+!B)+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_7_i347_3_lut_3_lut_3_lut_rep_597.init = 16'ha7a7;
    L6MUX21 i22166 (.D0(n860_adj_3517), .D1(n891_adj_3512), .SD(index_i[5]), 
            .Z(n24667));
    LUT4 mux_208_Mux_0_i985_3_lut_4_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[1]), .Z(n985)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_0_i985_3_lut_4_lut_4_lut_3_lut.init = 16'h1919;
    LUT4 mux_208_Mux_4_i142_3_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[3]), 
         .C(index_i[2]), .Z(n142_adj_3617)) /* synthesis lut_function=(A (B (C))+!A !(B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_4_i142_3_lut_4_lut_3_lut.init = 16'h9595;
    LUT4 mux_208_Mux_8_i93_3_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n93_adj_3647)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_8_i93_3_lut_3_lut_4_lut.init = 16'h0f85;
    LUT4 n53_bdd_3_lut_26927_3_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n27646)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C (D)))+!A (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n53_bdd_3_lut_26927_3_lut_4_lut.init = 16'h0fa7;
    LUT4 mux_208_Mux_4_i221_3_lut_3_lut (.A(index_i[0]), .B(index_i[4]), 
         .C(n205), .Z(n221_adj_3638)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_4_i221_3_lut_3_lut.init = 16'h7474;
    LUT4 mux_208_Mux_1_i890_4_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[3]), 
         .C(n29214), .D(index_i[4]), .Z(n890_adj_3524)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (D))+!A !((C+(D))+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_1_i890_4_lut_4_lut_4_lut_4_lut.init = 16'h55f3;
    LUT4 mux_208_Mux_3_i890_3_lut_4_lut (.A(n29223), .B(index_i[2]), .C(index_i[3]), 
         .D(n396), .Z(n890_adj_3510)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_3_i890_3_lut_4_lut.init = 16'h6f60;
    LUT4 i21066_3_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[0]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n23548)) /* synthesis lut_function=(A (B (C+(D))+!B !(D))+!A !(B (C+(D))+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21066_3_lut_4_lut_4_lut.init = 16'h99a7;
    LUT4 i13830_2_lut_3_lut_3_lut (.A(index_i[0]), .B(index_i[3]), .C(index_i[2]), 
         .Z(n16239)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i13830_2_lut_3_lut_3_lut.init = 16'h4040;
    LUT4 i21048_3_lut_4_lut_4_lut (.A(index_i[0]), .B(n29226), .C(index_i[3]), 
         .D(n29218), .Z(n23530)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21048_3_lut_4_lut_4_lut.init = 16'hc5c0;
    LUT4 mux_208_Mux_6_i332_3_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[1]), .Z(n332)) /* synthesis lut_function=(!(A (B)+!A !(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_6_i332_3_lut_4_lut_3_lut.init = 16'h6767;
    LUT4 n269_bdd_3_lut_24987_4_lut (.A(n29223), .B(index_i[2]), .C(index_i[3]), 
         .D(n32049), .Z(n26556)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n269_bdd_3_lut_24987_4_lut.init = 16'hf606;
    LUT4 i20959_3_lut_4_lut (.A(n29223), .B(index_i[2]), .C(index_i[3]), 
         .D(n32041), .Z(n23441)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20959_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_208_Mux_0_i762_3_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n762)) /* synthesis lut_function=(A (B+!(D))+!A !(B ((D)+!C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_0_i762_3_lut_4_lut_4_lut.init = 16'h98fa;
    LUT4 i13829_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(n29325), .C(index_i[4]), 
         .D(index_i[1]), .Z(n16238)) /* synthesis lut_function=(!(A (D)+!A !(B (C+!(D))+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i13829_3_lut_4_lut_4_lut_4_lut.init = 16'h40ff;
    LUT4 mux_208_Mux_5_i30_3_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n30)) /* synthesis lut_function=(A ((D)+!B)+!A !(B (D)+!B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_5_i30_3_lut_4_lut.init = 16'haa67;
    LUT4 mux_208_Mux_0_i348_3_lut_4_lut (.A(n29223), .B(index_i[2]), .C(index_i[3]), 
         .D(n32032), .Z(n348_adj_3620)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_0_i348_3_lut_4_lut.init = 16'h6f60;
    LUT4 i11185_3_lut_4_lut_4_lut (.A(index_i[0]), .B(n29229), .C(index_i[4]), 
         .D(index_i[3]), .Z(n605_adj_3629)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A !(B+(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11185_3_lut_4_lut_4_lut.init = 16'h555c;
    LUT4 i12936_3_lut_3_lut_3_lut (.A(index_i[0]), .B(index_i[2]), .C(index_i[1]), 
         .Z(n676)) /* synthesis lut_function=(!(A (C)+!A !(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12936_3_lut_3_lut_3_lut.init = 16'h4f4f;
    LUT4 i21030_3_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[0]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n23512)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21030_3_lut_4_lut_4_lut.init = 16'h5a58;
    LUT4 mux_208_Mux_4_i773_3_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[1]), .Z(n7)) /* synthesis lut_function=(!(A (B+(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_4_i773_3_lut_4_lut_3_lut.init = 16'h5656;
    LUT4 mux_208_Mux_5_i573_3_lut_3_lut (.A(index_i[0]), .B(index_i[4]), 
         .C(n572_adj_3607), .Z(n573_adj_3628)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_5_i573_3_lut_3_lut.init = 16'hd1d1;
    LUT4 mux_208_Mux_2_i507_3_lut_3_lut (.A(index_i[0]), .B(index_i[4]), 
         .C(n491_adj_3630), .Z(n507_adj_3666)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_2_i507_3_lut_3_lut.init = 16'h7474;
    L6MUX21 i25657 (.D0(n27406), .D1(n27404), .SD(index_i[5]), .Z(n27407));
    LUT4 n285_bdd_3_lut (.A(n32052), .B(n32043), .C(index_i[3]), .Z(n26558)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n285_bdd_3_lut.init = 16'hacac;
    LUT4 i11213_3_lut_4_lut_4_lut (.A(index_i[0]), .B(n7), .C(index_i[4]), 
         .D(n29218), .Z(n13509)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B ((D)+!C)+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11213_3_lut_4_lut_4_lut.init = 16'h5c0c;
    LUT4 mux_208_Mux_2_i859_3_lut_4_lut_4_lut (.A(index_i[0]), .B(n32052), 
         .C(index_i[3]), .D(n29218), .Z(n859_adj_3516)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B ((D)+!C)+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_2_i859_3_lut_4_lut_4_lut.init = 16'h5c0c;
    PFUMX i25655 (.BLUT(n27405), .ALUT(n285_adj_3664), .C0(index_i[4]), 
          .Z(n27406));
    LUT4 mux_208_Mux_2_i349_3_lut_3_lut (.A(index_i[0]), .B(index_i[4]), 
         .C(n348_adj_3669), .Z(n349_adj_3665)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_2_i349_3_lut_3_lut.init = 16'hd1d1;
    PFUMX i25653 (.BLUT(n78), .ALUT(n27403), .C0(index_i[4]), .Z(n27404));
    LUT4 mux_208_Mux_0_i684_3_lut_4_lut_4_lut (.A(index_i[0]), .B(n29255), 
         .C(index_i[3]), .D(n29218), .Z(n684_adj_3650)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B ((D)+!C)+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_0_i684_3_lut_4_lut_4_lut.init = 16'h5c0c;
    LUT4 mux_208_Mux_2_i763_4_lut_4_lut (.A(index_i[0]), .B(n13501), .C(index_i[4]), 
         .D(n157), .Z(n763_adj_3668)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_2_i763_4_lut_4_lut.init = 16'hdfd0;
    LUT4 mux_208_Mux_5_i564_3_lut_4_lut_3_lut_rep_752 (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[1]), .Z(n29412)) /* synthesis lut_function=(A (B (C))+!A !(B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_5_i564_3_lut_4_lut_3_lut_rep_752.init = 16'h9595;
    LUT4 mux_208_Mux_6_i156_3_lut_4_lut_4_lut_3_lut_rep_753 (.A(index_i[0]), 
         .B(index_i[2]), .C(index_i[1]), .Z(n29413)) /* synthesis lut_function=(!(A (B+(C))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_6_i156_3_lut_4_lut_4_lut_3_lut_rep_753.init = 16'h4646;
    PFUMX i22851 (.BLUT(n781_adj_3478), .ALUT(n796), .C0(index_i[4]), 
          .Z(n25352));
    LUT4 i21073_3_lut_4_lut (.A(index_i[0]), .B(index_i[2]), .C(index_i[1]), 
         .D(index_i[3]), .Z(n23555)) /* synthesis lut_function=(A (B+(D))+!A !(B (C+(D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21073_3_lut_4_lut.init = 16'haa9d;
    LUT4 mux_208_Mux_3_i444_3_lut_4_lut (.A(index_i[0]), .B(index_i[3]), 
         .C(n29349), .D(index_i[4]), .Z(n444_adj_3662)) /* synthesis lut_function=(!(A (B (D)+!B (C (D)))+!A !(B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_3_i444_3_lut_4_lut.init = 16'h46aa;
    LUT4 mux_208_Mux_4_i252_4_lut_4_lut (.A(index_i[0]), .B(index_i[3]), 
         .C(n29218), .D(index_i[4]), .Z(n252_adj_3639)) /* synthesis lut_function=(!(A (B (D)+!B !(D))+!A !(B ((D)+!C)+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_4_i252_4_lut_4_lut.init = 16'h669d;
    LUT4 mux_208_Mux_2_i348_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[1]), .D(index_i[3]), .Z(n348_adj_3669)) /* synthesis lut_function=(!(A (B (D)+!B (C+!(D)))+!A !(B (D)+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_2_i348_3_lut_4_lut_4_lut.init = 16'h4699;
    PFUMX i22852 (.BLUT(n812_adj_3624), .ALUT(n13515), .C0(index_i[4]), 
          .Z(n25353));
    LUT4 i20958_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[2]), .C(index_i[1]), 
         .D(index_i[3]), .Z(n23440)) /* synthesis lut_function=(!(A (B+!((D)+!C))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20958_3_lut_4_lut_4_lut.init = 16'h6646;
    LUT4 mux_208_Mux_4_i205_3_lut_4_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[1]), .D(index_i[3]), .Z(n205)) /* synthesis lut_function=(!(A (B (D)+!B (C (D)))+!A !(B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_4_i205_3_lut_4_lut.init = 16'h46aa;
    LUT4 mux_208_Mux_5_i572_3_lut_4_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[1]), .D(index_i[3]), .Z(n572_adj_3607)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A !(B (C+(D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_5_i572_3_lut_4_lut.init = 16'haa95;
    LUT4 mux_208_Mux_1_i93_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[1]), .D(index_i[3]), .Z(n93_adj_3667)) /* synthesis lut_function=(A (B (C (D))+!B !(D))+!A !(B (C (D))+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_1_i93_3_lut_4_lut_4_lut.init = 16'h9566;
    LUT4 mux_208_Mux_1_i62_3_lut_4_lut (.A(index_i[0]), .B(index_i[3]), 
         .C(index_i[2]), .D(index_i[4]), .Z(n62_adj_3661)) /* synthesis lut_function=(A (B (D)+!B ((D)+!C))+!A !(B (D)+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_1_i62_3_lut_4_lut.init = 16'haa56;
    PFUMX i22854 (.BLUT(n875_adj_3657), .ALUT(n890_adj_3480), .C0(index_i[4]), 
          .Z(n25355));
    LUT4 i24508_2_lut_rep_757 (.A(index_i[1]), .B(index_i[2]), .Z(n29417)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i24508_2_lut_rep_757.init = 16'h9999;
    LUT4 n442_bdd_2_lut_26997_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[3]), 
         .Z(n28936)) /* synthesis lut_function=(A (B+(C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n442_bdd_2_lut_26997_3_lut.init = 16'hf9f9;
    LUT4 mux_208_Mux_0_i93_3_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .Z(n93_adj_3567)) /* synthesis lut_function=(A (B)+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_0_i93_3_lut_3_lut.init = 16'h9c9c;
    LUT4 i8382_2_lut_rep_601 (.A(index_i[3]), .B(index_i[4]), .Z(n29261)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i8382_2_lut_rep_601.init = 16'heeee;
    LUT4 i1_3_lut_4_lut_adj_193 (.A(index_i[3]), .B(index_i[4]), .C(index_i[5]), 
         .D(n29349), .Z(n22204)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_3_lut_4_lut_adj_193.init = 16'hfffe;
    LUT4 mux_208_Mux_4_i262_3_lut_3_lut_rep_836 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n32037)) /* synthesis lut_function=(A (B+(C))+!A !(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_4_i262_3_lut_3_lut_rep_836.init = 16'ha9a9;
    LUT4 i14315_2_lut (.A(index_i[1]), .B(index_i[3]), .Z(n541)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i14315_2_lut.init = 16'h1111;
    LUT4 i21045_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n23527)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A !(B (D)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21045_3_lut_3_lut_4_lut.init = 16'ha955;
    LUT4 mux_208_Mux_0_i526_3_lut (.A(n29239), .B(n29229), .C(index_i[3]), 
         .Z(n526)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_0_i526_3_lut.init = 16'hcaca;
    PFUMX i22855 (.BLUT(n908), .ALUT(n923), .C0(index_i[4]), .Z(n25356));
    PFUMX i22856 (.BLUT(n939), .ALUT(n954_adj_3590), .C0(index_i[4]), 
          .Z(n25357));
    PFUMX i22857 (.BLUT(n971), .ALUT(n986), .C0(index_i[4]), .Z(n25358));
    PFUMX i22858 (.BLUT(n1002), .ALUT(n1017), .C0(index_i[4]), .Z(n25359));
    PFUMX i21083 (.BLUT(n23563), .ALUT(n23564), .C0(index_i[4]), .Z(n23565));
    LUT4 i24410_3_lut_rep_377_4_lut (.A(n29105), .B(index_i[5]), .C(index_i[8]), 
         .D(n1021), .Z(n29037)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i24410_3_lut_rep_377_4_lut.init = 16'hf808;
    LUT4 i24085_3_lut (.A(n286_adj_3504), .B(n317_adj_3555), .C(index_i[5]), 
         .Z(n25177)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24085_3_lut.init = 16'hcaca;
    LUT4 n23456_bdd_3_lut (.A(n32045), .B(n32044), .C(index_i[3]), .Z(n26561)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n23456_bdd_3_lut.init = 16'hcaca;
    LUT4 mux_208_Mux_1_i317_3_lut (.A(n301), .B(n908_adj_3578), .C(index_i[4]), 
         .Z(n317)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_208_Mux_1_i317_3_lut.init = 16'hcaca;
    PFUMX i17680 (.BLUT(n19992), .ALUT(n19993), .C0(index_i[4]), .Z(n19994));
    PFUMX i24965 (.BLUT(n26607), .ALUT(n26606), .C0(index_i[4]), .Z(n26608));
    PFUMX i21086 (.BLUT(n23566), .ALUT(n23567), .C0(index_i[4]), .Z(n23568));
    
endmodule
//
// Verilog Description of module \nco(OW=12) 
//

module \nco(OW=12)  (increment, GND_net, o_phase, dac_clk_p_c, i_sw0_c) /* synthesis syn_module_defined=1 */ ;
    input [30:0]increment;
    input GND_net;
    output [11:0]o_phase;
    input dac_clk_p_c;
    input i_sw0_c;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[29:38])
    
    wire n19891;
    wire [31:0]n233;
    wire [31:0]n133;
    
    wire n19892, n19890, n19889, n19888, n19887, n19886, n19885, 
        n19899, n19898, n19897, n19896, n19895, n19894, n19893;
    
    CCU2D phase_register_857_add_4_16 (.A0(increment[14]), .B0(n233[14]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[15]), .B1(n233[15]), 
          .C1(GND_net), .D1(GND_net), .CIN(n19891), .COUT(n19892), .S0(n133[14]), 
          .S1(n133[15]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_857_add_4_16.INIT0 = 16'h5666;
    defparam phase_register_857_add_4_16.INIT1 = 16'h5666;
    defparam phase_register_857_add_4_16.INJECT1_0 = "NO";
    defparam phase_register_857_add_4_16.INJECT1_1 = "NO";
    CCU2D phase_register_857_add_4_14 (.A0(increment[12]), .B0(n233[12]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[13]), .B1(n233[13]), 
          .C1(GND_net), .D1(GND_net), .CIN(n19890), .COUT(n19891), .S0(n133[12]), 
          .S1(n133[13]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_857_add_4_14.INIT0 = 16'h5666;
    defparam phase_register_857_add_4_14.INIT1 = 16'h5666;
    defparam phase_register_857_add_4_14.INJECT1_0 = "NO";
    defparam phase_register_857_add_4_14.INJECT1_1 = "NO";
    CCU2D phase_register_857_add_4_12 (.A0(increment[10]), .B0(n233[10]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[11]), .B1(n233[11]), 
          .C1(GND_net), .D1(GND_net), .CIN(n19889), .COUT(n19890), .S0(n133[10]), 
          .S1(n133[11]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_857_add_4_12.INIT0 = 16'h5666;
    defparam phase_register_857_add_4_12.INIT1 = 16'h5666;
    defparam phase_register_857_add_4_12.INJECT1_0 = "NO";
    defparam phase_register_857_add_4_12.INJECT1_1 = "NO";
    CCU2D phase_register_857_add_4_10 (.A0(increment[8]), .B0(n233[8]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[9]), .B1(n233[9]), 
          .C1(GND_net), .D1(GND_net), .CIN(n19888), .COUT(n19889), .S0(n133[8]), 
          .S1(n133[9]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_857_add_4_10.INIT0 = 16'h5666;
    defparam phase_register_857_add_4_10.INIT1 = 16'h5666;
    defparam phase_register_857_add_4_10.INJECT1_0 = "NO";
    defparam phase_register_857_add_4_10.INJECT1_1 = "NO";
    CCU2D phase_register_857_add_4_8 (.A0(increment[6]), .B0(n233[6]), .C0(GND_net), 
          .D0(GND_net), .A1(increment[7]), .B1(n233[7]), .C1(GND_net), 
          .D1(GND_net), .CIN(n19887), .COUT(n19888), .S0(n133[6]), .S1(n133[7]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_857_add_4_8.INIT0 = 16'h5666;
    defparam phase_register_857_add_4_8.INIT1 = 16'h5666;
    defparam phase_register_857_add_4_8.INJECT1_0 = "NO";
    defparam phase_register_857_add_4_8.INJECT1_1 = "NO";
    CCU2D phase_register_857_add_4_6 (.A0(increment[4]), .B0(n233[4]), .C0(GND_net), 
          .D0(GND_net), .A1(increment[5]), .B1(n233[5]), .C1(GND_net), 
          .D1(GND_net), .CIN(n19886), .COUT(n19887), .S0(n133[4]), .S1(n133[5]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_857_add_4_6.INIT0 = 16'h5666;
    defparam phase_register_857_add_4_6.INIT1 = 16'h5666;
    defparam phase_register_857_add_4_6.INJECT1_0 = "NO";
    defparam phase_register_857_add_4_6.INJECT1_1 = "NO";
    CCU2D phase_register_857_add_4_4 (.A0(increment[2]), .B0(n233[2]), .C0(GND_net), 
          .D0(GND_net), .A1(increment[3]), .B1(n233[3]), .C1(GND_net), 
          .D1(GND_net), .CIN(n19885), .COUT(n19886), .S0(n133[2]), .S1(n133[3]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_857_add_4_4.INIT0 = 16'h5666;
    defparam phase_register_857_add_4_4.INIT1 = 16'h5666;
    defparam phase_register_857_add_4_4.INJECT1_0 = "NO";
    defparam phase_register_857_add_4_4.INJECT1_1 = "NO";
    CCU2D phase_register_857_add_4_2 (.A0(increment[0]), .B0(n233[0]), .C0(GND_net), 
          .D0(GND_net), .A1(increment[1]), .B1(n233[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n19885), .S1(n133[1]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_857_add_4_2.INIT0 = 16'h7000;
    defparam phase_register_857_add_4_2.INIT1 = 16'h5666;
    defparam phase_register_857_add_4_2.INJECT1_0 = "NO";
    defparam phase_register_857_add_4_2.INJECT1_1 = "NO";
    FD1S3DX phase_register_857__i31 (.D(n133[31]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_phase[11])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_857__i31.GSR = "DISABLED";
    FD1S3DX phase_register_857__i30 (.D(n133[30]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_phase[10])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_857__i30.GSR = "DISABLED";
    FD1S3DX phase_register_857__i29 (.D(n133[29]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_phase[9])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_857__i29.GSR = "DISABLED";
    FD1S3DX phase_register_857__i28 (.D(n133[28]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_phase[8])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_857__i28.GSR = "DISABLED";
    FD1S3DX phase_register_857__i27 (.D(n133[27]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_phase[7])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_857__i27.GSR = "DISABLED";
    FD1S3DX phase_register_857__i26 (.D(n133[26]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_phase[6])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_857__i26.GSR = "DISABLED";
    FD1S3DX phase_register_857__i25 (.D(n133[25]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_phase[5])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_857__i25.GSR = "DISABLED";
    FD1S3DX phase_register_857__i24 (.D(n133[24]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_phase[4])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_857__i24.GSR = "DISABLED";
    FD1S3DX phase_register_857__i23 (.D(n133[23]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_phase[3])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_857__i23.GSR = "DISABLED";
    FD1S3DX phase_register_857__i22 (.D(n133[22]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_phase[2])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_857__i22.GSR = "DISABLED";
    FD1S3DX phase_register_857__i21 (.D(n133[21]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_phase[1])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_857__i21.GSR = "DISABLED";
    FD1S3DX phase_register_857__i20 (.D(n133[20]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_phase[0])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_857__i20.GSR = "DISABLED";
    FD1S3DX phase_register_857__i19 (.D(n133[19]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[19])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_857__i19.GSR = "DISABLED";
    FD1S3DX phase_register_857__i18 (.D(n133[18]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[18])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_857__i18.GSR = "DISABLED";
    FD1S3DX phase_register_857__i17 (.D(n133[17]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[17])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_857__i17.GSR = "DISABLED";
    FD1S3DX phase_register_857__i16 (.D(n133[16]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[16])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_857__i16.GSR = "DISABLED";
    FD1S3DX phase_register_857__i15 (.D(n133[15]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[15])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_857__i15.GSR = "DISABLED";
    FD1S3DX phase_register_857__i14 (.D(n133[14]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[14])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_857__i14.GSR = "DISABLED";
    FD1S3DX phase_register_857__i13 (.D(n133[13]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[13])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_857__i13.GSR = "DISABLED";
    FD1S3DX phase_register_857__i12 (.D(n133[12]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[12])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_857__i12.GSR = "DISABLED";
    FD1S3DX phase_register_857__i11 (.D(n133[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[11])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_857__i11.GSR = "DISABLED";
    FD1S3DX phase_register_857__i10 (.D(n133[10]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[10])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_857__i10.GSR = "DISABLED";
    FD1S3DX phase_register_857__i9 (.D(n133[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[9])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_857__i9.GSR = "DISABLED";
    FD1S3DX phase_register_857__i8 (.D(n133[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[8])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_857__i8.GSR = "DISABLED";
    FD1S3DX phase_register_857__i7 (.D(n133[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[7])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_857__i7.GSR = "DISABLED";
    FD1S3DX phase_register_857__i6 (.D(n133[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[6])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_857__i6.GSR = "DISABLED";
    FD1S3DX phase_register_857__i5 (.D(n133[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[5])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_857__i5.GSR = "DISABLED";
    FD1S3DX phase_register_857__i4 (.D(n133[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[4])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_857__i4.GSR = "DISABLED";
    FD1S3DX phase_register_857__i3 (.D(n133[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[3])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_857__i3.GSR = "DISABLED";
    FD1S3DX phase_register_857__i2 (.D(n133[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[2])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_857__i2.GSR = "DISABLED";
    FD1S3DX phase_register_857__i1 (.D(n133[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[1])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_857__i1.GSR = "DISABLED";
    LUT4 i17621_2_lut (.A(increment[0]), .B(n233[0]), .Z(n133[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i17621_2_lut.init = 16'h6666;
    CCU2D phase_register_857_add_4_32 (.A0(increment[30]), .B0(o_phase[10]), 
          .C0(GND_net), .D0(GND_net), .A1(o_phase[11]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n19899), .S0(n133[30]), .S1(n133[31]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_857_add_4_32.INIT0 = 16'h5666;
    defparam phase_register_857_add_4_32.INIT1 = 16'hfaaa;
    defparam phase_register_857_add_4_32.INJECT1_0 = "NO";
    defparam phase_register_857_add_4_32.INJECT1_1 = "NO";
    CCU2D phase_register_857_add_4_30 (.A0(increment[28]), .B0(o_phase[8]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[29]), .B1(o_phase[9]), 
          .C1(GND_net), .D1(GND_net), .CIN(n19898), .COUT(n19899), .S0(n133[28]), 
          .S1(n133[29]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_857_add_4_30.INIT0 = 16'h5666;
    defparam phase_register_857_add_4_30.INIT1 = 16'h5666;
    defparam phase_register_857_add_4_30.INJECT1_0 = "NO";
    defparam phase_register_857_add_4_30.INJECT1_1 = "NO";
    CCU2D phase_register_857_add_4_28 (.A0(increment[26]), .B0(o_phase[6]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[27]), .B1(o_phase[7]), 
          .C1(GND_net), .D1(GND_net), .CIN(n19897), .COUT(n19898), .S0(n133[26]), 
          .S1(n133[27]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_857_add_4_28.INIT0 = 16'h5666;
    defparam phase_register_857_add_4_28.INIT1 = 16'h5666;
    defparam phase_register_857_add_4_28.INJECT1_0 = "NO";
    defparam phase_register_857_add_4_28.INJECT1_1 = "NO";
    CCU2D phase_register_857_add_4_26 (.A0(increment[24]), .B0(o_phase[4]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[25]), .B1(o_phase[5]), 
          .C1(GND_net), .D1(GND_net), .CIN(n19896), .COUT(n19897), .S0(n133[24]), 
          .S1(n133[25]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_857_add_4_26.INIT0 = 16'h5666;
    defparam phase_register_857_add_4_26.INIT1 = 16'h5666;
    defparam phase_register_857_add_4_26.INJECT1_0 = "NO";
    defparam phase_register_857_add_4_26.INJECT1_1 = "NO";
    CCU2D phase_register_857_add_4_24 (.A0(increment[22]), .B0(o_phase[2]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[23]), .B1(o_phase[3]), 
          .C1(GND_net), .D1(GND_net), .CIN(n19895), .COUT(n19896), .S0(n133[22]), 
          .S1(n133[23]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_857_add_4_24.INIT0 = 16'h5666;
    defparam phase_register_857_add_4_24.INIT1 = 16'h5666;
    defparam phase_register_857_add_4_24.INJECT1_0 = "NO";
    defparam phase_register_857_add_4_24.INJECT1_1 = "NO";
    CCU2D phase_register_857_add_4_22 (.A0(increment[20]), .B0(o_phase[0]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[21]), .B1(o_phase[1]), 
          .C1(GND_net), .D1(GND_net), .CIN(n19894), .COUT(n19895), .S0(n133[20]), 
          .S1(n133[21]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_857_add_4_22.INIT0 = 16'h5666;
    defparam phase_register_857_add_4_22.INIT1 = 16'h5666;
    defparam phase_register_857_add_4_22.INJECT1_0 = "NO";
    defparam phase_register_857_add_4_22.INJECT1_1 = "NO";
    CCU2D phase_register_857_add_4_20 (.A0(increment[18]), .B0(n233[18]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[19]), .B1(n233[19]), 
          .C1(GND_net), .D1(GND_net), .CIN(n19893), .COUT(n19894), .S0(n133[18]), 
          .S1(n133[19]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_857_add_4_20.INIT0 = 16'h5666;
    defparam phase_register_857_add_4_20.INIT1 = 16'h5666;
    defparam phase_register_857_add_4_20.INJECT1_0 = "NO";
    defparam phase_register_857_add_4_20.INJECT1_1 = "NO";
    CCU2D phase_register_857_add_4_18 (.A0(increment[16]), .B0(n233[16]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[17]), .B1(n233[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n19892), .COUT(n19893), .S0(n133[16]), 
          .S1(n133[17]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_857_add_4_18.INIT0 = 16'h5666;
    defparam phase_register_857_add_4_18.INIT1 = 16'h5666;
    defparam phase_register_857_add_4_18.INJECT1_0 = "NO";
    defparam phase_register_857_add_4_18.INJECT1_1 = "NO";
    FD1S3DX phase_register_857__i0 (.D(n133[0]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[0])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_857__i0.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module sgnmpy_14x16_U25
//

module sgnmpy_14x16_U25 (dac_clk_p_c, i_sw0_c, \o_sample_dc_offset_i[7] , 
            u_s, \addr_space[3][13] , o_sample_i, GND_net, \u_s[12] , 
            \u_s[10] , \u_s[8] , \u_s[6] , \u_s[4] , \u_s[2] , \addr_space[3][12] , 
            \addr_space[3][10] , \addr_space[3][11] , \addr_space[3][8] , 
            \addr_space[3][9] , \addr_space[3][6] , \addr_space[3][7] , 
            \addr_space[3][4] , \addr_space[3][5] , \addr_space[3][2] , 
            \addr_space[3][3] , \addr_space[3][0] , \addr_space[3][1] , 
            \o_sample_dc_offset_i[15] , \o_sample_dc_offset_i[14] , \o_sample_dc_offset_i[13] , 
            \o_sample_dc_offset_i[12] , \o_sample_dc_offset_i[11] , \o_sample_dc_offset_i[10] , 
            \o_sample_dc_offset_i[9] , \o_sample_dc_offset_i[8] , n9490, 
            n9492, n9494, n9496, n9498, n9504, n9506) /* synthesis syn_module_defined=1 */ ;
    input dac_clk_p_c;
    input i_sw0_c;
    output \o_sample_dc_offset_i[7] ;
    output [13:0]u_s;
    input \addr_space[3][13] ;
    input [15:0]o_sample_i;
    input GND_net;
    output \u_s[12] ;
    output \u_s[10] ;
    output \u_s[8] ;
    output \u_s[6] ;
    output \u_s[4] ;
    output \u_s[2] ;
    input \addr_space[3][12] ;
    input \addr_space[3][10] ;
    input \addr_space[3][11] ;
    input \addr_space[3][8] ;
    input \addr_space[3][9] ;
    input \addr_space[3][6] ;
    input \addr_space[3][7] ;
    input \addr_space[3][4] ;
    input \addr_space[3][5] ;
    input \addr_space[3][2] ;
    input \addr_space[3][3] ;
    input \addr_space[3][0] ;
    input \addr_space[3][1] ;
    output \o_sample_dc_offset_i[15] ;
    output \o_sample_dc_offset_i[14] ;
    output \o_sample_dc_offset_i[13] ;
    output \o_sample_dc_offset_i[12] ;
    output \o_sample_dc_offset_i[11] ;
    output \o_sample_dc_offset_i[10] ;
    output \o_sample_dc_offset_i[9] ;
    output \o_sample_dc_offset_i[8] ;
    input n9490;
    input n9492;
    input n9494;
    input n9496;
    input n9498;
    input n9504;
    input n9506;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[29:38])
    wire [15:0]o_sample_i_c /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(30[39:49])
    wire [15:0]u_l;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(62[18:21])
    wire [15:0]u_l_15__N_1965;
    wire [4:0]u_sgn;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(63[19:24])
    wire [4:0]u_sgn_4__N_1981;
    wire [29:0]o_p_29__N_1986;
    wire [13:0]u_s_13__N_1951;
    wire [29:0]u_r;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(93[21:24])
    wire [29:0]n215;
    
    wire n14224, n19430, n19429, n19428, n19427, n19426, n19425, 
        n19424, n19423, n19422, n19421, n19420, n19419, n19418, 
        n19417;
    wire [13:0]u_s_c;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(61[18:21])
    
    wire n19586, n19585, n19584, n19583, n19582, n19581, n19580, 
        n19579, n19578, n19577, n19576, n19575, n19574, n19573, 
        n19572;
    
    FD1S3IX u_l__i0 (.D(u_l_15__N_1965[0]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_l[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=108, LSE_RLINE=108 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_l__i0.GSR = "DISABLED";
    FD1S3IX u_sgn__i0 (.D(u_sgn_4__N_1981[0]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_sgn[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=108, LSE_RLINE=108 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(87[9] 91[60])
    defparam u_sgn__i0.GSR = "DISABLED";
    FD1S3IX o_p__i1 (.D(o_p_29__N_1986[21]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_sample_dc_offset_i[7] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=108, LSE_RLINE=108 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(98[9] 102[36])
    defparam o_p__i1.GSR = "DISABLED";
    FD1S3IX u_s__i0 (.D(u_s_13__N_1951[0]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_s[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=108, LSE_RLINE=108 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_s__i0.GSR = "DISABLED";
    LUT4 i17_2_lut (.A(\addr_space[3][13] ), .B(o_sample_i[15]), .Z(u_sgn_4__N_1981[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(91[32:57])
    defparam i17_2_lut.init = 16'h6666;
    LUT4 mux_643_i1_3_lut (.A(u_r[21]), .B(n215[21]), .C(u_sgn[4]), .Z(o_p_29__N_1986[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[10:35])
    defparam mux_643_i1_3_lut.init = 16'hcaca;
    LUT4 i11848_1_lut (.A(u_l[0]), .Z(n14224)) /* synthesis lut_function=(!(A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam i11848_1_lut.init = 16'h5555;
    CCU2D add_536_29 (.A0(u_r[28]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(u_r[29]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19430), 
          .S0(n215[28]), .S1(n215[29]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[25:31])
    defparam add_536_29.INIT0 = 16'hf555;
    defparam add_536_29.INIT1 = 16'hf555;
    defparam add_536_29.INJECT1_0 = "NO";
    defparam add_536_29.INJECT1_1 = "NO";
    CCU2D add_536_27 (.A0(u_r[26]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(u_r[27]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19429), 
          .COUT(n19430), .S0(n215[26]), .S1(n215[27]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[25:31])
    defparam add_536_27.INIT0 = 16'hf555;
    defparam add_536_27.INIT1 = 16'hf555;
    defparam add_536_27.INJECT1_0 = "NO";
    defparam add_536_27.INJECT1_1 = "NO";
    CCU2D add_536_25 (.A0(u_r[24]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(u_r[25]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19428), 
          .COUT(n19429), .S0(n215[24]), .S1(n215[25]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[25:31])
    defparam add_536_25.INIT0 = 16'hf555;
    defparam add_536_25.INIT1 = 16'hf555;
    defparam add_536_25.INJECT1_0 = "NO";
    defparam add_536_25.INJECT1_1 = "NO";
    CCU2D add_536_23 (.A0(u_r[22]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(u_r[23]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19427), 
          .COUT(n19428), .S0(n215[22]), .S1(n215[23]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[25:31])
    defparam add_536_23.INIT0 = 16'hf555;
    defparam add_536_23.INIT1 = 16'hf555;
    defparam add_536_23.INJECT1_0 = "NO";
    defparam add_536_23.INJECT1_1 = "NO";
    CCU2D add_536_21 (.A0(u_r[20]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(u_r[21]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19426), 
          .COUT(n19427), .S1(n215[21]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[25:31])
    defparam add_536_21.INIT0 = 16'hf555;
    defparam add_536_21.INIT1 = 16'hf555;
    defparam add_536_21.INJECT1_0 = "NO";
    defparam add_536_21.INJECT1_1 = "NO";
    CCU2D add_536_19 (.A0(u_r[18]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(u_r[19]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19425), 
          .COUT(n19426));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[25:31])
    defparam add_536_19.INIT0 = 16'hf555;
    defparam add_536_19.INIT1 = 16'hf555;
    defparam add_536_19.INJECT1_0 = "NO";
    defparam add_536_19.INJECT1_1 = "NO";
    CCU2D add_536_17 (.A0(u_r[16]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(u_r[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19424), 
          .COUT(n19425));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[25:31])
    defparam add_536_17.INIT0 = 16'hf555;
    defparam add_536_17.INIT1 = 16'hf555;
    defparam add_536_17.INJECT1_0 = "NO";
    defparam add_536_17.INJECT1_1 = "NO";
    CCU2D add_536_15 (.A0(u_r[14]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(u_r[15]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19423), 
          .COUT(n19424));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[25:31])
    defparam add_536_15.INIT0 = 16'hf555;
    defparam add_536_15.INIT1 = 16'hf555;
    defparam add_536_15.INJECT1_0 = "NO";
    defparam add_536_15.INJECT1_1 = "NO";
    CCU2D add_536_13 (.A0(u_r[12]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(u_r[13]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19422), 
          .COUT(n19423));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[25:31])
    defparam add_536_13.INIT0 = 16'hf555;
    defparam add_536_13.INIT1 = 16'hf555;
    defparam add_536_13.INJECT1_0 = "NO";
    defparam add_536_13.INJECT1_1 = "NO";
    CCU2D add_536_11 (.A0(u_r[10]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(u_r[11]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19421), 
          .COUT(n19422));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[25:31])
    defparam add_536_11.INIT0 = 16'hf555;
    defparam add_536_11.INIT1 = 16'hf555;
    defparam add_536_11.INJECT1_0 = "NO";
    defparam add_536_11.INJECT1_1 = "NO";
    CCU2D add_536_9 (.A0(u_r[8]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(u_r[9]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19420), 
          .COUT(n19421));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[25:31])
    defparam add_536_9.INIT0 = 16'hf555;
    defparam add_536_9.INIT1 = 16'hf555;
    defparam add_536_9.INJECT1_0 = "NO";
    defparam add_536_9.INJECT1_1 = "NO";
    CCU2D add_536_7 (.A0(u_r[6]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(u_r[7]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19419), 
          .COUT(n19420));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[25:31])
    defparam add_536_7.INIT0 = 16'hf555;
    defparam add_536_7.INIT1 = 16'hf555;
    defparam add_536_7.INJECT1_0 = "NO";
    defparam add_536_7.INJECT1_1 = "NO";
    CCU2D add_536_5 (.A0(u_r[4]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(u_r[5]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19418), 
          .COUT(n19419));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[25:31])
    defparam add_536_5.INIT0 = 16'hf555;
    defparam add_536_5.INIT1 = 16'hf555;
    defparam add_536_5.INJECT1_0 = "NO";
    defparam add_536_5.INJECT1_1 = "NO";
    CCU2D add_536_3 (.A0(u_r[2]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(u_r[3]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19417), 
          .COUT(n19418));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[25:31])
    defparam add_536_3.INIT0 = 16'hf555;
    defparam add_536_3.INIT1 = 16'hf555;
    defparam add_536_3.INJECT1_0 = "NO";
    defparam add_536_3.INJECT1_1 = "NO";
    CCU2D add_536_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(u_r[0]), .B1(u_r[1]), .C1(GND_net), .D1(GND_net), .COUT(n19417));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[25:31])
    defparam add_536_1.INIT0 = 16'hF000;
    defparam add_536_1.INIT1 = 16'ha666;
    defparam add_536_1.INJECT1_0 = "NO";
    defparam add_536_1.INJECT1_1 = "NO";
    FD1S3IX u_s__i13 (.D(u_s_13__N_1951[13]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_s_c[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=108, LSE_RLINE=108 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_s__i13.GSR = "DISABLED";
    FD1S3IX u_s__i12 (.D(u_s_13__N_1951[12]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\u_s[12] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=108, LSE_RLINE=108 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_s__i12.GSR = "DISABLED";
    FD1S3IX u_s__i11 (.D(u_s_13__N_1951[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_s_c[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=108, LSE_RLINE=108 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_s__i11.GSR = "DISABLED";
    FD1S3IX u_s__i10 (.D(u_s_13__N_1951[10]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\u_s[10] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=108, LSE_RLINE=108 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_s__i10.GSR = "DISABLED";
    FD1S3IX u_s__i9 (.D(u_s_13__N_1951[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_s_c[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=108, LSE_RLINE=108 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_s__i9.GSR = "DISABLED";
    FD1S3IX u_s__i8 (.D(u_s_13__N_1951[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\u_s[8] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=108, LSE_RLINE=108 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_s__i8.GSR = "DISABLED";
    FD1S3IX u_s__i7 (.D(u_s_13__N_1951[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_s_c[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=108, LSE_RLINE=108 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_s__i7.GSR = "DISABLED";
    FD1S3IX u_s__i6 (.D(u_s_13__N_1951[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\u_s[6] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=108, LSE_RLINE=108 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_s__i6.GSR = "DISABLED";
    FD1S3IX u_s__i5 (.D(u_s_13__N_1951[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_s_c[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=108, LSE_RLINE=108 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_s__i5.GSR = "DISABLED";
    FD1S3IX u_s__i4 (.D(u_s_13__N_1951[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\u_s[4] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=108, LSE_RLINE=108 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_s__i4.GSR = "DISABLED";
    FD1S3IX u_s__i3 (.D(u_s_13__N_1951[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_s_c[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=108, LSE_RLINE=108 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_s__i3.GSR = "DISABLED";
    FD1S3IX u_s__i2 (.D(u_s_13__N_1951[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\u_s[2] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=108, LSE_RLINE=108 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_s__i2.GSR = "DISABLED";
    FD1S3IX u_s__i1 (.D(u_s_13__N_1951[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_s_c[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=108, LSE_RLINE=108 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_s__i1.GSR = "DISABLED";
    CCU2D unary_minus_8_add_3_17 (.A0(o_sample_i[14]), .B0(o_sample_i[15]), 
          .C0(GND_net), .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n19586), .S0(u_l_15__N_1965[15]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(83[22:28])
    defparam unary_minus_8_add_3_17.INIT0 = 16'hd111;
    defparam unary_minus_8_add_3_17.INIT1 = 16'h0000;
    defparam unary_minus_8_add_3_17.INJECT1_0 = "NO";
    defparam unary_minus_8_add_3_17.INJECT1_1 = "NO";
    CCU2D unary_minus_8_add_3_15 (.A0(o_sample_i[12]), .B0(o_sample_i[15]), 
          .C0(o_sample_i[13]), .D0(GND_net), .A1(o_sample_i[13]), .B1(o_sample_i[15]), 
          .C1(o_sample_i[14]), .D1(GND_net), .CIN(n19585), .COUT(n19586), 
          .S0(u_l_15__N_1965[13]), .S1(u_l_15__N_1965[14]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(83[22:28])
    defparam unary_minus_8_add_3_15.INIT0 = 16'hdd2d;
    defparam unary_minus_8_add_3_15.INIT1 = 16'hdd2d;
    defparam unary_minus_8_add_3_15.INJECT1_0 = "NO";
    defparam unary_minus_8_add_3_15.INJECT1_1 = "NO";
    CCU2D unary_minus_8_add_3_13 (.A0(o_sample_i[10]), .B0(o_sample_i[15]), 
          .C0(o_sample_i[11]), .D0(GND_net), .A1(o_sample_i[11]), .B1(o_sample_i[15]), 
          .C1(o_sample_i[12]), .D1(GND_net), .CIN(n19584), .COUT(n19585), 
          .S0(u_l_15__N_1965[11]), .S1(u_l_15__N_1965[12]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(83[22:28])
    defparam unary_minus_8_add_3_13.INIT0 = 16'hdd2d;
    defparam unary_minus_8_add_3_13.INIT1 = 16'hdd2d;
    defparam unary_minus_8_add_3_13.INJECT1_0 = "NO";
    defparam unary_minus_8_add_3_13.INJECT1_1 = "NO";
    CCU2D unary_minus_8_add_3_11 (.A0(o_sample_i[8]), .B0(o_sample_i[15]), 
          .C0(o_sample_i[9]), .D0(GND_net), .A1(o_sample_i[9]), .B1(o_sample_i[15]), 
          .C1(o_sample_i[10]), .D1(GND_net), .CIN(n19583), .COUT(n19584), 
          .S0(u_l_15__N_1965[9]), .S1(u_l_15__N_1965[10]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(83[22:28])
    defparam unary_minus_8_add_3_11.INIT0 = 16'hdd2d;
    defparam unary_minus_8_add_3_11.INIT1 = 16'hdd2d;
    defparam unary_minus_8_add_3_11.INJECT1_0 = "NO";
    defparam unary_minus_8_add_3_11.INJECT1_1 = "NO";
    CCU2D unary_minus_8_add_3_9 (.A0(o_sample_i[6]), .B0(o_sample_i[15]), 
          .C0(o_sample_i[7]), .D0(GND_net), .A1(o_sample_i[7]), .B1(o_sample_i[15]), 
          .C1(o_sample_i[8]), .D1(GND_net), .CIN(n19582), .COUT(n19583), 
          .S0(u_l_15__N_1965[7]), .S1(u_l_15__N_1965[8]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(83[22:28])
    defparam unary_minus_8_add_3_9.INIT0 = 16'hdd2d;
    defparam unary_minus_8_add_3_9.INIT1 = 16'hdd2d;
    defparam unary_minus_8_add_3_9.INJECT1_0 = "NO";
    defparam unary_minus_8_add_3_9.INJECT1_1 = "NO";
    CCU2D unary_minus_8_add_3_7 (.A0(o_sample_i[4]), .B0(o_sample_i[15]), 
          .C0(o_sample_i[5]), .D0(GND_net), .A1(o_sample_i[5]), .B1(o_sample_i[15]), 
          .C1(o_sample_i[6]), .D1(GND_net), .CIN(n19581), .COUT(n19582), 
          .S0(u_l_15__N_1965[5]), .S1(u_l_15__N_1965[6]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(83[22:28])
    defparam unary_minus_8_add_3_7.INIT0 = 16'hdd2d;
    defparam unary_minus_8_add_3_7.INIT1 = 16'hdd2d;
    defparam unary_minus_8_add_3_7.INJECT1_0 = "NO";
    defparam unary_minus_8_add_3_7.INJECT1_1 = "NO";
    CCU2D unary_minus_8_add_3_5 (.A0(o_sample_i[2]), .B0(o_sample_i[15]), 
          .C0(o_sample_i[3]), .D0(GND_net), .A1(o_sample_i[3]), .B1(o_sample_i[15]), 
          .C1(o_sample_i[4]), .D1(GND_net), .CIN(n19580), .COUT(n19581), 
          .S0(u_l_15__N_1965[3]), .S1(u_l_15__N_1965[4]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(83[22:28])
    defparam unary_minus_8_add_3_5.INIT0 = 16'hdd2d;
    defparam unary_minus_8_add_3_5.INIT1 = 16'hdd2d;
    defparam unary_minus_8_add_3_5.INJECT1_0 = "NO";
    defparam unary_minus_8_add_3_5.INJECT1_1 = "NO";
    CCU2D unary_minus_8_add_3_3 (.A0(o_sample_i[0]), .B0(o_sample_i[15]), 
          .C0(o_sample_i[1]), .D0(GND_net), .A1(o_sample_i[1]), .B1(o_sample_i[15]), 
          .C1(o_sample_i[2]), .D1(GND_net), .CIN(n19579), .COUT(n19580), 
          .S0(u_l_15__N_1965[1]), .S1(u_l_15__N_1965[2]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(83[22:28])
    defparam unary_minus_8_add_3_3.INIT0 = 16'hdd2d;
    defparam unary_minus_8_add_3_3.INIT1 = 16'hdd2d;
    defparam unary_minus_8_add_3_3.INJECT1_0 = "NO";
    defparam unary_minus_8_add_3_3.INJECT1_1 = "NO";
    CCU2D unary_minus_8_add_3_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(o_sample_i[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n19579), .S1(u_l_15__N_1965[0]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(83[22:28])
    defparam unary_minus_8_add_3_1.INIT0 = 16'hF000;
    defparam unary_minus_8_add_3_1.INIT1 = 16'h0aaa;
    defparam unary_minus_8_add_3_1.INJECT1_0 = "NO";
    defparam unary_minus_8_add_3_1.INJECT1_1 = "NO";
    CCU2D unary_minus_6_add_3_15 (.A0(\addr_space[3][12] ), .B0(\addr_space[3][13] ), 
          .C0(GND_net), .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n19578), .S0(u_s_13__N_1951[13]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(82[22:28])
    defparam unary_minus_6_add_3_15.INIT0 = 16'hd111;
    defparam unary_minus_6_add_3_15.INIT1 = 16'h0000;
    defparam unary_minus_6_add_3_15.INJECT1_0 = "NO";
    defparam unary_minus_6_add_3_15.INJECT1_1 = "NO";
    CCU2D unary_minus_6_add_3_13 (.A0(\addr_space[3][10] ), .B0(\addr_space[3][13] ), 
          .C0(\addr_space[3][11] ), .D0(GND_net), .A1(\addr_space[3][11] ), 
          .B1(\addr_space[3][13] ), .C1(\addr_space[3][12] ), .D1(GND_net), 
          .CIN(n19577), .COUT(n19578), .S0(u_s_13__N_1951[11]), .S1(u_s_13__N_1951[12]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(82[22:28])
    defparam unary_minus_6_add_3_13.INIT0 = 16'hdd2d;
    defparam unary_minus_6_add_3_13.INIT1 = 16'hdd2d;
    defparam unary_minus_6_add_3_13.INJECT1_0 = "NO";
    defparam unary_minus_6_add_3_13.INJECT1_1 = "NO";
    CCU2D unary_minus_6_add_3_11 (.A0(\addr_space[3][8] ), .B0(\addr_space[3][13] ), 
          .C0(\addr_space[3][9] ), .D0(GND_net), .A1(\addr_space[3][9] ), 
          .B1(\addr_space[3][13] ), .C1(\addr_space[3][10] ), .D1(GND_net), 
          .CIN(n19576), .COUT(n19577), .S0(u_s_13__N_1951[9]), .S1(u_s_13__N_1951[10]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(82[22:28])
    defparam unary_minus_6_add_3_11.INIT0 = 16'hdd2d;
    defparam unary_minus_6_add_3_11.INIT1 = 16'hdd2d;
    defparam unary_minus_6_add_3_11.INJECT1_0 = "NO";
    defparam unary_minus_6_add_3_11.INJECT1_1 = "NO";
    CCU2D unary_minus_6_add_3_9 (.A0(\addr_space[3][6] ), .B0(\addr_space[3][13] ), 
          .C0(\addr_space[3][7] ), .D0(GND_net), .A1(\addr_space[3][7] ), 
          .B1(\addr_space[3][13] ), .C1(\addr_space[3][8] ), .D1(GND_net), 
          .CIN(n19575), .COUT(n19576), .S0(u_s_13__N_1951[7]), .S1(u_s_13__N_1951[8]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(82[22:28])
    defparam unary_minus_6_add_3_9.INIT0 = 16'hdd2d;
    defparam unary_minus_6_add_3_9.INIT1 = 16'hdd2d;
    defparam unary_minus_6_add_3_9.INJECT1_0 = "NO";
    defparam unary_minus_6_add_3_9.INJECT1_1 = "NO";
    CCU2D unary_minus_6_add_3_7 (.A0(\addr_space[3][4] ), .B0(\addr_space[3][13] ), 
          .C0(\addr_space[3][5] ), .D0(GND_net), .A1(\addr_space[3][5] ), 
          .B1(\addr_space[3][13] ), .C1(\addr_space[3][6] ), .D1(GND_net), 
          .CIN(n19574), .COUT(n19575), .S0(u_s_13__N_1951[5]), .S1(u_s_13__N_1951[6]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(82[22:28])
    defparam unary_minus_6_add_3_7.INIT0 = 16'hdd2d;
    defparam unary_minus_6_add_3_7.INIT1 = 16'hdd2d;
    defparam unary_minus_6_add_3_7.INJECT1_0 = "NO";
    defparam unary_minus_6_add_3_7.INJECT1_1 = "NO";
    CCU2D unary_minus_6_add_3_5 (.A0(\addr_space[3][2] ), .B0(\addr_space[3][13] ), 
          .C0(\addr_space[3][3] ), .D0(GND_net), .A1(\addr_space[3][3] ), 
          .B1(\addr_space[3][13] ), .C1(\addr_space[3][4] ), .D1(GND_net), 
          .CIN(n19573), .COUT(n19574), .S0(u_s_13__N_1951[3]), .S1(u_s_13__N_1951[4]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(82[22:28])
    defparam unary_minus_6_add_3_5.INIT0 = 16'hdd2d;
    defparam unary_minus_6_add_3_5.INIT1 = 16'hdd2d;
    defparam unary_minus_6_add_3_5.INJECT1_0 = "NO";
    defparam unary_minus_6_add_3_5.INJECT1_1 = "NO";
    CCU2D unary_minus_6_add_3_3 (.A0(\addr_space[3][0] ), .B0(\addr_space[3][13] ), 
          .C0(\addr_space[3][1] ), .D0(GND_net), .A1(\addr_space[3][1] ), 
          .B1(\addr_space[3][13] ), .C1(\addr_space[3][2] ), .D1(GND_net), 
          .CIN(n19572), .COUT(n19573), .S0(u_s_13__N_1951[1]), .S1(u_s_13__N_1951[2]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(82[22:28])
    defparam unary_minus_6_add_3_3.INIT0 = 16'hdd2d;
    defparam unary_minus_6_add_3_3.INIT1 = 16'hdd2d;
    defparam unary_minus_6_add_3_3.INJECT1_0 = "NO";
    defparam unary_minus_6_add_3_3.INJECT1_1 = "NO";
    CCU2D unary_minus_6_add_3_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\addr_space[3][0] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n19572), .S1(u_s_13__N_1951[0]));   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(82[22:28])
    defparam unary_minus_6_add_3_1.INIT0 = 16'hF000;
    defparam unary_minus_6_add_3_1.INIT1 = 16'h0aaa;
    defparam unary_minus_6_add_3_1.INJECT1_0 = "NO";
    defparam unary_minus_6_add_3_1.INJECT1_1 = "NO";
    LUT4 mux_643_i9_3_lut (.A(u_r[29]), .B(n215[29]), .C(u_sgn[4]), .Z(o_p_29__N_1986[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[10:35])
    defparam mux_643_i9_3_lut.init = 16'hcaca;
    LUT4 mux_643_i8_3_lut (.A(u_r[28]), .B(n215[28]), .C(u_sgn[4]), .Z(o_p_29__N_1986[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[10:35])
    defparam mux_643_i8_3_lut.init = 16'hcaca;
    LUT4 mux_643_i7_3_lut (.A(u_r[27]), .B(n215[27]), .C(u_sgn[4]), .Z(o_p_29__N_1986[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[10:35])
    defparam mux_643_i7_3_lut.init = 16'hcaca;
    LUT4 mux_643_i6_3_lut (.A(u_r[26]), .B(n215[26]), .C(u_sgn[4]), .Z(o_p_29__N_1986[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[10:35])
    defparam mux_643_i6_3_lut.init = 16'hcaca;
    LUT4 mux_643_i5_3_lut (.A(u_r[25]), .B(n215[25]), .C(u_sgn[4]), .Z(o_p_29__N_1986[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[10:35])
    defparam mux_643_i5_3_lut.init = 16'hcaca;
    LUT4 mux_643_i4_3_lut (.A(u_r[24]), .B(n215[24]), .C(u_sgn[4]), .Z(o_p_29__N_1986[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[10:35])
    defparam mux_643_i4_3_lut.init = 16'hcaca;
    LUT4 mux_643_i3_3_lut (.A(u_r[23]), .B(n215[23]), .C(u_sgn[4]), .Z(o_p_29__N_1986[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[10:35])
    defparam mux_643_i3_3_lut.init = 16'hcaca;
    LUT4 mux_643_i2_3_lut (.A(u_r[22]), .B(n215[22]), .C(u_sgn[4]), .Z(o_p_29__N_1986[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(102[10:35])
    defparam mux_643_i2_3_lut.init = 16'hcaca;
    FD1S3IX o_p__i9 (.D(o_p_29__N_1986[29]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_sample_dc_offset_i[15] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=108, LSE_RLINE=108 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(98[9] 102[36])
    defparam o_p__i9.GSR = "DISABLED";
    FD1S3IX o_p__i8 (.D(o_p_29__N_1986[28]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_sample_dc_offset_i[14] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=108, LSE_RLINE=108 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(98[9] 102[36])
    defparam o_p__i8.GSR = "DISABLED";
    FD1S3IX o_p__i7 (.D(o_p_29__N_1986[27]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_sample_dc_offset_i[13] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=108, LSE_RLINE=108 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(98[9] 102[36])
    defparam o_p__i7.GSR = "DISABLED";
    FD1S3IX o_p__i6 (.D(o_p_29__N_1986[26]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_sample_dc_offset_i[12] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=108, LSE_RLINE=108 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(98[9] 102[36])
    defparam o_p__i6.GSR = "DISABLED";
    FD1S3IX o_p__i5 (.D(o_p_29__N_1986[25]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_sample_dc_offset_i[11] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=108, LSE_RLINE=108 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(98[9] 102[36])
    defparam o_p__i5.GSR = "DISABLED";
    FD1S3IX o_p__i4 (.D(o_p_29__N_1986[24]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_sample_dc_offset_i[10] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=108, LSE_RLINE=108 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(98[9] 102[36])
    defparam o_p__i4.GSR = "DISABLED";
    FD1S3IX o_p__i3 (.D(o_p_29__N_1986[23]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_sample_dc_offset_i[9] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=108, LSE_RLINE=108 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(98[9] 102[36])
    defparam o_p__i3.GSR = "DISABLED";
    FD1S3IX o_p__i2 (.D(o_p_29__N_1986[22]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_sample_dc_offset_i[8] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=108, LSE_RLINE=108 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(98[9] 102[36])
    defparam o_p__i2.GSR = "DISABLED";
    FD1S3IX u_sgn__i4 (.D(u_sgn[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(u_sgn[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=108, LSE_RLINE=108 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(87[9] 91[60])
    defparam u_sgn__i4.GSR = "DISABLED";
    FD1S3IX u_sgn__i3 (.D(u_sgn[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(u_sgn[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=108, LSE_RLINE=108 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(87[9] 91[60])
    defparam u_sgn__i3.GSR = "DISABLED";
    FD1S3IX u_sgn__i2 (.D(u_sgn[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(u_sgn[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=108, LSE_RLINE=108 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(87[9] 91[60])
    defparam u_sgn__i2.GSR = "DISABLED";
    FD1S3IX u_sgn__i1 (.D(u_sgn[0]), .CK(dac_clk_p_c), .CD(i_sw0_c), .Q(u_sgn[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=108, LSE_RLINE=108 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(87[9] 91[60])
    defparam u_sgn__i1.GSR = "DISABLED";
    FD1S3IX u_l__i15 (.D(u_l_15__N_1965[15]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_l[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=108, LSE_RLINE=108 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_l__i15.GSR = "DISABLED";
    FD1S3IX u_l__i14 (.D(u_l_15__N_1965[14]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_l[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=108, LSE_RLINE=108 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_l__i14.GSR = "DISABLED";
    FD1S3IX u_l__i13 (.D(u_l_15__N_1965[13]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_l[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=108, LSE_RLINE=108 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_l__i13.GSR = "DISABLED";
    FD1S3IX u_l__i12 (.D(u_l_15__N_1965[12]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_l[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=108, LSE_RLINE=108 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_l__i12.GSR = "DISABLED";
    FD1S3IX u_l__i11 (.D(u_l_15__N_1965[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_l[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=108, LSE_RLINE=108 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_l__i11.GSR = "DISABLED";
    FD1S3IX u_l__i10 (.D(u_l_15__N_1965[10]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_l[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=108, LSE_RLINE=108 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_l__i10.GSR = "DISABLED";
    FD1S3IX u_l__i9 (.D(u_l_15__N_1965[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_l[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=108, LSE_RLINE=108 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_l__i9.GSR = "DISABLED";
    FD1S3IX u_l__i8 (.D(u_l_15__N_1965[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_l[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=108, LSE_RLINE=108 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_l__i8.GSR = "DISABLED";
    FD1S3IX u_l__i7 (.D(u_l_15__N_1965[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_l[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=108, LSE_RLINE=108 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_l__i7.GSR = "DISABLED";
    FD1S3IX u_l__i6 (.D(u_l_15__N_1965[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_l[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=108, LSE_RLINE=108 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_l__i6.GSR = "DISABLED";
    FD1S3IX u_l__i5 (.D(u_l_15__N_1965[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_l[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=108, LSE_RLINE=108 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_l__i5.GSR = "DISABLED";
    FD1S3IX u_l__i4 (.D(u_l_15__N_1965[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_l[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=108, LSE_RLINE=108 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_l__i4.GSR = "DISABLED";
    FD1S3IX u_l__i3 (.D(u_l_15__N_1965[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_l[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=108, LSE_RLINE=108 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_l__i3.GSR = "DISABLED";
    FD1S3IX u_l__i2 (.D(u_l_15__N_1965[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_l[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=108, LSE_RLINE=108 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_l__i2.GSR = "DISABLED";
    FD1S3IX u_l__i1 (.D(u_l_15__N_1965[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_l[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=4, LSE_LCOL=14, LSE_RCOL=99, LSE_LLINE=108, LSE_RLINE=108 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(75[9] 84[5])
    defparam u_l__i1.GSR = "DISABLED";
    umpy_14x16_U21 umpy (.GND_net(GND_net), .dac_clk_p_c(dac_clk_p_c), .i_sw0_c(i_sw0_c), 
            .u_r({u_r}), .n14224(n14224), .n9490(n9490), .u_l({u_l}), 
            .u_s({u_s_c[13], \u_s[12] , u_s_c[11], \u_s[10] , u_s_c[9], 
            \u_s[8] , u_s_c[7], \u_s[6] , u_s_c[5], \u_s[4] , u_s_c[3], 
            \u_s[2] , u_s_c[1], u_s[0]}), .n9492(n9492), .n9494(n9494), 
            .n9496(n9496), .n9498(n9498), .n9504(n9504), .n9506(n9506)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/sgnmpy_14x16.v(95[13:68])
    
endmodule
//
// Verilog Description of module umpy_14x16_U21
//

module umpy_14x16_U21 (GND_net, dac_clk_p_c, i_sw0_c, u_r, n14224, 
            n9490, u_l, u_s, n9492, n9494, n9496, n9498, n9504, 
            n9506) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input dac_clk_p_c;
    input i_sw0_c;
    output [29:0]u_r;
    input n14224;
    input n9490;
    input [15:0]u_l;
    input [13:0]u_s;
    input n9492;
    input n9494;
    input n9496;
    input n9498;
    input n9504;
    input n9506;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[29:38])
    
    wire n19559;
    wire [17:0]S_0_00;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(71[14:20])
    wire [17:0]S_0_01;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(74[14:20])
    wire [20:0]S_1_00_20__N_2184;
    
    wire n19560, n19558, n19557, n19556, n19555, n19554, n19553;
    wire [20:0]S_1_00;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(103[17:23])
    wire [20:0]S_1_01;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(104[17:23])
    wire [17:0]S_0_02;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(77[14:20])
    wire [25:0]S_2_01_25__N_2294;
    wire [17:0]S_0_04;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(83[14:20])
    wire [20:0]S_1_03;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(106[17:23])
    wire [17:0]S_0_06;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(89[14:20])
    wire [29:0]o_p_29__N_2320;
    wire [25:0]S_2_01;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(140[17:23])
    
    wire n19340;
    wire [25:0]S_2_00_25__N_2268;
    
    wire n19682;
    wire [20:0]S_1_02_20__N_2226;
    
    wire n19681;
    wire [17:0]S_0_05;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(86[14:20])
    
    wire n19680, n19679, n19678, n19677, n19676, n19675, n19674, 
        n19374;
    wire [20:0]S_1_01_20__N_2205;
    
    wire n19373;
    wire [17:0]S_0_03;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(80[14:20])
    
    wire n19372, n19371, n19370, n19369, n19368, n19367, n19366, 
        n19339, n19338, n19337, n19336, n19331, n19332, n19333, 
        n19334, n19335, n19407;
    wire [20:0]S_1_02;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(105[17:23])
    
    wire n19406, n19405, n19404, n19403, n19597, n19596, n19595;
    wire [25:0]S_2_00;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(139[17:23])
    
    wire n19402, n19594, n19593, n19592, n19591, n19590, n19589, 
        n19588, n19401, n19400, n19561;
    
    CCU2D add_835_16 (.A0(S_0_00[16]), .B0(S_0_01[14]), .C0(GND_net), 
          .D0(GND_net), .A1(S_0_00[17]), .B1(S_0_01[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n19559), .COUT(n19560), .S0(S_1_00_20__N_2184[16]), 
          .S1(S_1_00_20__N_2184[17]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(122[13:48])
    defparam add_835_16.INIT0 = 16'h5666;
    defparam add_835_16.INIT1 = 16'h5666;
    defparam add_835_16.INJECT1_0 = "NO";
    defparam add_835_16.INJECT1_1 = "NO";
    CCU2D add_835_14 (.A0(S_0_00[14]), .B0(S_0_01[12]), .C0(GND_net), 
          .D0(GND_net), .A1(S_0_00[15]), .B1(S_0_01[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n19558), .COUT(n19559), .S0(S_1_00_20__N_2184[14]), 
          .S1(S_1_00_20__N_2184[15]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(122[13:48])
    defparam add_835_14.INIT0 = 16'h5666;
    defparam add_835_14.INIT1 = 16'h5666;
    defparam add_835_14.INJECT1_0 = "NO";
    defparam add_835_14.INJECT1_1 = "NO";
    CCU2D add_835_12 (.A0(S_0_00[12]), .B0(S_0_01[10]), .C0(GND_net), 
          .D0(GND_net), .A1(S_0_00[13]), .B1(S_0_01[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n19557), .COUT(n19558), .S0(S_1_00_20__N_2184[12]), 
          .S1(S_1_00_20__N_2184[13]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(122[13:48])
    defparam add_835_12.INIT0 = 16'h5666;
    defparam add_835_12.INIT1 = 16'h5666;
    defparam add_835_12.INJECT1_0 = "NO";
    defparam add_835_12.INJECT1_1 = "NO";
    CCU2D add_835_10 (.A0(S_0_00[10]), .B0(S_0_01[8]), .C0(GND_net), .D0(GND_net), 
          .A1(S_0_00[11]), .B1(S_0_01[9]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19556), .COUT(n19557), .S0(S_1_00_20__N_2184[10]), .S1(S_1_00_20__N_2184[11]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(122[13:48])
    defparam add_835_10.INIT0 = 16'h5666;
    defparam add_835_10.INIT1 = 16'h5666;
    defparam add_835_10.INJECT1_0 = "NO";
    defparam add_835_10.INJECT1_1 = "NO";
    CCU2D add_835_8 (.A0(S_0_00[8]), .B0(S_0_01[6]), .C0(GND_net), .D0(GND_net), 
          .A1(S_0_00[9]), .B1(S_0_01[7]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19555), .COUT(n19556), .S0(S_1_00_20__N_2184[8]), .S1(S_1_00_20__N_2184[9]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(122[13:48])
    defparam add_835_8.INIT0 = 16'h5666;
    defparam add_835_8.INIT1 = 16'h5666;
    defparam add_835_8.INJECT1_0 = "NO";
    defparam add_835_8.INJECT1_1 = "NO";
    CCU2D add_835_6 (.A0(S_0_00[6]), .B0(S_0_01[4]), .C0(GND_net), .D0(GND_net), 
          .A1(S_0_00[7]), .B1(S_0_01[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19554), .COUT(n19555), .S0(S_1_00_20__N_2184[6]), .S1(S_1_00_20__N_2184[7]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(122[13:48])
    defparam add_835_6.INIT0 = 16'h5666;
    defparam add_835_6.INIT1 = 16'h5666;
    defparam add_835_6.INJECT1_0 = "NO";
    defparam add_835_6.INJECT1_1 = "NO";
    CCU2D add_835_4 (.A0(S_0_00[4]), .B0(S_0_01[2]), .C0(GND_net), .D0(GND_net), 
          .A1(S_0_00[5]), .B1(S_0_01[3]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19553), .COUT(n19554), .S0(S_1_00_20__N_2184[4]), .S1(S_1_00_20__N_2184[5]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(122[13:48])
    defparam add_835_4.INIT0 = 16'h5666;
    defparam add_835_4.INIT1 = 16'h5666;
    defparam add_835_4.INJECT1_0 = "NO";
    defparam add_835_4.INJECT1_1 = "NO";
    FD1S3IX S_1_00__i0 (.D(S_0_00[0]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_00[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i0.GSR = "DISABLED";
    FD1S3IX S_1_01__i0 (.D(S_0_02[0]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i0.GSR = "DISABLED";
    FD1S3IX S_1_02__i1 (.D(S_0_04[0]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01_25__N_2294[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i1.GSR = "DISABLED";
    FD1S3IX S_1_03__i1 (.D(S_0_06[0]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_03[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_03__i1.GSR = "DISABLED";
    FD1S3IX S_2_00__i1 (.D(S_1_00[0]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_p_29__N_2320[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i1.GSR = "DISABLED";
    FD1S3IX S_2_01__i1 (.D(S_2_01_25__N_2294[0]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i1.GSR = "DISABLED";
    FD1S3IX S_3_00__i0 (.D(o_p_29__N_2320[0]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i0.GSR = "DISABLED";
    CCU2D add_835_2 (.A0(S_0_00[2]), .B0(S_0_01[0]), .C0(GND_net), .D0(GND_net), 
          .A1(S_0_00[3]), .B1(S_0_01[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n19553), .S1(S_1_00_20__N_2184[3]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(122[13:48])
    defparam add_835_2.INIT0 = 16'h7000;
    defparam add_835_2.INIT1 = 16'h5666;
    defparam add_835_2.INJECT1_0 = "NO";
    defparam add_835_2.INJECT1_1 = "NO";
    CCU2D add_815_22 (.A0(S_1_01[20]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19340), 
          .S0(S_2_00_25__N_2268[24]), .S1(S_2_00_25__N_2268[25]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(152[13:48])
    defparam add_815_22.INIT0 = 16'hfaaa;
    defparam add_815_22.INIT1 = 16'h0000;
    defparam add_815_22.INJECT1_0 = "NO";
    defparam add_815_22.INJECT1_1 = "NO";
    CCU2D add_837_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19682), 
          .S0(S_1_02_20__N_2226[20]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(124[13:48])
    defparam add_837_cout.INIT0 = 16'h0000;
    defparam add_837_cout.INIT1 = 16'h0000;
    defparam add_837_cout.INJECT1_0 = "NO";
    defparam add_837_cout.INJECT1_1 = "NO";
    CCU2D add_837_18 (.A0(S_0_05[16]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(S_0_05[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n19681), .COUT(n19682), .S0(S_1_02_20__N_2226[18]), .S1(S_1_02_20__N_2226[19]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(124[13:48])
    defparam add_837_18.INIT0 = 16'hfaaa;
    defparam add_837_18.INIT1 = 16'hfaaa;
    defparam add_837_18.INJECT1_0 = "NO";
    defparam add_837_18.INJECT1_1 = "NO";
    CCU2D add_837_16 (.A0(S_0_04[16]), .B0(S_0_05[14]), .C0(GND_net), 
          .D0(GND_net), .A1(S_0_04[17]), .B1(S_0_05[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n19680), .COUT(n19681), .S0(S_1_02_20__N_2226[16]), 
          .S1(S_1_02_20__N_2226[17]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(124[13:48])
    defparam add_837_16.INIT0 = 16'h5666;
    defparam add_837_16.INIT1 = 16'h5666;
    defparam add_837_16.INJECT1_0 = "NO";
    defparam add_837_16.INJECT1_1 = "NO";
    CCU2D add_837_14 (.A0(S_0_04[14]), .B0(S_0_05[12]), .C0(GND_net), 
          .D0(GND_net), .A1(S_0_04[15]), .B1(S_0_05[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n19679), .COUT(n19680), .S0(S_1_02_20__N_2226[14]), 
          .S1(S_1_02_20__N_2226[15]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(124[13:48])
    defparam add_837_14.INIT0 = 16'h5666;
    defparam add_837_14.INIT1 = 16'h5666;
    defparam add_837_14.INJECT1_0 = "NO";
    defparam add_837_14.INJECT1_1 = "NO";
    CCU2D add_837_12 (.A0(S_0_04[12]), .B0(S_0_05[10]), .C0(GND_net), 
          .D0(GND_net), .A1(S_0_04[13]), .B1(S_0_05[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n19678), .COUT(n19679), .S0(S_1_02_20__N_2226[12]), 
          .S1(S_1_02_20__N_2226[13]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(124[13:48])
    defparam add_837_12.INIT0 = 16'h5666;
    defparam add_837_12.INIT1 = 16'h5666;
    defparam add_837_12.INJECT1_0 = "NO";
    defparam add_837_12.INJECT1_1 = "NO";
    CCU2D add_837_10 (.A0(S_0_04[10]), .B0(S_0_05[8]), .C0(GND_net), .D0(GND_net), 
          .A1(S_0_04[11]), .B1(S_0_05[9]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19677), .COUT(n19678), .S0(S_1_02_20__N_2226[10]), .S1(S_1_02_20__N_2226[11]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(124[13:48])
    defparam add_837_10.INIT0 = 16'h5666;
    defparam add_837_10.INIT1 = 16'h5666;
    defparam add_837_10.INJECT1_0 = "NO";
    defparam add_837_10.INJECT1_1 = "NO";
    CCU2D add_837_8 (.A0(S_0_04[8]), .B0(S_0_05[6]), .C0(GND_net), .D0(GND_net), 
          .A1(S_0_04[9]), .B1(S_0_05[7]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19676), .COUT(n19677), .S0(S_1_02_20__N_2226[8]), .S1(S_1_02_20__N_2226[9]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(124[13:48])
    defparam add_837_8.INIT0 = 16'h5666;
    defparam add_837_8.INIT1 = 16'h5666;
    defparam add_837_8.INJECT1_0 = "NO";
    defparam add_837_8.INJECT1_1 = "NO";
    CCU2D add_837_6 (.A0(S_0_04[6]), .B0(S_0_05[4]), .C0(GND_net), .D0(GND_net), 
          .A1(S_0_04[7]), .B1(S_0_05[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19675), .COUT(n19676), .S0(S_1_02_20__N_2226[6]), .S1(S_1_02_20__N_2226[7]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(124[13:48])
    defparam add_837_6.INIT0 = 16'h5666;
    defparam add_837_6.INIT1 = 16'h5666;
    defparam add_837_6.INJECT1_0 = "NO";
    defparam add_837_6.INJECT1_1 = "NO";
    CCU2D add_837_4 (.A0(S_0_04[4]), .B0(S_0_05[2]), .C0(GND_net), .D0(GND_net), 
          .A1(S_0_04[5]), .B1(S_0_05[3]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19674), .COUT(n19675), .S0(S_1_02_20__N_2226[4]), .S1(S_1_02_20__N_2226[5]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(124[13:48])
    defparam add_837_4.INIT0 = 16'h5666;
    defparam add_837_4.INIT1 = 16'h5666;
    defparam add_837_4.INJECT1_0 = "NO";
    defparam add_837_4.INJECT1_1 = "NO";
    CCU2D add_837_2 (.A0(S_0_04[2]), .B0(S_0_05[0]), .C0(GND_net), .D0(GND_net), 
          .A1(S_0_04[3]), .B1(S_0_05[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n19674), .S1(S_1_02_20__N_2226[3]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(124[13:48])
    defparam add_837_2.INIT0 = 16'h7000;
    defparam add_837_2.INIT1 = 16'h5666;
    defparam add_837_2.INJECT1_0 = "NO";
    defparam add_837_2.INJECT1_1 = "NO";
    CCU2D add_814_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19374), 
          .S0(S_1_01_20__N_2205[20]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(123[13:48])
    defparam add_814_cout.INIT0 = 16'h0000;
    defparam add_814_cout.INIT1 = 16'h0000;
    defparam add_814_cout.INJECT1_0 = "NO";
    defparam add_814_cout.INJECT1_1 = "NO";
    CCU2D add_814_18 (.A0(S_0_03[16]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(S_0_03[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n19373), .COUT(n19374), .S0(S_1_01_20__N_2205[18]), .S1(S_1_01_20__N_2205[19]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(123[13:48])
    defparam add_814_18.INIT0 = 16'hfaaa;
    defparam add_814_18.INIT1 = 16'hfaaa;
    defparam add_814_18.INJECT1_0 = "NO";
    defparam add_814_18.INJECT1_1 = "NO";
    CCU2D add_814_16 (.A0(S_0_02[16]), .B0(S_0_03[14]), .C0(GND_net), 
          .D0(GND_net), .A1(S_0_02[17]), .B1(S_0_03[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n19372), .COUT(n19373), .S0(S_1_01_20__N_2205[16]), 
          .S1(S_1_01_20__N_2205[17]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(123[13:48])
    defparam add_814_16.INIT0 = 16'h5666;
    defparam add_814_16.INIT1 = 16'h5666;
    defparam add_814_16.INJECT1_0 = "NO";
    defparam add_814_16.INJECT1_1 = "NO";
    CCU2D add_814_14 (.A0(S_0_02[14]), .B0(S_0_03[12]), .C0(GND_net), 
          .D0(GND_net), .A1(S_0_02[15]), .B1(S_0_03[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n19371), .COUT(n19372), .S0(S_1_01_20__N_2205[14]), 
          .S1(S_1_01_20__N_2205[15]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(123[13:48])
    defparam add_814_14.INIT0 = 16'h5666;
    defparam add_814_14.INIT1 = 16'h5666;
    defparam add_814_14.INJECT1_0 = "NO";
    defparam add_814_14.INJECT1_1 = "NO";
    CCU2D add_814_12 (.A0(S_0_02[12]), .B0(S_0_03[10]), .C0(GND_net), 
          .D0(GND_net), .A1(S_0_02[13]), .B1(S_0_03[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n19370), .COUT(n19371), .S0(S_1_01_20__N_2205[12]), 
          .S1(S_1_01_20__N_2205[13]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(123[13:48])
    defparam add_814_12.INIT0 = 16'h5666;
    defparam add_814_12.INIT1 = 16'h5666;
    defparam add_814_12.INJECT1_0 = "NO";
    defparam add_814_12.INJECT1_1 = "NO";
    CCU2D add_814_10 (.A0(S_0_02[10]), .B0(S_0_03[8]), .C0(GND_net), .D0(GND_net), 
          .A1(S_0_02[11]), .B1(S_0_03[9]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19369), .COUT(n19370), .S0(S_1_01_20__N_2205[10]), .S1(S_1_01_20__N_2205[11]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(123[13:48])
    defparam add_814_10.INIT0 = 16'h5666;
    defparam add_814_10.INIT1 = 16'h5666;
    defparam add_814_10.INJECT1_0 = "NO";
    defparam add_814_10.INJECT1_1 = "NO";
    CCU2D add_814_8 (.A0(S_0_02[8]), .B0(S_0_03[6]), .C0(GND_net), .D0(GND_net), 
          .A1(S_0_02[9]), .B1(S_0_03[7]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19368), .COUT(n19369), .S0(S_1_01_20__N_2205[8]), .S1(S_1_01_20__N_2205[9]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(123[13:48])
    defparam add_814_8.INIT0 = 16'h5666;
    defparam add_814_8.INIT1 = 16'h5666;
    defparam add_814_8.INJECT1_0 = "NO";
    defparam add_814_8.INJECT1_1 = "NO";
    CCU2D add_814_6 (.A0(S_0_02[6]), .B0(S_0_03[4]), .C0(GND_net), .D0(GND_net), 
          .A1(S_0_02[7]), .B1(S_0_03[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19367), .COUT(n19368), .S0(S_1_01_20__N_2205[6]), .S1(S_1_01_20__N_2205[7]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(123[13:48])
    defparam add_814_6.INIT0 = 16'h5666;
    defparam add_814_6.INIT1 = 16'h5666;
    defparam add_814_6.INJECT1_0 = "NO";
    defparam add_814_6.INJECT1_1 = "NO";
    CCU2D add_814_4 (.A0(S_0_02[4]), .B0(S_0_03[2]), .C0(GND_net), .D0(GND_net), 
          .A1(S_0_02[5]), .B1(S_0_03[3]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19366), .COUT(n19367), .S0(S_1_01_20__N_2205[4]), .S1(S_1_01_20__N_2205[5]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(123[13:48])
    defparam add_814_4.INIT0 = 16'h5666;
    defparam add_814_4.INIT1 = 16'h5666;
    defparam add_814_4.INJECT1_0 = "NO";
    defparam add_814_4.INJECT1_1 = "NO";
    CCU2D add_814_2 (.A0(S_0_02[2]), .B0(S_0_03[0]), .C0(GND_net), .D0(GND_net), 
          .A1(S_0_02[3]), .B1(S_0_03[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n19366), .S1(S_1_01_20__N_2205[3]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(123[13:48])
    defparam add_814_2.INIT0 = 16'h7000;
    defparam add_814_2.INIT1 = 16'h5666;
    defparam add_814_2.INJECT1_0 = "NO";
    defparam add_814_2.INJECT1_1 = "NO";
    CCU2D add_815_20 (.A0(S_1_01[18]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(S_1_01[19]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n19339), .COUT(n19340), .S0(S_2_00_25__N_2268[22]), .S1(S_2_00_25__N_2268[23]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(152[13:48])
    defparam add_815_20.INIT0 = 16'hfaaa;
    defparam add_815_20.INIT1 = 16'hfaaa;
    defparam add_815_20.INJECT1_0 = "NO";
    defparam add_815_20.INJECT1_1 = "NO";
    CCU2D add_815_18 (.A0(S_1_00[20]), .B0(S_1_01[16]), .C0(GND_net), 
          .D0(GND_net), .A1(S_1_01[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n19338), .COUT(n19339), .S0(S_2_00_25__N_2268[20]), 
          .S1(S_2_00_25__N_2268[21]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(152[13:48])
    defparam add_815_18.INIT0 = 16'h5666;
    defparam add_815_18.INIT1 = 16'hfaaa;
    defparam add_815_18.INJECT1_0 = "NO";
    defparam add_815_18.INJECT1_1 = "NO";
    CCU2D add_815_16 (.A0(S_1_00[18]), .B0(S_1_01[14]), .C0(GND_net), 
          .D0(GND_net), .A1(S_1_00[19]), .B1(S_1_01[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n19337), .COUT(n19338), .S0(S_2_00_25__N_2268[18]), 
          .S1(S_2_00_25__N_2268[19]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(152[13:48])
    defparam add_815_16.INIT0 = 16'h5666;
    defparam add_815_16.INIT1 = 16'h5666;
    defparam add_815_16.INJECT1_0 = "NO";
    defparam add_815_16.INJECT1_1 = "NO";
    CCU2D add_815_14 (.A0(S_1_00[16]), .B0(S_1_01[12]), .C0(GND_net), 
          .D0(GND_net), .A1(S_1_00[17]), .B1(S_1_01[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n19336), .COUT(n19337), .S0(S_2_00_25__N_2268[16]), 
          .S1(S_2_00_25__N_2268[17]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(152[13:48])
    defparam add_815_14.INIT0 = 16'h5666;
    defparam add_815_14.INIT1 = 16'h5666;
    defparam add_815_14.INJECT1_0 = "NO";
    defparam add_815_14.INJECT1_1 = "NO";
    CCU2D add_815_4 (.A0(S_1_00[6]), .B0(S_1_01[2]), .C0(GND_net), .D0(GND_net), 
          .A1(S_1_00[7]), .B1(S_1_01[3]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19331), .COUT(n19332), .S0(S_2_00_25__N_2268[6]), .S1(S_2_00_25__N_2268[7]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(152[13:48])
    defparam add_815_4.INIT0 = 16'h5666;
    defparam add_815_4.INIT1 = 16'h5666;
    defparam add_815_4.INJECT1_0 = "NO";
    defparam add_815_4.INJECT1_1 = "NO";
    CCU2D add_815_8 (.A0(S_1_00[10]), .B0(S_1_01[6]), .C0(GND_net), .D0(GND_net), 
          .A1(S_1_00[11]), .B1(S_1_01[7]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19333), .COUT(n19334), .S0(S_2_00_25__N_2268[10]), .S1(S_2_00_25__N_2268[11]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(152[13:48])
    defparam add_815_8.INIT0 = 16'h5666;
    defparam add_815_8.INIT1 = 16'h5666;
    defparam add_815_8.INJECT1_0 = "NO";
    defparam add_815_8.INJECT1_1 = "NO";
    CCU2D add_815_2 (.A0(S_1_00[4]), .B0(S_1_01[0]), .C0(GND_net), .D0(GND_net), 
          .A1(S_1_00[5]), .B1(S_1_01[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n19331), .S1(S_2_00_25__N_2268[5]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(152[13:48])
    defparam add_815_2.INIT0 = 16'h7000;
    defparam add_815_2.INIT1 = 16'h5666;
    defparam add_815_2.INJECT1_0 = "NO";
    defparam add_815_2.INJECT1_1 = "NO";
    CCU2D add_815_12 (.A0(S_1_00[14]), .B0(S_1_01[10]), .C0(GND_net), 
          .D0(GND_net), .A1(S_1_00[15]), .B1(S_1_01[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n19335), .COUT(n19336), .S0(S_2_00_25__N_2268[14]), 
          .S1(S_2_00_25__N_2268[15]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(152[13:48])
    defparam add_815_12.INIT0 = 16'h5666;
    defparam add_815_12.INIT1 = 16'h5666;
    defparam add_815_12.INJECT1_0 = "NO";
    defparam add_815_12.INJECT1_1 = "NO";
    CCU2D add_410_18 (.A0(S_1_02[20]), .B0(S_1_03[16]), .C0(GND_net), 
          .D0(GND_net), .A1(S_1_03[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n19407), .S0(S_2_01_25__N_2294[20]), .S1(S_2_01_25__N_2294[21]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(153[13:48])
    defparam add_410_18.INIT0 = 16'h5666;
    defparam add_410_18.INIT1 = 16'hfaaa;
    defparam add_410_18.INJECT1_0 = "NO";
    defparam add_410_18.INJECT1_1 = "NO";
    CCU2D add_410_16 (.A0(S_1_02[18]), .B0(S_1_03[14]), .C0(GND_net), 
          .D0(GND_net), .A1(S_1_02[19]), .B1(S_1_03[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n19406), .COUT(n19407), .S0(S_2_01_25__N_2294[18]), 
          .S1(S_2_01_25__N_2294[19]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(153[13:48])
    defparam add_410_16.INIT0 = 16'h5666;
    defparam add_410_16.INIT1 = 16'h5666;
    defparam add_410_16.INJECT1_0 = "NO";
    defparam add_410_16.INJECT1_1 = "NO";
    CCU2D add_410_14 (.A0(S_1_02[16]), .B0(S_1_03[12]), .C0(GND_net), 
          .D0(GND_net), .A1(S_1_02[17]), .B1(S_1_03[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n19405), .COUT(n19406), .S0(S_2_01_25__N_2294[16]), 
          .S1(S_2_01_25__N_2294[17]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(153[13:48])
    defparam add_410_14.INIT0 = 16'h5666;
    defparam add_410_14.INIT1 = 16'h5666;
    defparam add_410_14.INJECT1_0 = "NO";
    defparam add_410_14.INJECT1_1 = "NO";
    CCU2D add_410_12 (.A0(S_1_02[14]), .B0(S_1_03[10]), .C0(GND_net), 
          .D0(GND_net), .A1(S_1_02[15]), .B1(S_1_03[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n19404), .COUT(n19405), .S0(S_2_01_25__N_2294[14]), 
          .S1(S_2_01_25__N_2294[15]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(153[13:48])
    defparam add_410_12.INIT0 = 16'h5666;
    defparam add_410_12.INIT1 = 16'h5666;
    defparam add_410_12.INJECT1_0 = "NO";
    defparam add_410_12.INJECT1_1 = "NO";
    CCU2D add_410_10 (.A0(S_1_02[12]), .B0(S_1_03[8]), .C0(GND_net), .D0(GND_net), 
          .A1(S_1_02[13]), .B1(S_1_03[9]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19403), .COUT(n19404), .S0(S_2_01_25__N_2294[12]), .S1(S_2_01_25__N_2294[13]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(153[13:48])
    defparam add_410_10.INIT0 = 16'h5666;
    defparam add_410_10.INIT1 = 16'h5666;
    defparam add_410_10.INJECT1_0 = "NO";
    defparam add_410_10.INJECT1_1 = "NO";
    CCU2D add_35_22 (.A0(S_2_01[20]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(S_2_01[21]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n19597), .S0(o_p_29__N_2320[28]), .S1(o_p_29__N_2320[29]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(177[13] 178[15])
    defparam add_35_22.INIT0 = 16'hfaaa;
    defparam add_35_22.INIT1 = 16'hfaaa;
    defparam add_35_22.INJECT1_0 = "NO";
    defparam add_35_22.INJECT1_1 = "NO";
    CCU2D add_35_20 (.A0(S_2_01[18]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(S_2_01[19]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n19596), .COUT(n19597), .S0(o_p_29__N_2320[26]), .S1(o_p_29__N_2320[27]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(177[13] 178[15])
    defparam add_35_20.INIT0 = 16'hfaaa;
    defparam add_35_20.INIT1 = 16'hfaaa;
    defparam add_35_20.INJECT1_0 = "NO";
    defparam add_35_20.INJECT1_1 = "NO";
    CCU2D add_815_6 (.A0(S_1_00[8]), .B0(S_1_01[4]), .C0(GND_net), .D0(GND_net), 
          .A1(S_1_00[9]), .B1(S_1_01[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19332), .COUT(n19333), .S0(S_2_00_25__N_2268[8]), .S1(S_2_00_25__N_2268[9]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(152[13:48])
    defparam add_815_6.INIT0 = 16'h5666;
    defparam add_815_6.INIT1 = 16'h5666;
    defparam add_815_6.INJECT1_0 = "NO";
    defparam add_815_6.INJECT1_1 = "NO";
    CCU2D add_35_18 (.A0(S_2_00[24]), .B0(S_2_01[16]), .C0(GND_net), .D0(GND_net), 
          .A1(S_2_00[25]), .B1(S_2_01[17]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19595), .COUT(n19596), .S0(o_p_29__N_2320[24]), .S1(o_p_29__N_2320[25]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(177[13] 178[15])
    defparam add_35_18.INIT0 = 16'h5666;
    defparam add_35_18.INIT1 = 16'h5666;
    defparam add_35_18.INJECT1_0 = "NO";
    defparam add_35_18.INJECT1_1 = "NO";
    CCU2D add_410_8 (.A0(S_1_02[10]), .B0(S_1_03[6]), .C0(GND_net), .D0(GND_net), 
          .A1(S_1_02[11]), .B1(S_1_03[7]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19402), .COUT(n19403), .S0(S_2_01_25__N_2294[10]), .S1(S_2_01_25__N_2294[11]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(153[13:48])
    defparam add_410_8.INIT0 = 16'h5666;
    defparam add_410_8.INIT1 = 16'h5666;
    defparam add_410_8.INJECT1_0 = "NO";
    defparam add_410_8.INJECT1_1 = "NO";
    CCU2D add_35_16 (.A0(S_2_00[22]), .B0(S_2_01[14]), .C0(GND_net), .D0(GND_net), 
          .A1(S_2_00[23]), .B1(S_2_01[15]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19594), .COUT(n19595), .S0(o_p_29__N_2320[22]), .S1(o_p_29__N_2320[23]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(177[13] 178[15])
    defparam add_35_16.INIT0 = 16'h5666;
    defparam add_35_16.INIT1 = 16'h5666;
    defparam add_35_16.INJECT1_0 = "NO";
    defparam add_35_16.INJECT1_1 = "NO";
    CCU2D add_35_14 (.A0(S_2_00[20]), .B0(S_2_01[12]), .C0(GND_net), .D0(GND_net), 
          .A1(S_2_00[21]), .B1(S_2_01[13]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19593), .COUT(n19594), .S0(o_p_29__N_2320[20]), .S1(o_p_29__N_2320[21]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(177[13] 178[15])
    defparam add_35_14.INIT0 = 16'h5666;
    defparam add_35_14.INIT1 = 16'h5666;
    defparam add_35_14.INJECT1_0 = "NO";
    defparam add_35_14.INJECT1_1 = "NO";
    CCU2D add_35_12 (.A0(S_2_00[18]), .B0(S_2_01[10]), .C0(GND_net), .D0(GND_net), 
          .A1(S_2_00[19]), .B1(S_2_01[11]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19592), .COUT(n19593), .S0(o_p_29__N_2320[18]), .S1(o_p_29__N_2320[19]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(177[13] 178[15])
    defparam add_35_12.INIT0 = 16'h5666;
    defparam add_35_12.INIT1 = 16'h5666;
    defparam add_35_12.INJECT1_0 = "NO";
    defparam add_35_12.INJECT1_1 = "NO";
    CCU2D add_35_10 (.A0(S_2_00[16]), .B0(S_2_01[8]), .C0(GND_net), .D0(GND_net), 
          .A1(S_2_00[17]), .B1(S_2_01[9]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19591), .COUT(n19592), .S0(o_p_29__N_2320[16]), .S1(o_p_29__N_2320[17]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(177[13] 178[15])
    defparam add_35_10.INIT0 = 16'h5666;
    defparam add_35_10.INIT1 = 16'h5666;
    defparam add_35_10.INJECT1_0 = "NO";
    defparam add_35_10.INJECT1_1 = "NO";
    CCU2D add_35_8 (.A0(S_2_00[14]), .B0(S_2_01[6]), .C0(GND_net), .D0(GND_net), 
          .A1(S_2_00[15]), .B1(S_2_01[7]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19590), .COUT(n19591), .S0(o_p_29__N_2320[14]), .S1(o_p_29__N_2320[15]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(177[13] 178[15])
    defparam add_35_8.INIT0 = 16'h5666;
    defparam add_35_8.INIT1 = 16'h5666;
    defparam add_35_8.INJECT1_0 = "NO";
    defparam add_35_8.INJECT1_1 = "NO";
    CCU2D add_35_6 (.A0(S_2_00[12]), .B0(S_2_01[4]), .C0(GND_net), .D0(GND_net), 
          .A1(S_2_00[13]), .B1(S_2_01[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19589), .COUT(n19590), .S0(o_p_29__N_2320[12]), .S1(o_p_29__N_2320[13]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(177[13] 178[15])
    defparam add_35_6.INIT0 = 16'h5666;
    defparam add_35_6.INIT1 = 16'h5666;
    defparam add_35_6.INJECT1_0 = "NO";
    defparam add_35_6.INJECT1_1 = "NO";
    CCU2D add_35_4 (.A0(S_2_00[10]), .B0(S_2_01[2]), .C0(GND_net), .D0(GND_net), 
          .A1(S_2_00[11]), .B1(S_2_01[3]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19588), .COUT(n19589), .S0(o_p_29__N_2320[10]), .S1(o_p_29__N_2320[11]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(177[13] 178[15])
    defparam add_35_4.INIT0 = 16'h5666;
    defparam add_35_4.INIT1 = 16'h5666;
    defparam add_35_4.INJECT1_0 = "NO";
    defparam add_35_4.INJECT1_1 = "NO";
    CCU2D add_410_6 (.A0(S_1_02[8]), .B0(S_1_03[4]), .C0(GND_net), .D0(GND_net), 
          .A1(S_1_02[9]), .B1(S_1_03[5]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19401), .COUT(n19402), .S0(S_2_01_25__N_2294[8]), .S1(S_2_01_25__N_2294[9]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(153[13:48])
    defparam add_410_6.INIT0 = 16'h5666;
    defparam add_410_6.INIT1 = 16'h5666;
    defparam add_410_6.INJECT1_0 = "NO";
    defparam add_410_6.INJECT1_1 = "NO";
    CCU2D add_35_2 (.A0(S_2_00[8]), .B0(S_2_01[0]), .C0(GND_net), .D0(GND_net), 
          .A1(S_2_00[9]), .B1(S_2_01[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n19588), .S1(o_p_29__N_2320[9]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(177[13] 178[15])
    defparam add_35_2.INIT0 = 16'h7000;
    defparam add_35_2.INIT1 = 16'h5666;
    defparam add_35_2.INJECT1_0 = "NO";
    defparam add_35_2.INJECT1_1 = "NO";
    CCU2D add_410_4 (.A0(S_1_02[6]), .B0(S_1_03[2]), .C0(GND_net), .D0(GND_net), 
          .A1(S_1_02[7]), .B1(S_1_03[3]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19400), .COUT(n19401), .S0(S_2_01_25__N_2294[6]), .S1(S_2_01_25__N_2294[7]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(153[13:48])
    defparam add_410_4.INIT0 = 16'h5666;
    defparam add_410_4.INIT1 = 16'h5666;
    defparam add_410_4.INJECT1_0 = "NO";
    defparam add_410_4.INJECT1_1 = "NO";
    CCU2D add_410_2 (.A0(S_1_02[4]), .B0(S_1_03[0]), .C0(GND_net), .D0(GND_net), 
          .A1(S_1_02[5]), .B1(S_1_03[1]), .C1(GND_net), .D1(GND_net), 
          .COUT(n19400), .S1(S_2_01_25__N_2294[5]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(153[13:48])
    defparam add_410_2.INIT0 = 16'h7000;
    defparam add_410_2.INIT1 = 16'h5666;
    defparam add_410_2.INJECT1_0 = "NO";
    defparam add_410_2.INJECT1_1 = "NO";
    LUT4 i17606_2_lut (.A(S_2_00[8]), .B(S_2_01[0]), .Z(o_p_29__N_2320[8])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i17606_2_lut.init = 16'h6666;
    LUT4 i17603_2_lut (.A(S_1_02[4]), .B(S_1_03[0]), .Z(S_2_01_25__N_2294[4])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i17603_2_lut.init = 16'h6666;
    LUT4 i17600_2_lut (.A(S_1_00[4]), .B(S_1_01[0]), .Z(S_2_00_25__N_2268[4])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i17600_2_lut.init = 16'h6666;
    LUT4 i17611_2_lut (.A(S_0_04[2]), .B(S_0_05[0]), .Z(S_1_02_20__N_2226[2])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i17611_2_lut.init = 16'h6666;
    CCU2D add_815_10 (.A0(S_1_00[12]), .B0(S_1_01[8]), .C0(GND_net), .D0(GND_net), 
          .A1(S_1_00[13]), .B1(S_1_01[9]), .C1(GND_net), .D1(GND_net), 
          .CIN(n19334), .COUT(n19335), .S0(S_2_00_25__N_2268[12]), .S1(S_2_00_25__N_2268[13]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(152[13:48])
    defparam add_815_10.INIT0 = 16'h5666;
    defparam add_815_10.INIT1 = 16'h5666;
    defparam add_815_10.INJECT1_0 = "NO";
    defparam add_815_10.INJECT1_1 = "NO";
    LUT4 i17601_2_lut (.A(S_0_02[2]), .B(S_0_03[0]), .Z(S_1_01_20__N_2205[2])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i17601_2_lut.init = 16'h6666;
    LUT4 i17604_2_lut (.A(S_0_00[2]), .B(S_0_01[0]), .Z(S_1_00_20__N_2184[2])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i17604_2_lut.init = 16'h6666;
    FD1S3IX S_3_00__i29 (.D(o_p_29__N_2320[29]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i29.GSR = "DISABLED";
    FD1S3IX S_3_00__i28 (.D(o_p_29__N_2320[28]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i28.GSR = "DISABLED";
    FD1S3IX S_3_00__i27 (.D(o_p_29__N_2320[27]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i27.GSR = "DISABLED";
    FD1S3IX S_3_00__i26 (.D(o_p_29__N_2320[26]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i26.GSR = "DISABLED";
    FD1S3IX S_3_00__i25 (.D(o_p_29__N_2320[25]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i25.GSR = "DISABLED";
    FD1S3IX S_3_00__i24 (.D(o_p_29__N_2320[24]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i24.GSR = "DISABLED";
    FD1S3IX S_3_00__i23 (.D(o_p_29__N_2320[23]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i23.GSR = "DISABLED";
    FD1S3IX S_3_00__i22 (.D(o_p_29__N_2320[22]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i22.GSR = "DISABLED";
    FD1S3IX S_3_00__i21 (.D(o_p_29__N_2320[21]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i21.GSR = "DISABLED";
    FD1S3IX S_3_00__i20 (.D(o_p_29__N_2320[20]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i20.GSR = "DISABLED";
    FD1S3IX S_3_00__i19 (.D(o_p_29__N_2320[19]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i19.GSR = "DISABLED";
    FD1S3IX S_3_00__i18 (.D(o_p_29__N_2320[18]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i18.GSR = "DISABLED";
    FD1S3IX S_3_00__i17 (.D(o_p_29__N_2320[17]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i17.GSR = "DISABLED";
    FD1S3IX S_3_00__i16 (.D(o_p_29__N_2320[16]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i16.GSR = "DISABLED";
    FD1S3IX S_3_00__i15 (.D(o_p_29__N_2320[15]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i15.GSR = "DISABLED";
    FD1S3IX S_3_00__i14 (.D(o_p_29__N_2320[14]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i14.GSR = "DISABLED";
    FD1S3IX S_3_00__i13 (.D(o_p_29__N_2320[13]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i13.GSR = "DISABLED";
    FD1S3IX S_3_00__i12 (.D(o_p_29__N_2320[12]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i12.GSR = "DISABLED";
    FD1S3IX S_3_00__i11 (.D(o_p_29__N_2320[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i11.GSR = "DISABLED";
    FD1S3IX S_3_00__i10 (.D(o_p_29__N_2320[10]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i10.GSR = "DISABLED";
    FD1S3IX S_3_00__i9 (.D(o_p_29__N_2320[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i9.GSR = "DISABLED";
    FD1S3IX S_3_00__i8 (.D(o_p_29__N_2320[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i8.GSR = "DISABLED";
    FD1S3IX S_3_00__i7 (.D(o_p_29__N_2320[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i7.GSR = "DISABLED";
    FD1S3IX S_3_00__i6 (.D(o_p_29__N_2320[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i6.GSR = "DISABLED";
    FD1S3IX S_3_00__i5 (.D(o_p_29__N_2320[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i5.GSR = "DISABLED";
    FD1S3IX S_3_00__i4 (.D(o_p_29__N_2320[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i4.GSR = "DISABLED";
    FD1S3IX S_3_00__i3 (.D(o_p_29__N_2320[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i3.GSR = "DISABLED";
    FD1S3IX S_3_00__i2 (.D(o_p_29__N_2320[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i2.GSR = "DISABLED";
    FD1S3IX S_3_00__i1 (.D(o_p_29__N_2320[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(u_r[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(171[9] 181[5])
    defparam S_3_00__i1.GSR = "DISABLED";
    FD1S3IX S_2_01__i22 (.D(S_2_01_25__N_2294[21]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i22.GSR = "DISABLED";
    FD1S3IX S_2_01__i21 (.D(S_2_01_25__N_2294[20]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i21.GSR = "DISABLED";
    FD1S3IX S_2_01__i20 (.D(S_2_01_25__N_2294[19]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i20.GSR = "DISABLED";
    FD1S3IX S_2_01__i19 (.D(S_2_01_25__N_2294[18]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i19.GSR = "DISABLED";
    FD1S3IX S_2_01__i18 (.D(S_2_01_25__N_2294[17]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i18.GSR = "DISABLED";
    FD1S3IX S_2_01__i17 (.D(S_2_01_25__N_2294[16]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i17.GSR = "DISABLED";
    FD1S3IX S_2_01__i16 (.D(S_2_01_25__N_2294[15]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i16.GSR = "DISABLED";
    FD1S3IX S_2_01__i15 (.D(S_2_01_25__N_2294[14]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i15.GSR = "DISABLED";
    FD1S3IX S_2_01__i14 (.D(S_2_01_25__N_2294[13]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i14.GSR = "DISABLED";
    FD1S3IX S_2_01__i13 (.D(S_2_01_25__N_2294[12]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i13.GSR = "DISABLED";
    FD1S3IX S_2_01__i12 (.D(S_2_01_25__N_2294[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i12.GSR = "DISABLED";
    FD1S3IX S_2_01__i11 (.D(S_2_01_25__N_2294[10]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i11.GSR = "DISABLED";
    FD1S3IX S_2_01__i10 (.D(S_2_01_25__N_2294[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i10.GSR = "DISABLED";
    FD1S3IX S_2_01__i9 (.D(S_2_01_25__N_2294[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i9.GSR = "DISABLED";
    FD1S3IX S_2_01__i8 (.D(S_2_01_25__N_2294[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i8.GSR = "DISABLED";
    FD1S3IX S_2_01__i7 (.D(S_2_01_25__N_2294[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i7.GSR = "DISABLED";
    FD1S3IX S_2_01__i6 (.D(S_2_01_25__N_2294[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i6.GSR = "DISABLED";
    FD1S3IX S_2_01__i5 (.D(S_2_01_25__N_2294[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i5.GSR = "DISABLED";
    FD1S3IX S_2_01__i4 (.D(S_2_01_25__N_2294[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i4.GSR = "DISABLED";
    FD1S3IX S_2_01__i3 (.D(S_2_01_25__N_2294[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i3.GSR = "DISABLED";
    FD1S3IX S_2_01__i2 (.D(S_2_01_25__N_2294[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_01__i2.GSR = "DISABLED";
    FD1S3IX S_2_00__i26 (.D(S_2_00_25__N_2268[25]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i26.GSR = "DISABLED";
    FD1S3IX S_2_00__i25 (.D(S_2_00_25__N_2268[24]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i25.GSR = "DISABLED";
    FD1S3IX S_2_00__i24 (.D(S_2_00_25__N_2268[23]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i24.GSR = "DISABLED";
    FD1S3IX S_2_00__i23 (.D(S_2_00_25__N_2268[22]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i23.GSR = "DISABLED";
    FD1S3IX S_2_00__i22 (.D(S_2_00_25__N_2268[21]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i22.GSR = "DISABLED";
    FD1S3IX S_2_00__i21 (.D(S_2_00_25__N_2268[20]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i21.GSR = "DISABLED";
    FD1S3IX S_2_00__i20 (.D(S_2_00_25__N_2268[19]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i20.GSR = "DISABLED";
    FD1S3IX S_2_00__i19 (.D(S_2_00_25__N_2268[18]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i19.GSR = "DISABLED";
    FD1S3IX S_2_00__i18 (.D(S_2_00_25__N_2268[17]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i18.GSR = "DISABLED";
    FD1S3IX S_2_00__i17 (.D(S_2_00_25__N_2268[16]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i17.GSR = "DISABLED";
    FD1S3IX S_2_00__i16 (.D(S_2_00_25__N_2268[15]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i16.GSR = "DISABLED";
    FD1S3IX S_2_00__i15 (.D(S_2_00_25__N_2268[14]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i15.GSR = "DISABLED";
    FD1S3IX S_2_00__i14 (.D(S_2_00_25__N_2268[13]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i14.GSR = "DISABLED";
    FD1S3IX S_2_00__i13 (.D(S_2_00_25__N_2268[12]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i13.GSR = "DISABLED";
    FD1S3IX S_2_00__i12 (.D(S_2_00_25__N_2268[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i12.GSR = "DISABLED";
    FD1S3IX S_2_00__i11 (.D(S_2_00_25__N_2268[10]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i11.GSR = "DISABLED";
    FD1S3IX S_2_00__i10 (.D(S_2_00_25__N_2268[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i10.GSR = "DISABLED";
    FD1S3IX S_2_00__i9 (.D(S_2_00_25__N_2268[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i9.GSR = "DISABLED";
    FD1S3IX S_2_00__i8 (.D(S_2_00_25__N_2268[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_p_29__N_2320[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i8.GSR = "DISABLED";
    FD1S3IX S_2_00__i7 (.D(S_2_00_25__N_2268[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_p_29__N_2320[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i7.GSR = "DISABLED";
    FD1S3IX S_2_00__i6 (.D(S_2_00_25__N_2268[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_p_29__N_2320[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i6.GSR = "DISABLED";
    FD1S3IX S_2_00__i5 (.D(S_2_00_25__N_2268[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_p_29__N_2320[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i5.GSR = "DISABLED";
    FD1S3IX S_2_00__i4 (.D(S_2_00_25__N_2268[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_p_29__N_2320[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i4.GSR = "DISABLED";
    FD1S3IX S_2_00__i3 (.D(S_2_00_25__N_2268[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_p_29__N_2320[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i3.GSR = "DISABLED";
    FD1S3IX S_2_00__i2 (.D(S_2_00_25__N_2268[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_p_29__N_2320[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(145[9] 154[5])
    defparam S_2_00__i2.GSR = "DISABLED";
    FD1S3IX S_1_03__i18 (.D(S_0_06[17]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_03[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_03__i18.GSR = "DISABLED";
    FD1S3IX S_1_03__i17 (.D(S_0_06[16]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_03[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_03__i17.GSR = "DISABLED";
    FD1S3IX S_1_03__i16 (.D(S_0_06[15]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_03[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_03__i16.GSR = "DISABLED";
    FD1S3IX S_1_03__i15 (.D(S_0_06[14]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_03[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_03__i15.GSR = "DISABLED";
    FD1S3IX S_1_03__i14 (.D(S_0_06[13]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_03[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_03__i14.GSR = "DISABLED";
    FD1S3IX S_1_03__i13 (.D(S_0_06[12]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_03[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_03__i13.GSR = "DISABLED";
    FD1S3IX S_1_03__i12 (.D(S_0_06[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_03[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_03__i12.GSR = "DISABLED";
    FD1S3IX S_1_03__i11 (.D(S_0_06[10]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_03[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_03__i11.GSR = "DISABLED";
    FD1S3IX S_1_03__i10 (.D(S_0_06[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_03[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_03__i10.GSR = "DISABLED";
    FD1S3IX S_1_03__i9 (.D(S_0_06[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_03[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_03__i9.GSR = "DISABLED";
    FD1S3IX S_1_03__i8 (.D(S_0_06[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_03[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_03__i8.GSR = "DISABLED";
    FD1S3IX S_1_03__i7 (.D(S_0_06[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_03[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_03__i7.GSR = "DISABLED";
    FD1S3IX S_1_03__i6 (.D(S_0_06[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_03[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_03__i6.GSR = "DISABLED";
    FD1S3IX S_1_03__i5 (.D(S_0_06[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_03[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_03__i5.GSR = "DISABLED";
    FD1S3IX S_1_03__i4 (.D(S_0_06[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_03[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_03__i4.GSR = "DISABLED";
    FD1S3IX S_1_03__i3 (.D(S_0_06[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_03[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_03__i3.GSR = "DISABLED";
    FD1S3IX S_1_03__i2 (.D(S_0_06[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_03[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_03__i2.GSR = "DISABLED";
    FD1S3IX S_1_02__i21 (.D(S_1_02_20__N_2226[20]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_02[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i21.GSR = "DISABLED";
    FD1S3IX S_1_02__i20 (.D(S_1_02_20__N_2226[19]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_02[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i20.GSR = "DISABLED";
    FD1S3IX S_1_02__i19 (.D(S_1_02_20__N_2226[18]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_02[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i19.GSR = "DISABLED";
    FD1S3IX S_1_02__i18 (.D(S_1_02_20__N_2226[17]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_02[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i18.GSR = "DISABLED";
    FD1S3IX S_1_02__i17 (.D(S_1_02_20__N_2226[16]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_02[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i17.GSR = "DISABLED";
    FD1S3IX S_1_02__i16 (.D(S_1_02_20__N_2226[15]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_02[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i16.GSR = "DISABLED";
    FD1S3IX S_1_02__i15 (.D(S_1_02_20__N_2226[14]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_02[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i15.GSR = "DISABLED";
    FD1S3IX S_1_02__i14 (.D(S_1_02_20__N_2226[13]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_02[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i14.GSR = "DISABLED";
    FD1S3IX S_1_02__i13 (.D(S_1_02_20__N_2226[12]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_02[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i13.GSR = "DISABLED";
    FD1S3IX S_1_02__i12 (.D(S_1_02_20__N_2226[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_02[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i12.GSR = "DISABLED";
    FD1S3IX S_1_02__i11 (.D(S_1_02_20__N_2226[10]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_02[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i11.GSR = "DISABLED";
    FD1S3IX S_1_02__i10 (.D(S_1_02_20__N_2226[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_02[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i10.GSR = "DISABLED";
    FD1S3IX S_1_02__i9 (.D(S_1_02_20__N_2226[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_02[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i9.GSR = "DISABLED";
    FD1S3IX S_1_02__i8 (.D(S_1_02_20__N_2226[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_02[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i8.GSR = "DISABLED";
    FD1S3IX S_1_02__i7 (.D(S_1_02_20__N_2226[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_02[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i7.GSR = "DISABLED";
    FD1S3IX S_1_02__i6 (.D(S_1_02_20__N_2226[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_02[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i6.GSR = "DISABLED";
    FD1S3IX S_1_02__i5 (.D(S_1_02_20__N_2226[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_02[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i5.GSR = "DISABLED";
    FD1S3IX S_1_02__i4 (.D(S_1_02_20__N_2226[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01_25__N_2294[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i4.GSR = "DISABLED";
    FD1S3IX S_1_02__i3 (.D(S_1_02_20__N_2226[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01_25__N_2294[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i3.GSR = "DISABLED";
    FD1S3IX S_1_02__i2 (.D(S_1_02_20__N_2226[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_01_25__N_2294[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_02__i2.GSR = "DISABLED";
    CCU2D add_835_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19561), 
          .S0(S_1_00_20__N_2184[20]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(122[13:48])
    defparam add_835_cout.INIT0 = 16'h0000;
    defparam add_835_cout.INIT1 = 16'h0000;
    defparam add_835_cout.INJECT1_0 = "NO";
    defparam add_835_cout.INJECT1_1 = "NO";
    CCU2D add_835_18 (.A0(S_0_01[16]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(S_0_01[17]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n19560), .COUT(n19561), .S0(S_1_00_20__N_2184[18]), .S1(S_1_00_20__N_2184[19]));   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(122[13:48])
    defparam add_835_18.INIT0 = 16'hfaaa;
    defparam add_835_18.INIT1 = 16'hfaaa;
    defparam add_835_18.INJECT1_0 = "NO";
    defparam add_835_18.INJECT1_1 = "NO";
    FD1S3IX S_1_01__i20 (.D(S_1_01_20__N_2205[20]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i20.GSR = "DISABLED";
    FD1S3IX S_1_01__i19 (.D(S_1_01_20__N_2205[19]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i19.GSR = "DISABLED";
    FD1S3IX S_1_01__i18 (.D(S_1_01_20__N_2205[18]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i18.GSR = "DISABLED";
    FD1S3IX S_1_01__i17 (.D(S_1_01_20__N_2205[17]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i17.GSR = "DISABLED";
    FD1S3IX S_1_01__i16 (.D(S_1_01_20__N_2205[16]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i16.GSR = "DISABLED";
    FD1S3IX S_1_01__i15 (.D(S_1_01_20__N_2205[15]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i15.GSR = "DISABLED";
    FD1S3IX S_1_01__i14 (.D(S_1_01_20__N_2205[14]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i14.GSR = "DISABLED";
    FD1S3IX S_1_01__i13 (.D(S_1_01_20__N_2205[13]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i13.GSR = "DISABLED";
    FD1S3IX S_1_01__i12 (.D(S_1_01_20__N_2205[12]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i12.GSR = "DISABLED";
    FD1S3IX S_1_01__i11 (.D(S_1_01_20__N_2205[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i11.GSR = "DISABLED";
    FD1S3IX S_1_01__i10 (.D(S_1_01_20__N_2205[10]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i10.GSR = "DISABLED";
    FD1S3IX S_1_01__i9 (.D(S_1_01_20__N_2205[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i9.GSR = "DISABLED";
    FD1S3IX S_1_01__i8 (.D(S_1_01_20__N_2205[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i8.GSR = "DISABLED";
    FD1S3IX S_1_01__i7 (.D(S_1_01_20__N_2205[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i7.GSR = "DISABLED";
    FD1S3IX S_1_01__i6 (.D(S_1_01_20__N_2205[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i6.GSR = "DISABLED";
    FD1S3IX S_1_01__i5 (.D(S_1_01_20__N_2205[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i5.GSR = "DISABLED";
    FD1S3IX S_1_01__i4 (.D(S_1_01_20__N_2205[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i4.GSR = "DISABLED";
    FD1S3IX S_1_01__i3 (.D(S_1_01_20__N_2205[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i3.GSR = "DISABLED";
    FD1S3IX S_1_01__i2 (.D(S_1_01_20__N_2205[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i2.GSR = "DISABLED";
    FD1S3IX S_1_01__i1 (.D(S_1_01_20__N_2205[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_01[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_01__i1.GSR = "DISABLED";
    FD1S3IX S_1_00__i20 (.D(S_1_00_20__N_2184[20]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_00[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i20.GSR = "DISABLED";
    FD1S3IX S_1_00__i19 (.D(S_1_00_20__N_2184[19]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_00[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i19.GSR = "DISABLED";
    FD1S3IX S_1_00__i18 (.D(S_1_00_20__N_2184[18]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_00[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i18.GSR = "DISABLED";
    FD1S3IX S_1_00__i17 (.D(S_1_00_20__N_2184[17]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_00[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i17.GSR = "DISABLED";
    FD1S3IX S_1_00__i16 (.D(S_1_00_20__N_2184[16]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_00[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i16.GSR = "DISABLED";
    FD1S3IX S_1_00__i15 (.D(S_1_00_20__N_2184[15]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_00[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i15.GSR = "DISABLED";
    FD1S3IX S_1_00__i14 (.D(S_1_00_20__N_2184[14]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_00[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i14.GSR = "DISABLED";
    FD1S3IX S_1_00__i13 (.D(S_1_00_20__N_2184[13]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_00[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i13.GSR = "DISABLED";
    FD1S3IX S_1_00__i12 (.D(S_1_00_20__N_2184[12]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_00[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i12.GSR = "DISABLED";
    FD1S3IX S_1_00__i11 (.D(S_1_00_20__N_2184[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_00[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i11.GSR = "DISABLED";
    FD1S3IX S_1_00__i10 (.D(S_1_00_20__N_2184[10]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_00[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i10.GSR = "DISABLED";
    FD1S3IX S_1_00__i9 (.D(S_1_00_20__N_2184[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_00[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i9.GSR = "DISABLED";
    FD1S3IX S_1_00__i8 (.D(S_1_00_20__N_2184[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_00[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i8.GSR = "DISABLED";
    FD1S3IX S_1_00__i7 (.D(S_1_00_20__N_2184[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_00[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i7.GSR = "DISABLED";
    FD1S3IX S_1_00__i6 (.D(S_1_00_20__N_2184[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_00[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i6.GSR = "DISABLED";
    FD1S3IX S_1_00__i5 (.D(S_1_00_20__N_2184[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_00[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i5.GSR = "DISABLED";
    FD1S3IX S_1_00__i4 (.D(S_1_00_20__N_2184[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_1_00[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i4.GSR = "DISABLED";
    FD1S3IX S_1_00__i3 (.D(S_1_00_20__N_2184[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00_25__N_2268[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i3.GSR = "DISABLED";
    FD1S3IX S_1_00__i2 (.D(S_1_00_20__N_2184[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00_25__N_2268[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i2.GSR = "DISABLED";
    FD1S3IX S_1_00__i1 (.D(S_1_00_20__N_2184[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_2_00_25__N_2268[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=28, LSE_LCOL=13, LSE_RCOL=68, LSE_LLINE=95, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(113[9] 126[5])
    defparam S_1_00__i1.GSR = "DISABLED";
    \bimpy(BW=16)_U13  initialmpy_6_0 (.S_0_06({S_0_06}), .dac_clk_p_c(dac_clk_p_c), 
            .n14224(n14224), .n9490(n9490), .GND_net(GND_net), .u_l({u_l}), 
            .\u_s[13] (u_s[13]), .\u_s[12] (u_s[12]), .i_sw0_c(i_sw0_c)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(90[14:75])
    \bimpy(BW=16)_U14  initialmpy_5_0 (.S_0_05({S_0_05}), .dac_clk_p_c(dac_clk_p_c), 
            .n14224(n14224), .n9492(n9492), .GND_net(GND_net), .u_l({u_l}), 
            .\u_s[11] (u_s[11]), .\u_s[10] (u_s[10]), .i_sw0_c(i_sw0_c)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(87[14:75])
    \bimpy(BW=16)_U15  initialmpy_4_0 (.\S_0_04[0] (S_0_04[0]), .dac_clk_p_c(dac_clk_p_c), 
            .n14224(n14224), .n9494(n9494), .GND_net(GND_net), .u_l({u_l}), 
            .\u_s[9] (u_s[9]), .\u_s[8] (u_s[8]), .\S_0_04[17] (S_0_04[17]), 
            .i_sw0_c(i_sw0_c), .\S_0_04[16] (S_0_04[16]), .\S_0_04[15] (S_0_04[15]), 
            .\S_0_04[14] (S_0_04[14]), .\S_0_04[13] (S_0_04[13]), .\S_0_04[12] (S_0_04[12]), 
            .\S_0_04[11] (S_0_04[11]), .\S_0_04[10] (S_0_04[10]), .\S_0_04[9] (S_0_04[9]), 
            .\S_0_04[8] (S_0_04[8]), .\S_0_04[7] (S_0_04[7]), .\S_0_04[6] (S_0_04[6]), 
            .\S_0_04[5] (S_0_04[5]), .\S_0_04[4] (S_0_04[4]), .\S_0_04[3] (S_0_04[3]), 
            .\S_0_04[2] (S_0_04[2]), .\S_1_02_20__N_2226[1] (S_1_02_20__N_2226[1])) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(84[14:73])
    \bimpy(BW=16)_U16  initialmpy_3_0 (.S_0_03({S_0_03}), .dac_clk_p_c(dac_clk_p_c), 
            .n14224(n14224), .n9496(n9496), .u_l({u_l}), .\u_s[6] (u_s[6]), 
            .\u_s[7] (u_s[7]), .i_sw0_c(i_sw0_c), .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(81[14:73])
    \bimpy(BW=16)_U17  initialmpy_2_0 (.\S_0_02[0] (S_0_02[0]), .dac_clk_p_c(dac_clk_p_c), 
            .n14224(n14224), .n9498(n9498), .GND_net(GND_net), .u_l({u_l}), 
            .\u_s[5] (u_s[5]), .\u_s[4] (u_s[4]), .\S_0_02[17] (S_0_02[17]), 
            .i_sw0_c(i_sw0_c), .\S_0_02[16] (S_0_02[16]), .\S_0_02[15] (S_0_02[15]), 
            .\S_0_02[14] (S_0_02[14]), .\S_0_02[13] (S_0_02[13]), .\S_0_02[12] (S_0_02[12]), 
            .\S_0_02[11] (S_0_02[11]), .\S_0_02[10] (S_0_02[10]), .\S_0_02[9] (S_0_02[9]), 
            .\S_0_02[8] (S_0_02[8]), .\S_0_02[7] (S_0_02[7]), .\S_0_02[6] (S_0_02[6]), 
            .\S_0_02[5] (S_0_02[5]), .\S_0_02[4] (S_0_02[4]), .\S_0_02[3] (S_0_02[3]), 
            .\S_0_02[2] (S_0_02[2]), .\S_1_01_20__N_2205[1] (S_1_01_20__N_2205[1])) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(78[14:73])
    \bimpy(BW=16)_U18  initialmpy_1_0 (.S_0_01({S_0_01}), .dac_clk_p_c(dac_clk_p_c), 
            .n14224(n14224), .n9504(n9504), .GND_net(GND_net), .u_l({u_l}), 
            .\u_s[3] (u_s[3]), .\u_s[2] (u_s[2]), .i_sw0_c(i_sw0_c)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(75[14:73])
    \bimpy(BW=16)_U19  initialmpy_0_0 (.u_l({u_l}), .\u_s[1] (u_s[1]), .\u_s[0] (u_s[0]), 
            .\S_0_00[0] (S_0_00[0]), .dac_clk_p_c(dac_clk_p_c), .n14224(n14224), 
            .n9506(n9506), .GND_net(GND_net), .\S_0_00[17] (S_0_00[17]), 
            .i_sw0_c(i_sw0_c), .\S_0_00[16] (S_0_00[16]), .\S_0_00[15] (S_0_00[15]), 
            .\S_0_00[14] (S_0_00[14]), .\S_0_00[13] (S_0_00[13]), .\S_0_00[12] (S_0_00[12]), 
            .\S_0_00[11] (S_0_00[11]), .\S_0_00[10] (S_0_00[10]), .\S_0_00[9] (S_0_00[9]), 
            .\S_0_00[8] (S_0_00[8]), .\S_0_00[7] (S_0_00[7]), .\S_0_00[6] (S_0_00[6]), 
            .\S_0_00[5] (S_0_00[5]), .\S_0_00[4] (S_0_00[4]), .\S_0_00[3] (S_0_00[3]), 
            .\S_0_00[2] (S_0_00[2]), .\S_1_00_20__N_2184[1] (S_1_00_20__N_2184[1])) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/umpy_14x16.v(72[14:73])
    
endmodule
//
// Verilog Description of module \bimpy(BW=16)_U13 
//

module \bimpy(BW=16)_U13  (S_0_06, dac_clk_p_c, n14224, n9490, GND_net, 
            u_l, \u_s[13] , \u_s[12] , i_sw0_c) /* synthesis syn_module_defined=1 */ ;
    output [17:0]S_0_06;
    input dac_clk_p_c;
    input n14224;
    input n9490;
    input GND_net;
    input [15:0]u_l;
    input \u_s[13] ;
    input \u_s[12] ;
    input i_sw0_c;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[29:38])
    
    wire n19535;
    wire [17:0]o_r_17__N_2438;
    
    wire n19534;
    wire [14:0]c_15__N_2408;
    wire [14:0]c_15__N_2423;
    
    wire n19533, n19532, n19531, n19530, n19529, n19528, n29297, 
        n29296;
    
    FD1S3IX o_r__i0 (.D(n9490), .CK(dac_clk_p_c), .CD(n14224), .Q(S_0_06[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=90, LSE_RLINE=90 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i0.GSR = "DISABLED";
    CCU2D add_832_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19535), 
          .S0(o_r_17__N_2438[17]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_832_cout.INIT0 = 16'h0000;
    defparam add_832_cout.INIT1 = 16'h0000;
    defparam add_832_cout.INJECT1_0 = "NO";
    defparam add_832_cout.INJECT1_1 = "NO";
    CCU2D add_832_15 (.A0(c_15__N_2408[14]), .B0(c_15__N_2423[14]), .C0(c_15__N_2408[13]), 
          .D0(c_15__N_2423[13]), .A1(u_l[15]), .B1(\u_s[13] ), .C1(c_15__N_2408[14]), 
          .D1(c_15__N_2423[14]), .CIN(n19534), .COUT(n19535), .S0(o_r_17__N_2438[15]), 
          .S1(o_r_17__N_2438[16]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_832_15.INIT0 = 16'h9666;
    defparam add_832_15.INIT1 = 16'h7888;
    defparam add_832_15.INJECT1_0 = "NO";
    defparam add_832_15.INJECT1_1 = "NO";
    CCU2D add_832_13 (.A0(c_15__N_2408[12]), .B0(c_15__N_2423[12]), .C0(c_15__N_2408[11]), 
          .D0(c_15__N_2423[11]), .A1(c_15__N_2408[13]), .B1(c_15__N_2423[13]), 
          .C1(c_15__N_2408[12]), .D1(c_15__N_2423[12]), .CIN(n19533), 
          .COUT(n19534), .S0(o_r_17__N_2438[13]), .S1(o_r_17__N_2438[14]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_832_13.INIT0 = 16'h9666;
    defparam add_832_13.INIT1 = 16'h9666;
    defparam add_832_13.INJECT1_0 = "NO";
    defparam add_832_13.INJECT1_1 = "NO";
    CCU2D add_832_11 (.A0(c_15__N_2408[10]), .B0(c_15__N_2423[10]), .C0(c_15__N_2408[9]), 
          .D0(c_15__N_2423[9]), .A1(c_15__N_2408[11]), .B1(c_15__N_2423[11]), 
          .C1(c_15__N_2408[10]), .D1(c_15__N_2423[10]), .CIN(n19532), 
          .COUT(n19533), .S0(o_r_17__N_2438[11]), .S1(o_r_17__N_2438[12]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_832_11.INIT0 = 16'h9666;
    defparam add_832_11.INIT1 = 16'h9666;
    defparam add_832_11.INJECT1_0 = "NO";
    defparam add_832_11.INJECT1_1 = "NO";
    CCU2D add_832_9 (.A0(c_15__N_2408[8]), .B0(c_15__N_2423[8]), .C0(c_15__N_2408[7]), 
          .D0(c_15__N_2423[7]), .A1(c_15__N_2408[9]), .B1(c_15__N_2423[9]), 
          .C1(c_15__N_2408[8]), .D1(c_15__N_2423[8]), .CIN(n19531), .COUT(n19532), 
          .S0(o_r_17__N_2438[9]), .S1(o_r_17__N_2438[10]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_832_9.INIT0 = 16'h9666;
    defparam add_832_9.INIT1 = 16'h9666;
    defparam add_832_9.INJECT1_0 = "NO";
    defparam add_832_9.INJECT1_1 = "NO";
    CCU2D add_832_7 (.A0(c_15__N_2408[6]), .B0(c_15__N_2423[6]), .C0(c_15__N_2408[5]), 
          .D0(c_15__N_2423[5]), .A1(c_15__N_2408[7]), .B1(c_15__N_2423[7]), 
          .C1(c_15__N_2408[6]), .D1(c_15__N_2423[6]), .CIN(n19530), .COUT(n19531), 
          .S0(o_r_17__N_2438[7]), .S1(o_r_17__N_2438[8]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_832_7.INIT0 = 16'h9666;
    defparam add_832_7.INIT1 = 16'h9666;
    defparam add_832_7.INJECT1_0 = "NO";
    defparam add_832_7.INJECT1_1 = "NO";
    CCU2D add_832_5 (.A0(c_15__N_2408[4]), .B0(c_15__N_2423[4]), .C0(c_15__N_2408[3]), 
          .D0(c_15__N_2423[3]), .A1(c_15__N_2408[5]), .B1(c_15__N_2423[5]), 
          .C1(c_15__N_2408[4]), .D1(c_15__N_2423[4]), .CIN(n19529), .COUT(n19530), 
          .S0(o_r_17__N_2438[5]), .S1(o_r_17__N_2438[6]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_832_5.INIT0 = 16'h9666;
    defparam add_832_5.INIT1 = 16'h9666;
    defparam add_832_5.INJECT1_0 = "NO";
    defparam add_832_5.INJECT1_1 = "NO";
    CCU2D add_832_3 (.A0(c_15__N_2408[2]), .B0(c_15__N_2423[2]), .C0(c_15__N_2408[1]), 
          .D0(c_15__N_2423[1]), .A1(c_15__N_2408[3]), .B1(c_15__N_2423[3]), 
          .C1(c_15__N_2408[2]), .D1(c_15__N_2423[2]), .CIN(n19528), .COUT(n19529), 
          .S0(o_r_17__N_2438[3]), .S1(o_r_17__N_2438[4]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_832_3.INIT0 = 16'h9666;
    defparam add_832_3.INIT1 = 16'h9666;
    defparam add_832_3.INJECT1_0 = "NO";
    defparam add_832_3.INJECT1_1 = "NO";
    CCU2D add_832_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(c_15__N_2408[1]), .B1(c_15__N_2423[1]), .C1(n29297), .D1(n29296), 
          .COUT(n19528), .S1(o_r_17__N_2438[2]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_832_1.INIT0 = 16'hF000;
    defparam add_832_1.INIT1 = 16'h9666;
    defparam add_832_1.INJECT1_0 = "NO";
    defparam add_832_1.INJECT1_1 = "NO";
    LUT4 i13627_2_lut (.A(u_l[14]), .B(\u_s[13] ), .Z(c_15__N_2408[14])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13627_2_lut.init = 16'h8888;
    LUT4 i13613_2_lut (.A(u_l[15]), .B(\u_s[12] ), .Z(c_15__N_2423[14])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13613_2_lut.init = 16'h8888;
    LUT4 i13628_2_lut (.A(u_l[13]), .B(\u_s[13] ), .Z(c_15__N_2408[13])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13628_2_lut.init = 16'h8888;
    LUT4 i13614_2_lut (.A(u_l[14]), .B(\u_s[12] ), .Z(c_15__N_2423[13])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13614_2_lut.init = 16'h8888;
    LUT4 i13629_2_lut (.A(u_l[12]), .B(\u_s[13] ), .Z(c_15__N_2408[12])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13629_2_lut.init = 16'h8888;
    LUT4 i13615_2_lut (.A(u_l[13]), .B(\u_s[12] ), .Z(c_15__N_2423[12])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13615_2_lut.init = 16'h8888;
    LUT4 i13630_2_lut (.A(u_l[11]), .B(\u_s[13] ), .Z(c_15__N_2408[11])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13630_2_lut.init = 16'h8888;
    LUT4 i13616_2_lut (.A(u_l[12]), .B(\u_s[12] ), .Z(c_15__N_2423[11])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13616_2_lut.init = 16'h8888;
    LUT4 i13631_2_lut (.A(u_l[10]), .B(\u_s[13] ), .Z(c_15__N_2408[10])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13631_2_lut.init = 16'h8888;
    LUT4 i13617_2_lut (.A(u_l[11]), .B(\u_s[12] ), .Z(c_15__N_2423[10])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13617_2_lut.init = 16'h8888;
    LUT4 i13632_2_lut (.A(u_l[9]), .B(\u_s[13] ), .Z(c_15__N_2408[9])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13632_2_lut.init = 16'h8888;
    LUT4 i13618_2_lut (.A(u_l[10]), .B(\u_s[12] ), .Z(c_15__N_2423[9])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13618_2_lut.init = 16'h8888;
    LUT4 i13633_2_lut (.A(u_l[8]), .B(\u_s[13] ), .Z(c_15__N_2408[8])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13633_2_lut.init = 16'h8888;
    LUT4 i13619_2_lut (.A(u_l[9]), .B(\u_s[12] ), .Z(c_15__N_2423[8])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13619_2_lut.init = 16'h8888;
    LUT4 i13634_2_lut (.A(u_l[7]), .B(\u_s[13] ), .Z(c_15__N_2408[7])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13634_2_lut.init = 16'h8888;
    LUT4 i13620_2_lut (.A(u_l[8]), .B(\u_s[12] ), .Z(c_15__N_2423[7])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13620_2_lut.init = 16'h8888;
    LUT4 i13635_2_lut (.A(u_l[6]), .B(\u_s[13] ), .Z(c_15__N_2408[6])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13635_2_lut.init = 16'h8888;
    LUT4 i13621_2_lut (.A(u_l[7]), .B(\u_s[12] ), .Z(c_15__N_2423[6])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13621_2_lut.init = 16'h8888;
    LUT4 i13636_2_lut (.A(u_l[5]), .B(\u_s[13] ), .Z(c_15__N_2408[5])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13636_2_lut.init = 16'h8888;
    LUT4 i13622_2_lut (.A(u_l[6]), .B(\u_s[12] ), .Z(c_15__N_2423[5])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13622_2_lut.init = 16'h8888;
    LUT4 i13637_2_lut (.A(u_l[4]), .B(\u_s[13] ), .Z(c_15__N_2408[4])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13637_2_lut.init = 16'h8888;
    LUT4 i13623_2_lut (.A(u_l[5]), .B(\u_s[12] ), .Z(c_15__N_2423[4])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13623_2_lut.init = 16'h8888;
    LUT4 i13638_2_lut (.A(u_l[3]), .B(\u_s[13] ), .Z(c_15__N_2408[3])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13638_2_lut.init = 16'h8888;
    LUT4 i13624_2_lut (.A(u_l[4]), .B(\u_s[12] ), .Z(c_15__N_2423[3])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13624_2_lut.init = 16'h8888;
    LUT4 i13639_2_lut (.A(u_l[2]), .B(\u_s[13] ), .Z(c_15__N_2408[2])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13639_2_lut.init = 16'h8888;
    LUT4 i13625_2_lut (.A(u_l[3]), .B(\u_s[12] ), .Z(c_15__N_2423[2])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13625_2_lut.init = 16'h8888;
    LUT4 i13640_2_lut (.A(u_l[1]), .B(\u_s[13] ), .Z(c_15__N_2408[1])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13640_2_lut.init = 16'h8888;
    LUT4 i13626_2_lut (.A(u_l[2]), .B(\u_s[12] ), .Z(c_15__N_2423[1])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13626_2_lut.init = 16'h8888;
    LUT4 i12483_2_lut_rep_636 (.A(u_l[1]), .B(\u_s[12] ), .Z(n29296)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i12483_2_lut_rep_636.init = 16'h8888;
    LUT4 i12482_2_lut_rep_637 (.A(u_l[0]), .B(\u_s[13] ), .Z(n29297)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(51[18:45])
    defparam i12482_2_lut_rep_637.init = 16'h8888;
    LUT4 w_r_16__I_0_i2_2_lut_3_lut_4_lut (.A(u_l[0]), .B(\u_s[13] ), .C(\u_s[12] ), 
         .D(u_l[1]), .Z(o_r_17__N_2438[1])) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(51[18:45])
    defparam w_r_16__I_0_i2_2_lut_3_lut_4_lut.init = 16'h7888;
    FD1S3IX o_r__i17 (.D(o_r_17__N_2438[17]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_06[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=90, LSE_RLINE=90 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i17.GSR = "DISABLED";
    FD1S3IX o_r__i16 (.D(o_r_17__N_2438[16]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_06[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=90, LSE_RLINE=90 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i16.GSR = "DISABLED";
    FD1S3IX o_r__i15 (.D(o_r_17__N_2438[15]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_06[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=90, LSE_RLINE=90 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i15.GSR = "DISABLED";
    FD1S3IX o_r__i14 (.D(o_r_17__N_2438[14]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_06[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=90, LSE_RLINE=90 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i14.GSR = "DISABLED";
    FD1S3IX o_r__i13 (.D(o_r_17__N_2438[13]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_06[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=90, LSE_RLINE=90 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i13.GSR = "DISABLED";
    FD1S3IX o_r__i12 (.D(o_r_17__N_2438[12]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_06[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=90, LSE_RLINE=90 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i12.GSR = "DISABLED";
    FD1S3IX o_r__i11 (.D(o_r_17__N_2438[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_06[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=90, LSE_RLINE=90 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i11.GSR = "DISABLED";
    FD1S3IX o_r__i10 (.D(o_r_17__N_2438[10]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_06[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=90, LSE_RLINE=90 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i10.GSR = "DISABLED";
    FD1S3IX o_r__i9 (.D(o_r_17__N_2438[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_06[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=90, LSE_RLINE=90 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i9.GSR = "DISABLED";
    FD1S3IX o_r__i8 (.D(o_r_17__N_2438[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_06[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=90, LSE_RLINE=90 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i8.GSR = "DISABLED";
    FD1S3IX o_r__i7 (.D(o_r_17__N_2438[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_06[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=90, LSE_RLINE=90 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i7.GSR = "DISABLED";
    FD1S3IX o_r__i6 (.D(o_r_17__N_2438[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_06[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=90, LSE_RLINE=90 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i6.GSR = "DISABLED";
    FD1S3IX o_r__i5 (.D(o_r_17__N_2438[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_06[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=90, LSE_RLINE=90 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i5.GSR = "DISABLED";
    FD1S3IX o_r__i4 (.D(o_r_17__N_2438[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_06[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=90, LSE_RLINE=90 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i4.GSR = "DISABLED";
    FD1S3IX o_r__i3 (.D(o_r_17__N_2438[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_06[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=90, LSE_RLINE=90 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i3.GSR = "DISABLED";
    FD1S3IX o_r__i2 (.D(o_r_17__N_2438[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_06[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=90, LSE_RLINE=90 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i2.GSR = "DISABLED";
    FD1S3IX o_r__i1 (.D(o_r_17__N_2438[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_06[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=90, LSE_RLINE=90 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i1.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module \bimpy(BW=16)_U14 
//

module \bimpy(BW=16)_U14  (S_0_05, dac_clk_p_c, n14224, n9492, GND_net, 
            u_l, \u_s[11] , \u_s[10] , i_sw0_c) /* synthesis syn_module_defined=1 */ ;
    output [17:0]S_0_05;
    input dac_clk_p_c;
    input n14224;
    input n9492;
    input GND_net;
    input [15:0]u_l;
    input \u_s[11] ;
    input \u_s[10] ;
    input i_sw0_c;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[29:38])
    
    wire n19543;
    wire [17:0]o_r_17__N_2438;
    
    wire n19542;
    wire [14:0]c_15__N_2408;
    wire [14:0]c_15__N_2423;
    
    wire n19541, n19540, n19539, n19538, n19537, n19536, n29299, 
        n29298;
    
    FD1S3IX o_r__i0 (.D(n9492), .CK(dac_clk_p_c), .CD(n14224), .Q(S_0_05[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=87, LSE_RLINE=87 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i0.GSR = "DISABLED";
    CCU2D add_833_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19543), 
          .S0(o_r_17__N_2438[17]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_833_cout.INIT0 = 16'h0000;
    defparam add_833_cout.INIT1 = 16'h0000;
    defparam add_833_cout.INJECT1_0 = "NO";
    defparam add_833_cout.INJECT1_1 = "NO";
    CCU2D add_833_15 (.A0(c_15__N_2408[14]), .B0(c_15__N_2423[14]), .C0(c_15__N_2408[13]), 
          .D0(c_15__N_2423[13]), .A1(u_l[15]), .B1(\u_s[11] ), .C1(c_15__N_2408[14]), 
          .D1(c_15__N_2423[14]), .CIN(n19542), .COUT(n19543), .S0(o_r_17__N_2438[15]), 
          .S1(o_r_17__N_2438[16]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_833_15.INIT0 = 16'h9666;
    defparam add_833_15.INIT1 = 16'h7888;
    defparam add_833_15.INJECT1_0 = "NO";
    defparam add_833_15.INJECT1_1 = "NO";
    CCU2D add_833_13 (.A0(c_15__N_2408[12]), .B0(c_15__N_2423[12]), .C0(c_15__N_2408[11]), 
          .D0(c_15__N_2423[11]), .A1(c_15__N_2408[13]), .B1(c_15__N_2423[13]), 
          .C1(c_15__N_2408[12]), .D1(c_15__N_2423[12]), .CIN(n19541), 
          .COUT(n19542), .S0(o_r_17__N_2438[13]), .S1(o_r_17__N_2438[14]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_833_13.INIT0 = 16'h9666;
    defparam add_833_13.INIT1 = 16'h9666;
    defparam add_833_13.INJECT1_0 = "NO";
    defparam add_833_13.INJECT1_1 = "NO";
    CCU2D add_833_11 (.A0(c_15__N_2408[10]), .B0(c_15__N_2423[10]), .C0(c_15__N_2408[9]), 
          .D0(c_15__N_2423[9]), .A1(c_15__N_2408[11]), .B1(c_15__N_2423[11]), 
          .C1(c_15__N_2408[10]), .D1(c_15__N_2423[10]), .CIN(n19540), 
          .COUT(n19541), .S0(o_r_17__N_2438[11]), .S1(o_r_17__N_2438[12]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_833_11.INIT0 = 16'h9666;
    defparam add_833_11.INIT1 = 16'h9666;
    defparam add_833_11.INJECT1_0 = "NO";
    defparam add_833_11.INJECT1_1 = "NO";
    CCU2D add_833_9 (.A0(c_15__N_2408[8]), .B0(c_15__N_2423[8]), .C0(c_15__N_2408[7]), 
          .D0(c_15__N_2423[7]), .A1(c_15__N_2408[9]), .B1(c_15__N_2423[9]), 
          .C1(c_15__N_2408[8]), .D1(c_15__N_2423[8]), .CIN(n19539), .COUT(n19540), 
          .S0(o_r_17__N_2438[9]), .S1(o_r_17__N_2438[10]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_833_9.INIT0 = 16'h9666;
    defparam add_833_9.INIT1 = 16'h9666;
    defparam add_833_9.INJECT1_0 = "NO";
    defparam add_833_9.INJECT1_1 = "NO";
    CCU2D add_833_7 (.A0(c_15__N_2408[6]), .B0(c_15__N_2423[6]), .C0(c_15__N_2408[5]), 
          .D0(c_15__N_2423[5]), .A1(c_15__N_2408[7]), .B1(c_15__N_2423[7]), 
          .C1(c_15__N_2408[6]), .D1(c_15__N_2423[6]), .CIN(n19538), .COUT(n19539), 
          .S0(o_r_17__N_2438[7]), .S1(o_r_17__N_2438[8]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_833_7.INIT0 = 16'h9666;
    defparam add_833_7.INIT1 = 16'h9666;
    defparam add_833_7.INJECT1_0 = "NO";
    defparam add_833_7.INJECT1_1 = "NO";
    CCU2D add_833_5 (.A0(c_15__N_2408[4]), .B0(c_15__N_2423[4]), .C0(c_15__N_2408[3]), 
          .D0(c_15__N_2423[3]), .A1(c_15__N_2408[5]), .B1(c_15__N_2423[5]), 
          .C1(c_15__N_2408[4]), .D1(c_15__N_2423[4]), .CIN(n19537), .COUT(n19538), 
          .S0(o_r_17__N_2438[5]), .S1(o_r_17__N_2438[6]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_833_5.INIT0 = 16'h9666;
    defparam add_833_5.INIT1 = 16'h9666;
    defparam add_833_5.INJECT1_0 = "NO";
    defparam add_833_5.INJECT1_1 = "NO";
    CCU2D add_833_3 (.A0(c_15__N_2408[2]), .B0(c_15__N_2423[2]), .C0(c_15__N_2408[1]), 
          .D0(c_15__N_2423[1]), .A1(c_15__N_2408[3]), .B1(c_15__N_2423[3]), 
          .C1(c_15__N_2408[2]), .D1(c_15__N_2423[2]), .CIN(n19536), .COUT(n19537), 
          .S0(o_r_17__N_2438[3]), .S1(o_r_17__N_2438[4]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_833_3.INIT0 = 16'h9666;
    defparam add_833_3.INIT1 = 16'h9666;
    defparam add_833_3.INJECT1_0 = "NO";
    defparam add_833_3.INJECT1_1 = "NO";
    CCU2D add_833_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(c_15__N_2408[1]), .B1(c_15__N_2423[1]), .C1(n29299), .D1(n29298), 
          .COUT(n19536), .S1(o_r_17__N_2438[2]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_833_1.INIT0 = 16'hF000;
    defparam add_833_1.INIT1 = 16'h9666;
    defparam add_833_1.INJECT1_0 = "NO";
    defparam add_833_1.INJECT1_1 = "NO";
    LUT4 i13657_2_lut (.A(u_l[14]), .B(\u_s[11] ), .Z(c_15__N_2408[14])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13657_2_lut.init = 16'h8888;
    LUT4 i13643_2_lut (.A(u_l[15]), .B(\u_s[10] ), .Z(c_15__N_2423[14])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13643_2_lut.init = 16'h8888;
    LUT4 i13658_2_lut (.A(u_l[13]), .B(\u_s[11] ), .Z(c_15__N_2408[13])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13658_2_lut.init = 16'h8888;
    LUT4 i13644_2_lut (.A(u_l[14]), .B(\u_s[10] ), .Z(c_15__N_2423[13])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13644_2_lut.init = 16'h8888;
    LUT4 i13659_2_lut (.A(u_l[12]), .B(\u_s[11] ), .Z(c_15__N_2408[12])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13659_2_lut.init = 16'h8888;
    LUT4 i13645_2_lut (.A(u_l[13]), .B(\u_s[10] ), .Z(c_15__N_2423[12])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13645_2_lut.init = 16'h8888;
    LUT4 i13660_2_lut (.A(u_l[11]), .B(\u_s[11] ), .Z(c_15__N_2408[11])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13660_2_lut.init = 16'h8888;
    LUT4 i13646_2_lut (.A(u_l[12]), .B(\u_s[10] ), .Z(c_15__N_2423[11])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13646_2_lut.init = 16'h8888;
    LUT4 i13661_2_lut (.A(u_l[10]), .B(\u_s[11] ), .Z(c_15__N_2408[10])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13661_2_lut.init = 16'h8888;
    LUT4 i13647_2_lut (.A(u_l[11]), .B(\u_s[10] ), .Z(c_15__N_2423[10])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13647_2_lut.init = 16'h8888;
    LUT4 i13662_2_lut (.A(u_l[9]), .B(\u_s[11] ), .Z(c_15__N_2408[9])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13662_2_lut.init = 16'h8888;
    LUT4 i13648_2_lut (.A(u_l[10]), .B(\u_s[10] ), .Z(c_15__N_2423[9])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13648_2_lut.init = 16'h8888;
    LUT4 i13663_2_lut (.A(u_l[8]), .B(\u_s[11] ), .Z(c_15__N_2408[8])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13663_2_lut.init = 16'h8888;
    LUT4 i13649_2_lut (.A(u_l[9]), .B(\u_s[10] ), .Z(c_15__N_2423[8])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13649_2_lut.init = 16'h8888;
    LUT4 i13664_2_lut (.A(u_l[7]), .B(\u_s[11] ), .Z(c_15__N_2408[7])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13664_2_lut.init = 16'h8888;
    LUT4 i13650_2_lut (.A(u_l[8]), .B(\u_s[10] ), .Z(c_15__N_2423[7])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13650_2_lut.init = 16'h8888;
    LUT4 i13665_2_lut (.A(u_l[6]), .B(\u_s[11] ), .Z(c_15__N_2408[6])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13665_2_lut.init = 16'h8888;
    LUT4 i13651_2_lut (.A(u_l[7]), .B(\u_s[10] ), .Z(c_15__N_2423[6])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13651_2_lut.init = 16'h8888;
    LUT4 i13666_2_lut (.A(u_l[5]), .B(\u_s[11] ), .Z(c_15__N_2408[5])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13666_2_lut.init = 16'h8888;
    LUT4 i13652_2_lut (.A(u_l[6]), .B(\u_s[10] ), .Z(c_15__N_2423[5])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13652_2_lut.init = 16'h8888;
    LUT4 i13667_2_lut (.A(u_l[4]), .B(\u_s[11] ), .Z(c_15__N_2408[4])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13667_2_lut.init = 16'h8888;
    LUT4 i13653_2_lut (.A(u_l[5]), .B(\u_s[10] ), .Z(c_15__N_2423[4])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13653_2_lut.init = 16'h8888;
    LUT4 i13668_2_lut (.A(u_l[3]), .B(\u_s[11] ), .Z(c_15__N_2408[3])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13668_2_lut.init = 16'h8888;
    LUT4 i13654_2_lut (.A(u_l[4]), .B(\u_s[10] ), .Z(c_15__N_2423[3])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13654_2_lut.init = 16'h8888;
    LUT4 i13669_2_lut (.A(u_l[2]), .B(\u_s[11] ), .Z(c_15__N_2408[2])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13669_2_lut.init = 16'h8888;
    LUT4 i13655_2_lut (.A(u_l[3]), .B(\u_s[10] ), .Z(c_15__N_2423[2])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13655_2_lut.init = 16'h8888;
    LUT4 i13670_2_lut (.A(u_l[1]), .B(\u_s[11] ), .Z(c_15__N_2408[1])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13670_2_lut.init = 16'h8888;
    LUT4 i13656_2_lut (.A(u_l[2]), .B(\u_s[10] ), .Z(c_15__N_2423[1])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13656_2_lut.init = 16'h8888;
    LUT4 i12481_2_lut_rep_638 (.A(u_l[1]), .B(\u_s[10] ), .Z(n29298)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i12481_2_lut_rep_638.init = 16'h8888;
    LUT4 i12480_2_lut_rep_639 (.A(u_l[0]), .B(\u_s[11] ), .Z(n29299)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(51[18:45])
    defparam i12480_2_lut_rep_639.init = 16'h8888;
    LUT4 w_r_16__I_0_i2_2_lut_3_lut_4_lut (.A(u_l[0]), .B(\u_s[11] ), .C(\u_s[10] ), 
         .D(u_l[1]), .Z(o_r_17__N_2438[1])) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(51[18:45])
    defparam w_r_16__I_0_i2_2_lut_3_lut_4_lut.init = 16'h7888;
    FD1S3IX o_r__i17 (.D(o_r_17__N_2438[17]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_05[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=87, LSE_RLINE=87 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i17.GSR = "DISABLED";
    FD1S3IX o_r__i16 (.D(o_r_17__N_2438[16]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_05[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=87, LSE_RLINE=87 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i16.GSR = "DISABLED";
    FD1S3IX o_r__i15 (.D(o_r_17__N_2438[15]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_05[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=87, LSE_RLINE=87 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i15.GSR = "DISABLED";
    FD1S3IX o_r__i14 (.D(o_r_17__N_2438[14]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_05[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=87, LSE_RLINE=87 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i14.GSR = "DISABLED";
    FD1S3IX o_r__i13 (.D(o_r_17__N_2438[13]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_05[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=87, LSE_RLINE=87 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i13.GSR = "DISABLED";
    FD1S3IX o_r__i12 (.D(o_r_17__N_2438[12]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_05[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=87, LSE_RLINE=87 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i12.GSR = "DISABLED";
    FD1S3IX o_r__i11 (.D(o_r_17__N_2438[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_05[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=87, LSE_RLINE=87 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i11.GSR = "DISABLED";
    FD1S3IX o_r__i10 (.D(o_r_17__N_2438[10]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_05[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=87, LSE_RLINE=87 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i10.GSR = "DISABLED";
    FD1S3IX o_r__i9 (.D(o_r_17__N_2438[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_05[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=87, LSE_RLINE=87 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i9.GSR = "DISABLED";
    FD1S3IX o_r__i8 (.D(o_r_17__N_2438[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_05[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=87, LSE_RLINE=87 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i8.GSR = "DISABLED";
    FD1S3IX o_r__i7 (.D(o_r_17__N_2438[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_05[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=87, LSE_RLINE=87 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i7.GSR = "DISABLED";
    FD1S3IX o_r__i6 (.D(o_r_17__N_2438[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_05[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=87, LSE_RLINE=87 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i6.GSR = "DISABLED";
    FD1S3IX o_r__i5 (.D(o_r_17__N_2438[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_05[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=87, LSE_RLINE=87 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i5.GSR = "DISABLED";
    FD1S3IX o_r__i4 (.D(o_r_17__N_2438[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_05[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=87, LSE_RLINE=87 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i4.GSR = "DISABLED";
    FD1S3IX o_r__i3 (.D(o_r_17__N_2438[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_05[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=87, LSE_RLINE=87 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i3.GSR = "DISABLED";
    FD1S3IX o_r__i2 (.D(o_r_17__N_2438[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_05[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=87, LSE_RLINE=87 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i2.GSR = "DISABLED";
    FD1S3IX o_r__i1 (.D(o_r_17__N_2438[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_05[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=75, LSE_LLINE=87, LSE_RLINE=87 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i1.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module \bimpy(BW=16)_U15 
//

module \bimpy(BW=16)_U15  (\S_0_04[0] , dac_clk_p_c, n14224, n9494, 
            GND_net, u_l, \u_s[9] , \u_s[8] , \S_0_04[17] , i_sw0_c, 
            \S_0_04[16] , \S_0_04[15] , \S_0_04[14] , \S_0_04[13] , 
            \S_0_04[12] , \S_0_04[11] , \S_0_04[10] , \S_0_04[9] , \S_0_04[8] , 
            \S_0_04[7] , \S_0_04[6] , \S_0_04[5] , \S_0_04[4] , \S_0_04[3] , 
            \S_0_04[2] , \S_1_02_20__N_2226[1] ) /* synthesis syn_module_defined=1 */ ;
    output \S_0_04[0] ;
    input dac_clk_p_c;
    input n14224;
    input n9494;
    input GND_net;
    input [15:0]u_l;
    input \u_s[9] ;
    input \u_s[8] ;
    output \S_0_04[17] ;
    input i_sw0_c;
    output \S_0_04[16] ;
    output \S_0_04[15] ;
    output \S_0_04[14] ;
    output \S_0_04[13] ;
    output \S_0_04[12] ;
    output \S_0_04[11] ;
    output \S_0_04[10] ;
    output \S_0_04[9] ;
    output \S_0_04[8] ;
    output \S_0_04[7] ;
    output \S_0_04[6] ;
    output \S_0_04[5] ;
    output \S_0_04[4] ;
    output \S_0_04[3] ;
    output \S_0_04[2] ;
    output \S_1_02_20__N_2226[1] ;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[29:38])
    
    wire n19551;
    wire [17:0]o_r_17__N_2438;
    
    wire n19550;
    wire [14:0]c_15__N_2408;
    wire [14:0]c_15__N_2423;
    
    wire n19549, n19548, n19547, n19546, n19545, n19544, n29308, 
        n29307;
    
    FD1S3IX o_r__i0 (.D(n9494), .CK(dac_clk_p_c), .CD(n14224), .Q(\S_0_04[0] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=84, LSE_RLINE=84 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i0.GSR = "DISABLED";
    CCU2D add_834_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19551), 
          .S0(o_r_17__N_2438[17]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_834_cout.INIT0 = 16'h0000;
    defparam add_834_cout.INIT1 = 16'h0000;
    defparam add_834_cout.INJECT1_0 = "NO";
    defparam add_834_cout.INJECT1_1 = "NO";
    CCU2D add_834_15 (.A0(c_15__N_2408[14]), .B0(c_15__N_2423[14]), .C0(c_15__N_2408[13]), 
          .D0(c_15__N_2423[13]), .A1(u_l[15]), .B1(\u_s[9] ), .C1(c_15__N_2408[14]), 
          .D1(c_15__N_2423[14]), .CIN(n19550), .COUT(n19551), .S0(o_r_17__N_2438[15]), 
          .S1(o_r_17__N_2438[16]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_834_15.INIT0 = 16'h9666;
    defparam add_834_15.INIT1 = 16'h7888;
    defparam add_834_15.INJECT1_0 = "NO";
    defparam add_834_15.INJECT1_1 = "NO";
    CCU2D add_834_13 (.A0(c_15__N_2408[12]), .B0(c_15__N_2423[12]), .C0(c_15__N_2408[11]), 
          .D0(c_15__N_2423[11]), .A1(c_15__N_2408[13]), .B1(c_15__N_2423[13]), 
          .C1(c_15__N_2408[12]), .D1(c_15__N_2423[12]), .CIN(n19549), 
          .COUT(n19550), .S0(o_r_17__N_2438[13]), .S1(o_r_17__N_2438[14]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_834_13.INIT0 = 16'h9666;
    defparam add_834_13.INIT1 = 16'h9666;
    defparam add_834_13.INJECT1_0 = "NO";
    defparam add_834_13.INJECT1_1 = "NO";
    CCU2D add_834_11 (.A0(c_15__N_2408[10]), .B0(c_15__N_2423[10]), .C0(c_15__N_2408[9]), 
          .D0(c_15__N_2423[9]), .A1(c_15__N_2408[11]), .B1(c_15__N_2423[11]), 
          .C1(c_15__N_2408[10]), .D1(c_15__N_2423[10]), .CIN(n19548), 
          .COUT(n19549), .S0(o_r_17__N_2438[11]), .S1(o_r_17__N_2438[12]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_834_11.INIT0 = 16'h9666;
    defparam add_834_11.INIT1 = 16'h9666;
    defparam add_834_11.INJECT1_0 = "NO";
    defparam add_834_11.INJECT1_1 = "NO";
    CCU2D add_834_9 (.A0(c_15__N_2408[8]), .B0(c_15__N_2423[8]), .C0(c_15__N_2408[7]), 
          .D0(c_15__N_2423[7]), .A1(c_15__N_2408[9]), .B1(c_15__N_2423[9]), 
          .C1(c_15__N_2408[8]), .D1(c_15__N_2423[8]), .CIN(n19547), .COUT(n19548), 
          .S0(o_r_17__N_2438[9]), .S1(o_r_17__N_2438[10]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_834_9.INIT0 = 16'h9666;
    defparam add_834_9.INIT1 = 16'h9666;
    defparam add_834_9.INJECT1_0 = "NO";
    defparam add_834_9.INJECT1_1 = "NO";
    CCU2D add_834_7 (.A0(c_15__N_2408[6]), .B0(c_15__N_2423[6]), .C0(c_15__N_2408[5]), 
          .D0(c_15__N_2423[5]), .A1(c_15__N_2408[7]), .B1(c_15__N_2423[7]), 
          .C1(c_15__N_2408[6]), .D1(c_15__N_2423[6]), .CIN(n19546), .COUT(n19547), 
          .S0(o_r_17__N_2438[7]), .S1(o_r_17__N_2438[8]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_834_7.INIT0 = 16'h9666;
    defparam add_834_7.INIT1 = 16'h9666;
    defparam add_834_7.INJECT1_0 = "NO";
    defparam add_834_7.INJECT1_1 = "NO";
    CCU2D add_834_5 (.A0(c_15__N_2408[4]), .B0(c_15__N_2423[4]), .C0(c_15__N_2408[3]), 
          .D0(c_15__N_2423[3]), .A1(c_15__N_2408[5]), .B1(c_15__N_2423[5]), 
          .C1(c_15__N_2408[4]), .D1(c_15__N_2423[4]), .CIN(n19545), .COUT(n19546), 
          .S0(o_r_17__N_2438[5]), .S1(o_r_17__N_2438[6]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_834_5.INIT0 = 16'h9666;
    defparam add_834_5.INIT1 = 16'h9666;
    defparam add_834_5.INJECT1_0 = "NO";
    defparam add_834_5.INJECT1_1 = "NO";
    CCU2D add_834_3 (.A0(c_15__N_2408[2]), .B0(c_15__N_2423[2]), .C0(c_15__N_2408[1]), 
          .D0(c_15__N_2423[1]), .A1(c_15__N_2408[3]), .B1(c_15__N_2423[3]), 
          .C1(c_15__N_2408[2]), .D1(c_15__N_2423[2]), .CIN(n19544), .COUT(n19545), 
          .S0(o_r_17__N_2438[3]), .S1(o_r_17__N_2438[4]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_834_3.INIT0 = 16'h9666;
    defparam add_834_3.INIT1 = 16'h9666;
    defparam add_834_3.INJECT1_0 = "NO";
    defparam add_834_3.INJECT1_1 = "NO";
    CCU2D add_834_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(c_15__N_2408[1]), .B1(c_15__N_2423[1]), .C1(n29308), .D1(n29307), 
          .COUT(n19544), .S1(o_r_17__N_2438[2]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_834_1.INIT0 = 16'hF000;
    defparam add_834_1.INIT1 = 16'h9666;
    defparam add_834_1.INJECT1_0 = "NO";
    defparam add_834_1.INJECT1_1 = "NO";
    LUT4 i13686_2_lut (.A(u_l[14]), .B(\u_s[9] ), .Z(c_15__N_2408[14])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13686_2_lut.init = 16'h8888;
    LUT4 i13672_2_lut (.A(u_l[15]), .B(\u_s[8] ), .Z(c_15__N_2423[14])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13672_2_lut.init = 16'h8888;
    LUT4 i13687_2_lut (.A(u_l[13]), .B(\u_s[9] ), .Z(c_15__N_2408[13])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13687_2_lut.init = 16'h8888;
    LUT4 i13673_2_lut (.A(u_l[14]), .B(\u_s[8] ), .Z(c_15__N_2423[13])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13673_2_lut.init = 16'h8888;
    LUT4 i13688_2_lut (.A(u_l[12]), .B(\u_s[9] ), .Z(c_15__N_2408[12])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13688_2_lut.init = 16'h8888;
    LUT4 i13674_2_lut (.A(u_l[13]), .B(\u_s[8] ), .Z(c_15__N_2423[12])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13674_2_lut.init = 16'h8888;
    LUT4 i13689_2_lut (.A(u_l[11]), .B(\u_s[9] ), .Z(c_15__N_2408[11])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13689_2_lut.init = 16'h8888;
    LUT4 i13675_2_lut (.A(u_l[12]), .B(\u_s[8] ), .Z(c_15__N_2423[11])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13675_2_lut.init = 16'h8888;
    LUT4 i13690_2_lut (.A(u_l[10]), .B(\u_s[9] ), .Z(c_15__N_2408[10])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13690_2_lut.init = 16'h8888;
    LUT4 i13676_2_lut (.A(u_l[11]), .B(\u_s[8] ), .Z(c_15__N_2423[10])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13676_2_lut.init = 16'h8888;
    LUT4 i13691_2_lut (.A(u_l[9]), .B(\u_s[9] ), .Z(c_15__N_2408[9])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13691_2_lut.init = 16'h8888;
    LUT4 i13677_2_lut (.A(u_l[10]), .B(\u_s[8] ), .Z(c_15__N_2423[9])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13677_2_lut.init = 16'h8888;
    LUT4 i13692_2_lut (.A(u_l[8]), .B(\u_s[9] ), .Z(c_15__N_2408[8])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13692_2_lut.init = 16'h8888;
    LUT4 i13678_2_lut (.A(u_l[9]), .B(\u_s[8] ), .Z(c_15__N_2423[8])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13678_2_lut.init = 16'h8888;
    LUT4 i13693_2_lut (.A(u_l[7]), .B(\u_s[9] ), .Z(c_15__N_2408[7])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13693_2_lut.init = 16'h8888;
    LUT4 i13679_2_lut (.A(u_l[8]), .B(\u_s[8] ), .Z(c_15__N_2423[7])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13679_2_lut.init = 16'h8888;
    LUT4 i13694_2_lut (.A(u_l[6]), .B(\u_s[9] ), .Z(c_15__N_2408[6])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13694_2_lut.init = 16'h8888;
    LUT4 i13680_2_lut (.A(u_l[7]), .B(\u_s[8] ), .Z(c_15__N_2423[6])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13680_2_lut.init = 16'h8888;
    LUT4 i13695_2_lut (.A(u_l[5]), .B(\u_s[9] ), .Z(c_15__N_2408[5])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13695_2_lut.init = 16'h8888;
    LUT4 i13681_2_lut (.A(u_l[6]), .B(\u_s[8] ), .Z(c_15__N_2423[5])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13681_2_lut.init = 16'h8888;
    LUT4 i13696_2_lut (.A(u_l[4]), .B(\u_s[9] ), .Z(c_15__N_2408[4])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13696_2_lut.init = 16'h8888;
    LUT4 i13682_2_lut (.A(u_l[5]), .B(\u_s[8] ), .Z(c_15__N_2423[4])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13682_2_lut.init = 16'h8888;
    LUT4 i13697_2_lut (.A(u_l[3]), .B(\u_s[9] ), .Z(c_15__N_2408[3])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13697_2_lut.init = 16'h8888;
    LUT4 i13683_2_lut (.A(u_l[4]), .B(\u_s[8] ), .Z(c_15__N_2423[3])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13683_2_lut.init = 16'h8888;
    LUT4 i13698_2_lut (.A(u_l[2]), .B(\u_s[9] ), .Z(c_15__N_2408[2])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13698_2_lut.init = 16'h8888;
    LUT4 i13684_2_lut (.A(u_l[3]), .B(\u_s[8] ), .Z(c_15__N_2423[2])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13684_2_lut.init = 16'h8888;
    LUT4 i13699_2_lut (.A(u_l[1]), .B(\u_s[9] ), .Z(c_15__N_2408[1])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13699_2_lut.init = 16'h8888;
    LUT4 i13685_2_lut (.A(u_l[2]), .B(\u_s[8] ), .Z(c_15__N_2423[1])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13685_2_lut.init = 16'h8888;
    LUT4 i12479_2_lut_rep_647 (.A(u_l[1]), .B(\u_s[8] ), .Z(n29307)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i12479_2_lut_rep_647.init = 16'h8888;
    LUT4 i12477_2_lut_rep_648 (.A(u_l[0]), .B(\u_s[9] ), .Z(n29308)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(51[18:45])
    defparam i12477_2_lut_rep_648.init = 16'h8888;
    LUT4 w_r_16__I_0_i2_2_lut_3_lut_4_lut (.A(u_l[0]), .B(\u_s[9] ), .C(\u_s[8] ), 
         .D(u_l[1]), .Z(o_r_17__N_2438[1])) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(51[18:45])
    defparam w_r_16__I_0_i2_2_lut_3_lut_4_lut.init = 16'h7888;
    FD1S3IX o_r__i17 (.D(o_r_17__N_2438[17]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_04[17] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=84, LSE_RLINE=84 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i17.GSR = "DISABLED";
    FD1S3IX o_r__i16 (.D(o_r_17__N_2438[16]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_04[16] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=84, LSE_RLINE=84 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i16.GSR = "DISABLED";
    FD1S3IX o_r__i15 (.D(o_r_17__N_2438[15]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_04[15] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=84, LSE_RLINE=84 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i15.GSR = "DISABLED";
    FD1S3IX o_r__i14 (.D(o_r_17__N_2438[14]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_04[14] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=84, LSE_RLINE=84 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i14.GSR = "DISABLED";
    FD1S3IX o_r__i13 (.D(o_r_17__N_2438[13]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_04[13] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=84, LSE_RLINE=84 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i13.GSR = "DISABLED";
    FD1S3IX o_r__i12 (.D(o_r_17__N_2438[12]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_04[12] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=84, LSE_RLINE=84 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i12.GSR = "DISABLED";
    FD1S3IX o_r__i11 (.D(o_r_17__N_2438[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_04[11] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=84, LSE_RLINE=84 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i11.GSR = "DISABLED";
    FD1S3IX o_r__i10 (.D(o_r_17__N_2438[10]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_04[10] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=84, LSE_RLINE=84 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i10.GSR = "DISABLED";
    FD1S3IX o_r__i9 (.D(o_r_17__N_2438[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_04[9] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=84, LSE_RLINE=84 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i9.GSR = "DISABLED";
    FD1S3IX o_r__i8 (.D(o_r_17__N_2438[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_04[8] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=84, LSE_RLINE=84 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i8.GSR = "DISABLED";
    FD1S3IX o_r__i7 (.D(o_r_17__N_2438[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_04[7] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=84, LSE_RLINE=84 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i7.GSR = "DISABLED";
    FD1S3IX o_r__i6 (.D(o_r_17__N_2438[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_04[6] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=84, LSE_RLINE=84 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i6.GSR = "DISABLED";
    FD1S3IX o_r__i5 (.D(o_r_17__N_2438[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_04[5] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=84, LSE_RLINE=84 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i5.GSR = "DISABLED";
    FD1S3IX o_r__i4 (.D(o_r_17__N_2438[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_04[4] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=84, LSE_RLINE=84 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i4.GSR = "DISABLED";
    FD1S3IX o_r__i3 (.D(o_r_17__N_2438[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_04[3] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=84, LSE_RLINE=84 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i3.GSR = "DISABLED";
    FD1S3IX o_r__i2 (.D(o_r_17__N_2438[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_04[2] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=84, LSE_RLINE=84 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i2.GSR = "DISABLED";
    FD1S3IX o_r__i1 (.D(o_r_17__N_2438[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_1_02_20__N_2226[1] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=84, LSE_RLINE=84 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i1.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module \bimpy(BW=16)_U16 
//

module \bimpy(BW=16)_U16  (S_0_03, dac_clk_p_c, n14224, n9496, u_l, 
            \u_s[6] , \u_s[7] , i_sw0_c, GND_net) /* synthesis syn_module_defined=1 */ ;
    output [17:0]S_0_03;
    input dac_clk_p_c;
    input n14224;
    input n9496;
    input [15:0]u_l;
    input \u_s[6] ;
    input \u_s[7] ;
    input i_sw0_c;
    input GND_net;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[29:38])
    
    wire n29243, n29244;
    wire [17:0]o_r_17__N_2438;
    wire [14:0]c_15__N_2408;
    wire [14:0]c_15__N_2423;
    
    wire n19721, n19720, n19719, n19718, n19717, n19716, n19715, 
        n19714;
    
    FD1S3IX o_r__i0 (.D(n9496), .CK(dac_clk_p_c), .CD(n14224), .Q(S_0_03[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=81, LSE_RLINE=81 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i0.GSR = "DISABLED";
    LUT4 i12476_2_lut_rep_583 (.A(u_l[1]), .B(\u_s[6] ), .Z(n29243)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i12476_2_lut_rep_583.init = 16'h8888;
    LUT4 i12475_2_lut_rep_584 (.A(u_l[0]), .B(\u_s[7] ), .Z(n29244)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(51[18:45])
    defparam i12475_2_lut_rep_584.init = 16'h8888;
    LUT4 w_r_16__I_0_i2_2_lut_3_lut_4_lut (.A(u_l[0]), .B(\u_s[7] ), .C(\u_s[6] ), 
         .D(u_l[1]), .Z(o_r_17__N_2438[1])) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(51[18:45])
    defparam w_r_16__I_0_i2_2_lut_3_lut_4_lut.init = 16'h7888;
    LUT4 i13716_2_lut (.A(u_l[14]), .B(\u_s[7] ), .Z(c_15__N_2408[14])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13716_2_lut.init = 16'h8888;
    LUT4 i13702_2_lut (.A(u_l[15]), .B(\u_s[6] ), .Z(c_15__N_2423[14])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13702_2_lut.init = 16'h8888;
    LUT4 i13717_2_lut (.A(u_l[13]), .B(\u_s[7] ), .Z(c_15__N_2408[13])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13717_2_lut.init = 16'h8888;
    LUT4 i13703_2_lut (.A(u_l[14]), .B(\u_s[6] ), .Z(c_15__N_2423[13])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13703_2_lut.init = 16'h8888;
    LUT4 i13718_2_lut (.A(u_l[12]), .B(\u_s[7] ), .Z(c_15__N_2408[12])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13718_2_lut.init = 16'h8888;
    LUT4 i13704_2_lut (.A(u_l[13]), .B(\u_s[6] ), .Z(c_15__N_2423[12])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13704_2_lut.init = 16'h8888;
    LUT4 i13719_2_lut (.A(u_l[11]), .B(\u_s[7] ), .Z(c_15__N_2408[11])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13719_2_lut.init = 16'h8888;
    LUT4 i13705_2_lut (.A(u_l[12]), .B(\u_s[6] ), .Z(c_15__N_2423[11])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13705_2_lut.init = 16'h8888;
    LUT4 i13720_2_lut (.A(u_l[10]), .B(\u_s[7] ), .Z(c_15__N_2408[10])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13720_2_lut.init = 16'h8888;
    LUT4 i13706_2_lut (.A(u_l[11]), .B(\u_s[6] ), .Z(c_15__N_2423[10])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13706_2_lut.init = 16'h8888;
    LUT4 i13721_2_lut (.A(u_l[9]), .B(\u_s[7] ), .Z(c_15__N_2408[9])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13721_2_lut.init = 16'h8888;
    LUT4 i13707_2_lut (.A(u_l[10]), .B(\u_s[6] ), .Z(c_15__N_2423[9])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13707_2_lut.init = 16'h8888;
    LUT4 i13722_2_lut (.A(u_l[8]), .B(\u_s[7] ), .Z(c_15__N_2408[8])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13722_2_lut.init = 16'h8888;
    LUT4 i13708_2_lut (.A(u_l[9]), .B(\u_s[6] ), .Z(c_15__N_2423[8])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13708_2_lut.init = 16'h8888;
    LUT4 i13723_2_lut (.A(u_l[7]), .B(\u_s[7] ), .Z(c_15__N_2408[7])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13723_2_lut.init = 16'h8888;
    LUT4 i13709_2_lut (.A(u_l[8]), .B(\u_s[6] ), .Z(c_15__N_2423[7])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13709_2_lut.init = 16'h8888;
    LUT4 i13724_2_lut (.A(u_l[6]), .B(\u_s[7] ), .Z(c_15__N_2408[6])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13724_2_lut.init = 16'h8888;
    LUT4 i13710_2_lut (.A(u_l[7]), .B(\u_s[6] ), .Z(c_15__N_2423[6])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13710_2_lut.init = 16'h8888;
    LUT4 i13725_2_lut (.A(u_l[5]), .B(\u_s[7] ), .Z(c_15__N_2408[5])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13725_2_lut.init = 16'h8888;
    LUT4 i13711_2_lut (.A(u_l[6]), .B(\u_s[6] ), .Z(c_15__N_2423[5])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13711_2_lut.init = 16'h8888;
    LUT4 i13726_2_lut (.A(u_l[4]), .B(\u_s[7] ), .Z(c_15__N_2408[4])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13726_2_lut.init = 16'h8888;
    LUT4 i13712_2_lut (.A(u_l[5]), .B(\u_s[6] ), .Z(c_15__N_2423[4])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13712_2_lut.init = 16'h8888;
    LUT4 i13727_2_lut (.A(u_l[3]), .B(\u_s[7] ), .Z(c_15__N_2408[3])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13727_2_lut.init = 16'h8888;
    LUT4 i13713_2_lut (.A(u_l[4]), .B(\u_s[6] ), .Z(c_15__N_2423[3])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13713_2_lut.init = 16'h8888;
    LUT4 i13728_2_lut (.A(u_l[2]), .B(\u_s[7] ), .Z(c_15__N_2408[2])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13728_2_lut.init = 16'h8888;
    LUT4 i13714_2_lut (.A(u_l[3]), .B(\u_s[6] ), .Z(c_15__N_2423[2])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13714_2_lut.init = 16'h8888;
    LUT4 i13729_2_lut (.A(u_l[1]), .B(\u_s[7] ), .Z(c_15__N_2408[1])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13729_2_lut.init = 16'h8888;
    LUT4 i13715_2_lut (.A(u_l[2]), .B(\u_s[6] ), .Z(c_15__N_2423[1])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13715_2_lut.init = 16'h8888;
    FD1S3IX o_r__i17 (.D(o_r_17__N_2438[17]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_03[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=81, LSE_RLINE=81 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i17.GSR = "DISABLED";
    FD1S3IX o_r__i16 (.D(o_r_17__N_2438[16]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_03[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=81, LSE_RLINE=81 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i16.GSR = "DISABLED";
    FD1S3IX o_r__i15 (.D(o_r_17__N_2438[15]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_03[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=81, LSE_RLINE=81 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i15.GSR = "DISABLED";
    FD1S3IX o_r__i14 (.D(o_r_17__N_2438[14]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_03[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=81, LSE_RLINE=81 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i14.GSR = "DISABLED";
    FD1S3IX o_r__i13 (.D(o_r_17__N_2438[13]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_03[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=81, LSE_RLINE=81 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i13.GSR = "DISABLED";
    FD1S3IX o_r__i12 (.D(o_r_17__N_2438[12]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_03[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=81, LSE_RLINE=81 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i12.GSR = "DISABLED";
    FD1S3IX o_r__i11 (.D(o_r_17__N_2438[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_03[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=81, LSE_RLINE=81 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i11.GSR = "DISABLED";
    FD1S3IX o_r__i10 (.D(o_r_17__N_2438[10]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_03[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=81, LSE_RLINE=81 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i10.GSR = "DISABLED";
    FD1S3IX o_r__i9 (.D(o_r_17__N_2438[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_03[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=81, LSE_RLINE=81 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i9.GSR = "DISABLED";
    FD1S3IX o_r__i8 (.D(o_r_17__N_2438[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_03[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=81, LSE_RLINE=81 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i8.GSR = "DISABLED";
    FD1S3IX o_r__i7 (.D(o_r_17__N_2438[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_03[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=81, LSE_RLINE=81 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i7.GSR = "DISABLED";
    FD1S3IX o_r__i6 (.D(o_r_17__N_2438[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_03[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=81, LSE_RLINE=81 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i6.GSR = "DISABLED";
    FD1S3IX o_r__i5 (.D(o_r_17__N_2438[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_03[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=81, LSE_RLINE=81 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i5.GSR = "DISABLED";
    FD1S3IX o_r__i4 (.D(o_r_17__N_2438[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_03[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=81, LSE_RLINE=81 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i4.GSR = "DISABLED";
    FD1S3IX o_r__i3 (.D(o_r_17__N_2438[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_03[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=81, LSE_RLINE=81 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i3.GSR = "DISABLED";
    FD1S3IX o_r__i2 (.D(o_r_17__N_2438[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_03[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=81, LSE_RLINE=81 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i2.GSR = "DISABLED";
    FD1S3IX o_r__i1 (.D(o_r_17__N_2438[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_03[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=81, LSE_RLINE=81 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i1.GSR = "DISABLED";
    CCU2D add_838_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19721), 
          .S0(o_r_17__N_2438[17]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_838_cout.INIT0 = 16'h0000;
    defparam add_838_cout.INIT1 = 16'h0000;
    defparam add_838_cout.INJECT1_0 = "NO";
    defparam add_838_cout.INJECT1_1 = "NO";
    CCU2D add_838_15 (.A0(c_15__N_2408[14]), .B0(c_15__N_2423[14]), .C0(c_15__N_2408[13]), 
          .D0(c_15__N_2423[13]), .A1(u_l[15]), .B1(\u_s[7] ), .C1(c_15__N_2408[14]), 
          .D1(c_15__N_2423[14]), .CIN(n19720), .COUT(n19721), .S0(o_r_17__N_2438[15]), 
          .S1(o_r_17__N_2438[16]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_838_15.INIT0 = 16'h9666;
    defparam add_838_15.INIT1 = 16'h7888;
    defparam add_838_15.INJECT1_0 = "NO";
    defparam add_838_15.INJECT1_1 = "NO";
    CCU2D add_838_13 (.A0(c_15__N_2408[12]), .B0(c_15__N_2423[12]), .C0(c_15__N_2408[11]), 
          .D0(c_15__N_2423[11]), .A1(c_15__N_2408[13]), .B1(c_15__N_2423[13]), 
          .C1(c_15__N_2408[12]), .D1(c_15__N_2423[12]), .CIN(n19719), 
          .COUT(n19720), .S0(o_r_17__N_2438[13]), .S1(o_r_17__N_2438[14]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_838_13.INIT0 = 16'h9666;
    defparam add_838_13.INIT1 = 16'h9666;
    defparam add_838_13.INJECT1_0 = "NO";
    defparam add_838_13.INJECT1_1 = "NO";
    CCU2D add_838_11 (.A0(c_15__N_2408[10]), .B0(c_15__N_2423[10]), .C0(c_15__N_2408[9]), 
          .D0(c_15__N_2423[9]), .A1(c_15__N_2408[11]), .B1(c_15__N_2423[11]), 
          .C1(c_15__N_2408[10]), .D1(c_15__N_2423[10]), .CIN(n19718), 
          .COUT(n19719), .S0(o_r_17__N_2438[11]), .S1(o_r_17__N_2438[12]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_838_11.INIT0 = 16'h9666;
    defparam add_838_11.INIT1 = 16'h9666;
    defparam add_838_11.INJECT1_0 = "NO";
    defparam add_838_11.INJECT1_1 = "NO";
    CCU2D add_838_9 (.A0(c_15__N_2408[8]), .B0(c_15__N_2423[8]), .C0(c_15__N_2408[7]), 
          .D0(c_15__N_2423[7]), .A1(c_15__N_2408[9]), .B1(c_15__N_2423[9]), 
          .C1(c_15__N_2408[8]), .D1(c_15__N_2423[8]), .CIN(n19717), .COUT(n19718), 
          .S0(o_r_17__N_2438[9]), .S1(o_r_17__N_2438[10]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_838_9.INIT0 = 16'h9666;
    defparam add_838_9.INIT1 = 16'h9666;
    defparam add_838_9.INJECT1_0 = "NO";
    defparam add_838_9.INJECT1_1 = "NO";
    CCU2D add_838_7 (.A0(c_15__N_2408[6]), .B0(c_15__N_2423[6]), .C0(c_15__N_2408[5]), 
          .D0(c_15__N_2423[5]), .A1(c_15__N_2408[7]), .B1(c_15__N_2423[7]), 
          .C1(c_15__N_2408[6]), .D1(c_15__N_2423[6]), .CIN(n19716), .COUT(n19717), 
          .S0(o_r_17__N_2438[7]), .S1(o_r_17__N_2438[8]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_838_7.INIT0 = 16'h9666;
    defparam add_838_7.INIT1 = 16'h9666;
    defparam add_838_7.INJECT1_0 = "NO";
    defparam add_838_7.INJECT1_1 = "NO";
    CCU2D add_838_5 (.A0(c_15__N_2408[4]), .B0(c_15__N_2423[4]), .C0(c_15__N_2408[3]), 
          .D0(c_15__N_2423[3]), .A1(c_15__N_2408[5]), .B1(c_15__N_2423[5]), 
          .C1(c_15__N_2408[4]), .D1(c_15__N_2423[4]), .CIN(n19715), .COUT(n19716), 
          .S0(o_r_17__N_2438[5]), .S1(o_r_17__N_2438[6]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_838_5.INIT0 = 16'h9666;
    defparam add_838_5.INIT1 = 16'h9666;
    defparam add_838_5.INJECT1_0 = "NO";
    defparam add_838_5.INJECT1_1 = "NO";
    CCU2D add_838_3 (.A0(c_15__N_2408[2]), .B0(c_15__N_2423[2]), .C0(c_15__N_2408[1]), 
          .D0(c_15__N_2423[1]), .A1(c_15__N_2408[3]), .B1(c_15__N_2423[3]), 
          .C1(c_15__N_2408[2]), .D1(c_15__N_2423[2]), .CIN(n19714), .COUT(n19715), 
          .S0(o_r_17__N_2438[3]), .S1(o_r_17__N_2438[4]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_838_3.INIT0 = 16'h9666;
    defparam add_838_3.INIT1 = 16'h9666;
    defparam add_838_3.INJECT1_0 = "NO";
    defparam add_838_3.INJECT1_1 = "NO";
    CCU2D add_838_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(c_15__N_2408[1]), .B1(c_15__N_2423[1]), .C1(n29244), .D1(n29243), 
          .COUT(n19714), .S1(o_r_17__N_2438[2]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_838_1.INIT0 = 16'hF000;
    defparam add_838_1.INIT1 = 16'h9666;
    defparam add_838_1.INJECT1_0 = "NO";
    defparam add_838_1.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module \bimpy(BW=16)_U17 
//

module \bimpy(BW=16)_U17  (\S_0_02[0] , dac_clk_p_c, n14224, n9498, 
            GND_net, u_l, \u_s[5] , \u_s[4] , \S_0_02[17] , i_sw0_c, 
            \S_0_02[16] , \S_0_02[15] , \S_0_02[14] , \S_0_02[13] , 
            \S_0_02[12] , \S_0_02[11] , \S_0_02[10] , \S_0_02[9] , \S_0_02[8] , 
            \S_0_02[7] , \S_0_02[6] , \S_0_02[5] , \S_0_02[4] , \S_0_02[3] , 
            \S_0_02[2] , \S_1_01_20__N_2205[1] ) /* synthesis syn_module_defined=1 */ ;
    output \S_0_02[0] ;
    input dac_clk_p_c;
    input n14224;
    input n9498;
    input GND_net;
    input [15:0]u_l;
    input \u_s[5] ;
    input \u_s[4] ;
    output \S_0_02[17] ;
    input i_sw0_c;
    output \S_0_02[16] ;
    output \S_0_02[15] ;
    output \S_0_02[14] ;
    output \S_0_02[13] ;
    output \S_0_02[12] ;
    output \S_0_02[11] ;
    output \S_0_02[10] ;
    output \S_0_02[9] ;
    output \S_0_02[8] ;
    output \S_0_02[7] ;
    output \S_0_02[6] ;
    output \S_0_02[5] ;
    output \S_0_02[4] ;
    output \S_0_02[3] ;
    output \S_0_02[2] ;
    output \S_1_01_20__N_2205[1] ;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[29:38])
    
    wire n19729;
    wire [17:0]o_r_17__N_2438;
    
    wire n19728;
    wire [14:0]c_15__N_2408;
    wire [14:0]c_15__N_2423;
    
    wire n19727, n19726, n19725, n19724, n29245, n29246, n19723, 
        n19722;
    
    FD1S3IX o_r__i0 (.D(n9498), .CK(dac_clk_p_c), .CD(n14224), .Q(\S_0_02[0] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i0.GSR = "DISABLED";
    CCU2D add_839_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19729), 
          .S0(o_r_17__N_2438[17]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_839_cout.INIT0 = 16'h0000;
    defparam add_839_cout.INIT1 = 16'h0000;
    defparam add_839_cout.INJECT1_0 = "NO";
    defparam add_839_cout.INJECT1_1 = "NO";
    CCU2D add_839_15 (.A0(c_15__N_2408[14]), .B0(c_15__N_2423[14]), .C0(c_15__N_2408[13]), 
          .D0(c_15__N_2423[13]), .A1(u_l[15]), .B1(\u_s[5] ), .C1(c_15__N_2408[14]), 
          .D1(c_15__N_2423[14]), .CIN(n19728), .COUT(n19729), .S0(o_r_17__N_2438[15]), 
          .S1(o_r_17__N_2438[16]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_839_15.INIT0 = 16'h9666;
    defparam add_839_15.INIT1 = 16'h7888;
    defparam add_839_15.INJECT1_0 = "NO";
    defparam add_839_15.INJECT1_1 = "NO";
    CCU2D add_839_13 (.A0(c_15__N_2408[12]), .B0(c_15__N_2423[12]), .C0(c_15__N_2408[11]), 
          .D0(c_15__N_2423[11]), .A1(c_15__N_2408[13]), .B1(c_15__N_2423[13]), 
          .C1(c_15__N_2408[12]), .D1(c_15__N_2423[12]), .CIN(n19727), 
          .COUT(n19728), .S0(o_r_17__N_2438[13]), .S1(o_r_17__N_2438[14]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_839_13.INIT0 = 16'h9666;
    defparam add_839_13.INIT1 = 16'h9666;
    defparam add_839_13.INJECT1_0 = "NO";
    defparam add_839_13.INJECT1_1 = "NO";
    CCU2D add_839_11 (.A0(c_15__N_2408[10]), .B0(c_15__N_2423[10]), .C0(c_15__N_2408[9]), 
          .D0(c_15__N_2423[9]), .A1(c_15__N_2408[11]), .B1(c_15__N_2423[11]), 
          .C1(c_15__N_2408[10]), .D1(c_15__N_2423[10]), .CIN(n19726), 
          .COUT(n19727), .S0(o_r_17__N_2438[11]), .S1(o_r_17__N_2438[12]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_839_11.INIT0 = 16'h9666;
    defparam add_839_11.INIT1 = 16'h9666;
    defparam add_839_11.INJECT1_0 = "NO";
    defparam add_839_11.INJECT1_1 = "NO";
    CCU2D add_839_9 (.A0(c_15__N_2408[8]), .B0(c_15__N_2423[8]), .C0(c_15__N_2408[7]), 
          .D0(c_15__N_2423[7]), .A1(c_15__N_2408[9]), .B1(c_15__N_2423[9]), 
          .C1(c_15__N_2408[8]), .D1(c_15__N_2423[8]), .CIN(n19725), .COUT(n19726), 
          .S0(o_r_17__N_2438[9]), .S1(o_r_17__N_2438[10]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_839_9.INIT0 = 16'h9666;
    defparam add_839_9.INIT1 = 16'h9666;
    defparam add_839_9.INJECT1_0 = "NO";
    defparam add_839_9.INJECT1_1 = "NO";
    CCU2D add_839_7 (.A0(c_15__N_2408[6]), .B0(c_15__N_2423[6]), .C0(c_15__N_2408[5]), 
          .D0(c_15__N_2423[5]), .A1(c_15__N_2408[7]), .B1(c_15__N_2423[7]), 
          .C1(c_15__N_2408[6]), .D1(c_15__N_2423[6]), .CIN(n19724), .COUT(n19725), 
          .S0(o_r_17__N_2438[7]), .S1(o_r_17__N_2438[8]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_839_7.INIT0 = 16'h9666;
    defparam add_839_7.INIT1 = 16'h9666;
    defparam add_839_7.INJECT1_0 = "NO";
    defparam add_839_7.INJECT1_1 = "NO";
    LUT4 i13745_2_lut (.A(u_l[14]), .B(\u_s[5] ), .Z(c_15__N_2408[14])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13745_2_lut.init = 16'h8888;
    LUT4 i13731_2_lut (.A(u_l[15]), .B(\u_s[4] ), .Z(c_15__N_2423[14])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13731_2_lut.init = 16'h8888;
    LUT4 i13746_2_lut (.A(u_l[13]), .B(\u_s[5] ), .Z(c_15__N_2408[13])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13746_2_lut.init = 16'h8888;
    LUT4 i13732_2_lut (.A(u_l[14]), .B(\u_s[4] ), .Z(c_15__N_2423[13])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13732_2_lut.init = 16'h8888;
    LUT4 i13747_2_lut (.A(u_l[12]), .B(\u_s[5] ), .Z(c_15__N_2408[12])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13747_2_lut.init = 16'h8888;
    LUT4 i13733_2_lut (.A(u_l[13]), .B(\u_s[4] ), .Z(c_15__N_2423[12])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13733_2_lut.init = 16'h8888;
    LUT4 i13748_2_lut (.A(u_l[11]), .B(\u_s[5] ), .Z(c_15__N_2408[11])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13748_2_lut.init = 16'h8888;
    LUT4 i13734_2_lut (.A(u_l[12]), .B(\u_s[4] ), .Z(c_15__N_2423[11])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13734_2_lut.init = 16'h8888;
    LUT4 i13749_2_lut (.A(u_l[10]), .B(\u_s[5] ), .Z(c_15__N_2408[10])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13749_2_lut.init = 16'h8888;
    LUT4 i13735_2_lut (.A(u_l[11]), .B(\u_s[4] ), .Z(c_15__N_2423[10])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13735_2_lut.init = 16'h8888;
    LUT4 i13750_2_lut (.A(u_l[9]), .B(\u_s[5] ), .Z(c_15__N_2408[9])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13750_2_lut.init = 16'h8888;
    LUT4 i13736_2_lut (.A(u_l[10]), .B(\u_s[4] ), .Z(c_15__N_2423[9])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13736_2_lut.init = 16'h8888;
    LUT4 i13751_2_lut (.A(u_l[8]), .B(\u_s[5] ), .Z(c_15__N_2408[8])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13751_2_lut.init = 16'h8888;
    LUT4 i13737_2_lut (.A(u_l[9]), .B(\u_s[4] ), .Z(c_15__N_2423[8])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13737_2_lut.init = 16'h8888;
    LUT4 i13752_2_lut (.A(u_l[7]), .B(\u_s[5] ), .Z(c_15__N_2408[7])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13752_2_lut.init = 16'h8888;
    LUT4 i13738_2_lut (.A(u_l[8]), .B(\u_s[4] ), .Z(c_15__N_2423[7])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13738_2_lut.init = 16'h8888;
    LUT4 i12474_2_lut_rep_585 (.A(u_l[1]), .B(\u_s[4] ), .Z(n29245)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i12474_2_lut_rep_585.init = 16'h8888;
    LUT4 i12473_2_lut_rep_586 (.A(u_l[0]), .B(\u_s[5] ), .Z(n29246)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(51[18:45])
    defparam i12473_2_lut_rep_586.init = 16'h8888;
    LUT4 i13753_2_lut (.A(u_l[6]), .B(\u_s[5] ), .Z(c_15__N_2408[6])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13753_2_lut.init = 16'h8888;
    LUT4 i13739_2_lut (.A(u_l[7]), .B(\u_s[4] ), .Z(c_15__N_2423[6])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13739_2_lut.init = 16'h8888;
    LUT4 i13754_2_lut (.A(u_l[5]), .B(\u_s[5] ), .Z(c_15__N_2408[5])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13754_2_lut.init = 16'h8888;
    LUT4 i13740_2_lut (.A(u_l[6]), .B(\u_s[4] ), .Z(c_15__N_2423[5])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13740_2_lut.init = 16'h8888;
    LUT4 w_r_16__I_0_i2_2_lut_3_lut_4_lut (.A(u_l[0]), .B(\u_s[5] ), .C(\u_s[4] ), 
         .D(u_l[1]), .Z(o_r_17__N_2438[1])) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(51[18:45])
    defparam w_r_16__I_0_i2_2_lut_3_lut_4_lut.init = 16'h7888;
    CCU2D add_839_5 (.A0(c_15__N_2408[4]), .B0(c_15__N_2423[4]), .C0(c_15__N_2408[3]), 
          .D0(c_15__N_2423[3]), .A1(c_15__N_2408[5]), .B1(c_15__N_2423[5]), 
          .C1(c_15__N_2408[4]), .D1(c_15__N_2423[4]), .CIN(n19723), .COUT(n19724), 
          .S0(o_r_17__N_2438[5]), .S1(o_r_17__N_2438[6]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_839_5.INIT0 = 16'h9666;
    defparam add_839_5.INIT1 = 16'h9666;
    defparam add_839_5.INJECT1_0 = "NO";
    defparam add_839_5.INJECT1_1 = "NO";
    LUT4 i13755_2_lut (.A(u_l[4]), .B(\u_s[5] ), .Z(c_15__N_2408[4])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13755_2_lut.init = 16'h8888;
    LUT4 i13741_2_lut (.A(u_l[5]), .B(\u_s[4] ), .Z(c_15__N_2423[4])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13741_2_lut.init = 16'h8888;
    LUT4 i13756_2_lut (.A(u_l[3]), .B(\u_s[5] ), .Z(c_15__N_2408[3])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13756_2_lut.init = 16'h8888;
    LUT4 i13742_2_lut (.A(u_l[4]), .B(\u_s[4] ), .Z(c_15__N_2423[3])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13742_2_lut.init = 16'h8888;
    LUT4 i13757_2_lut (.A(u_l[2]), .B(\u_s[5] ), .Z(c_15__N_2408[2])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13757_2_lut.init = 16'h8888;
    LUT4 i13743_2_lut (.A(u_l[3]), .B(\u_s[4] ), .Z(c_15__N_2423[2])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13743_2_lut.init = 16'h8888;
    LUT4 i13758_2_lut (.A(u_l[1]), .B(\u_s[5] ), .Z(c_15__N_2408[1])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13758_2_lut.init = 16'h8888;
    LUT4 i13744_2_lut (.A(u_l[2]), .B(\u_s[4] ), .Z(c_15__N_2423[1])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13744_2_lut.init = 16'h8888;
    CCU2D add_839_3 (.A0(c_15__N_2408[2]), .B0(c_15__N_2423[2]), .C0(c_15__N_2408[1]), 
          .D0(c_15__N_2423[1]), .A1(c_15__N_2408[3]), .B1(c_15__N_2423[3]), 
          .C1(c_15__N_2408[2]), .D1(c_15__N_2423[2]), .CIN(n19722), .COUT(n19723), 
          .S0(o_r_17__N_2438[3]), .S1(o_r_17__N_2438[4]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_839_3.INIT0 = 16'h9666;
    defparam add_839_3.INIT1 = 16'h9666;
    defparam add_839_3.INJECT1_0 = "NO";
    defparam add_839_3.INJECT1_1 = "NO";
    CCU2D add_839_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(c_15__N_2408[1]), .B1(c_15__N_2423[1]), .C1(n29246), .D1(n29245), 
          .COUT(n19722), .S1(o_r_17__N_2438[2]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_839_1.INIT0 = 16'hF000;
    defparam add_839_1.INIT1 = 16'h9666;
    defparam add_839_1.INJECT1_0 = "NO";
    defparam add_839_1.INJECT1_1 = "NO";
    FD1S3IX o_r__i17 (.D(o_r_17__N_2438[17]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_02[17] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i17.GSR = "DISABLED";
    FD1S3IX o_r__i16 (.D(o_r_17__N_2438[16]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_02[16] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i16.GSR = "DISABLED";
    FD1S3IX o_r__i15 (.D(o_r_17__N_2438[15]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_02[15] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i15.GSR = "DISABLED";
    FD1S3IX o_r__i14 (.D(o_r_17__N_2438[14]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_02[14] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i14.GSR = "DISABLED";
    FD1S3IX o_r__i13 (.D(o_r_17__N_2438[13]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_02[13] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i13.GSR = "DISABLED";
    FD1S3IX o_r__i12 (.D(o_r_17__N_2438[12]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_02[12] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i12.GSR = "DISABLED";
    FD1S3IX o_r__i11 (.D(o_r_17__N_2438[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_02[11] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i11.GSR = "DISABLED";
    FD1S3IX o_r__i10 (.D(o_r_17__N_2438[10]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_02[10] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i10.GSR = "DISABLED";
    FD1S3IX o_r__i9 (.D(o_r_17__N_2438[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_02[9] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i9.GSR = "DISABLED";
    FD1S3IX o_r__i8 (.D(o_r_17__N_2438[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_02[8] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i8.GSR = "DISABLED";
    FD1S3IX o_r__i7 (.D(o_r_17__N_2438[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_02[7] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i7.GSR = "DISABLED";
    FD1S3IX o_r__i6 (.D(o_r_17__N_2438[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_02[6] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i6.GSR = "DISABLED";
    FD1S3IX o_r__i5 (.D(o_r_17__N_2438[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_02[5] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i5.GSR = "DISABLED";
    FD1S3IX o_r__i4 (.D(o_r_17__N_2438[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_02[4] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i4.GSR = "DISABLED";
    FD1S3IX o_r__i3 (.D(o_r_17__N_2438[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_02[3] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i3.GSR = "DISABLED";
    FD1S3IX o_r__i2 (.D(o_r_17__N_2438[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_02[2] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i2.GSR = "DISABLED";
    FD1S3IX o_r__i1 (.D(o_r_17__N_2438[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_1_01_20__N_2205[1] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i1.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module \bimpy(BW=16)_U18 
//

module \bimpy(BW=16)_U18  (S_0_01, dac_clk_p_c, n14224, n9504, GND_net, 
            u_l, \u_s[3] , \u_s[2] , i_sw0_c) /* synthesis syn_module_defined=1 */ ;
    output [17:0]S_0_01;
    input dac_clk_p_c;
    input n14224;
    input n9504;
    input GND_net;
    input [15:0]u_l;
    input \u_s[3] ;
    input \u_s[2] ;
    input i_sw0_c;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[29:38])
    
    wire n19737;
    wire [17:0]o_r_17__N_2438;
    
    wire n19736;
    wire [14:0]c_15__N_2408;
    wire [14:0]c_15__N_2423;
    
    wire n19735, n19734, n19733, n19732, n19731, n19730, n29260, 
        n29259;
    
    FD1S3IX o_r__i0 (.D(n9504), .CK(dac_clk_p_c), .CD(n14224), .Q(S_0_01[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=75, LSE_RLINE=75 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i0.GSR = "DISABLED";
    CCU2D add_840_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19737), 
          .S0(o_r_17__N_2438[17]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_840_cout.INIT0 = 16'h0000;
    defparam add_840_cout.INIT1 = 16'h0000;
    defparam add_840_cout.INJECT1_0 = "NO";
    defparam add_840_cout.INJECT1_1 = "NO";
    CCU2D add_840_15 (.A0(c_15__N_2408[14]), .B0(c_15__N_2423[14]), .C0(c_15__N_2408[13]), 
          .D0(c_15__N_2423[13]), .A1(u_l[15]), .B1(\u_s[3] ), .C1(c_15__N_2408[14]), 
          .D1(c_15__N_2423[14]), .CIN(n19736), .COUT(n19737), .S0(o_r_17__N_2438[15]), 
          .S1(o_r_17__N_2438[16]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_840_15.INIT0 = 16'h9666;
    defparam add_840_15.INIT1 = 16'h7888;
    defparam add_840_15.INJECT1_0 = "NO";
    defparam add_840_15.INJECT1_1 = "NO";
    CCU2D add_840_13 (.A0(c_15__N_2408[12]), .B0(c_15__N_2423[12]), .C0(c_15__N_2408[11]), 
          .D0(c_15__N_2423[11]), .A1(c_15__N_2408[13]), .B1(c_15__N_2423[13]), 
          .C1(c_15__N_2408[12]), .D1(c_15__N_2423[12]), .CIN(n19735), 
          .COUT(n19736), .S0(o_r_17__N_2438[13]), .S1(o_r_17__N_2438[14]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_840_13.INIT0 = 16'h9666;
    defparam add_840_13.INIT1 = 16'h9666;
    defparam add_840_13.INJECT1_0 = "NO";
    defparam add_840_13.INJECT1_1 = "NO";
    CCU2D add_840_11 (.A0(c_15__N_2408[10]), .B0(c_15__N_2423[10]), .C0(c_15__N_2408[9]), 
          .D0(c_15__N_2423[9]), .A1(c_15__N_2408[11]), .B1(c_15__N_2423[11]), 
          .C1(c_15__N_2408[10]), .D1(c_15__N_2423[10]), .CIN(n19734), 
          .COUT(n19735), .S0(o_r_17__N_2438[11]), .S1(o_r_17__N_2438[12]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_840_11.INIT0 = 16'h9666;
    defparam add_840_11.INIT1 = 16'h9666;
    defparam add_840_11.INJECT1_0 = "NO";
    defparam add_840_11.INJECT1_1 = "NO";
    CCU2D add_840_9 (.A0(c_15__N_2408[8]), .B0(c_15__N_2423[8]), .C0(c_15__N_2408[7]), 
          .D0(c_15__N_2423[7]), .A1(c_15__N_2408[9]), .B1(c_15__N_2423[9]), 
          .C1(c_15__N_2408[8]), .D1(c_15__N_2423[8]), .CIN(n19733), .COUT(n19734), 
          .S0(o_r_17__N_2438[9]), .S1(o_r_17__N_2438[10]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_840_9.INIT0 = 16'h9666;
    defparam add_840_9.INIT1 = 16'h9666;
    defparam add_840_9.INJECT1_0 = "NO";
    defparam add_840_9.INJECT1_1 = "NO";
    CCU2D add_840_7 (.A0(c_15__N_2408[6]), .B0(c_15__N_2423[6]), .C0(c_15__N_2408[5]), 
          .D0(c_15__N_2423[5]), .A1(c_15__N_2408[7]), .B1(c_15__N_2423[7]), 
          .C1(c_15__N_2408[6]), .D1(c_15__N_2423[6]), .CIN(n19732), .COUT(n19733), 
          .S0(o_r_17__N_2438[7]), .S1(o_r_17__N_2438[8]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_840_7.INIT0 = 16'h9666;
    defparam add_840_7.INIT1 = 16'h9666;
    defparam add_840_7.INJECT1_0 = "NO";
    defparam add_840_7.INJECT1_1 = "NO";
    CCU2D add_840_5 (.A0(c_15__N_2408[4]), .B0(c_15__N_2423[4]), .C0(c_15__N_2408[3]), 
          .D0(c_15__N_2423[3]), .A1(c_15__N_2408[5]), .B1(c_15__N_2423[5]), 
          .C1(c_15__N_2408[4]), .D1(c_15__N_2423[4]), .CIN(n19731), .COUT(n19732), 
          .S0(o_r_17__N_2438[5]), .S1(o_r_17__N_2438[6]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_840_5.INIT0 = 16'h9666;
    defparam add_840_5.INIT1 = 16'h9666;
    defparam add_840_5.INJECT1_0 = "NO";
    defparam add_840_5.INJECT1_1 = "NO";
    CCU2D add_840_3 (.A0(c_15__N_2408[2]), .B0(c_15__N_2423[2]), .C0(c_15__N_2408[1]), 
          .D0(c_15__N_2423[1]), .A1(c_15__N_2408[3]), .B1(c_15__N_2423[3]), 
          .C1(c_15__N_2408[2]), .D1(c_15__N_2423[2]), .CIN(n19730), .COUT(n19731), 
          .S0(o_r_17__N_2438[3]), .S1(o_r_17__N_2438[4]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_840_3.INIT0 = 16'h9666;
    defparam add_840_3.INIT1 = 16'h9666;
    defparam add_840_3.INJECT1_0 = "NO";
    defparam add_840_3.INJECT1_1 = "NO";
    LUT4 i13774_2_lut (.A(u_l[14]), .B(\u_s[3] ), .Z(c_15__N_2408[14])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13774_2_lut.init = 16'h8888;
    CCU2D add_840_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(c_15__N_2408[1]), .B1(c_15__N_2423[1]), .C1(n29260), .D1(n29259), 
          .COUT(n19730), .S1(o_r_17__N_2438[2]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_840_1.INIT0 = 16'hF000;
    defparam add_840_1.INIT1 = 16'h9666;
    defparam add_840_1.INJECT1_0 = "NO";
    defparam add_840_1.INJECT1_1 = "NO";
    LUT4 i13760_2_lut (.A(u_l[15]), .B(\u_s[2] ), .Z(c_15__N_2423[14])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13760_2_lut.init = 16'h8888;
    LUT4 i13775_2_lut (.A(u_l[13]), .B(\u_s[3] ), .Z(c_15__N_2408[13])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13775_2_lut.init = 16'h8888;
    LUT4 i13761_2_lut (.A(u_l[14]), .B(\u_s[2] ), .Z(c_15__N_2423[13])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13761_2_lut.init = 16'h8888;
    LUT4 i13776_2_lut (.A(u_l[12]), .B(\u_s[3] ), .Z(c_15__N_2408[12])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13776_2_lut.init = 16'h8888;
    LUT4 i13762_2_lut (.A(u_l[13]), .B(\u_s[2] ), .Z(c_15__N_2423[12])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13762_2_lut.init = 16'h8888;
    LUT4 i13777_2_lut (.A(u_l[11]), .B(\u_s[3] ), .Z(c_15__N_2408[11])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13777_2_lut.init = 16'h8888;
    LUT4 i13763_2_lut (.A(u_l[12]), .B(\u_s[2] ), .Z(c_15__N_2423[11])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13763_2_lut.init = 16'h8888;
    LUT4 i13778_2_lut (.A(u_l[10]), .B(\u_s[3] ), .Z(c_15__N_2408[10])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13778_2_lut.init = 16'h8888;
    LUT4 i13764_2_lut (.A(u_l[11]), .B(\u_s[2] ), .Z(c_15__N_2423[10])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13764_2_lut.init = 16'h8888;
    LUT4 i13779_2_lut (.A(u_l[9]), .B(\u_s[3] ), .Z(c_15__N_2408[9])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13779_2_lut.init = 16'h8888;
    LUT4 i13765_2_lut (.A(u_l[10]), .B(\u_s[2] ), .Z(c_15__N_2423[9])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13765_2_lut.init = 16'h8888;
    LUT4 i13780_2_lut (.A(u_l[8]), .B(\u_s[3] ), .Z(c_15__N_2408[8])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13780_2_lut.init = 16'h8888;
    LUT4 i13766_2_lut (.A(u_l[9]), .B(\u_s[2] ), .Z(c_15__N_2423[8])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13766_2_lut.init = 16'h8888;
    LUT4 i13781_2_lut (.A(u_l[7]), .B(\u_s[3] ), .Z(c_15__N_2408[7])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13781_2_lut.init = 16'h8888;
    LUT4 i13767_2_lut (.A(u_l[8]), .B(\u_s[2] ), .Z(c_15__N_2423[7])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13767_2_lut.init = 16'h8888;
    LUT4 i13782_2_lut (.A(u_l[6]), .B(\u_s[3] ), .Z(c_15__N_2408[6])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13782_2_lut.init = 16'h8888;
    LUT4 i13768_2_lut (.A(u_l[7]), .B(\u_s[2] ), .Z(c_15__N_2423[6])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13768_2_lut.init = 16'h8888;
    LUT4 i13783_2_lut (.A(u_l[5]), .B(\u_s[3] ), .Z(c_15__N_2408[5])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13783_2_lut.init = 16'h8888;
    LUT4 i13769_2_lut (.A(u_l[6]), .B(\u_s[2] ), .Z(c_15__N_2423[5])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13769_2_lut.init = 16'h8888;
    LUT4 i13784_2_lut (.A(u_l[4]), .B(\u_s[3] ), .Z(c_15__N_2408[4])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13784_2_lut.init = 16'h8888;
    LUT4 i13770_2_lut (.A(u_l[5]), .B(\u_s[2] ), .Z(c_15__N_2423[4])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13770_2_lut.init = 16'h8888;
    LUT4 i13785_2_lut (.A(u_l[3]), .B(\u_s[3] ), .Z(c_15__N_2408[3])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13785_2_lut.init = 16'h8888;
    LUT4 i13771_2_lut (.A(u_l[4]), .B(\u_s[2] ), .Z(c_15__N_2423[3])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13771_2_lut.init = 16'h8888;
    LUT4 i13786_2_lut (.A(u_l[2]), .B(\u_s[3] ), .Z(c_15__N_2408[2])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13786_2_lut.init = 16'h8888;
    LUT4 i13772_2_lut (.A(u_l[3]), .B(\u_s[2] ), .Z(c_15__N_2423[2])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13772_2_lut.init = 16'h8888;
    LUT4 i13787_2_lut (.A(u_l[1]), .B(\u_s[3] ), .Z(c_15__N_2408[1])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13787_2_lut.init = 16'h8888;
    LUT4 i13773_2_lut (.A(u_l[2]), .B(\u_s[2] ), .Z(c_15__N_2423[1])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13773_2_lut.init = 16'h8888;
    FD1S3IX o_r__i17 (.D(o_r_17__N_2438[17]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_01[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=75, LSE_RLINE=75 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i17.GSR = "DISABLED";
    FD1S3IX o_r__i16 (.D(o_r_17__N_2438[16]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_01[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=75, LSE_RLINE=75 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i16.GSR = "DISABLED";
    FD1S3IX o_r__i15 (.D(o_r_17__N_2438[15]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_01[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=75, LSE_RLINE=75 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i15.GSR = "DISABLED";
    FD1S3IX o_r__i14 (.D(o_r_17__N_2438[14]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_01[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=75, LSE_RLINE=75 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i14.GSR = "DISABLED";
    FD1S3IX o_r__i13 (.D(o_r_17__N_2438[13]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_01[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=75, LSE_RLINE=75 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i13.GSR = "DISABLED";
    FD1S3IX o_r__i12 (.D(o_r_17__N_2438[12]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_01[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=75, LSE_RLINE=75 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i12.GSR = "DISABLED";
    FD1S3IX o_r__i11 (.D(o_r_17__N_2438[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_01[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=75, LSE_RLINE=75 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i11.GSR = "DISABLED";
    FD1S3IX o_r__i10 (.D(o_r_17__N_2438[10]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_01[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=75, LSE_RLINE=75 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i10.GSR = "DISABLED";
    FD1S3IX o_r__i9 (.D(o_r_17__N_2438[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_01[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=75, LSE_RLINE=75 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i9.GSR = "DISABLED";
    FD1S3IX o_r__i8 (.D(o_r_17__N_2438[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_01[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=75, LSE_RLINE=75 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i8.GSR = "DISABLED";
    FD1S3IX o_r__i7 (.D(o_r_17__N_2438[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_01[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=75, LSE_RLINE=75 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i7.GSR = "DISABLED";
    FD1S3IX o_r__i6 (.D(o_r_17__N_2438[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_01[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=75, LSE_RLINE=75 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i6.GSR = "DISABLED";
    FD1S3IX o_r__i5 (.D(o_r_17__N_2438[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_01[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=75, LSE_RLINE=75 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i5.GSR = "DISABLED";
    FD1S3IX o_r__i4 (.D(o_r_17__N_2438[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_01[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=75, LSE_RLINE=75 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i4.GSR = "DISABLED";
    FD1S3IX o_r__i3 (.D(o_r_17__N_2438[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_01[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=75, LSE_RLINE=75 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i3.GSR = "DISABLED";
    FD1S3IX o_r__i2 (.D(o_r_17__N_2438[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_01[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=75, LSE_RLINE=75 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i2.GSR = "DISABLED";
    FD1S3IX o_r__i1 (.D(o_r_17__N_2438[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(S_0_01[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=75, LSE_RLINE=75 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i1.GSR = "DISABLED";
    LUT4 i12472_2_lut_rep_599 (.A(u_l[1]), .B(\u_s[2] ), .Z(n29259)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i12472_2_lut_rep_599.init = 16'h8888;
    LUT4 i12471_2_lut_rep_600 (.A(u_l[0]), .B(\u_s[3] ), .Z(n29260)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(51[18:45])
    defparam i12471_2_lut_rep_600.init = 16'h8888;
    LUT4 w_r_16__I_0_i2_2_lut_3_lut_4_lut (.A(u_l[0]), .B(\u_s[3] ), .C(\u_s[2] ), 
         .D(u_l[1]), .Z(o_r_17__N_2438[1])) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(51[18:45])
    defparam w_r_16__I_0_i2_2_lut_3_lut_4_lut.init = 16'h7888;
    
endmodule
//
// Verilog Description of module \bimpy(BW=16)_U19 
//

module \bimpy(BW=16)_U19  (u_l, \u_s[1] , \u_s[0] , \S_0_00[0] , dac_clk_p_c, 
            n14224, n9506, GND_net, \S_0_00[17] , i_sw0_c, \S_0_00[16] , 
            \S_0_00[15] , \S_0_00[14] , \S_0_00[13] , \S_0_00[12] , 
            \S_0_00[11] , \S_0_00[10] , \S_0_00[9] , \S_0_00[8] , \S_0_00[7] , 
            \S_0_00[6] , \S_0_00[5] , \S_0_00[4] , \S_0_00[3] , \S_0_00[2] , 
            \S_1_00_20__N_2184[1] ) /* synthesis syn_module_defined=1 */ ;
    input [15:0]u_l;
    input \u_s[1] ;
    input \u_s[0] ;
    output \S_0_00[0] ;
    input dac_clk_p_c;
    input n14224;
    input n9506;
    input GND_net;
    output \S_0_00[17] ;
    input i_sw0_c;
    output \S_0_00[16] ;
    output \S_0_00[15] ;
    output \S_0_00[14] ;
    output \S_0_00[13] ;
    output \S_0_00[12] ;
    output \S_0_00[11] ;
    output \S_0_00[10] ;
    output \S_0_00[9] ;
    output \S_0_00[8] ;
    output \S_0_00[7] ;
    output \S_0_00[6] ;
    output \S_0_00[5] ;
    output \S_0_00[4] ;
    output \S_0_00[3] ;
    output \S_0_00[2] ;
    output \S_1_00_20__N_2184[1] ;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[29:38])
    wire [14:0]c_15__N_2408;
    wire [14:0]c_15__N_2423;
    
    wire n19753;
    wire [17:0]o_r_17__N_2438;
    
    wire n19752, n19751, n19750, n19749, n19748, n19747, n19746, 
        n29265, n29264;
    
    LUT4 i13813_2_lut (.A(u_l[4]), .B(\u_s[1] ), .Z(c_15__N_2408[4])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13813_2_lut.init = 16'h8888;
    LUT4 i13799_2_lut (.A(u_l[5]), .B(\u_s[0] ), .Z(c_15__N_2423[4])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13799_2_lut.init = 16'h8888;
    LUT4 i13814_2_lut (.A(u_l[3]), .B(\u_s[1] ), .Z(c_15__N_2408[3])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13814_2_lut.init = 16'h8888;
    LUT4 i13800_2_lut (.A(u_l[4]), .B(\u_s[0] ), .Z(c_15__N_2423[3])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13800_2_lut.init = 16'h8888;
    LUT4 i13815_2_lut (.A(u_l[2]), .B(\u_s[1] ), .Z(c_15__N_2408[2])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13815_2_lut.init = 16'h8888;
    LUT4 i13801_2_lut (.A(u_l[3]), .B(\u_s[0] ), .Z(c_15__N_2423[2])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13801_2_lut.init = 16'h8888;
    LUT4 i13816_2_lut (.A(u_l[1]), .B(\u_s[1] ), .Z(c_15__N_2408[1])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13816_2_lut.init = 16'h8888;
    LUT4 i13802_2_lut (.A(u_l[2]), .B(\u_s[0] ), .Z(c_15__N_2423[1])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13802_2_lut.init = 16'h8888;
    FD1S3IX o_r__i0 (.D(n9506), .CK(dac_clk_p_c), .CD(n14224), .Q(\S_0_00[0] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i0.GSR = "DISABLED";
    CCU2D add_841_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19753), 
          .S0(o_r_17__N_2438[17]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_841_cout.INIT0 = 16'h0000;
    defparam add_841_cout.INIT1 = 16'h0000;
    defparam add_841_cout.INJECT1_0 = "NO";
    defparam add_841_cout.INJECT1_1 = "NO";
    CCU2D add_841_15 (.A0(c_15__N_2408[14]), .B0(c_15__N_2423[14]), .C0(c_15__N_2408[13]), 
          .D0(c_15__N_2423[13]), .A1(u_l[15]), .B1(\u_s[1] ), .C1(c_15__N_2408[14]), 
          .D1(c_15__N_2423[14]), .CIN(n19752), .COUT(n19753), .S0(o_r_17__N_2438[15]), 
          .S1(o_r_17__N_2438[16]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_841_15.INIT0 = 16'h9666;
    defparam add_841_15.INIT1 = 16'h7888;
    defparam add_841_15.INJECT1_0 = "NO";
    defparam add_841_15.INJECT1_1 = "NO";
    CCU2D add_841_13 (.A0(c_15__N_2408[12]), .B0(c_15__N_2423[12]), .C0(c_15__N_2408[11]), 
          .D0(c_15__N_2423[11]), .A1(c_15__N_2408[13]), .B1(c_15__N_2423[13]), 
          .C1(c_15__N_2408[12]), .D1(c_15__N_2423[12]), .CIN(n19751), 
          .COUT(n19752), .S0(o_r_17__N_2438[13]), .S1(o_r_17__N_2438[14]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_841_13.INIT0 = 16'h9666;
    defparam add_841_13.INIT1 = 16'h9666;
    defparam add_841_13.INJECT1_0 = "NO";
    defparam add_841_13.INJECT1_1 = "NO";
    CCU2D add_841_11 (.A0(c_15__N_2408[10]), .B0(c_15__N_2423[10]), .C0(c_15__N_2408[9]), 
          .D0(c_15__N_2423[9]), .A1(c_15__N_2408[11]), .B1(c_15__N_2423[11]), 
          .C1(c_15__N_2408[10]), .D1(c_15__N_2423[10]), .CIN(n19750), 
          .COUT(n19751), .S0(o_r_17__N_2438[11]), .S1(o_r_17__N_2438[12]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_841_11.INIT0 = 16'h9666;
    defparam add_841_11.INIT1 = 16'h9666;
    defparam add_841_11.INJECT1_0 = "NO";
    defparam add_841_11.INJECT1_1 = "NO";
    CCU2D add_841_9 (.A0(c_15__N_2408[8]), .B0(c_15__N_2423[8]), .C0(c_15__N_2408[7]), 
          .D0(c_15__N_2423[7]), .A1(c_15__N_2408[9]), .B1(c_15__N_2423[9]), 
          .C1(c_15__N_2408[8]), .D1(c_15__N_2423[8]), .CIN(n19749), .COUT(n19750), 
          .S0(o_r_17__N_2438[9]), .S1(o_r_17__N_2438[10]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_841_9.INIT0 = 16'h9666;
    defparam add_841_9.INIT1 = 16'h9666;
    defparam add_841_9.INJECT1_0 = "NO";
    defparam add_841_9.INJECT1_1 = "NO";
    CCU2D add_841_7 (.A0(c_15__N_2408[6]), .B0(c_15__N_2423[6]), .C0(c_15__N_2408[5]), 
          .D0(c_15__N_2423[5]), .A1(c_15__N_2408[7]), .B1(c_15__N_2423[7]), 
          .C1(c_15__N_2408[6]), .D1(c_15__N_2423[6]), .CIN(n19748), .COUT(n19749), 
          .S0(o_r_17__N_2438[7]), .S1(o_r_17__N_2438[8]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_841_7.INIT0 = 16'h9666;
    defparam add_841_7.INIT1 = 16'h9666;
    defparam add_841_7.INJECT1_0 = "NO";
    defparam add_841_7.INJECT1_1 = "NO";
    CCU2D add_841_5 (.A0(c_15__N_2408[4]), .B0(c_15__N_2423[4]), .C0(c_15__N_2408[3]), 
          .D0(c_15__N_2423[3]), .A1(c_15__N_2408[5]), .B1(c_15__N_2423[5]), 
          .C1(c_15__N_2408[4]), .D1(c_15__N_2423[4]), .CIN(n19747), .COUT(n19748), 
          .S0(o_r_17__N_2438[5]), .S1(o_r_17__N_2438[6]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_841_5.INIT0 = 16'h9666;
    defparam add_841_5.INIT1 = 16'h9666;
    defparam add_841_5.INJECT1_0 = "NO";
    defparam add_841_5.INJECT1_1 = "NO";
    CCU2D add_841_3 (.A0(c_15__N_2408[2]), .B0(c_15__N_2423[2]), .C0(c_15__N_2408[1]), 
          .D0(c_15__N_2423[1]), .A1(c_15__N_2408[3]), .B1(c_15__N_2423[3]), 
          .C1(c_15__N_2408[2]), .D1(c_15__N_2423[2]), .CIN(n19746), .COUT(n19747), 
          .S0(o_r_17__N_2438[3]), .S1(o_r_17__N_2438[4]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_841_3.INIT0 = 16'h9666;
    defparam add_841_3.INIT1 = 16'h9666;
    defparam add_841_3.INJECT1_0 = "NO";
    defparam add_841_3.INJECT1_1 = "NO";
    CCU2D add_841_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(c_15__N_2408[1]), .B1(c_15__N_2423[1]), .C1(n29265), .D1(n29264), 
          .COUT(n19746), .S1(o_r_17__N_2438[2]));   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(61[10:27])
    defparam add_841_1.INIT0 = 16'hF000;
    defparam add_841_1.INIT1 = 16'h9666;
    defparam add_841_1.INJECT1_0 = "NO";
    defparam add_841_1.INJECT1_1 = "NO";
    LUT4 i13803_2_lut (.A(u_l[14]), .B(\u_s[1] ), .Z(c_15__N_2408[14])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13803_2_lut.init = 16'h8888;
    LUT4 i13789_2_lut (.A(u_l[15]), .B(\u_s[0] ), .Z(c_15__N_2423[14])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13789_2_lut.init = 16'h8888;
    LUT4 i13804_2_lut (.A(u_l[13]), .B(\u_s[1] ), .Z(c_15__N_2408[13])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13804_2_lut.init = 16'h8888;
    LUT4 i13790_2_lut (.A(u_l[14]), .B(\u_s[0] ), .Z(c_15__N_2423[13])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13790_2_lut.init = 16'h8888;
    LUT4 i13805_2_lut (.A(u_l[12]), .B(\u_s[1] ), .Z(c_15__N_2408[12])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13805_2_lut.init = 16'h8888;
    LUT4 i13791_2_lut (.A(u_l[13]), .B(\u_s[0] ), .Z(c_15__N_2423[12])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13791_2_lut.init = 16'h8888;
    LUT4 i13806_2_lut (.A(u_l[11]), .B(\u_s[1] ), .Z(c_15__N_2408[11])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13806_2_lut.init = 16'h8888;
    LUT4 i13792_2_lut (.A(u_l[12]), .B(\u_s[0] ), .Z(c_15__N_2423[11])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13792_2_lut.init = 16'h8888;
    LUT4 i13807_2_lut (.A(u_l[10]), .B(\u_s[1] ), .Z(c_15__N_2408[10])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13807_2_lut.init = 16'h8888;
    LUT4 i13793_2_lut (.A(u_l[11]), .B(\u_s[0] ), .Z(c_15__N_2423[10])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13793_2_lut.init = 16'h8888;
    LUT4 i13808_2_lut (.A(u_l[9]), .B(\u_s[1] ), .Z(c_15__N_2408[9])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13808_2_lut.init = 16'h8888;
    LUT4 i13794_2_lut (.A(u_l[10]), .B(\u_s[0] ), .Z(c_15__N_2423[9])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13794_2_lut.init = 16'h8888;
    LUT4 i13809_2_lut (.A(u_l[8]), .B(\u_s[1] ), .Z(c_15__N_2408[8])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13809_2_lut.init = 16'h8888;
    LUT4 i13795_2_lut (.A(u_l[9]), .B(\u_s[0] ), .Z(c_15__N_2423[8])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13795_2_lut.init = 16'h8888;
    LUT4 i13810_2_lut (.A(u_l[7]), .B(\u_s[1] ), .Z(c_15__N_2408[7])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13810_2_lut.init = 16'h8888;
    LUT4 i13796_2_lut (.A(u_l[8]), .B(\u_s[0] ), .Z(c_15__N_2423[7])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13796_2_lut.init = 16'h8888;
    LUT4 i13811_2_lut (.A(u_l[6]), .B(\u_s[1] ), .Z(c_15__N_2408[6])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13811_2_lut.init = 16'h8888;
    LUT4 i13797_2_lut (.A(u_l[7]), .B(\u_s[0] ), .Z(c_15__N_2423[6])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13797_2_lut.init = 16'h8888;
    LUT4 i13812_2_lut (.A(u_l[5]), .B(\u_s[1] ), .Z(c_15__N_2408[5])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(53[15:54])
    defparam i13812_2_lut.init = 16'h8888;
    LUT4 i13798_2_lut (.A(u_l[6]), .B(\u_s[0] ), .Z(c_15__N_2423[5])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i13798_2_lut.init = 16'h8888;
    FD1S3IX o_r__i17 (.D(o_r_17__N_2438[17]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_00[17] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i17.GSR = "DISABLED";
    FD1S3IX o_r__i16 (.D(o_r_17__N_2438[16]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_00[16] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i16.GSR = "DISABLED";
    FD1S3IX o_r__i15 (.D(o_r_17__N_2438[15]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_00[15] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i15.GSR = "DISABLED";
    FD1S3IX o_r__i14 (.D(o_r_17__N_2438[14]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_00[14] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i14.GSR = "DISABLED";
    FD1S3IX o_r__i13 (.D(o_r_17__N_2438[13]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_00[13] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i13.GSR = "DISABLED";
    FD1S3IX o_r__i12 (.D(o_r_17__N_2438[12]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_00[12] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i12.GSR = "DISABLED";
    FD1S3IX o_r__i11 (.D(o_r_17__N_2438[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_00[11] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i11.GSR = "DISABLED";
    FD1S3IX o_r__i10 (.D(o_r_17__N_2438[10]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_00[10] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i10.GSR = "DISABLED";
    FD1S3IX o_r__i9 (.D(o_r_17__N_2438[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_00[9] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i9.GSR = "DISABLED";
    FD1S3IX o_r__i8 (.D(o_r_17__N_2438[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_00[8] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i8.GSR = "DISABLED";
    FD1S3IX o_r__i7 (.D(o_r_17__N_2438[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_00[7] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i7.GSR = "DISABLED";
    FD1S3IX o_r__i6 (.D(o_r_17__N_2438[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_00[6] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i6.GSR = "DISABLED";
    FD1S3IX o_r__i5 (.D(o_r_17__N_2438[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_00[5] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i5.GSR = "DISABLED";
    FD1S3IX o_r__i4 (.D(o_r_17__N_2438[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_00[4] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i4.GSR = "DISABLED";
    FD1S3IX o_r__i3 (.D(o_r_17__N_2438[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_00[3] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i3.GSR = "DISABLED";
    FD1S3IX o_r__i2 (.D(o_r_17__N_2438[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_0_00[2] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i2.GSR = "DISABLED";
    FD1S3IX o_r__i1 (.D(o_r_17__N_2438[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\S_1_00_20__N_2184[1] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=27, LSE_LCOL=14, LSE_RCOL=73, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(57[9] 61[28])
    defparam o_r__i1.GSR = "DISABLED";
    LUT4 i12470_2_lut_rep_604 (.A(u_l[1]), .B(\u_s[0] ), .Z(n29264)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(54[6:45])
    defparam i12470_2_lut_rep_604.init = 16'h8888;
    LUT4 i12460_2_lut_rep_605 (.A(u_l[0]), .B(\u_s[1] ), .Z(n29265)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(51[18:45])
    defparam i12460_2_lut_rep_605.init = 16'h8888;
    LUT4 w_r_16__I_0_i2_2_lut_3_lut_4_lut (.A(u_l[0]), .B(\u_s[1] ), .C(\u_s[0] ), 
         .D(u_l[1]), .Z(o_r_17__N_2438[1])) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/bimpy.v(51[18:45])
    defparam w_r_16__I_0_i2_2_lut_3_lut_4_lut.init = 16'h7888;
    
endmodule
//
// Verilog Description of module dds_U26
//

module dds_U26 (dac_clk_p_c, i_sw0_c, carrier_increment, GND_net, dac_clk_p_c_enable_630, 
            o_sample_q, o_sample_i, \quarter_wave_sample_register_i[15] , 
            n32066) /* synthesis syn_module_defined=1 */ ;
    input dac_clk_p_c;
    input i_sw0_c;
    input [30:0]carrier_increment;
    input GND_net;
    input dac_clk_p_c_enable_630;
    output [15:0]o_sample_q;
    output [15:0]o_sample_i;
    output \quarter_wave_sample_register_i[15] ;
    input n32066;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[29:38])
    wire [15:0]o_sample_q_c /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(30[51:61])
    wire [15:0]o_sample_i_c /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(30[39:49])
    wire [30:0]increment;   // d:/documents/git_local/fm_modulator/rtl/dds.v(14[31:40])
    wire [11:0]o_phase;   // d:/documents/git_local/fm_modulator/rtl/dds.v(18[26:33])
    
    FD1S3DX increment_i0 (.D(carrier_increment[0]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[0])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=91, LSE_RLINE=91 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i0.GSR = "DISABLED";
    FD1S3DX increment_i30 (.D(carrier_increment[30]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(increment[30])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=91, LSE_RLINE=91 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i30.GSR = "DISABLED";
    FD1S3DX increment_i29 (.D(carrier_increment[29]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(increment[29])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=91, LSE_RLINE=91 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i29.GSR = "DISABLED";
    FD1S3DX increment_i28 (.D(carrier_increment[28]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(increment[28])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=91, LSE_RLINE=91 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i28.GSR = "DISABLED";
    FD1S3DX increment_i27 (.D(carrier_increment[27]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(increment[27])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=91, LSE_RLINE=91 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i27.GSR = "DISABLED";
    FD1S3DX increment_i26 (.D(carrier_increment[26]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(increment[26])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=91, LSE_RLINE=91 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i26.GSR = "DISABLED";
    FD1S3DX increment_i25 (.D(carrier_increment[25]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(increment[25])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=91, LSE_RLINE=91 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i25.GSR = "DISABLED";
    FD1S3DX increment_i24 (.D(carrier_increment[24]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(increment[24])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=91, LSE_RLINE=91 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i24.GSR = "DISABLED";
    FD1S3DX increment_i23 (.D(carrier_increment[23]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(increment[23])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=91, LSE_RLINE=91 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i23.GSR = "DISABLED";
    FD1S3DX increment_i22 (.D(carrier_increment[22]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(increment[22])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=91, LSE_RLINE=91 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i22.GSR = "DISABLED";
    FD1S3DX increment_i21 (.D(carrier_increment[21]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(increment[21])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=91, LSE_RLINE=91 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i21.GSR = "DISABLED";
    FD1S3DX increment_i20 (.D(carrier_increment[20]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(increment[20])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=91, LSE_RLINE=91 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i20.GSR = "DISABLED";
    FD1S3DX increment_i19 (.D(carrier_increment[19]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(increment[19])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=91, LSE_RLINE=91 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i19.GSR = "DISABLED";
    FD1S3DX increment_i18 (.D(carrier_increment[18]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(increment[18])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=91, LSE_RLINE=91 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i18.GSR = "DISABLED";
    FD1S3DX increment_i17 (.D(carrier_increment[17]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(increment[17])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=91, LSE_RLINE=91 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i17.GSR = "DISABLED";
    FD1S3DX increment_i16 (.D(carrier_increment[16]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(increment[16])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=91, LSE_RLINE=91 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i16.GSR = "DISABLED";
    FD1S3DX increment_i15 (.D(carrier_increment[15]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(increment[15])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=91, LSE_RLINE=91 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i15.GSR = "DISABLED";
    FD1S3DX increment_i14 (.D(carrier_increment[14]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(increment[14])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=91, LSE_RLINE=91 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i14.GSR = "DISABLED";
    FD1S3DX increment_i13 (.D(carrier_increment[13]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(increment[13])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=91, LSE_RLINE=91 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i13.GSR = "DISABLED";
    FD1S3DX increment_i12 (.D(carrier_increment[12]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(increment[12])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=91, LSE_RLINE=91 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i12.GSR = "DISABLED";
    FD1S3DX increment_i11 (.D(carrier_increment[11]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(increment[11])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=91, LSE_RLINE=91 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i11.GSR = "DISABLED";
    FD1S3DX increment_i10 (.D(carrier_increment[10]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(increment[10])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=91, LSE_RLINE=91 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i10.GSR = "DISABLED";
    FD1S3DX increment_i9 (.D(carrier_increment[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[9])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=91, LSE_RLINE=91 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i9.GSR = "DISABLED";
    FD1S3DX increment_i8 (.D(carrier_increment[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[8])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=91, LSE_RLINE=91 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i8.GSR = "DISABLED";
    FD1S3DX increment_i7 (.D(carrier_increment[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[7])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=91, LSE_RLINE=91 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i7.GSR = "DISABLED";
    FD1S3DX increment_i6 (.D(carrier_increment[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[6])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=91, LSE_RLINE=91 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i6.GSR = "DISABLED";
    FD1S3DX increment_i5 (.D(carrier_increment[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[5])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=91, LSE_RLINE=91 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i5.GSR = "DISABLED";
    FD1S3DX increment_i4 (.D(carrier_increment[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[4])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=91, LSE_RLINE=91 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i4.GSR = "DISABLED";
    FD1S3DX increment_i3 (.D(carrier_increment[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[3])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=91, LSE_RLINE=91 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i3.GSR = "DISABLED";
    FD1S3DX increment_i2 (.D(carrier_increment[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[2])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=91, LSE_RLINE=91 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i2.GSR = "DISABLED";
    FD1S3DX increment_i1 (.D(carrier_increment[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(increment[1])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=91, LSE_RLINE=91 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i1.GSR = "DISABLED";
    quarter_wave_sine_lookup_U22 qtr_inst (.GND_net(GND_net), .dac_clk_p_c(dac_clk_p_c), 
            .dac_clk_p_c_enable_630(dac_clk_p_c_enable_630), .o_phase({o_phase}), 
            .o_sample_q({o_sample_q}), .i_sw0_c(i_sw0_c), .o_sample_i({o_sample_i}), 
            .\quarter_wave_sample_register_i[15] (\quarter_wave_sample_register_i[15] ), 
            .n32066(n32066)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(21[70:134])
    \nco(OW=12)_U23  nco_inst (.o_phase({o_phase}), .dac_clk_p_c(dac_clk_p_c), 
            .i_sw0_c(i_sw0_c), .increment({increment}), .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(20[49:100])
    
endmodule
//
// Verilog Description of module quarter_wave_sine_lookup_U22
//

module quarter_wave_sine_lookup_U22 (GND_net, dac_clk_p_c, dac_clk_p_c_enable_630, 
            o_phase, o_sample_q, i_sw0_c, o_sample_i, \quarter_wave_sample_register_i[15] , 
            n32066) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input dac_clk_p_c;
    input dac_clk_p_c_enable_630;
    input [11:0]o_phase;
    output [15:0]o_sample_q;
    input i_sw0_c;
    output [15:0]o_sample_i;
    output \quarter_wave_sample_register_i[15] ;
    input n32066;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[29:38])
    wire [15:0]o_sample_q_c /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(30[51:61])
    wire [15:0]\o_val_pipeline_q[0]  /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(16[24:40])
    wire [15:0]o_sample_i_c /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(30[39:49])
    wire [15:0]\o_val_pipeline_i[0]  /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(15[24:40])
    
    wire n27193, n25146;
    wire [9:0]index_i;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(31[17:24])
    
    wire n27194, n27192, n27191;
    wire [9:0]index_q;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(31[26:33])
    
    wire n101, n19707;
    wire [15:0]quarter_wave_sample_register_q;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(22[56:86])
    wire [15:0]o_val_pipeline_q_0__15__N_1831;
    
    wire n19708, n29392, n325, n32029, n23071, n27189, n27186, 
        n27190, n29406, n32019, n27188, n27187, n797, n828, n24956, 
        n24944, n24945, n24960, n24946, n24947, n24961, n24948, 
        n24949, n24962, n24950, n24951, n24963, n27185, n27184, 
        n24952, n24953, n24964, n19706, n24958, n24959, n24967, 
        n23242, n23204, n24991, n24992, n24999;
    wire [11:0]phase_i;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(11[17:24])
    
    wire n24997, n24998, n25002, n29371, n25022, n25023, n25030, 
        n29512, n29513, n29514, n25028, n25029, n25033, n25058, 
        n25059, n25074, n25060, n25061, n25075, n23218, n23219, 
        n23220, n25062, n25063, n25076, n25064, n25065, n25077, 
        n25066, n25067, n25078, n25068, n25069, n25079, n318, 
        n381, n23284, n29581, n29389, n763, n23221, n23222, n23223;
    wire [1:0]phase_negation_i;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(23[12:28])
    wire [1:0]phase_negation_q;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(23[30:46])
    wire [11:0]phase_q;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(12[17:24])
    wire [9:0]index_i_9__N_1748;
    wire [9:0]index_q_9__N_1758;
    wire [14:0]quarter_wave_sample_register_q_15__N_1783;
    wire [15:0]quarter_wave_sample_register_i;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(22[24:54])
    wire [14:0]quarter_wave_sample_register_i_15__N_1768;
    
    wire n318_adj_2938, n381_adj_2939, n23266, n23125, n23126, n476, 
        n28141, n62, n23105, n29509, n29510, n29511, n13548, n13549, 
        n24318, n13335, n28139, n526, n29167, n13556, n13557, 
        n24310, n13394, n29393, n23131, n19705;
    wire [15:0]o_val_pipeline_i_0__15__N_1799;
    
    wire n19704, n27072, n29459, n19703, n29394, n23227, n23228, 
        n23229, n29506, n29507, n29508, n716, n25163, n25164, 
        n25167, n173, n221, n252, n24334, n25165, n25166, n25168, 
        n23974, n29041, n23396, n23230, n23231, n23232, n28659, 
        n572, n954, n19702, n29079, n23236, n23237, n23238, n285, 
        n29386, n20016, n29503, n29504, n29505, n348, n349, n23243, 
        n23244, n46, n158, n189, n24364, n24801, n24802, n24805, 
        n557, n24803, n24804, n24806, n19701, n19700, n526_adj_2940, 
        n541, n25313, n24808, n24809, n24812, n25199, n25200, 
        n25211, n25201, n25202, n25212, n32018, n851, n23615, 
        n25203, n25204, n25213, n24810, n24811, n24813, n25205, 
        n25206, n25214, n13382, n23325, n25223, n29054, n285_adj_2941, 
        n23331, n23334, n25225, n574, n23337, n25226, n23340, 
        n764, n25227, n93, n94, n25237, n25238, n25241, n25239, 
        n25240, n25242, n890, n13357, n29335, n173_adj_2942, n844, 
        n13320, n25260, n25261, n25268, n32034, n620, n25262, 
        n25263, n25269, n404, n23966, n25264, n25265, n25270, 
        n882, n25266, n25267, n25271, n29181, n20015, n13317, 
        n29423, n173_adj_2943, n635, n27538, n23401, n28140, n747, 
        n29095, n29395, n25290, n25291, n25302, n25292, n25293, 
        n25303, n25294, n25295, n25304, n25296, n25297, n25305, 
        n27389, n23134, n444, n25329, n25330, n25337, n25331, 
        n25332, n25338, n25333, n25334, n25339, n29326, n892, 
        n23150, n25335, n25336, n25340, n731, n796, n27071, n491, 
        n29460, n32054, n29070, n251, n25089, n348_adj_2944, n109, 
        n1017, n716_adj_2945, n716_adj_2946, n32036, n23423, n29147, 
        n29086, n29499, n29500, n29501, n27460, n908, n23207, 
        n27462, n460, n316, n29148, n29064, n812, n62_adj_2947, 
        n29376, n731_adj_2948, n32022, n23930, n931, n29429, n23068, 
        n13328, n13331, n875, n13565, n29370, n29396, n23390, 
        n762, n252_adj_2949, n812_adj_2950, n443, n604, n428, n443_adj_2951, 
        n23393, n29518, n32039, n23174, n29405, n29447, n20013, 
        n27073, n29372, n29063, n251_adj_2952, n29441, n20012, n15, 
        n844_adj_2953, n24815, n24816, n24819, n588, n23932, n23216, 
        n956, n22180, n24730, n109_adj_2954, n25092, n251_adj_2955, 
        n460_adj_2956, n23111, n25090, n13554, n526_adj_2957, n23613, 
        n173_adj_2958, n190, n491_adj_2959, n507, n29058, n379, 
        n32035, n908_adj_2960, n23387, n109_adj_2961, n27619, n24738, 
        n24739, n24742, n443_adj_2962, n24740, n24741, n24743, n25091, 
        n557_adj_2963, n428_adj_2964, n716_adj_2965, n732, n24303, 
        n764_adj_2966, n29354, n29390, n26642, n24745, n24746, n24749, 
        n109_adj_2967, n460_adj_2968, n443_adj_2969, n24747, n24748, 
        n24750, n379_adj_2970, n542, n13528, n574_adj_2971, n19699, 
        n23180, n19698, n29176, n445, n900, n684, n32025, n26726, 
        n325_adj_2972, n890_adj_2973, n684_adj_2974, n32056, n348_adj_2975, 
        n29437, n23918, n29301, n29436, n491_adj_2976, n29519, n29180, 
        n475, n604_adj_2977, n29204, n445_adj_2978, n29357, n26646, 
        n890_adj_2979, n412, n29388, n26649, n684_adj_2980, n23422, 
        n699, n699_adj_2981, n29356, n29353, n19982, n23921, n716_adj_2982, 
        n19981, n29521, n29402, n29433, n26718, n668, n890_adj_2983, 
        n747_adj_2984, n763_adj_2985, n27373, n29385, n1001, n27372, 
        n412_adj_2986, n29520, n29475, n653, n23198, n23351, n29177, 
        n29146, n317, n32020, n301, n32021, n29391, n29387, n26652, 
        n29470, n475_adj_2987, n25072, n28680, n25081, n747_adj_2988, 
        n844_adj_2989, n860, n29355, n32033, n26655, n645, n23612, 
        n23353, n221_adj_2990, n28839, n46_adj_2991, n29168, n29903, 
        n23999, n204, n29901, n29900, n29400, n29439, n908_adj_2992, 
        n29523, n31, n23976, n24331, n23318, n348_adj_2993, n349_adj_2994, 
        n716_adj_2995, n29446, n23117, n26659, n157, n26660, n94_adj_2996, 
        n125, n24332, n27400, n23116, n23118, n29336, n653_adj_2997, 
        n29465, n29461, n731_adj_2998, n844_adj_2999, n860_adj_3000, 
        n23867, n23420, n620_adj_3001, n29315, n20003, n16258, n24333, 
        n24817, n24818, n24820, n23985, n23988, n24335, n23991, 
        n23994, n24336, n413, n444_adj_3002, n24337, n29432, n27414, 
        n589, n23203, n29316, n731_adj_3003, n27416, n29578, n23201, 
        n23202, n29585, n29586, n29587, n29444, n23114, n29418, 
        n635_adj_3004, n23885, n526_adj_3005, n189_adj_3006, n508, 
        n476_adj_3007, n507_adj_3008, n24338, n29361, n29133, n16858, 
        n475_adj_3009, n619, n27466, n27483, n29379, n23135, n23900, 
        n684_adj_3010, n29088, n28360, n29026, n475_adj_3011, n23954, 
        n29377, n653_adj_3012, n29424, n28281, n29028, n20017, n573, 
        n24339, n23902, n604_adj_3013, n605, n636, n24340, n23997, 
        n700, n24341, n29367, n557_adj_3014, n573_adj_3015, n125_adj_3016, 
        n24004, n29438, n27511, n732_adj_3017, n24000, n24342, n797_adj_3018, 
        n828_adj_3019, n24343, n124, n28488, n573_adj_3020, n573_adj_3021, 
        n860_adj_3022, n891, n24344, n812_adj_3023, n25322, n30203, 
        n23362, n30204, n29067, n29066, n25229, n23197, n23199, 
        n24780, n24781, n24784, n29136, n29068, n24782, n24783, 
        n24785, n29330, n460_adj_3024, n285_adj_3025, n29384, n23611, 
        n23381, n23072, n29329, n16898, n875_adj_3026, n25324, n29420, 
        n285_adj_3027, n23993, n364, n460_adj_3028, n29324, n700_adj_3029, 
        n27572, n23195, n29178, n25172, n29165, n23338, n94_adj_3030, 
        n24003, n24363, n23192, n23191, n908_adj_3031, n923, n25325, 
        n28340, n16900, n124_adj_3032, n875_adj_3033, n890_adj_3034, 
        n891_adj_3035, n189_adj_3036, n29467, n29331, n27586, n508_adj_3037, 
        n23110, n23112, n29369, n254, n14983, n828_adj_3038, n653_adj_3039, 
        n797_adj_3040, n221_adj_3041, n252_adj_3042, n24365, n29309, 
        n22131, n285_adj_3043, n124_adj_3044, n28534, n573_adj_3045, 
        n573_adj_3046, n653_adj_3047, n668_adj_3048, n669, n286, n24006, 
        n24366, n125_adj_3049, n573_adj_3050, n859, n24009, n24367, 
        n32023, n124_adj_3051, n94_adj_3052, n15_adj_3053, n29486, 
        n24975, n29463, n32055, n668_adj_3054, n29034, n29477, n16844, 
        n364_adj_3055, n29373, n30466, n30467, n29080, n574_adj_3056, 
        n23215, n23217, n23728, n23729, n23730, n29464, n23189, 
        n812_adj_3057, n541_adj_3058, n542_adj_3059, n29404, n26721, 
        n669_adj_3060, n700_adj_3061, n24372, n23212, n762_adj_3062, 
        n29534, n379_adj_3063, n85, n23188, n23190, n23186, n332, 
        n23185, n23102, n23101, n251_adj_3064, n12265, n252_adj_3065, 
        n23103, n28840, n25285, n30579, n30580, n30581, n506, 
        n985, n986, n29382, n971, n29403, n29440, n26725, n30578, 
        n29100, n30577, n30582, n32024, n30583, n30584, n23064, 
        n24373, n29185, n939, n23147, n29334, n29360, n444_adj_3066, 
        n29409, n923_adj_3067, n23416, n747_adj_3068, n23070, n828_adj_3069, 
        n24374, n251_adj_3070, n301_adj_3071, n890_adj_3072, n891_adj_3073, 
        n29351, n26639, n812_adj_3074, n15114, n828_adj_3075, n781, 
        n29039, n797_adj_3076, n26728, n860_adj_3077, n23076, n24375, 
        n29533, n29471, n27747, n30637, n30638, n30636, n30635, 
        n653_adj_3078, n668_adj_3079, n669_adj_3080, n30639, n30640, 
        n30641, n30642, n668_adj_3081, n763_adj_3082, n29430, n29445, 
        n716_adj_3083, n541_adj_3084, n542_adj_3085, n29036, n701, 
        n27756, n12338, n252_adj_3086, n24807, n28803, n25194, n32028, 
        n653_adj_3087, n31750, n25243, n27760, n125_adj_3088, n24394, 
        n29442, n620_adj_3089, n23959, n589_adj_3090, n23090, n541_adj_3091, 
        n526_adj_3092, n158_adj_3093, n189_adj_3094, n24395, n29038, 
        n701_adj_3095, n27781, n491_adj_3096, n507_adj_3097, n860_adj_3098, 
        n31713, n25169, n27785, n443_adj_3099, n684_adj_3100, n700_adj_3101, 
        n221_adj_3102, n252_adj_3103, n24396, n27805, n21714, n1018, 
        n653_adj_3104, n29374, n254_adj_3105, n286_adj_3106, n23088, 
        n24397, n29559, n27806, n27811, n286_adj_3107, n349_adj_3108, 
        n23097, n24398, n413_adj_3109, n444_adj_3110, n24399, n29166, 
        n637, n24814, n476_adj_3111, n507_adj_3112, n24400, n16828, 
        n28143, n29029, n23106, n24401, n15_adj_3113, n24823, n27836, 
        n29346, n348_adj_3114, n13369, n24402, n29553, n27837, n27842, 
        n24822, n24826, n108, n29375, n173_adj_3115, n620_adj_3116, 
        n669_adj_3117, n700_adj_3118, n24403, n638, n23316, n27860, 
        n23115, n763_adj_3119, n24404, n498, n23984, n860_adj_3120, 
        n891_adj_3121, n24406, n23099, n24824, n24825, n24827, n382, 
        n509, n27862, n23098, n23100, n26741, n924, n24407, n23121, 
        n1018_adj_3122, n24408, n890_adj_3123, n23074, n26744, n28082, 
        n29032, n24821, n29127, n61, n62_adj_3124, n15_adj_3125, 
        n29190, n31_adj_3126, n158_adj_3127, n24426, n142, n221_adj_3128, 
        n23136, n24427, n23310, n27863, n29537, n23398, n24380, 
        n24381, n27878, n286_adj_3129, n317_adj_3130, n24428, n21712, 
        n29040, n24382, n24383, n27876, n23356, n397, n24379, 
        n24378, n27879, n28285, n349_adj_3131, n23139, n24429, n638_adj_3132, 
        n23298, n27897, n413_adj_3133, n23142, n24430, n30, n28491, 
        n382_adj_3134, n509_adj_3135, n27899, n13386, n29904, n30_adj_3136, 
        n31_adj_3137, n23145, n507_adj_3138, n24431, n939_adj_3139, 
        n954_adj_3140, n25326, n16860, n252_adj_3141, n13403, n13404, 
        n13444, n13445, n23809, n23810, n23811, n475_adj_3142, n24847, 
        n23148, n24432, n23292, n27900, n28284, n572_adj_3143, n29579, 
        n29580, n364_adj_3144, n605_adj_3145, n23151, n24433, n24894, 
        n24893, n27924, n24892, n24891, n27925, n62_adj_3146, n22572, 
        n13385, n24895, n24896, n27922, n23335, n23143, n955, 
        n669_adj_3147, n700_adj_3148, n24434, n23096, n16668, n23095, 
        n605_adj_3149, n29089, n574_adj_3150, n24828, n732_adj_3151, 
        n763_adj_3152, n24435, n29049, n29536, n25277, n23917, n860_adj_3153, 
        n23960, n29130, n189_adj_3154, n25144, n26651, n25196, n27977, 
        n971_adj_3155, n986_adj_3156, n25327, n1002, n25197, n26657, 
        n27976, n26645, n25192, n27979, n828_adj_3157, n93_adj_3158, 
        n29540, n491_adj_3159, n25143, n908_adj_3160, n716_adj_3161, 
        n732_adj_3162, n27575, n16798, n28079, n29031, n29078, n638_adj_3163, 
        n29407, n25137, n653_adj_3164, n475_adj_3165, n669_adj_3166, 
        n1017_adj_3167, n25328, n660, n25136, n142_adj_3168, n605_adj_3169, 
        n29134, n221_adj_3170, n23405, n23919, n25135, n23372, n23373, 
        n29443, n25134, n23368, n23369, n23370, n507_adj_3171, n23953, 
        n29408, n27386, n859_adj_3172, n443_adj_3173, n21706, n21704, 
        n28073, n157_adj_3174, n29571, n24889, n542_adj_3175, n24883, 
        n860_adj_3176, n891_adj_3177, n24437, n29574, n24881, n491_adj_3178, 
        n732_adj_3179, n29539, n924_adj_3180, n28075, n28076, n29161, 
        n23239, n29042, n316_adj_3181, n285_adj_3182, n28100, n28103, 
        n28102, n28104, n317_adj_3183, n397_adj_3184, n413_adj_3185, 
        n731_adj_3186, n732_adj_3187, n684_adj_3188, n700_adj_3189, 
        n24976, n93_adj_3190, n24977, n23267, n1021, n316_adj_3191, 
        n317_adj_3192, n270, n653_adj_3193, n286_adj_3194, n27418, 
        n28106, n23920, n23922, n29522, n28107, n491_adj_3195, n732_adj_3196, 
        n188, n23073, n29179, n16610, n27387, n29380, n27391, 
        n23816, n23817, n22201, n21709, n24458, n732_adj_3197, n28108, 
        n28109, n28110, n28111, n511, n364_adj_3198, n28074, n29173, 
        n29143, n29047, n27467, n24376, n23926, n23927, n23928, 
        n542_adj_3199, n24370, n444_adj_3200, n24368, n31_adj_3201, 
        n62_adj_3202, n142_adj_3203, n28344, n32031, n796_adj_3204, 
        n23929, n23931, n29099, n28170, n890_adj_3205, n924_adj_3206, 
        n28172, n28173, n23140, n684_adj_3207, n700_adj_3208, n23092, 
        n23093, n23094, n15165, n158_adj_3209, n30_adj_3210, n28537, 
        n27539, n23912, n23913, n29365, n21737, n24719, n13387, 
        n892_adj_3211, n25228, n29250, n22031, n28364, n13529, n475_adj_3212, 
        n572_adj_3213, n22576, n28363, n23884, n29053, n23933, n23934, 
        n23962, n28664, n25071, n25080, n29101, n124_adj_3214, n23935, 
        n23936, n23937, n1002_adj_3215, n29549, n29087, n638_adj_3216, 
        n23428, n23429, n23430, n23206, n25099, n25098, n23285, 
        n27465, n25096, n333, n13530, n892_adj_3217, n24835, n23425, 
        n29548, n23426, n23427, n236, n25013, n29102, n1021_adj_3218, 
        n25342, n25341, n25309, n25288, n26746, n25301, n26730, 
        n25287, n25300, n26724, n25283, n25298, n25273, n25272, 
        n25224, n25231, n25222, n25230, n158_adj_3219, n189_adj_3220, 
        n24877, n94_adj_3221, n125_adj_3222, n24845, n25232, n25233, 
        n25235, n25218, n20006, n16248, n24846, n29552, n27757, 
        n27758, n29551, n25032, n25035, n25031, n25034, n25001, 
        n25004, n25000, n25003, n24897, n24898, n24902, n24464, 
        n24465, n24471, n31_adj_3223, n62_adj_3224, n24875, n24462, 
        n24463, n24470, n26753, n157_adj_3225, n26754, n24831, n24832, 
        n24838, n24829, n24830, n24837, n24839, n24840, n24842, 
        n29251, n22033, n24384, n24385, n24389, n511_adj_3226, n16882, 
        n766, n27195, n24726, n24732, n24723, n24724, n24731, 
        n23866, n23868, n31711, n252_adj_3227, n31708, n62_adj_3228, 
        n31710, n16930, n766_adj_3229, n25234, n956_adj_3230, n22170, 
        n24469, n15_adj_3231, n30_adj_3232, n25006, n23417, n25084, 
        n25085, n25087, n25082, n25083, n25086, n31747, n24866, 
        n28174, n24871, n24864, n24865, n24870, n24873, n252_adj_3233, 
        n31745, n31748, n24841, n23967, n23970, n24848, n24450, 
        n24453, n24448, n24449, n24452, n23869, n23870, n23871, 
        n1022, n1022_adj_3234, n28148, n23286, n23248, n23995, n24353, 
        n28077, n24358, n24351, n24352, n24357, n24360, n29558, 
        n731_adj_3235, n28084, n23268, n23209, n24970, n24971, n24973, 
        n24968, n24969, n24972, n24534, n24535, n24537, n24532, 
        n24533, n24536, n24868, n24869, n24872, n24503, n24504, 
        n24506, n24501, n24502, n24505, n24419, n24420, n24422, 
        n24417, n24418, n24421, n29575, n29576, n29577, n637_adj_3236, 
        n23287, n23213, n24355, n24356, n24359, n23973, n24849, 
        n23269, n29557, n413_adj_3237, n24850, n285_adj_3238, n23963, 
        n23964, n557_adj_3239, n699_adj_3240, n23419, n23957, n413_adj_3241, 
        n348_adj_3242, n26901, n26899, n26902, n23399, n491_adj_3243, 
        n29132, n28442, n476_adj_3244, n28443, n23878, n23879, n23880, 
        n23965, n94_adj_3245, n24478, n316_adj_3246, n27559, n23205, 
        n23208, n24479, n13553, n526_adj_3247, n157_adj_3248, n828_adj_3249, 
        n1002_adj_3250, n29541, n28444, n28447, n26900, n732_adj_3251, 
        n526_adj_3252, n27390, n23968, n23969, n23089, n476_adj_3253, 
        n507_adj_3254, n24851, n28502, n635_adj_3255, n23971, n23972, 
        n24311, n27573, n29479, n27557, n23881, n23882, n23883, 
        n29057, n747_adj_3256, n23404, n26898, n15110, n141, n124_adj_3257, 
        n23155, n23156, n23157, n29472, n29478, n716_adj_3258, n23886, 
        n30_adj_3259, n23384, n526_adj_3260, n27748, n620_adj_3261, 
        n93_adj_3262, n23173, n23956, n762_adj_3263, n29476, n716_adj_3264, 
        n28501, n28504, n23214, n24481, n23983, n23413, n29317, 
        n13422, n28171, n29045, n19977, n573_adj_3265, n24852, n860_adj_3266, 
        n28575, n23887, n23888, n23889, n28578, n28146, n955_adj_3267, 
        n23080, n93_adj_3268, n25008, n636_adj_3269, n15097, n23893, 
        n23894, n23895, n46_adj_3270, n25007, n220, n25012, n23896, 
        n23897, n23898, n23899, n23901, n23980, n29502, n23982, 
        n28343, n747_adj_3271, n29333, n28662, n924_adj_3272, n27782, 
        n27783, n890_adj_3273, n891_adj_3274, n23903, n23904, n23986, 
        n23987, n23402, n349_adj_3275, n24482, n24483, n24484, n605_adj_3276, 
        n636_adj_3277, n24853, n93_adj_3278, n15_adj_3279, n29435, 
        n669_adj_3280, n29427, n124_adj_3281, n985_adj_3282, n23082, 
        n700_adj_3283, n24854, n875_adj_3284, n890_adj_3285, n891_adj_3286, 
        n732_adj_3287, n23091, n24855, n397_adj_3288, n797_adj_3289, 
        n24856, n13432, n28676, n23905, n23906, n23907, n859_adj_3290, 
        n860_adj_3291, n23908, n23909, n23910, n28678, n506_adj_3292, 
        n636_adj_3293, n24486, n188_adj_3294, n23241, n24487, n23158, 
        n23159, n23160, n23958, n860_adj_3295, n891_adj_3296, n24857, 
        n476_adj_3297, n23395, n397_adj_3298, n29281, n413_adj_3299, 
        n29481, n16645, n286_adj_3300, n24489, n924_adj_3301, n23940, 
        n24491, n158_adj_3302, n29572, n29573, n125_adj_3303, n397_adj_3304, 
        n23392, n23394, n859_adj_3305, n987, n23943, n24492, n875_adj_3306, 
        n29483, n301_adj_3307, n31_adj_3308, n908_adj_3309, n317_adj_3310, 
        n30_adj_3311, n29516, n23317, n23319, n29482, n94_adj_3312, 
        n24876, n187, n188_adj_3313, n94_adj_3314, n23382, n24509, 
        n270_adj_3315, n762_adj_3316, n23320, n23321, n23322, n25009, 
        n747_adj_3317, n763_adj_3318, n29426, n900_adj_3319, n23383, 
        n221_adj_3320, n252_adj_3321, n24878, n668_adj_3322, n23989, 
        n23990, n684_adj_3323, n23992, n286_adj_3324, n24879, n349_adj_3325, 
        n24880, n23385, n23388, n24510, n23998, n23391, n24512, 
        n27620, n124_adj_3326, n24978, n23087, n23086, n23350, n349_adj_3327, 
        n24513, n23397, n23400, n24514, n397_adj_3328, n23347, n23374, 
        n23403, n23406, n24515, n23375, n23376, n348_adj_3329, n23345, 
        n23344, n23342, n333_adj_3330, n23341, n23168, n23329, n23330, 
        n23167, n23169, n29569, n29570, n15092, n348_adj_3331, n669_adj_3332, 
        n700_adj_3333, n24885, n23164, n316_adj_3334, n412_adj_3335, 
        n924_adj_3336, n23175, n24890, n29431, n908_adj_3337, n506_adj_3338, 
        n15_adj_3339, n860_adj_3340, n23133, n24886, n731_adj_3341, 
        n23165, n23166, n23412, n24517, n23415, n700_adj_3342, n24518, 
        n270_adj_3343, n316_adj_3344, n23332, n23333, n491_adj_3345, 
        n506_adj_3346, n397_adj_3347, n23414, n23132, n23418, n23421, 
        n24520, n684_adj_3348, n828_adj_3349, n24887, n16626, n29480, 
        n24884, n24888, n24008, n24007, n635_adj_3350, n23336, n24005, 
        n24522, n987_adj_3351, n24523, n23389, n23339, n24001, n24002, 
        n23343, n23346, n23348, n23349, n24093, n13389, n890_adj_3352, 
        n891_adj_3353, n24882, n94_adj_3354, n460_adj_3355, n23352, 
        n270_adj_3356, n15_adj_3357, n23354, n23355, n29422, n93_adj_3358, 
        n13436, n763_adj_3359, n859_adj_3360, n61_adj_3361, n29283, 
        n23363, n23364, n23360, n142_adj_3362, n157_adj_3363, n25010, 
        n29484, n28802, n23359, n23361, n23386, n25011, n23357, 
        n23358, n25097, n142_adj_3364, n157_adj_3365, n24979, n29419, 
        n205, n62_adj_3366, n891_adj_3367, n892_adj_3368, n875_adj_3369, 
        n859_adj_3370, n491_adj_3371, n507_adj_3372, n23410, n23240, 
        n23977, n16744, n93_adj_3373, n173_adj_3374, n23952, n24844, 
        n23081, n333_adj_3375, n25016, n157_adj_3376, n29112, n444_adj_3377, 
        n25017, n882_adj_3378, n890_adj_3379, n29311, n891_adj_3380, 
        n29285, n25018, n541_adj_3381, n25019, n28675, n526_adj_3382, 
        n397_adj_3383, n25020, n397_adj_3384, n348_adj_3385, n491_adj_3386, 
        n12581, n25021, n349_adj_3387, n23949, n635_adj_3388, n16249, 
        n636_adj_3389, n19975, n19976, n348_adj_3390, n24980, n28679, 
        n28677, n23978, n23979, n491_adj_3391, n23975, n23063, n460_adj_3392, 
        n475_adj_3393, n23961, n506_adj_3394, n93_adj_3395, n28663, 
        n28660, n700_adj_3396, n24954, n29352, n28661, n986_adj_3397, 
        n24955, n24957, n763_adj_3398, n205_adj_3399, n23872, n23874, 
        n348_adj_3400, n23955, n23951, n23950, n16637, n23948, n986_adj_3401, 
        n29368, n29059, n23947, n23945, n413_adj_3402, n142_adj_3403, 
        n20004, n20005, n23941, n62_adj_3404, n23942, n812_adj_3405, 
        n684_adj_3406, n28577, n28576, n796_adj_3407, n797_adj_3408, 
        n16591, n23938, n23939, n24296, n13566, n13520, n28538, 
        n28536, n28535, n684_adj_3409, n844_adj_3410, n23075, n23411, 
        n29538, n253, n28503, n190_adj_3411, n28492, n28490, n62_adj_3412, 
        n572_adj_3413, n573_adj_3414, n28489, n29434, n605_adj_3415, 
        n620_adj_3416, n16308, n924_adj_3417, n27486, n891_adj_3418, 
        n892_adj_3419, n29276, n731_adj_3420, n24091, n29318, n348_adj_3421, 
        n28448, n542_adj_3422, n491_adj_3423, n653_adj_3424, n11112, 
        n13373, n684_adj_3425, n205_adj_3426, n142_adj_3427, n604_adj_3428, 
        n23210, n142_adj_3429, n572_adj_3430, n23249, n23144, n25036, 
        n25274, n25005, n25343, n31749, n31746, n24985, n24986, 
        n24996, n24987, n24988, n954_adj_3431, n25093, n24989, n24990, 
        n31712, n31709, n25306, n25307, n25310, n25094, n26755, 
        n28365, n24735, n23119, n24733, n24734, n24736, n24415, 
        n24416, n28345, n28342, n27413, n23149, n24413, n24414, 
        n24474, n24472, n24473, n24475, n24499, n24500, n24530, 
        n24531, n24493, n24494, n27488, n24497, n24498, n27513, 
        n24966, n24524, n24525, n27577, n25024, n25025, n24528, 
        n24529, n27588, n26752, n781_adj_3432, n25321, n23104, n28341, 
        n24965, n23424, n397_adj_3433, n29322, n25299, n9850, n24727, 
        n24728, n24729, n24347, n24348, n24349, n24350, n24405, 
        n24409, n24410, n24411, n24412, n747_adj_3434, n24833, n24834, 
        n286_adj_3435, n24442, n24443, n24441, n24444, n24445, n25027, 
        n24836, n25100, n28286, n25101, n29517, n1002_adj_3436, 
        n24377, n26722, n924_adj_3437, n221_adj_3438, n12256, n23069, 
        n27464, n25095, n24466, n24467, n24468, n29074, n29069, 
        n668_adj_3439, n24488, n24490, n24860, n24861, n24862, n24863, 
        n24495, n24496, n24519, n27537, n24521, n24526, n24527, 
        n23996, n24993, n29906, n27750, n28105, n23062, n27561, 
        n25217, n25308, n25102, n25140, n30_adj_3440, n28147, n635_adj_3441, 
        n317_adj_3442, n93_adj_3443, n24362, n24369, n24371, n27388, 
        n24393, n16259, n26745, n26742, n20002, n924_adj_3444, n924_adj_3445, 
        n29319, n24477, n699_adj_3446, n109_adj_3447, n875_adj_3448, 
        n28101, n28083, n24508, n26658, n23179, n25138, n635_adj_3449, 
        n25139, n668_adj_3450, n20001, n26640, n572_adj_3451, n573_adj_3452, 
        n27980, n27978, n27981, n25208, n23176, n23177, n23178, 
        n29145, n157_adj_3453, n29186, n844_adj_3454, n27926, n27923, 
        n27745, n27901, n27898, n62_adj_3455, n475_adj_3456, n364_adj_3457, 
        n27880, n27877, n27864, n27861, n23181, n25311;
    wire [15:0]n670;
    
    wire n254_adj_3458, n29515, n475_adj_3459, n25220, n254_adj_3460, 
        n25244, n557_adj_3461, n25245;
    wire [15:0]n671;
    
    wire n25246, n635_adj_3462, n25247, n27484, n25248, n491_adj_3463;
    wire [11:0]phase_q_11__N_1874;
    
    wire n23187, n19983, n25249, n23193, n27583, n25250, n27749, 
        n27746, n26729, n26727, n762_adj_3464, n25251, n781_adj_3465, 
        n796_adj_3466, n25252, n812_adj_3467, n25253, n22328, n25255, 
        n25256, n954_adj_3468, n25257, n25258, n25254, n25259, n26723, 
        n26720, n20014, n27585, n26719, n636_adj_3469, n22332, n19713, 
        n26647, n27587, n27584, n23141, n27576, n27574, n19712, 
        n19711, n19710, n27560, n27558, n19709, n27512, n27509, 
        n27510, n27508, n25314, n27487, n27485, n23113, n27463, 
        n27461, n23137, n27417, n27415, n25315, n25316, n25317, 
        n25318, n25319, n25320, n25323, n23138, n26661, n29902, 
        n29905, n26656, n26653, n26650, n26648, n26644, n26641;
    
    L6MUX21 i25486 (.D0(n27193), .D1(n25146), .SD(index_i[5]), .Z(n27194));
    PFUMX i25484 (.BLUT(n27192), .ALUT(n27191), .C0(index_i[4]), .Z(n27193));
    LUT4 mux_207_Mux_8_i101_3_lut_3_lut_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n101)) /* synthesis lut_function=(!(A (B (C))+!A (B (C)+!B !(C)))) */ ;
    defparam mux_207_Mux_8_i101_3_lut_3_lut_3_lut.init = 16'h3e3e;
    CCU2D unary_minus_27_add_3_5 (.A0(quarter_wave_sample_register_q[3]), 
          .B0(GND_net), .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_q[4]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19707), .COUT(n19708), 
          .S0(o_val_pipeline_q_0__15__N_1831[3]), .S1(o_val_pipeline_q_0__15__N_1831[4]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(81[29:60])
    defparam unary_minus_27_add_3_5.INIT0 = 16'hf555;
    defparam unary_minus_27_add_3_5.INIT1 = 16'hf555;
    defparam unary_minus_27_add_3_5.INJECT1_0 = "NO";
    defparam unary_minus_27_add_3_5.INJECT1_1 = "NO";
    LUT4 mux_207_Mux_6_i134_3_lut_4_lut_3_lut_rep_732 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29392)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_6_i134_3_lut_4_lut_3_lut_rep_732.init = 16'h9696;
    LUT4 i20589_3_lut (.A(n325), .B(n32029), .C(index_q[3]), .Z(n23071)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20589_3_lut.init = 16'hcaca;
    L6MUX21 i25481 (.D0(n27189), .D1(n27186), .SD(index_i[4]), .Z(n27190));
    LUT4 n459_bdd_3_lut (.A(n29406), .B(n32019), .C(index_i[3]), .Z(n27192)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n459_bdd_3_lut.init = 16'hcaca;
    PFUMX i25479 (.BLUT(n27188), .ALUT(n27187), .C0(index_i[3]), .Z(n27189));
    PFUMX i22455 (.BLUT(n797), .ALUT(n828), .C0(index_q[5]), .Z(n24956));
    L6MUX21 i22459 (.D0(n24944), .D1(n24945), .SD(index_q[6]), .Z(n24960));
    L6MUX21 i22460 (.D0(n24946), .D1(n24947), .SD(index_q[6]), .Z(n24961));
    L6MUX21 i22461 (.D0(n24948), .D1(n24949), .SD(index_q[6]), .Z(n24962));
    L6MUX21 i22462 (.D0(n24950), .D1(n24951), .SD(index_q[6]), .Z(n24963));
    PFUMX i25477 (.BLUT(n27185), .ALUT(n27184), .C0(index_i[5]), .Z(n27186));
    L6MUX21 i22463 (.D0(n24952), .D1(n24953), .SD(index_q[6]), .Z(n24964));
    CCU2D unary_minus_27_add_3_3 (.A0(quarter_wave_sample_register_q[1]), 
          .B0(GND_net), .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_q[2]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19706), .COUT(n19707), 
          .S0(o_val_pipeline_q_0__15__N_1831[1]), .S1(o_val_pipeline_q_0__15__N_1831[2]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(81[29:60])
    defparam unary_minus_27_add_3_3.INIT0 = 16'hf555;
    defparam unary_minus_27_add_3_3.INIT1 = 16'hf555;
    defparam unary_minus_27_add_3_3.INJECT1_0 = "NO";
    defparam unary_minus_27_add_3_3.INJECT1_1 = "NO";
    L6MUX21 i22466 (.D0(n24958), .D1(n24959), .SD(index_q[6]), .Z(n24967));
    LUT4 i20760_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n23242)) /* synthesis lut_function=(A (B (C)+!B (C (D)+!C !(D)))+!A !(B (C+!(D))+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20760_3_lut_4_lut_4_lut.init = 16'ha593;
    LUT4 i20722_3_lut_4_lut (.A(index_i[1]), .B(index_i[0]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n23204)) /* synthesis lut_function=(!(A (B (C (D))+!B (D))+!A (B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20722_3_lut_4_lut.init = 16'h18aa;
    L6MUX21 i22498 (.D0(n24991), .D1(n24992), .SD(index_q[6]), .Z(n24999));
    FD1P3AX phase_i_i0_i0 (.D(o_phase[0]), .SP(dac_clk_p_c_enable_630), 
            .CK(dac_clk_p_c), .Q(phase_i[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam phase_i_i0_i0.GSR = "DISABLED";
    L6MUX21 i22501 (.D0(n24997), .D1(n24998), .SD(index_q[6]), .Z(n25002));
    LUT4 i14377_2_lut_rep_711 (.A(index_q[2]), .B(index_q[0]), .Z(n29371)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14377_2_lut_rep_711.init = 16'heeee;
    L6MUX21 i22529 (.D0(n25022), .D1(n25023), .SD(index_i[6]), .Z(n25030));
    PFUMX i27092 (.BLUT(n29512), .ALUT(n29513), .C0(index_q[0]), .Z(n29514));
    L6MUX21 i22532 (.D0(n25028), .D1(n25029), .SD(index_i[6]), .Z(n25033));
    PFUMX i22573 (.BLUT(n25058), .ALUT(n25059), .C0(index_q[6]), .Z(n25074));
    L6MUX21 i22574 (.D0(n25060), .D1(n25061), .SD(index_q[6]), .Z(n25075));
    PFUMX i20738 (.BLUT(n23218), .ALUT(n23219), .C0(index_i[4]), .Z(n23220));
    L6MUX21 i22575 (.D0(n25062), .D1(n25063), .SD(index_q[6]), .Z(n25076));
    L6MUX21 i22576 (.D0(n25064), .D1(n25065), .SD(index_q[6]), .Z(n25077));
    L6MUX21 i22577 (.D0(n25066), .D1(n25067), .SD(index_q[6]), .Z(n25078));
    L6MUX21 i22578 (.D0(n25068), .D1(n25069), .SD(index_q[6]), .Z(n25079));
    PFUMX i20802 (.BLUT(n318), .ALUT(n381), .C0(index_i[6]), .Z(n23284));
    LUT4 mux_207_Mux_1_i763_3_lut_4_lut (.A(index_q[4]), .B(index_q[3]), 
         .C(n29581), .D(n29389), .Z(n763)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_1_i763_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i20741 (.BLUT(n23221), .ALUT(n23222), .C0(index_i[4]), .Z(n23223));
    FD1S3DX o_val_pipeline_q_1__i1 (.D(\o_val_pipeline_q[0] [0]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(o_sample_q[0])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_q_1__i1.GSR = "DISABLED";
    FD1S3DX phase_negation_i_i0 (.D(phase_i[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(phase_negation_i[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam phase_negation_i_i0.GSR = "DISABLED";
    FD1S3DX phase_negation_q_i0 (.D(phase_q[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(phase_negation_q[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam phase_negation_q_i0.GSR = "DISABLED";
    FD1S3DX index_i_i0 (.D(index_i_9__N_1748[0]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(index_i[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam index_i_i0.GSR = "DISABLED";
    FD1S3DX index_q_i0 (.D(index_q_9__N_1758[0]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(index_q[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam index_q_i0.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i0 (.D(quarter_wave_sample_register_q_15__N_1783[0]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_q[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_q_i0.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i1 (.D(\o_val_pipeline_i[0] [0]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(o_sample_i[0])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i1.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i0 (.D(quarter_wave_sample_register_i_15__N_1768[0]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_i[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_i_i0.GSR = "DISABLED";
    PFUMX i20784 (.BLUT(n318_adj_2938), .ALUT(n381_adj_2939), .C0(index_q[6]), 
          .Z(n23266));
    PFUMX i20645 (.BLUT(n23125), .ALUT(n23126), .C0(index_q[4]), .Z(n476));
    CCU2D unary_minus_27_add_3_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(quarter_wave_sample_register_q[0]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .COUT(n19706), .S1(o_val_pipeline_q_0__15__N_1831[0]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(81[29:60])
    defparam unary_minus_27_add_3_1.INIT0 = 16'hF000;
    defparam unary_minus_27_add_3_1.INIT1 = 16'h0aaa;
    defparam unary_minus_27_add_3_1.INJECT1_0 = "NO";
    defparam unary_minus_27_add_3_1.INJECT1_1 = "NO";
    LUT4 i24132_3_lut (.A(n28141), .B(n62), .C(index_q[5]), .Z(n25058)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24132_3_lut.init = 16'hcaca;
    LUT4 i20623_3_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[0]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n23105)) /* synthesis lut_function=(!(A (C)+!A (B (C+!(D))+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20623_3_lut_3_lut_4_lut.init = 16'h0f1a;
    PFUMX i27090 (.BLUT(n29509), .ALUT(n29510), .C0(index_q[1]), .Z(n29511));
    PFUMX i11039 (.BLUT(n13548), .ALUT(n13549), .C0(n24318), .Z(n13335));
    LUT4 n262_bdd_3_lut_26278_4_lut (.A(index_q[2]), .B(index_q[0]), .C(index_q[1]), 
         .D(index_q[4]), .Z(n28139)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B (D))) */ ;
    defparam n262_bdd_3_lut_26278_4_lut.init = 16'hf10e;
    LUT4 mux_206_Mux_4_i526_3_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n526)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A !(B ((D)+!C)+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_4_i526_3_lut_3_lut_4_lut.init = 16'h7e0f;
    LUT4 i1_2_lut_rep_507_3_lut (.A(index_q[2]), .B(index_q[0]), .C(index_q[1]), 
         .Z(n29167)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_507_3_lut.init = 16'hfefe;
    PFUMX i11098 (.BLUT(n13556), .ALUT(n13557), .C0(n24310), .Z(n13394));
    LUT4 mux_207_Mux_5_i459_3_lut_4_lut_3_lut_rep_733 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29393)) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_5_i459_3_lut_4_lut_3_lut_rep_733.init = 16'h6b6b;
    LUT4 i20649_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n23131)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i20649_3_lut_4_lut.init = 16'h64cc;
    CCU2D unary_minus_10_add_3_17 (.A0(\quarter_wave_sample_register_i[15] ), 
          .B0(GND_net), .C0(GND_net), .D0(GND_net), .A1(GND_net), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n19705), .S0(o_val_pipeline_i_0__15__N_1799[15]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam unary_minus_10_add_3_17.INIT0 = 16'hf555;
    defparam unary_minus_10_add_3_17.INIT1 = 16'h0000;
    defparam unary_minus_10_add_3_17.INJECT1_0 = "NO";
    defparam unary_minus_10_add_3_17.INJECT1_1 = "NO";
    CCU2D unary_minus_10_add_3_15 (.A0(quarter_wave_sample_register_i[13]), 
          .B0(GND_net), .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[14]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19704), .COUT(n19705), 
          .S0(o_val_pipeline_i_0__15__N_1799[13]), .S1(o_val_pipeline_i_0__15__N_1799[14]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam unary_minus_10_add_3_15.INIT0 = 16'hf555;
    defparam unary_minus_10_add_3_15.INIT1 = 16'hf555;
    defparam unary_minus_10_add_3_15.INJECT1_0 = "NO";
    defparam unary_minus_10_add_3_15.INJECT1_1 = "NO";
    LUT4 n966_bdd_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[4]), .Z(n27072)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !((D)+!C))+!A !(B (D)+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n966_bdd_3_lut_4_lut_4_lut.init = 16'h6693;
    LUT4 i14284_2_lut_rep_799 (.A(index_q[0]), .B(index_q[1]), .Z(n29459)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14284_2_lut_rep_799.init = 16'heeee;
    CCU2D unary_minus_10_add_3_13 (.A0(quarter_wave_sample_register_i[11]), 
          .B0(GND_net), .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[12]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19703), .COUT(n19704), 
          .S0(o_val_pipeline_i_0__15__N_1799[11]), .S1(o_val_pipeline_i_0__15__N_1799[12]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam unary_minus_10_add_3_13.INIT0 = 16'hf555;
    defparam unary_minus_10_add_3_13.INIT1 = 16'hf555;
    defparam unary_minus_10_add_3_13.INJECT1_0 = "NO";
    defparam unary_minus_10_add_3_13.INJECT1_1 = "NO";
    LUT4 mux_207_Mux_5_i754_3_lut_4_lut_3_lut_rep_734 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29394)) /* synthesis lut_function=(!(A (B)+!A ((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_5_i754_3_lut_4_lut_3_lut_rep_734.init = 16'h2626;
    PFUMX i20747 (.BLUT(n23227), .ALUT(n23228), .C0(index_i[4]), .Z(n23229));
    PFUMX i27088 (.BLUT(n29506), .ALUT(n29507), .C0(index_q[0]), .Z(n29508));
    LUT4 mux_206_Mux_7_i716_3_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n716)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C+!(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_7_i716_3_lut_3_lut_4_lut.init = 16'h0f81;
    PFUMX i22666 (.BLUT(n25163), .ALUT(n25164), .C0(index_i[6]), .Z(n25167));
    LUT4 mux_207_Mux_2_i173_3_lut_4_lut_4_lut_4_lut (.A(index_q[2]), .B(index_q[0]), 
         .C(index_q[3]), .D(index_q[1]), .Z(n173)) /* synthesis lut_function=(!(A (C)+!A (B (C+!(D))+!B (C (D)+!C !(D))))) */ ;
    defparam mux_207_Mux_2_i173_3_lut_4_lut_4_lut_4_lut.init = 16'h0f1a;
    PFUMX i21833 (.BLUT(n221), .ALUT(n252), .C0(index_i[5]), .Z(n24334));
    PFUMX i22667 (.BLUT(n25165), .ALUT(n25166), .C0(index_i[6]), .Z(n25168));
    LUT4 i21492_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n23974)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(D))+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21492_3_lut_3_lut_4_lut.init = 16'h3319;
    LUT4 mux_206_Mux_6_i796_3_lut_rep_381_3_lut_3_lut_4_lut (.A(index_i[1]), 
         .B(index_i[0]), .C(index_i[3]), .D(index_i[2]), .Z(n29041)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_6_i796_3_lut_rep_381_3_lut_3_lut_4_lut.init = 16'hfe01;
    LUT4 i20914_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n23396)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B ((D)+!C)+!B (C))) */ ;
    defparam i20914_3_lut_4_lut_4_lut.init = 16'hfc1c;
    PFUMX i20750 (.BLUT(n23230), .ALUT(n23231), .C0(index_i[4]), .Z(n23232));
    LUT4 n348_bdd_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n28659)) /* synthesis lut_function=(A (B (D)+!B (C+(D)))+!A (B (D)+!B !(C (D)+!C !(D)))) */ ;
    defparam n348_bdd_3_lut_4_lut_4_lut.init = 16'hef30;
    LUT4 mux_207_Mux_5_i572_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n572)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A !(B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_5_i572_3_lut_4_lut_4_lut.init = 16'ha9a5;
    LUT4 mux_207_Mux_5_i954_3_lut_3_lut_4_lut_4_lut (.A(index_q[2]), .B(index_q[0]), 
         .C(index_q[3]), .D(index_q[1]), .Z(n954)) /* synthesis lut_function=(!(A (C)+!A (B+((D)+!C)))) */ ;
    defparam mux_207_Mux_5_i954_3_lut_3_lut_4_lut_4_lut.init = 16'h0a1a;
    CCU2D unary_minus_10_add_3_11 (.A0(quarter_wave_sample_register_i[9]), 
          .B0(GND_net), .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[10]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19702), .COUT(n19703), 
          .S0(o_val_pipeline_i_0__15__N_1799[9]), .S1(o_val_pipeline_i_0__15__N_1799[10]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam unary_minus_10_add_3_11.INIT0 = 16'hf555;
    defparam unary_minus_10_add_3_11.INIT1 = 16'hf555;
    defparam unary_minus_10_add_3_11.INJECT1_0 = "NO";
    defparam unary_minus_10_add_3_11.INJECT1_1 = "NO";
    LUT4 i12545_2_lut_rep_419_3_lut_4_lut (.A(index_q[2]), .B(index_q[0]), 
         .C(index_q[3]), .D(index_q[1]), .Z(n29079)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;
    defparam i12545_2_lut_rep_419_3_lut_4_lut.init = 16'hf0e0;
    PFUMX i20756 (.BLUT(n23236), .ALUT(n23237), .C0(index_i[4]), .Z(n23238));
    LUT4 mux_206_Mux_8_i285_3_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n285)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C+!(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_8_i285_3_lut_3_lut_4_lut.init = 16'h0fa1;
    LUT4 i5082_2_lut_rep_726 (.A(index_q[0]), .B(index_q[1]), .Z(n29386)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i5082_2_lut_rep_726.init = 16'h6666;
    LUT4 i17702_3_lut_3_lut (.A(index_i[0]), .B(index_i[2]), .C(index_i[3]), 
         .Z(n20016)) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i17702_3_lut_3_lut.init = 16'h6a6a;
    PFUMX i27086 (.BLUT(n29503), .ALUT(n29504), .C0(index_q[1]), .Z(n29505));
    LUT4 mux_206_Mux_4_i349_3_lut_4_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[4]), .D(n348), .Z(n349)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_4_i349_3_lut_4_lut.init = 16'hf606;
    PFUMX i20762 (.BLUT(n23242), .ALUT(n23243), .C0(index_i[4]), .Z(n23244));
    LUT4 mux_207_Mux_0_i46_3_lut_4_lut_4_lut_4_lut (.A(index_q[2]), .B(index_q[0]), 
         .C(index_q[1]), .D(index_q[3]), .Z(n46)) /* synthesis lut_function=(A (D)+!A (B+(C+!(D)))) */ ;
    defparam mux_207_Mux_0_i46_3_lut_4_lut_4_lut_4_lut.init = 16'hfe55;
    PFUMX i21863 (.BLUT(n158), .ALUT(n189), .C0(index_i[5]), .Z(n24364));
    PFUMX i22304 (.BLUT(n24801), .ALUT(n24802), .C0(index_q[4]), .Z(n24805));
    LUT4 mux_206_Mux_3_i557_3_lut_3_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n557)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_3_i557_3_lut_3_lut_3_lut_4_lut.init = 16'hf10f;
    PFUMX i22305 (.BLUT(n24803), .ALUT(n24804), .C0(index_q[4]), .Z(n24806));
    CCU2D unary_minus_10_add_3_9 (.A0(quarter_wave_sample_register_i[7]), 
          .B0(GND_net), .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[8]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19701), .COUT(n19702), 
          .S0(o_val_pipeline_i_0__15__N_1799[7]), .S1(o_val_pipeline_i_0__15__N_1799[8]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam unary_minus_10_add_3_9.INIT0 = 16'hf555;
    defparam unary_minus_10_add_3_9.INIT1 = 16'hf555;
    defparam unary_minus_10_add_3_9.INJECT1_0 = "NO";
    defparam unary_minus_10_add_3_9.INJECT1_1 = "NO";
    CCU2D unary_minus_10_add_3_7 (.A0(quarter_wave_sample_register_i[5]), 
          .B0(GND_net), .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[6]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19700), .COUT(n19701), 
          .S0(o_val_pipeline_i_0__15__N_1799[5]), .S1(o_val_pipeline_i_0__15__N_1799[6]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam unary_minus_10_add_3_7.INIT0 = 16'hf555;
    defparam unary_minus_10_add_3_7.INIT1 = 16'hf555;
    defparam unary_minus_10_add_3_7.INJECT1_0 = "NO";
    defparam unary_minus_10_add_3_7.INJECT1_1 = "NO";
    PFUMX i22812 (.BLUT(n526_adj_2940), .ALUT(n541), .C0(index_q[4]), 
          .Z(n25313));
    PFUMX i22311 (.BLUT(n24808), .ALUT(n24809), .C0(index_q[4]), .Z(n24812));
    L6MUX21 i22710 (.D0(n25199), .D1(n25200), .SD(index_q[6]), .Z(n25211));
    L6MUX21 i22711 (.D0(n25201), .D1(n25202), .SD(index_q[6]), .Z(n25212));
    LUT4 i21133_3_lut (.A(n32018), .B(n851), .C(index_i[3]), .Z(n23615)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21133_3_lut.init = 16'hcaca;
    L6MUX21 i22712 (.D0(n25203), .D1(n25204), .SD(index_q[6]), .Z(n25213));
    PFUMX i22312 (.BLUT(n24810), .ALUT(n24811), .C0(index_q[4]), .Z(n24813));
    PFUMX i22713 (.BLUT(n25205), .ALUT(n25206), .C0(index_q[6]), .Z(n25214));
    PFUMX i22722 (.BLUT(n13382), .ALUT(n23325), .C0(index_q[6]), .Z(n25223));
    LUT4 i14171_1_lut_rep_394_2_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n29054)) /* synthesis lut_function=(!(A (C+(D))+!A (B (C+(D))+!B (C)))) */ ;
    defparam i14171_1_lut_rep_394_2_lut_3_lut_4_lut.init = 16'h010f;
    LUT4 mux_207_Mux_9_i285_3_lut_4_lut_4_lut (.A(index_q[2]), .B(index_q[0]), 
         .C(index_q[3]), .D(index_q[1]), .Z(n285_adj_2941)) /* synthesis lut_function=(A (C)+!A !(B+(C+(D)))) */ ;
    defparam mux_207_Mux_9_i285_3_lut_4_lut_4_lut.init = 16'ha0a1;
    L6MUX21 i22724 (.D0(n23331), .D1(n23334), .SD(index_q[6]), .Z(n25225));
    L6MUX21 i22725 (.D0(n574), .D1(n23337), .SD(index_q[6]), .Z(n25226));
    L6MUX21 i22726 (.D0(n23340), .D1(n764), .SD(index_q[6]), .Z(n25227));
    LUT4 mux_206_Mux_3_i94_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[4]), .D(n93), .Z(n94)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_3_i94_3_lut_4_lut.init = 16'hf606;
    PFUMX i22740 (.BLUT(n25237), .ALUT(n25238), .C0(index_q[6]), .Z(n25241));
    PFUMX i22741 (.BLUT(n25239), .ALUT(n25240), .C0(index_q[6]), .Z(n25242));
    LUT4 mux_206_Mux_2_i890_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n890)) /* synthesis lut_function=(A (B (C)+!B !(C+!(D)))+!A !(B (C+(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_2_i890_3_lut_4_lut_4_lut.init = 16'h9394;
    LUT4 i11061_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n13357)) /* synthesis lut_function=(!(A (B (C)+!B ((D)+!C))+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11061_3_lut_4_lut_4_lut.init = 16'h4969;
    LUT4 mux_207_Mux_0_i173_3_lut_4_lut (.A(n29371), .B(index_q[1]), .C(index_q[3]), 
         .D(n29335), .Z(n173_adj_2942)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_0_i173_3_lut_4_lut.init = 16'hdfd0;
    LUT4 i11080_3_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[3]), .C(index_i[0]), 
         .D(index_i[1]), .Z(n844)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11080_3_lut_4_lut_4_lut.init = 16'hf00e;
    LUT4 i11024_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n13320)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))+!A !(B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11024_3_lut_4_lut_4_lut.init = 16'hb5b3;
    L6MUX21 i22767 (.D0(n25260), .D1(n25261), .SD(index_i[6]), .Z(n25268));
    LUT4 mux_207_Mux_1_i620_3_lut_4_lut (.A(n29371), .B(index_q[1]), .C(index_q[3]), 
         .D(n32034), .Z(n620)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_1_i620_3_lut_4_lut.init = 16'hdfd0;
    L6MUX21 i22768 (.D0(n25262), .D1(n25263), .SD(index_i[6]), .Z(n25269));
    LUT4 i21484_3_lut_4_lut (.A(n29371), .B(index_q[1]), .C(index_q[3]), 
         .D(n404), .Z(n23966)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i21484_3_lut_4_lut.init = 16'hdfd0;
    L6MUX21 i22769 (.D0(n25264), .D1(n25265), .SD(index_i[6]), .Z(n25270));
    LUT4 mux_206_Mux_5_i252_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[4]), .Z(n252)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+(D)))+!A (B (C (D))+!B !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_5_i252_3_lut_4_lut.init = 16'hc993;
    LUT4 mux_207_Mux_1_i882_3_lut_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n882)) /* synthesis lut_function=(A ((C)+!B)+!A !((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_1_i882_3_lut_3_lut.init = 16'ha6a6;
    L6MUX21 i22770 (.D0(n25266), .D1(n25267), .SD(index_i[6]), .Z(n25271));
    LUT4 mux_207_Mux_0_i645_3_lut_rep_521_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29181)) /* synthesis lut_function=(!(A (B)+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_0_i645_3_lut_rep_521_3_lut.init = 16'h6363;
    LUT4 i20755_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[2]), .C(index_i[3]), 
         .D(index_i[1]), .Z(n23237)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+!(D)))+!A !(B+!(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20755_3_lut_4_lut_4_lut.init = 16'h6c67;
    LUT4 i17701_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[1]), .Z(n20015)) /* synthesis lut_function=(A (B (C (D))+!B !(C))+!A (B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i17701_3_lut_4_lut_4_lut_4_lut.init = 16'hd656;
    LUT4 i11021_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n13317)) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B ((D)+!C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11021_3_lut_4_lut_4_lut.init = 16'hcdad;
    LUT4 i12716_2_lut_rep_763 (.A(index_i[0]), .B(index_i[1]), .Z(n29423)) /* synthesis lut_function=(A+!(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12716_2_lut_rep_763.init = 16'hbbbb;
    LUT4 mux_206_Mux_2_i173_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), 
         .B(index_i[2]), .C(index_i[3]), .D(index_i[0]), .Z(n173_adj_2943)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B ((D)+!C)))) */ ;
    defparam mux_206_Mux_2_i173_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h0e1e;
    LUT4 i12777_2_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n635)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A (B (C+!(D))+!B (C+(D)))) */ ;
    defparam i12777_2_lut_4_lut_4_lut.init = 16'hf1fc;
    LUT4 i20749_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n23231)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B (C+!(D))+!B !(C)))) */ ;
    defparam i20749_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h1c18;
    LUT4 n45_bdd_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n27538)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B !(C)))) */ ;
    defparam n45_bdd_3_lut_4_lut_4_lut_4_lut.init = 16'h1e1c;
    LUT4 i20919_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n23401)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !(B (C+!(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i20919_3_lut_4_lut_4_lut.init = 16'ha5a9;
    LUT4 n262_bdd_3_lut_26735_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[4]), .Z(n28140)) /* synthesis lut_function=(A (B (D)+!B !((D)+!C))+!A !(B (D)+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam n262_bdd_3_lut_26735_4_lut_4_lut.init = 16'h9964;
    LUT4 mux_206_Mux_7_i747_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), 
         .B(index_i[2]), .C(index_i[3]), .D(index_i[0]), .Z(n747)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))+!A (B (C)+!B !(C))) */ ;
    defparam mux_206_Mux_7_i747_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'he1e3;
    LUT4 i12656_2_lut_rep_435_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n29095)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i12656_2_lut_rep_435_3_lut_4_lut.init = 16'hfef0;
    LUT4 mux_207_Mux_0_i525_3_lut_3_lut_rep_735 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29395)) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_0_i525_3_lut_3_lut_rep_735.init = 16'h6a6a;
    L6MUX21 i22801 (.D0(n25290), .D1(n25291), .SD(index_i[6]), .Z(n25302));
    L6MUX21 i22802 (.D0(n25292), .D1(n25293), .SD(index_i[6]), .Z(n25303));
    L6MUX21 i22803 (.D0(n25294), .D1(n25295), .SD(index_i[6]), .Z(n25304));
    PFUMX i22804 (.BLUT(n25296), .ALUT(n25297), .C0(index_i[6]), .Z(n25305));
    LUT4 n172_bdd_2_lut_3_lut_3_lut_4_lut (.A(index_q[2]), .B(index_q[0]), 
         .C(index_q[1]), .D(index_q[3]), .Z(n27389)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B ((D)+!C)))) */ ;
    defparam n172_bdd_2_lut_3_lut_3_lut_4_lut.init = 16'h00fe;
    LUT4 i20652_3_lut_3_lut_4_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n23134)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20652_3_lut_3_lut_4_lut_3_lut_4_lut.init = 16'h11ef;
    LUT4 i11134_3_lut_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[4]), .D(index_q[3]), .Z(n444)) /* synthesis lut_function=(!(A (B)+!A !(B (C (D))+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i11134_3_lut_3_lut_4_lut_4_lut.init = 16'h6333;
    L6MUX21 i22836 (.D0(n25329), .D1(n25330), .SD(index_q[6]), .Z(n25337));
    L6MUX21 i22837 (.D0(n25331), .D1(n25332), .SD(index_q[6]), .Z(n25338));
    L6MUX21 i22838 (.D0(n25333), .D1(n25334), .SD(index_q[6]), .Z(n25339));
    LUT4 i12669_3_lut_4_lut (.A(index_q[4]), .B(n29326), .C(index_q[5]), 
         .D(n29459), .Z(n892)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i12669_3_lut_4_lut.init = 16'hf8f0;
    LUT4 i20668_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n23150)) /* synthesis lut_function=(A (C+(D))+!A !(B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20668_3_lut_4_lut_4_lut.init = 16'haba5;
    L6MUX21 i22839 (.D0(n25335), .D1(n25336), .SD(index_q[6]), .Z(n25340));
    LUT4 mux_207_Mux_3_i796_3_lut (.A(index_q[2]), .B(n731), .C(index_q[4]), 
         .Z(n796)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_3_i796_3_lut.init = 16'hacac;
    LUT4 n966_bdd_4_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[0]), 
         .D(index_i[4]), .Z(n27071)) /* synthesis lut_function=(!(A (D)+!A !(B (D)+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n966_bdd_4_lut_3_lut_4_lut.init = 16'h54ab;
    LUT4 i20740_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[3]), 
         .C(index_i[2]), .D(index_i[0]), .Z(n23222)) /* synthesis lut_function=(!(A (B+!((D)+!C))+!A !(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20740_3_lut_4_lut_4_lut_4_lut.init = 16'h6747;
    LUT4 mux_206_Mux_7_i491_3_lut_4_lut_4_lut_4_lut_4_lut (.A(index_i[1]), 
         .B(index_i[3]), .C(index_i[2]), .D(index_i[0]), .Z(n491)) /* synthesis lut_function=(!(A (B (C+!(D))+!B ((D)+!C))+!A !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_7_i491_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'h5870;
    LUT4 mux_207_Mux_6_i731_3_lut (.A(n29460), .B(n32054), .C(index_q[3]), 
         .Z(n731)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_6_i731_3_lut.init = 16'hcaca;
    LUT4 i12710_2_lut_rep_410_4_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n29070)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12710_2_lut_rep_410_4_lut_4_lut_4_lut_4_lut.init = 16'h0058;
    LUT4 mux_206_Mux_0_i251_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n251)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A !(B ((D)+!C)+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i251_3_lut_4_lut_4_lut_4_lut.init = 16'h543c;
    LUT4 i22588_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[3]), 
         .C(index_i[2]), .D(index_i[0]), .Z(n25089)) /* synthesis lut_function=(A (B (C (D))+!B (C))+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i22588_3_lut_4_lut_4_lut_4_lut.init = 16'hb434;
    LUT4 mux_206_Mux_1_i348_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[3]), 
         .C(index_i[2]), .D(index_i[0]), .Z(n348_adj_2944)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_1_i348_3_lut_4_lut_4_lut_4_lut.init = 16'h7870;
    LUT4 mux_207_Mux_5_i109_3_lut_3_lut_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .Z(n109)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_5_i109_3_lut_3_lut_3_lut.init = 16'h3939;
    LUT4 mux_206_Mux_0_i1017_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n1017)) /* synthesis lut_function=(A (B (C)+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i1017_4_lut_4_lut_4_lut.init = 16'hd7d0;
    LUT4 mux_207_Mux_1_i716_3_lut_3_lut_4_lut_4_lut (.A(index_q[2]), .B(index_q[0]), 
         .C(index_q[1]), .D(index_q[3]), .Z(n716_adj_2945)) /* synthesis lut_function=(!(A (B (D)+!B !(C))+!A !(B (C (D))+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_1_i716_3_lut_3_lut_4_lut_4_lut.init = 16'h70a9;
    LUT4 mux_207_Mux_8_i716_3_lut_4_lut_4_lut_4_lut (.A(index_q[2]), .B(index_q[0]), 
         .C(index_q[1]), .D(index_q[3]), .Z(n716_adj_2946)) /* synthesis lut_function=(!(A (D)+!A !(B+(C+(D))))) */ ;
    defparam mux_207_Mux_8_i716_3_lut_4_lut_4_lut_4_lut.init = 16'h55fe;
    LUT4 i20941_3_lut_4_lut (.A(n29459), .B(index_q[2]), .C(index_q[3]), 
         .D(n32036), .Z(n23423)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i20941_3_lut_4_lut.init = 16'hdfd0;
    LUT4 i22663_3_lut_4_lut_4_lut (.A(n29147), .B(index_i[4]), .C(index_i[5]), 
         .D(n29086), .Z(n25164)) /* synthesis lut_function=(A ((C+!(D))+!B)+!A (B (C+!(D))+!B !(C))) */ ;
    defparam i22663_3_lut_4_lut_4_lut.init = 16'he3ef;
    PFUMX i27084 (.BLUT(n29499), .ALUT(n29500), .C0(index_i[1]), .Z(n29501));
    LUT4 n875_bdd_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n27460)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A !((C)+!B))) */ ;
    defparam n875_bdd_3_lut_4_lut_4_lut_4_lut.init = 16'h7173;
    LUT4 mux_206_Mux_6_i908_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), 
         .B(index_i[2]), .C(index_i[3]), .D(index_i[0]), .Z(n908)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B ((D)+!C)+!B !(C)))) */ ;
    defparam mux_206_Mux_6_i908_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h3878;
    LUT4 i20725_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n23207)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B (C+(D))+!B (C)))) */ ;
    defparam i20725_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h7c78;
    LUT4 n285_bdd_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n27462)) /* synthesis lut_function=(A (B (C)+!B ((D)+!C))+!A (B+!(C))) */ ;
    defparam n285_bdd_3_lut_4_lut_4_lut_4_lut.init = 16'he7c7;
    LUT4 mux_207_Mux_8_i460_3_lut_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n460)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B ((D)+!C))) */ ;
    defparam mux_207_Mux_8_i460_3_lut_3_lut_3_lut_4_lut.init = 16'hf10f;
    LUT4 mux_206_Mux_9_i316_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n316)) /* synthesis lut_function=(!(A (B (C)+!B !(C+(D)))+!A !(B+(C)))) */ ;
    defparam mux_206_Mux_9_i316_3_lut_4_lut_4_lut_4_lut.init = 16'h7e7c;
    LUT4 i22796_3_lut_4_lut_4_lut (.A(n29148), .B(index_i[5]), .C(index_i[4]), 
         .D(n29064), .Z(n25297)) /* synthesis lut_function=(A (B+(C (D)))+!A (B+((D)+!C))) */ ;
    defparam i22796_3_lut_4_lut_4_lut.init = 16'hfdcd;
    LUT4 mux_206_Mux_3_i62_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[4]), .D(n812), .Z(n62_adj_2947)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_3_i62_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_206_Mux_0_i731_3_lut_4_lut (.A(n29376), .B(index_i[2]), .C(index_i[3]), 
         .D(n32018), .Z(n731_adj_2948)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i731_3_lut_4_lut.init = 16'h4f40;
    LUT4 i21448_3_lut_4_lut (.A(n29376), .B(index_i[2]), .C(index_i[3]), 
         .D(n32022), .Z(n23930)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21448_3_lut_4_lut.init = 16'hf404;
    LUT4 i20586_3_lut (.A(n931), .B(n29429), .C(index_i[3]), .Z(n23068)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20586_3_lut.init = 16'hcaca;
    LUT4 i11032_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n13328)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))+!A !(B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i11032_3_lut_4_lut_4_lut.init = 16'hb5b3;
    LUT4 i11035_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n13331)) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B ((D)+!C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i11035_3_lut_4_lut_4_lut.init = 16'hcdad;
    LUT4 i11082_3_lut_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n875)) /* synthesis lut_function=(A (C (D))+!A !(B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11082_3_lut_3_lut_4_lut_4_lut.init = 16'hb555;
    LUT4 i11266_3_lut_3_lut_4_lut_4_lut_4_lut_4_lut (.A(index_i[3]), .B(index_i[1]), 
         .C(index_i[0]), .D(index_i[2]), .Z(n13565)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A !(B (D)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11266_3_lut_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'habd5;
    LUT4 i20908_3_lut_4_lut_4_lut (.A(n29370), .B(n29396), .C(index_q[3]), 
         .D(index_q[0]), .Z(n23390)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C))) */ ;
    defparam i20908_3_lut_4_lut_4_lut.init = 16'hcfc5;
    LUT4 i11075_3_lut_3_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[0]), .D(index_i[1]), .Z(n762)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C (D)+!C !(D)))+!A !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11075_3_lut_3_lut_4_lut_4_lut.init = 16'h700f;
    LUT4 mux_207_Mux_5_i252_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[4]), .Z(n252_adj_2949)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+(D)))+!A (B (C (D))+!B !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_5_i252_3_lut_4_lut.init = 16'hc993;
    LUT4 mux_206_Mux_4_i812_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[4]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n812_adj_2950)) /* synthesis lut_function=(A (B (C+(D)))+!A !(B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_4_i812_3_lut_3_lut_4_lut.init = 16'h9995;
    LUT4 mux_206_Mux_0_i443_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n443)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (D))+!A !(B (D)+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i443_3_lut_4_lut_4_lut_4_lut.init = 16'h54b3;
    LUT4 mux_207_Mux_0_i604_3_lut_4_lut_4_lut_4_lut (.A(index_q[2]), .B(index_q[0]), 
         .C(index_q[1]), .D(index_q[3]), .Z(n604)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A !(B (D)+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_0_i604_3_lut_4_lut_4_lut_4_lut.init = 16'h5439;
    LUT4 mux_207_Mux_0_i428_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_q[2]), 
         .B(index_q[0]), .C(index_q[1]), .D(index_q[3]), .Z(n428)) /* synthesis lut_function=(A (B (C+!(D))+!B !((D)+!C))+!A (B (D)+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_0_i428_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hd5a9;
    LUT4 mux_207_Mux_0_i443_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[0]), .D(index_q[3]), .Z(n443_adj_2951)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C (D))+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_0_i443_3_lut_4_lut_4_lut_4_lut.init = 16'h0ed5;
    LUT4 i20911_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n23393)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(D))+!A (B (D)+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i20911_3_lut_4_lut_4_lut_4_lut.init = 16'hd52b;
    LUT4 i20842_3_lut_else_4_lut (.A(index_q[4]), .B(index_q[1]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n29512)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A !(B (C+!(D))+!B ((D)+!C)))) */ ;
    defparam i20842_3_lut_else_4_lut.init = 16'h59e5;
    LUT4 index_q_0__bdd_4_lut_27767 (.A(index_q[0]), .B(index_q[3]), .C(index_q[1]), 
         .D(index_q[2]), .Z(n29518)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C (D)))+!A !(B (C+!(D))+!B !(C+(D))))) */ ;
    defparam index_q_0__bdd_4_lut_27767.init = 16'h4ae7;
    LUT4 i14149_3_lut_3_lut_rep_838 (.A(index_i[2]), .B(index_i[0]), .C(index_i[1]), 
         .Z(n32039)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i14149_3_lut_3_lut_rep_838.init = 16'hd0d0;
    LUT4 i20692_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n23174)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C))+!A (B (C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i20692_3_lut_4_lut_4_lut_4_lut.init = 16'he078;
    LUT4 i17699_3_lut (.A(n29405), .B(n29447), .C(index_i[3]), .Z(n20013)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17699_3_lut.init = 16'hcaca;
    LUT4 i22302_3_lut_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n24803)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C+!(D))+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i22302_3_lut_3_lut_4_lut_4_lut.init = 16'h1f81;
    PFUMX i25365 (.BLUT(n27072), .ALUT(n27071), .C0(index_i[3]), .Z(n27073));
    LUT4 i12852_2_lut_rep_712 (.A(index_i[2]), .B(index_i[3]), .Z(n29372)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12852_2_lut_rep_712.init = 16'heeee;
    LUT4 mux_207_Mux_8_i61_3_lut_rep_403_4_lut_4_lut_4_lut (.A(index_q[0]), 
         .B(index_q[1]), .C(index_q[2]), .D(index_q[3]), .Z(n29063)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A (B (C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_8_i61_3_lut_rep_403_4_lut_4_lut_4_lut.init = 16'he0f8;
    LUT4 mux_207_Mux_8_i251_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), 
         .B(index_q[1]), .C(index_q[2]), .D(index_q[3]), .Z(n251_adj_2952)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_8_i251_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h07e0;
    LUT4 i17698_3_lut (.A(n29447), .B(n29441), .C(index_i[3]), .Z(n20012)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17698_3_lut.init = 16'hcaca;
    LUT4 i22301_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n24802)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i22301_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hf81f;
    LUT4 mux_207_Mux_8_i157_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n15)) /* synthesis lut_function=(A (B (C)+!B !(C (D)+!C !(D)))+!A !(B ((D)+!C)+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_8_i157_3_lut_4_lut_4_lut.init = 16'h83e0;
    LUT4 i11143_3_lut_4_lut_3_lut_4_lut (.A(index_q[1]), .B(index_q[0]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n844_adj_2953)) /* synthesis lut_function=(A (B)+!A !(B+!(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i11143_3_lut_4_lut_3_lut_4_lut.init = 16'h9998;
    PFUMX i22318 (.BLUT(n24815), .ALUT(n24816), .C0(index_q[4]), .Z(n24819));
    LUT4 mux_207_Mux_0_i588_3_lut_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n588)) /* synthesis lut_function=(!(A (B+(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_0_i588_3_lut_3_lut.init = 16'h5656;
    LUT4 i21450_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n23932)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B+(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21450_3_lut_4_lut_4_lut_4_lut.init = 16'h2aab;
    LUT4 i20734_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n23216)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(D))+!A (B (D)+!B ((D)+!C))) */ ;
    defparam i20734_3_lut_4_lut_4_lut.init = 16'hd52b;
    PFUMX i22229 (.BLUT(n956), .ALUT(n22180), .C0(index_i[6]), .Z(n24730));
    LUT4 mux_206_Mux_8_i109_3_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n109_adj_2954)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (B (C+!(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_8_i109_3_lut_4_lut_4_lut.init = 16'hf85e;
    LUT4 i22591_3_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[0]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n25092)) /* synthesis lut_function=(A (B (C+!(D))+!B !((D)+!C))+!A !(B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i22591_3_lut_4_lut_4_lut.init = 16'h81f8;
    LUT4 mux_206_Mux_8_i251_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), 
         .B(index_i[0]), .C(index_i[2]), .D(index_i[3]), .Z(n251_adj_2955)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_8_i251_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h07e0;
    LUT4 mux_206_Mux_0_i460_3_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n460_adj_2956)) /* synthesis lut_function=(A (B+(C))+!A (C (D)+!C !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i460_3_lut_4_lut_4_lut.init = 16'hf8ad;
    LUT4 i20629_3_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[0]), .C(index_i[1]), 
         .D(index_i[3]), .Z(n23111)) /* synthesis lut_function=(A (B (C)+!B !(C+!(D)))+!A (B (C)+!B !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20629_3_lut_4_lut_4_lut.init = 16'hc3d0;
    LUT4 i22589_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n25090)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i22589_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hf81f;
    LUT4 i11255_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n13554)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B ((D)+!C)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i11255_3_lut_4_lut_4_lut.init = 16'h6c3c;
    LUT4 i11100_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n526_adj_2957)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+(D)))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i11100_3_lut_4_lut_4_lut.init = 16'h666c;
    PFUMX mux_206_Mux_7_i190 (.BLUT(n23613), .ALUT(n173_adj_2958), .C0(index_i[5]), 
          .Z(n190)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 mux_207_Mux_3_i507_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[4]), .D(n491_adj_2959), .Z(n507)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_3_i507_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_206_Mux_6_i859_3_lut_rep_398_4_lut_4_lut_4_lut (.A(index_i[1]), 
         .B(index_i[0]), .C(index_i[2]), .D(index_i[3]), .Z(n29058)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A (B (C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_6_i859_3_lut_rep_398_4_lut_4_lut_4_lut.init = 16'he0f8;
    LUT4 mux_206_Mux_0_i379_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n379)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !((D)+!C))+!A !(B ((D)+!C)+!B (D))) */ ;
    defparam mux_206_Mux_0_i379_3_lut_4_lut_4_lut.init = 16'h8079;
    LUT4 mux_207_Mux_3_i908_3_lut (.A(n29393), .B(n32035), .C(index_q[3]), 
         .Z(n908_adj_2960)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_3_i908_3_lut.init = 16'hcaca;
    LUT4 i20905_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n23387)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C+(D)))+!A (B (C (D)+!C !(D))+!B !(C)))) */ ;
    defparam i20905_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h3ef0;
    LUT4 mux_206_Mux_3_i109_3_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n109_adj_2961)) /* synthesis lut_function=(A (D)+!A !(B (C+!(D))+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_3_i109_3_lut_4_lut_4_lut.init = 16'haf10;
    LUT4 n273_bdd_3_lut_4_lut_3_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .Z(n27619)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)+!B !(C)))) */ ;
    defparam n273_bdd_3_lut_4_lut_3_lut.init = 16'h6161;
    PFUMX i22241 (.BLUT(n24738), .ALUT(n24739), .C0(index_q[5]), .Z(n24742));
    LUT4 mux_206_Mux_8_i443_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n443_adj_2962)) /* synthesis lut_function=(A (B (C+!(D))+!B !((D)+!C))+!A !(B (D)+!B ((D)+!C))) */ ;
    defparam mux_206_Mux_8_i443_3_lut_4_lut_4_lut.init = 16'h80fc;
    PFUMX i22242 (.BLUT(n24740), .ALUT(n24741), .C0(index_q[5]), .Z(n24743));
    LUT4 i22590_3_lut_3_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n25091)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C+!(D))+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i22590_3_lut_3_lut_4_lut_4_lut.init = 16'h1f81;
    LUT4 mux_206_Mux_2_i557_3_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n557_adj_2963)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C+!(D))+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_2_i557_3_lut_4_lut_4_lut.init = 16'h0f18;
    LUT4 mux_206_Mux_0_i428_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), 
         .B(index_i[0]), .C(index_i[2]), .D(index_i[3]), .Z(n428_adj_2964)) /* synthesis lut_function=(A (B (C+(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i428_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h8fe1;
    PFUMX mux_206_Mux_8_i764 (.BLUT(n716_adj_2965), .ALUT(n732), .C0(n24303), 
          .Z(n764_adj_2966)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 mux_207_Mux_2_i955_else_4_lut (.A(index_q[4]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n29506)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+(D)))+!A !(B (C+!(D))+!B !(C+!(D))))) */ ;
    defparam mux_207_Mux_2_i955_else_4_lut.init = 16'h49c6;
    LUT4 n22_bdd_3_lut_24997 (.A(n29354), .B(n29390), .C(index_q[3]), 
         .Z(n26642)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n22_bdd_3_lut_24997.init = 16'hcaca;
    LUT4 i22303_3_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[0]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n24804)) /* synthesis lut_function=(A (B (C+!(D))+!B !((D)+!C))+!A !(B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i22303_3_lut_4_lut_4_lut.init = 16'h81f8;
    PFUMX i22248 (.BLUT(n24745), .ALUT(n24746), .C0(index_q[5]), .Z(n24749));
    LUT4 mux_207_Mux_8_i109_3_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[0]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n109_adj_2967)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (B (C+!(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_8_i109_3_lut_4_lut_4_lut.init = 16'hf85e;
    LUT4 mux_207_Mux_0_i460_3_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[0]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n460_adj_2968)) /* synthesis lut_function=(A (B+(C))+!A (C (D)+!C !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_0_i460_3_lut_4_lut_4_lut.init = 16'hf8ad;
    LUT4 mux_207_Mux_8_i443_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n443_adj_2969)) /* synthesis lut_function=(A (B (C+!(D))+!B !((D)+!C))+!A !(B (D)+!B ((D)+!C))) */ ;
    defparam mux_207_Mux_8_i443_3_lut_4_lut_4_lut.init = 16'h80fc;
    PFUMX i22249 (.BLUT(n24747), .ALUT(n24748), .C0(index_q[5]), .Z(n24750));
    LUT4 mux_207_Mux_0_i379_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n379_adj_2970)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !((D)+!C))+!A !(B ((D)+!C)+!B (D))) */ ;
    defparam mux_207_Mux_0_i379_3_lut_4_lut_4_lut.init = 16'h8079;
    PFUMX mux_206_Mux_8_i574 (.BLUT(n542), .ALUT(n13528), .C0(index_i[5]), 
          .Z(n574_adj_2971)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    CCU2D unary_minus_10_add_3_5 (.A0(quarter_wave_sample_register_i[3]), 
          .B0(GND_net), .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[4]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19699), .COUT(n19700), 
          .S0(o_val_pipeline_i_0__15__N_1799[3]), .S1(o_val_pipeline_i_0__15__N_1799[4]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam unary_minus_10_add_3_5.INIT0 = 16'hf555;
    defparam unary_minus_10_add_3_5.INIT1 = 16'hf555;
    defparam unary_minus_10_add_3_5.INJECT1_0 = "NO";
    defparam unary_minus_10_add_3_5.INJECT1_1 = "NO";
    LUT4 i20698_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n23180)) /* synthesis lut_function=(A (C)+!A !(B (C)+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i20698_3_lut_4_lut_4_lut.init = 16'hb4b5;
    CCU2D unary_minus_10_add_3_3 (.A0(quarter_wave_sample_register_i[1]), 
          .B0(GND_net), .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[2]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19698), .COUT(n19699), 
          .S0(o_val_pipeline_i_0__15__N_1799[1]), .S1(o_val_pipeline_i_0__15__N_1799[2]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam unary_minus_10_add_3_3.INIT0 = 16'hf555;
    defparam unary_minus_10_add_3_3.INIT1 = 16'hf555;
    defparam unary_minus_10_add_3_3.INJECT1_0 = "NO";
    defparam unary_minus_10_add_3_3.INJECT1_1 = "NO";
    LUT4 mux_206_Mux_11_i445_3_lut_4_lut_4_lut_4_lut (.A(index_i[3]), .B(index_i[4]), 
         .C(index_i[5]), .D(n29176), .Z(n445)) /* synthesis lut_function=(!(A (B (C))+!A !(B+(C+(D))))) */ ;
    defparam mux_206_Mux_11_i445_3_lut_4_lut_4_lut_4_lut.init = 16'h7f7e;
    LUT4 mux_206_Mux_4_i900_3_lut_4_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n900)) /* synthesis lut_function=(A ((C)+!B)+!A !(B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_4_i900_3_lut_4_lut_4_lut_3_lut.init = 16'hb2b2;
    LUT4 index_i_5__bdd_2_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[2]), .D(index_i[5]), .Z(n27188)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam index_i_5__bdd_2_lut_4_lut_4_lut.init = 16'h718e;
    LUT4 mux_206_Mux_1_i684_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n684)) /* synthesis lut_function=(A (B ((D)+!C)+!B !((D)+!C))+!A !(B (C+(D))+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_1_i684_3_lut_4_lut_4_lut.init = 16'h992d;
    LUT4 n953_bdd_3_lut_25659_4_lut (.A(n29423), .B(index_i[2]), .C(index_i[3]), 
         .D(n32025), .Z(n26726)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n953_bdd_3_lut_25659_4_lut.init = 16'hf606;
    LUT4 mux_206_Mux_3_i890_3_lut_4_lut (.A(n29423), .B(index_i[2]), .C(index_i[3]), 
         .D(n325_adj_2972), .Z(n890_adj_2973)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_3_i890_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_207_Mux_1_i684_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n684_adj_2974)) /* synthesis lut_function=(A (B ((D)+!C)+!B !((D)+!C))+!A !(B (C+(D))+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_1_i684_3_lut_4_lut_4_lut.init = 16'h992d;
    LUT4 mux_206_Mux_0_i348_3_lut_4_lut (.A(n29423), .B(index_i[2]), .C(index_i[3]), 
         .D(n32056), .Z(n348_adj_2975)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i348_3_lut_4_lut.init = 16'h6f60;
    LUT4 i21436_3_lut_4_lut (.A(n29423), .B(index_i[2]), .C(index_i[3]), 
         .D(n29437), .Z(n23918)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21436_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_206_Mux_3_i491_3_lut_4_lut (.A(n29301), .B(index_i[1]), .C(index_i[3]), 
         .D(n29436), .Z(n491_adj_2976)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_3_i491_3_lut_4_lut.init = 16'h4f40;
    LUT4 index_q_1__bdd_4_lut_27802 (.A(index_q[1]), .B(index_q[0]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n29519)) /* synthesis lut_function=(!(A (B (D)+!B (C+!(D)))+!A !(B (C (D)+!C !(D))+!B !((D)+!C)))) */ ;
    defparam index_q_1__bdd_4_lut_27802.init = 16'h429c;
    LUT4 mux_206_Mux_0_i475_3_lut_4_lut (.A(n29301), .B(index_i[1]), .C(index_i[3]), 
         .D(n29180), .Z(n475)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i475_3_lut_4_lut.init = 16'h4f40;
    LUT4 mux_206_Mux_0_i604_3_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n604_adj_2977)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)))+!A (B (C (D)+!C !(D))+!B (C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i604_3_lut_4_lut_4_lut.init = 16'h0e63;
    LUT4 mux_207_Mux_11_i445_3_lut_4_lut_4_lut_4_lut (.A(index_q[3]), .B(index_q[4]), 
         .C(index_q[5]), .D(n29204), .Z(n445_adj_2978)) /* synthesis lut_function=(!(A (B (C))+!A !(B+(C+(D))))) */ ;
    defparam mux_207_Mux_11_i445_3_lut_4_lut_4_lut_4_lut.init = 16'h7f7e;
    LUT4 n953_bdd_3_lut_25002 (.A(n29357), .B(index_q[3]), .C(n29392), 
         .Z(n26646)) /* synthesis lut_function=(A (B+(C))+!A !(B+!(C))) */ ;
    defparam n953_bdd_3_lut_25002.init = 16'hb8b8;
    LUT4 mux_207_Mux_0_i890_3_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[0]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n890_adj_2979)) /* synthesis lut_function=(!(A (B (D)+!B !(C))+!A !(B (C (D)+!C !(D))+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_0_i890_3_lut_4_lut_4_lut.init = 16'h70ac;
    LUT4 mux_206_Mux_0_i412_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n412)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(D))+!A (B (D)+!B !(C+!(D)))) */ ;
    defparam mux_206_Mux_0_i412_3_lut_4_lut_4_lut.init = 16'hcd2a;
    LUT4 n285_bdd_3_lut (.A(n29357), .B(n29388), .C(index_q[3]), .Z(n26649)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n285_bdd_3_lut.init = 16'hacac;
    LUT4 mux_207_Mux_0_i684_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n684_adj_2980)) /* synthesis lut_function=(!(A ((D)+!B)+!A !(B (D)+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_0_i684_3_lut_4_lut_4_lut_4_lut.init = 16'h5498;
    LUT4 i20940_3_lut_4_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n23422)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B+(C+(D))))) */ ;
    defparam i20940_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'h2aab;
    LUT4 mux_206_Mux_7_i699_3_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n699)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C+!(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_7_i699_3_lut_4_lut_4_lut.init = 16'hf07e;
    LUT4 mux_207_Mux_7_i699_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n699_adj_2981)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C+!(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_7_i699_3_lut_4_lut_4_lut.init = 16'hf07e;
    LUT4 i17668_3_lut (.A(n29356), .B(n29353), .C(index_q[3]), .Z(n19982)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17668_3_lut.init = 16'hcaca;
    LUT4 i21439_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n23921)) /* synthesis lut_function=(A (C)+!A !(B (C)+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21439_3_lut_4_lut_4_lut.init = 16'hb4b5;
    LUT4 mux_206_Mux_1_i716_3_lut_3_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[1]), .D(index_i[3]), .Z(n716_adj_2982)) /* synthesis lut_function=(!(A (B (D)+!B !(C))+!A !(B (C (D))+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_1_i716_3_lut_3_lut_4_lut_4_lut.init = 16'h70a9;
    LUT4 i17667_3_lut (.A(n29353), .B(n29335), .C(index_q[3]), .Z(n19981)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17667_3_lut.init = 16'hcaca;
    LUT4 mux_206_Mux_2_i955_then_4_lut (.A(index_i[4]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n29521)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C (D)+!C !(D)))+!A (C+!(D))) */ ;
    defparam mux_206_Mux_2_i955_then_4_lut.init = 16'hda7d;
    LUT4 n773_bdd_3_lut_25068_4_lut (.A(n29402), .B(index_i[2]), .C(n29433), 
         .D(index_i[3]), .Z(n26718)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n773_bdd_3_lut_25068_4_lut.init = 16'hf066;
    LUT4 mux_206_Mux_3_i668_3_lut_4_lut (.A(n29402), .B(index_i[2]), .C(index_i[3]), 
         .D(n29441), .Z(n668)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_3_i668_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_206_Mux_0_i890_3_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n890_adj_2983)) /* synthesis lut_function=(!(A (B (D)+!B !(C))+!A !(B (C (D)+!C !(D))+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i890_3_lut_4_lut_4_lut.init = 16'h70ac;
    LUT4 mux_206_Mux_4_i763_3_lut_4_lut (.A(n29402), .B(index_i[2]), .C(index_i[4]), 
         .D(n747_adj_2984), .Z(n763_adj_2985)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_4_i763_3_lut_4_lut.init = 16'h6f60;
    LUT4 n698_bdd_3_lut_25715 (.A(n32039), .B(n32056), .C(index_i[3]), 
         .Z(n27373)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n698_bdd_3_lut_25715.init = 16'hcaca;
    LUT4 n698_bdd_3_lut_25625 (.A(n29385), .B(n1001), .C(index_i[3]), 
         .Z(n27372)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B+(C)))) */ ;
    defparam n698_bdd_3_lut_25625.init = 16'h5c5c;
    LUT4 mux_207_Mux_0_i412_3_lut_4_lut_4_lut (.A(index_q[2]), .B(index_q[0]), 
         .C(index_q[1]), .D(index_q[3]), .Z(n412_adj_2986)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C (D)))+!A (B (C+!(D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_0_i412_3_lut_4_lut_4_lut.init = 16'hf14c;
    LUT4 mux_206_Mux_2_i955_else_4_lut (.A(index_i[4]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n29520)) /* synthesis lut_function=(A (B (C (D))+!B !(C+(D)))+!A !(B (C (D))+!B (C+!(D)))) */ ;
    defparam mux_206_Mux_2_i955_else_4_lut.init = 16'h8546;
    LUT4 mux_207_Mux_7_i653_3_lut_4_lut (.A(n29459), .B(index_q[2]), .C(index_q[3]), 
         .D(n29475), .Z(n653)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_7_i653_3_lut_4_lut.init = 16'hf606;
    LUT4 i20716_3_lut_4_lut (.A(n29459), .B(index_q[2]), .C(index_q[3]), 
         .D(n32054), .Z(n23198)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i20716_3_lut_4_lut.init = 16'h6f60;
    LUT4 i20869_3_lut_4_lut_4_lut_4_lut (.A(n29459), .B(index_q[2]), .C(index_q[3]), 
         .D(index_q[4]), .Z(n23351)) /* synthesis lut_function=(A (B)+!A (B (C (D))+!B !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i20869_3_lut_4_lut_4_lut_4_lut.init = 16'hc999;
    CCU2D unary_minus_10_add_3_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(quarter_wave_sample_register_i[0]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .COUT(n19698), .S1(o_val_pipeline_i_0__15__N_1799[0]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam unary_minus_10_add_3_1.INIT0 = 16'hF000;
    defparam unary_minus_10_add_3_1.INIT1 = 16'h0aaa;
    defparam unary_minus_10_add_3_1.INJECT1_0 = "NO";
    defparam unary_minus_10_add_3_1.INJECT1_1 = "NO";
    LUT4 mux_206_Mux_10_i317_3_lut_3_lut_4_lut (.A(n29177), .B(index_i[3]), 
         .C(n29146), .D(index_i[4]), .Z(n317)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_10_i317_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 mux_206_Mux_0_i396_3_lut_4_lut_3_lut_rep_819 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n32020)) /* synthesis lut_function=(A ((C)+!B)+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i396_3_lut_4_lut_3_lut_rep_819.init = 16'hb6b6;
    LUT4 mux_206_Mux_1_i301_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n301)) /* synthesis lut_function=(A (B (C+(D))+!B !(D))+!A !(B (C+(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_1_i301_3_lut_4_lut_4_lut.init = 16'h99b6;
    LUT4 mux_206_Mux_0_i963_3_lut_3_lut_3_lut_rep_820 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n32021)) /* synthesis lut_function=(!(A (B)+!A (B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i963_3_lut_3_lut_3_lut_rep_820.init = 16'h3636;
    LUT4 n23195_bdd_3_lut_27008 (.A(n29391), .B(n29387), .C(index_q[3]), 
         .Z(n26652)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n23195_bdd_3_lut_27008.init = 16'hcaca;
    LUT4 mux_207_Mux_7_i475_3_lut_4_lut (.A(n29459), .B(index_q[2]), .C(index_q[3]), 
         .D(n29470), .Z(n475_adj_2987)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_7_i475_3_lut_4_lut.init = 16'h9f90;
    LUT4 i24310_3_lut (.A(n25072), .B(n28680), .C(index_q[6]), .Z(n25081)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24310_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_0_i747_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n747_adj_2988)) /* synthesis lut_function=(!(A (B+!(C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_0_i747_3_lut_4_lut_4_lut_4_lut.init = 16'h6556;
    LUT4 mux_207_Mux_6_i860_3_lut_3_lut (.A(n29063), .B(index_q[4]), .C(n844_adj_2989), 
         .Z(n860)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam mux_207_Mux_6_i860_3_lut_3_lut.init = 16'h7474;
    LUT4 n308_bdd_3_lut_27011 (.A(n29355), .B(n32033), .C(index_q[3]), 
         .Z(n26655)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n308_bdd_3_lut_27011.init = 16'hacac;
    LUT4 i21130_3_lut (.A(n32018), .B(n645), .C(index_i[3]), .Z(n23612)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21130_3_lut.init = 16'hcaca;
    LUT4 i20871_4_lut_4_lut_4_lut (.A(n29459), .B(index_q[2]), .C(index_q[4]), 
         .D(index_q[3]), .Z(n23353)) /* synthesis lut_function=(A (B)+!A !(B (C+(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i20871_4_lut_4_lut_4_lut.init = 16'h999c;
    LUT4 i11118_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(n29326), .D(index_q[4]), .Z(n221_adj_2990)) /* synthesis lut_function=(!(A (B)+!A (B (C+(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i11118_3_lut_4_lut_4_lut_4_lut.init = 16'h3336;
    LUT4 n201_bdd_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n28839)) /* synthesis lut_function=(!(A (D)+!A !(B (D)+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n201_bdd_4_lut_4_lut_4_lut.init = 16'h54bb;
    LUT4 mux_207_Mux_8_i46_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n46_adj_2991)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (D)+!B !(C (D)+!C !(D)))) */ ;
    defparam mux_207_Mux_8_i46_3_lut_4_lut_4_lut.init = 16'hcf10;
    LUT4 n29468_bdd_3_lut_27558 (.A(n29168), .B(n32033), .C(index_q[4]), 
         .Z(n29903)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n29468_bdd_3_lut_27558.init = 16'hcaca;
    LUT4 i21517_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n23999)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A (B (C (D)+!C !(D))+!B (D))) */ ;
    defparam i21517_3_lut_4_lut.init = 16'hd926;
    LUT4 mux_206_Mux_6_i204_3_lut_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n204)) /* synthesis lut_function=(!(A (C)+!A !((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_6_i204_3_lut_3_lut_3_lut.init = 16'h5b5b;
    LUT4 index_q_2__bdd_3_lut_27761 (.A(index_q[2]), .B(index_q[0]), .C(index_q[4]), 
         .Z(n29901)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B (C)+!B !(C)))) */ ;
    defparam index_q_2__bdd_3_lut_27761.init = 16'h6969;
    LUT4 index_q_2__bdd_4_lut_27760 (.A(index_q[2]), .B(index_q[0]), .C(index_q[4]), 
         .D(index_q[1]), .Z(n29900)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((C (D))+!B))) */ ;
    defparam index_q_2__bdd_4_lut_27760.init = 16'h0cec;
    LUT4 mux_206_Mux_0_i908_3_lut_4_lut (.A(index_i[0]), .B(n29400), .C(index_i[3]), 
         .D(n29439), .Z(n908_adj_2992)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (C+!(D)))) */ ;
    defparam mux_206_Mux_0_i908_3_lut_4_lut.init = 16'h2f20;
    LUT4 index_i_0__bdd_4_lut_27455 (.A(index_i[0]), .B(index_i[3]), .C(index_i[1]), 
         .D(index_i[2]), .Z(n29523)) /* synthesis lut_function=(A (B (C)+!B !(C+!(D)))+!A !(B ((D)+!C)+!B !(C (D)+!C !(D)))) */ ;
    defparam index_i_0__bdd_4_lut_27455.init = 16'h92c1;
    PFUMX i21830 (.BLUT(n31), .ALUT(n23976), .C0(index_i[5]), .Z(n24331));
    LUT4 i20836_3_lut_3_lut (.A(n29063), .B(index_q[4]), .C(n46_adj_2991), 
         .Z(n23318)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam i20836_3_lut_3_lut.init = 16'h7474;
    FD1P3AX phase_i_i0_i11 (.D(o_phase[11]), .SP(dac_clk_p_c_enable_630), 
            .CK(dac_clk_p_c), .Q(phase_i[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam phase_i_i0_i11.GSR = "DISABLED";
    LUT4 mux_207_Mux_2_i349_3_lut_3_lut (.A(index_q[0]), .B(index_q[4]), 
         .C(n348_adj_2993), .Z(n349_adj_2994)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_2_i349_3_lut_3_lut.init = 16'hd1d1;
    LUT4 mux_207_Mux_0_i716_3_lut (.A(n29394), .B(n32035), .C(index_q[3]), 
         .Z(n716_adj_2995)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_0_i716_3_lut.init = 16'hcaca;
    LUT4 i20635_3_lut (.A(n325_adj_2972), .B(n29446), .C(index_i[3]), 
         .Z(n23117)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20635_3_lut.init = 16'hcaca;
    LUT4 n26659_bdd_3_lut (.A(n26659), .B(n157), .C(index_q[4]), .Z(n26660)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n26659_bdd_3_lut.init = 16'hcaca;
    PFUMX i21831 (.BLUT(n94_adj_2996), .ALUT(n125), .C0(index_i[5]), .Z(n24332));
    LUT4 n557_bdd_3_lut_26430 (.A(n32025), .B(n32021), .C(index_i[3]), 
         .Z(n27400)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n557_bdd_3_lut_26430.init = 16'hcaca;
    LUT4 i23911_3_lut (.A(n23116), .B(n23117), .C(index_i[4]), .Z(n23118)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23911_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_0_i653_3_lut (.A(n29181), .B(n29336), .C(index_q[3]), 
         .Z(n653_adj_2997)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_0_i653_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_0_i731_3_lut_4_lut (.A(n29465), .B(index_q[2]), .C(index_q[3]), 
         .D(n29461), .Z(n731_adj_2998)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_0_i731_3_lut_4_lut.init = 16'h4f40;
    LUT4 mux_206_Mux_6_i860_3_lut_3_lut (.A(n29058), .B(index_i[4]), .C(n844_adj_2999), 
         .Z(n860_adj_3000)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam mux_206_Mux_6_i860_3_lut_3_lut.init = 16'h7474;
    LUT4 i21385_3_lut_3_lut (.A(n29058), .B(index_i[4]), .C(n109_adj_2961), 
         .Z(n23867)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam i21385_3_lut_3_lut.init = 16'h7474;
    LUT4 i20938_3_lut_4_lut (.A(n29465), .B(index_q[2]), .C(index_q[3]), 
         .D(n29391), .Z(n23420)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i20938_3_lut_4_lut.init = 16'hf404;
    LUT4 mux_207_Mux_0_i620_3_lut (.A(n29461), .B(n32034), .C(index_q[3]), 
         .Z(n620_adj_3001)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_0_i620_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_7_i77_3_lut_3_lut_rep_655 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29315)) /* synthesis lut_function=(A (B)+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_7_i77_3_lut_3_lut_rep_655.init = 16'h9c9c;
    PFUMX i21832 (.BLUT(n20003), .ALUT(n16258), .C0(index_i[5]), .Z(n24333));
    PFUMX i22319 (.BLUT(n24817), .ALUT(n24818), .C0(index_q[4]), .Z(n24820));
    L6MUX21 i21834 (.D0(n23985), .D1(n23988), .SD(index_i[5]), .Z(n24335));
    L6MUX21 i21835 (.D0(n23991), .D1(n23994), .SD(index_i[5]), .Z(n24336));
    PFUMX i21836 (.BLUT(n413), .ALUT(n444_adj_3002), .C0(index_i[5]), 
          .Z(n24337));
    FD1P3AX phase_i_i0_i10 (.D(o_phase[10]), .SP(dac_clk_p_c_enable_630), 
            .CK(dac_clk_p_c), .Q(phase_i[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam phase_i_i0_i10.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i9 (.D(o_phase[9]), .SP(dac_clk_p_c_enable_630), 
            .CK(dac_clk_p_c), .Q(phase_i[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam phase_i_i0_i9.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i8 (.D(o_phase[8]), .SP(dac_clk_p_c_enable_630), 
            .CK(dac_clk_p_c), .Q(phase_i[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam phase_i_i0_i8.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i7 (.D(o_phase[7]), .SP(dac_clk_p_c_enable_630), 
            .CK(dac_clk_p_c), .Q(phase_i[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam phase_i_i0_i7.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i6 (.D(o_phase[6]), .SP(dac_clk_p_c_enable_630), 
            .CK(dac_clk_p_c), .Q(phase_i[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam phase_i_i0_i6.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i5 (.D(o_phase[5]), .SP(dac_clk_p_c_enable_630), 
            .CK(dac_clk_p_c), .Q(phase_i[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam phase_i_i0_i5.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i4 (.D(o_phase[4]), .SP(dac_clk_p_c_enable_630), 
            .CK(dac_clk_p_c), .Q(phase_i[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam phase_i_i0_i4.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i3 (.D(o_phase[3]), .SP(dac_clk_p_c_enable_630), 
            .CK(dac_clk_p_c), .Q(phase_i[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam phase_i_i0_i3.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i2 (.D(o_phase[2]), .SP(dac_clk_p_c_enable_630), 
            .CK(dac_clk_p_c), .Q(phase_i[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam phase_i_i0_i2.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i1 (.D(o_phase[1]), .SP(dac_clk_p_c_enable_630), 
            .CK(dac_clk_p_c), .Q(phase_i[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam phase_i_i0_i1.GSR = "DISABLED";
    LUT4 n442_bdd_3_lut_25676 (.A(n29432), .B(n32039), .C(index_i[3]), 
         .Z(n27414)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n442_bdd_3_lut_25676.init = 16'hcaca;
    LUT4 mux_207_Mux_0_i589_3_lut (.A(n29470), .B(n588), .C(index_q[3]), 
         .Z(n589)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_0_i589_3_lut.init = 16'hcaca;
    LUT4 i20721_3_lut (.A(n900), .B(n29446), .C(index_i[3]), .Z(n23203)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20721_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_7_i45_3_lut_3_lut_rep_656 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29316)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_7_i45_3_lut_3_lut_rep_656.init = 16'h3939;
    LUT4 mux_207_Mux_2_i731_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n731_adj_3003)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_2_i731_3_lut_4_lut_4_lut.init = 16'h6cc6;
    LUT4 n340_bdd_3_lut (.A(n32025), .B(n931), .C(index_i[3]), .Z(n27416)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n340_bdd_3_lut.init = 16'hacac;
    LUT4 i23836_3_lut (.A(n29578), .B(n23201), .C(index_i[4]), .Z(n23202)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23836_3_lut.init = 16'hcaca;
    PFUMX i27141 (.BLUT(n29585), .ALUT(n29586), .C0(index_i[0]), .Z(n29587));
    LUT4 i20632_3_lut (.A(n29444), .B(n32020), .C(index_i[3]), .Z(n23114)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20632_3_lut.init = 16'hcaca;
    LUT4 i21403_3_lut_4_lut (.A(n29418), .B(index_i[3]), .C(index_i[4]), 
         .D(n635_adj_3004), .Z(n23885)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21403_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_206_Mux_8_i542_3_lut_4_lut (.A(n29418), .B(index_i[3]), .C(index_i[4]), 
         .D(n526_adj_3005), .Z(n542)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_8_i542_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_207_Mux_2_i189_3_lut_3_lut_4_lut (.A(index_q[1]), .B(n29326), 
         .C(n173), .D(index_q[4]), .Z(n189_adj_3006)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(C+(D)))) */ ;
    defparam mux_207_Mux_2_i189_3_lut_3_lut_4_lut.init = 16'h77f0;
    LUT4 i12587_2_lut_3_lut_4_lut (.A(index_q[1]), .B(n29326), .C(index_q[5]), 
         .D(index_q[4]), .Z(n508)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;
    defparam i12587_2_lut_3_lut_4_lut.init = 16'hf080;
    PFUMX i21837 (.BLUT(n476_adj_3007), .ALUT(n507_adj_3008), .C0(index_i[5]), 
          .Z(n24338));
    LUT4 mux_207_Mux_8_i763_3_lut_4_lut (.A(n29465), .B(n29361), .C(index_q[4]), 
         .D(n29133), .Z(n16858)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam mux_207_Mux_8_i763_3_lut_4_lut.init = 16'hfe0e;
    LUT4 mux_206_Mux_6_i475_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n475_adj_3009)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A !(B (C+(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_6_i475_3_lut_4_lut_4_lut.init = 16'h9936;
    LUT4 n698_bdd_3_lut_25743 (.A(n29439), .B(n619), .C(index_i[3]), .Z(n27466)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n698_bdd_3_lut_25743.init = 16'hcaca;
    LUT4 n994_bdd_3_lut_25732 (.A(n29437), .B(n32021), .C(index_i[3]), 
         .Z(n27483)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n994_bdd_3_lut_25732.init = 16'hacac;
    LUT4 i20653_3_lut_4_lut (.A(n29379), .B(index_i[2]), .C(index_i[3]), 
         .D(n851), .Z(n23135)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20653_3_lut_4_lut.init = 16'hf202;
    LUT4 i21418_3_lut_4_lut_4_lut_4_lut (.A(index_i[2]), .B(n29379), .C(index_i[3]), 
         .D(index_i[4]), .Z(n23900)) /* synthesis lut_function=(A (B+(C (D)))+!A !(B+(C (D)))) */ ;
    defparam i21418_3_lut_4_lut_4_lut_4_lut.init = 16'ha999;
    LUT4 mux_206_Mux_2_i684_3_lut_4_lut (.A(index_i[2]), .B(n29379), .C(index_i[3]), 
         .D(n32056), .Z(n684_adj_3010)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;
    defparam mux_206_Mux_2_i684_3_lut_4_lut.init = 16'h6f60;
    LUT4 n236_bdd_4_lut (.A(n29088), .B(index_i[4]), .C(n28360), .D(index_i[5]), 
         .Z(n29026)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (B (C (D))+!B (C+!(D)))) */ ;
    defparam n236_bdd_4_lut.init = 16'hf099;
    LUT4 mux_206_Mux_7_i475_3_lut_4_lut (.A(index_i[2]), .B(n29379), .C(index_i[3]), 
         .D(n32019), .Z(n475_adj_3011)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+(D)))) */ ;
    defparam mux_206_Mux_7_i475_3_lut_4_lut.init = 16'h9f90;
    LUT4 i21472_3_lut_4_lut (.A(index_i[2]), .B(n29379), .C(index_i[3]), 
         .D(n29406), .Z(n23954)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;
    defparam i21472_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_206_Mux_7_i653_3_lut_4_lut (.A(index_i[2]), .B(n29379), .C(index_i[3]), 
         .D(n29377), .Z(n653_adj_3012)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam mux_206_Mux_7_i653_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_206_Mux_6_i435_3_lut_4_lut_3_lut_rep_764 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29424)) /* synthesis lut_function=(A (B+!(C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_6_i435_3_lut_4_lut_3_lut_rep_764.init = 16'hdbdb;
    LUT4 n557_bdd_4_lut (.A(n29079), .B(index_q[4]), .C(n28281), .D(index_q[5]), 
         .Z(n29028)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (B (C (D))+!B (C+!(D)))) */ ;
    defparam n557_bdd_4_lut.init = 16'hf099;
    PFUMX i21838 (.BLUT(n20017), .ALUT(n573), .C0(index_i[5]), .Z(n24339));
    LUT4 i21420_4_lut_4_lut_4_lut (.A(index_i[2]), .B(n29379), .C(index_i[4]), 
         .D(index_i[3]), .Z(n23902)) /* synthesis lut_function=(A (B+!(C+(D)))+!A !(B+!(C+(D)))) */ ;
    defparam i21420_4_lut_4_lut_4_lut.init = 16'h999a;
    LUT4 mux_207_Mux_2_i604_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n604_adj_3013)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)+!C !(D)))+!A (B (D)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_2_i604_3_lut_4_lut_4_lut_4_lut.init = 16'h39cf;
    PFUMX i21839 (.BLUT(n605), .ALUT(n636), .C0(index_i[5]), .Z(n24340));
    PFUMX i21840 (.BLUT(n23997), .ALUT(n700), .C0(index_i[5]), .Z(n24341));
    LUT4 mux_207_Mux_2_i573_3_lut_3_lut_4_lut (.A(n29367), .B(index_q[3]), 
         .C(n557_adj_3014), .D(index_q[4]), .Z(n573_adj_3015)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_2_i573_3_lut_3_lut_4_lut.init = 16'h11f0;
    LUT4 i22237_3_lut_4_lut (.A(n29367), .B(index_q[3]), .C(index_q[4]), 
         .D(n285_adj_2941), .Z(n24738)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i22237_3_lut_4_lut.init = 16'hfe0e;
    LUT4 mux_207_Mux_10_i125_3_lut_4_lut_4_lut (.A(n29367), .B(index_q[3]), 
         .C(index_q[4]), .D(n29168), .Z(n125_adj_3016)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B (C (D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_10_i125_3_lut_4_lut_4_lut.init = 16'h3efe;
    LUT4 i21522_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n24004)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A !(B (C+!(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21522_3_lut_4_lut_4_lut.init = 16'ha52b;
    LUT4 n698_bdd_3_lut_26959 (.A(n29385), .B(n29438), .C(index_i[3]), 
         .Z(n27511)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n698_bdd_3_lut_26959.init = 16'hcaca;
    L6MUX21 i21841 (.D0(n732_adj_3017), .D1(n24000), .SD(index_i[5]), 
            .Z(n24342));
    PFUMX i21842 (.BLUT(n797_adj_3018), .ALUT(n828_adj_3019), .C0(index_i[5]), 
          .Z(n24343));
    LUT4 n124_bdd_3_lut_26558_4_lut (.A(n29367), .B(index_q[3]), .C(index_q[4]), 
         .D(n124), .Z(n28488)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam n124_bdd_3_lut_26558_4_lut.init = 16'hf101;
    LUT4 mux_207_Mux_4_i573_3_lut_3_lut_4_lut_4_lut (.A(n29367), .B(index_q[3]), 
         .C(index_q[4]), .D(n29204), .Z(n573_adj_3020)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_4_i573_3_lut_3_lut_4_lut_4_lut.init = 16'h1f1c;
    LUT4 mux_207_Mux_3_i573_3_lut_3_lut_4_lut (.A(n29367), .B(index_q[3]), 
         .C(n460), .D(index_q[4]), .Z(n573_adj_3021)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_3_i573_3_lut_3_lut_4_lut.init = 16'h11f0;
    PFUMX i21843 (.BLUT(n860_adj_3022), .ALUT(n891), .C0(index_i[5]), 
          .Z(n24344));
    PFUMX i22821 (.BLUT(n812_adj_3023), .ALUT(n13328), .C0(index_q[4]), 
          .Z(n25322));
    LUT4 index_i_1__bdd_4_lut_28653 (.A(index_i[1]), .B(index_i[3]), .C(index_i[0]), 
         .D(index_i[2]), .Z(n30203)) /* synthesis lut_function=(A (B (C+(D))+!B (C (D)))+!A !(B (C)+!B !(C+(D)))) */ ;
    defparam index_i_1__bdd_4_lut_28653.init = 16'hbd94;
    LUT4 i20880_3_lut_3_lut_4_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n23362)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B !((D)+!C)))) */ ;
    defparam i20880_3_lut_3_lut_4_lut_3_lut_4_lut.init = 16'h11ef;
    LUT4 n30203_bdd_3_lut (.A(n30203), .B(index_i[1]), .C(index_i[4]), 
         .Z(n30204)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n30203_bdd_3_lut.init = 16'hcaca;
    LUT4 i22728_3_lut_4_lut (.A(n29067), .B(n29066), .C(index_q[5]), .D(index_q[6]), 
         .Z(n25229)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (B+((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i22728_3_lut_4_lut.init = 16'hffc5;
    LUT4 i23547_3_lut (.A(n23197), .B(n23198), .C(index_q[4]), .Z(n23199)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23547_3_lut.init = 16'hcaca;
    PFUMX i22283 (.BLUT(n24780), .ALUT(n24781), .C0(index_i[5]), .Z(n24784));
    LUT4 i22705_3_lut_4_lut (.A(n29136), .B(n29068), .C(index_q[4]), .D(index_q[5]), 
         .Z(n25206)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (B+((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i22705_3_lut_4_lut.init = 16'hffc5;
    PFUMX i22284 (.BLUT(n24782), .ALUT(n24783), .C0(index_i[5]), .Z(n24785));
    LUT4 mux_207_Mux_3_i460_3_lut_4_lut (.A(n29330), .B(index_q[2]), .C(index_q[3]), 
         .D(n29395), .Z(n460_adj_3024)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_3_i460_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_207_Mux_6_i285_3_lut_4_lut (.A(n29330), .B(index_q[2]), .C(index_q[3]), 
         .D(n29390), .Z(n285_adj_3025)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_6_i285_3_lut_4_lut.init = 16'hf606;
    LUT4 i21129_3_lut (.A(n29384), .B(n851), .C(index_i[3]), .Z(n23611)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21129_3_lut.init = 16'hcaca;
    LUT4 i20899_3_lut_4_lut (.A(n29330), .B(index_q[2]), .C(index_q[3]), 
         .D(n29353), .Z(n23381)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i20899_3_lut_4_lut.init = 16'hf606;
    LUT4 i20590_3_lut_4_lut (.A(n29330), .B(index_q[2]), .C(index_q[3]), 
         .D(n29388), .Z(n23072)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i20590_3_lut_4_lut.init = 16'h6f60;
    LUT4 i14463_3_lut_4_lut (.A(n29329), .B(index_i[4]), .C(index_i[5]), 
         .D(n29379), .Z(n16898)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i14463_3_lut_4_lut.init = 16'hf8f0;
    PFUMX i22823 (.BLUT(n875_adj_3026), .ALUT(n890_adj_2979), .C0(index_q[4]), 
          .Z(n25324));
    LUT4 mux_206_Mux_6_i285_3_lut_4_lut (.A(n29420), .B(index_i[2]), .C(index_i[3]), 
         .D(n29437), .Z(n285_adj_3027)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_6_i285_3_lut_4_lut.init = 16'hf606;
    LUT4 i21511_3_lut_4_lut (.A(n29420), .B(index_i[2]), .C(index_i[3]), 
         .D(n32020), .Z(n23993)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21511_3_lut_4_lut.init = 16'h6f60;
    LUT4 i20719_3_lut_4_lut (.A(n29420), .B(index_i[2]), .C(index_i[3]), 
         .D(n29447), .Z(n23201)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20719_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_206_Mux_0_i364_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n364)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A ((C+!(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i364_3_lut_3_lut_4_lut.init = 16'hdb55;
    LUT4 mux_206_Mux_3_i460_3_lut_4_lut (.A(n29420), .B(index_i[2]), .C(index_i[3]), 
         .D(n29429), .Z(n460_adj_3028)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_3_i460_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_206_Mux_1_i700_3_lut_4_lut (.A(n29324), .B(index_i[3]), .C(index_i[4]), 
         .D(n684), .Z(n700_adj_3029)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_1_i700_3_lut_4_lut.init = 16'hefe0;
    LUT4 n77_bdd_3_lut_25818 (.A(n29390), .B(n29387), .C(index_q[3]), 
         .Z(n27572)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n77_bdd_3_lut_25818.init = 16'hacac;
    LUT4 i20713_3_lut (.A(n404), .B(n32036), .C(index_q[3]), .Z(n23195)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20713_3_lut.init = 16'hcaca;
    LUT4 i22671_4_lut_4_lut (.A(n29086), .B(n29178), .C(index_i[5]), .D(index_i[4]), 
         .Z(n25172)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C+(D))+!B !(C (D)+!C !(D)))) */ ;
    defparam i22671_4_lut_4_lut.init = 16'hcf50;
    LUT4 i20856_3_lut_4_lut_4_lut (.A(n29165), .B(index_q[4]), .C(index_q[3]), 
         .D(n29204), .Z(n23338)) /* synthesis lut_function=(A (B (C)+!B !(C+!(D)))+!A (B (C)+!B (C+(D)))) */ ;
    defparam i20856_3_lut_4_lut_4_lut.init = 16'hd3d0;
    PFUMX i21862 (.BLUT(n94_adj_3030), .ALUT(n24003), .C0(index_i[5]), 
          .Z(n24363));
    LUT4 i20710_3_lut (.A(n404), .B(n29356), .C(index_q[3]), .Z(n23192)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20710_3_lut.init = 16'hcaca;
    LUT4 i20709_3_lut (.A(n29335), .B(n325), .C(index_q[3]), .Z(n23191)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20709_3_lut.init = 16'hcaca;
    LUT4 mux_206_Mux_0_i978_3_lut_3_lut_rep_821 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n32022)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i978_3_lut_3_lut_rep_821.init = 16'h6c6c;
    PFUMX i22824 (.BLUT(n908_adj_3031), .ALUT(n923), .C0(index_q[4]), 
          .Z(n25325));
    LUT4 n16806_bdd_3_lut_26427_4_lut (.A(n29376), .B(n29372), .C(index_i[5]), 
         .D(n29329), .Z(n28340)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;
    defparam n16806_bdd_3_lut_26427_4_lut.init = 16'hf101;
    LUT4 mux_206_Mux_8_i763_3_lut_4_lut (.A(n29376), .B(n29372), .C(index_i[4]), 
         .D(n29147), .Z(n16900)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam mux_206_Mux_8_i763_3_lut_4_lut.init = 16'hfe0e;
    LUT4 mux_206_Mux_0_i124_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n124_adj_3032)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A !(B (D)+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i124_3_lut_4_lut_4_lut.init = 16'h6c99;
    LUT4 mux_206_Mux_6_i891_3_lut (.A(n875_adj_3033), .B(n890_adj_3034), 
         .C(index_i[4]), .Z(n891_adj_3035)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_6_i891_3_lut.init = 16'hcaca;
    LUT4 mux_206_Mux_2_i189_3_lut_3_lut_4_lut (.A(index_i[1]), .B(n29329), 
         .C(n173_adj_2943), .D(index_i[4]), .Z(n189_adj_3036)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(C+(D)))) */ ;
    defparam mux_206_Mux_2_i189_3_lut_3_lut_4_lut.init = 16'h77f0;
    LUT4 n284_bdd_3_lut_25851 (.A(n29467), .B(n29331), .C(index_q[3]), 
         .Z(n27586)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n284_bdd_3_lut_25851.init = 16'hcaca;
    LUT4 i12840_2_lut_3_lut_4_lut (.A(index_i[1]), .B(n29329), .C(index_i[5]), 
         .D(index_i[4]), .Z(n508_adj_3037)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;
    defparam i12840_2_lut_3_lut_4_lut.init = 16'hf080;
    LUT4 i23916_3_lut (.A(n23110), .B(n23111), .C(index_i[4]), .Z(n23112)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23916_3_lut.init = 16'hcaca;
    LUT4 i12537_2_lut_3_lut_4_lut (.A(n29204), .B(n29369), .C(index_q[6]), 
         .D(index_q[5]), .Z(n254)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i12537_2_lut_3_lut_4_lut.init = 16'hfef0;
    LUT4 mux_206_Mux_6_i828_4_lut (.A(n812), .B(n14983), .C(index_i[4]), 
         .D(index_i[2]), .Z(n828_adj_3038)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_6_i828_4_lut.init = 16'hfaca;
    LUT4 mux_206_Mux_6_i797_3_lut (.A(n653_adj_3039), .B(n29041), .C(index_i[4]), 
         .Z(n797_adj_3040)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_6_i797_3_lut.init = 16'hcaca;
    PFUMX i21864 (.BLUT(n221_adj_3041), .ALUT(n252_adj_3042), .C0(index_i[5]), 
          .Z(n24365));
    LUT4 i1_3_lut_4_lut (.A(n29379), .B(n29329), .C(index_i[6]), .D(n29309), 
         .Z(n22131)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;
    defparam i1_3_lut_4_lut.init = 16'hfff8;
    LUT4 i22279_3_lut_4_lut (.A(n29400), .B(index_i[3]), .C(index_i[4]), 
         .D(n285_adj_3043), .Z(n24780)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i22279_3_lut_4_lut.init = 16'hfe0e;
    LUT4 n124_bdd_3_lut_26598_4_lut (.A(n29400), .B(index_i[3]), .C(index_i[4]), 
         .D(n124_adj_3044), .Z(n28534)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n124_bdd_3_lut_26598_4_lut.init = 16'hf101;
    LUT4 mux_206_Mux_2_i573_3_lut_3_lut_4_lut (.A(n29400), .B(index_i[3]), 
         .C(n557_adj_2963), .D(index_i[4]), .Z(n573_adj_3045)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_2_i573_3_lut_3_lut_4_lut.init = 16'h11f0;
    LUT4 mux_206_Mux_3_i573_3_lut_3_lut_4_lut (.A(n29400), .B(index_i[3]), 
         .C(n557), .D(index_i[4]), .Z(n573_adj_3046)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_3_i573_3_lut_3_lut_4_lut.init = 16'h11f0;
    LUT4 mux_206_Mux_6_i669_3_lut (.A(n653_adj_3047), .B(n668_adj_3048), 
         .C(index_i[4]), .Z(n669)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_6_i669_3_lut.init = 16'hcaca;
    PFUMX i21865 (.BLUT(n286), .ALUT(n24006), .C0(index_i[5]), .Z(n24366));
    LUT4 mux_206_Mux_10_i125_3_lut_4_lut_4_lut (.A(n29400), .B(index_i[3]), 
         .C(index_i[4]), .D(n29180), .Z(n125_adj_3049)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B (C (D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_10_i125_3_lut_4_lut_4_lut.init = 16'h3efe;
    LUT4 mux_206_Mux_4_i573_3_lut_3_lut_4_lut_4_lut (.A(n29400), .B(index_i[3]), 
         .C(index_i[4]), .D(n29176), .Z(n573_adj_3050)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_4_i573_3_lut_3_lut_4_lut_4_lut.init = 16'h1f1c;
    LUT4 mux_207_Mux_3_i859_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n859)) /* synthesis lut_function=(!(A (B (D)+!B !(D))+!A (B (C+(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_3_i859_3_lut_3_lut_4_lut.init = 16'h339c;
    PFUMX i21866 (.BLUT(n349), .ALUT(n24009), .C0(index_i[5]), .Z(n24367));
    LUT4 mux_206_Mux_0_i795_3_lut_3_lut_rep_822 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n32023)) /* synthesis lut_function=(A (B+(C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i795_3_lut_3_lut_rep_822.init = 16'hadad;
    LUT4 mux_207_Mux_2_i94_3_lut (.A(index_q[1]), .B(n124_adj_3051), .C(index_q[4]), 
         .Z(n94_adj_3052)) /* synthesis lut_function=(A (B (C))+!A (B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_2_i94_3_lut.init = 16'hc5c5;
    LUT4 i22474_3_lut (.A(n15_adj_3053), .B(n29486), .C(index_q[4]), .Z(n24975)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22474_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_5_i124_3_lut (.A(n29181), .B(n29463), .C(index_q[3]), 
         .Z(n124_adj_3051)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_5_i124_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_4_i668_3_lut_3_lut (.A(n29467), .B(index_q[3]), .C(n32055), 
         .Z(n668_adj_3054)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;
    defparam mux_207_Mux_4_i668_3_lut_3_lut.init = 16'hd1d1;
    LUT4 i14490_2_lut_rep_374_3_lut_4_lut (.A(n29095), .B(index_q[4]), .C(index_q[6]), 
         .D(index_q[5]), .Z(n29034)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i14490_2_lut_rep_374_3_lut_4_lut.init = 16'hf080;
    LUT4 index_i_0__bdd_4_lut_27073 (.A(index_i[0]), .B(index_i[3]), .C(index_i[1]), 
         .D(index_i[2]), .Z(n29477)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C))+!A (B (C (D)+!C !(D))+!B !(C+!(D))))) */ ;
    defparam index_i_0__bdd_4_lut_27073.init = 16'h16d3;
    LUT4 i14416_2_lut_3_lut_4_lut (.A(n29079), .B(index_q[4]), .C(index_q[6]), 
         .D(index_q[5]), .Z(n16844)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i14416_2_lut_3_lut_4_lut.init = 16'hfef0;
    LUT4 mux_207_Mux_7_i364_3_lut_3_lut (.A(n29467), .B(index_q[3]), .C(n29461), 
         .Z(n364_adj_3055)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;
    defparam mux_207_Mux_7_i364_3_lut_3_lut.init = 16'hd1d1;
    LUT4 i20644_3_lut_3_lut (.A(n29467), .B(index_q[3]), .C(n29373), .Z(n23126)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam i20644_3_lut_3_lut.init = 16'h7474;
    LUT4 index_q_1__bdd_4_lut_27850 (.A(index_q[1]), .B(index_q[3]), .C(index_q[0]), 
         .D(index_q[2]), .Z(n30466)) /* synthesis lut_function=(A (B (C+(D))+!B (C (D)))+!A !(B (C)+!B !(C+(D)))) */ ;
    defparam index_q_1__bdd_4_lut_27850.init = 16'hbd94;
    LUT4 n30466_bdd_3_lut (.A(n30466), .B(index_q[1]), .C(index_q[4]), 
         .Z(n30467)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n30466_bdd_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_10_i574_4_lut_4_lut (.A(n29079), .B(index_q[4]), .C(index_q[5]), 
         .D(n29080), .Z(n574_adj_3056)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_10_i574_4_lut_4_lut.init = 16'h1f1c;
    LUT4 i23814_3_lut (.A(n23215), .B(n23216), .C(index_i[4]), .Z(n23217)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23814_3_lut.init = 16'hcaca;
    PFUMX i21248 (.BLUT(n23728), .ALUT(n23729), .C0(index_q[5]), .Z(n23730));
    LUT4 mux_207_Mux_6_i844_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n844_adj_2989)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (B (C)+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_6_i844_3_lut_4_lut_4_lut.init = 16'hc1e0;
    LUT4 i20707_3_lut (.A(n32055), .B(n29464), .C(index_q[3]), .Z(n23189)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20707_3_lut.init = 16'hcaca;
    LUT4 mux_206_Mux_6_i542_3_lut (.A(n812_adj_3057), .B(n541_adj_3058), 
         .C(index_i[4]), .Z(n542_adj_3059)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_6_i542_3_lut.init = 16'hcaca;
    LUT4 n22_bdd_3_lut_25071 (.A(n29404), .B(n29437), .C(index_i[3]), 
         .Z(n26721)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n22_bdd_3_lut_25071.init = 16'hcaca;
    PFUMX i21871 (.BLUT(n669_adj_3060), .ALUT(n700_adj_3061), .C0(index_i[5]), 
          .Z(n24372));
    LUT4 i20730_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n23212)) /* synthesis lut_function=(!(A (B (C (D))+!B (C (D)+!C !(D)))+!A !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20730_3_lut_4_lut_4_lut.init = 16'h5aad;
    LUT4 i11138_3_lut_3_lut_4_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n762_adj_3062)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A (B))) */ ;
    defparam i11138_3_lut_3_lut_4_lut_3_lut_4_lut.init = 16'h1999;
    LUT4 mux_206_Mux_9_i62_3_lut_3_lut_4_lut_then_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[1]), .D(index_i[4]), .Z(n29534)) /* synthesis lut_function=(!(A (B+(C+!(D)))+!A !(B (D)+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_9_i62_3_lut_3_lut_4_lut_then_4_lut.init = 16'h5701;
    LUT4 mux_207_Mux_7_i379_3_lut_3_lut (.A(n29467), .B(index_q[3]), .C(n29470), 
         .Z(n379_adj_3063)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam mux_207_Mux_7_i379_3_lut_3_lut.init = 16'h7474;
    LUT4 i20706_3_lut (.A(n29467), .B(n85), .C(index_q[3]), .Z(n23188)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20706_3_lut.init = 16'hcaca;
    LUT4 i23692_3_lut (.A(n23188), .B(n23189), .C(index_q[4]), .Z(n23190)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23692_3_lut.init = 16'hcaca;
    LUT4 i20704_3_lut (.A(n29335), .B(n29356), .C(index_q[3]), .Z(n23186)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20704_3_lut.init = 16'hcaca;
    LUT4 i20703_3_lut (.A(n325), .B(n332), .C(index_q[3]), .Z(n23185)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20703_3_lut.init = 16'hcaca;
    LUT4 i20620_3_lut (.A(n29335), .B(n29389), .C(index_q[3]), .Z(n23102)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20620_3_lut.init = 16'hcaca;
    LUT4 i20619_3_lut (.A(n29357), .B(n325), .C(index_q[3]), .Z(n23101)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20619_3_lut.init = 16'hcaca;
    LUT4 mux_206_Mux_6_i252_4_lut (.A(index_i[2]), .B(n251_adj_3064), .C(index_i[4]), 
         .D(n12265), .Z(n252_adj_3065)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_6_i252_4_lut.init = 16'hc5ca;
    LUT4 i23774_3_lut (.A(n23101), .B(n23102), .C(index_q[4]), .Z(n23103)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23774_3_lut.init = 16'hcaca;
    LUT4 i24040_3_lut (.A(n28840), .B(n252_adj_3065), .C(index_i[5]), 
         .Z(n25285)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24040_3_lut.init = 16'hcaca;
    LUT4 index_i_5__bdd_3_lut_28422 (.A(index_i[5]), .B(n30579), .C(index_i[3]), 
         .Z(n30580)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam index_i_5__bdd_3_lut_28422.init = 16'hcaca;
    LUT4 n29379_bdd_3_lut_28489 (.A(n29177), .B(index_i[6]), .C(index_i[5]), 
         .Z(n30581)) /* synthesis lut_function=(!(A (B)+!A (C))) */ ;
    defparam n29379_bdd_3_lut_28489.init = 16'h2727;
    LUT4 mux_206_Mux_7_i506_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n506)) /* synthesis lut_function=(!(A (D)+!A (B ((D)+!C)+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_7_i506_3_lut_4_lut_4_lut_4_lut.init = 16'h01ea;
    LUT4 mux_206_Mux_0_i986_3_lut (.A(n32022), .B(n985), .C(index_i[3]), 
         .Z(n986)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i986_3_lut.init = 16'hcaca;
    LUT4 mux_206_Mux_0_i971_3_lut (.A(n32021), .B(n29382), .C(index_i[3]), 
         .Z(n971)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i971_3_lut.init = 16'hcaca;
    LUT4 n953_bdd_3_lut_25076 (.A(n29403), .B(index_i[3]), .C(n29440), 
         .Z(n26725)) /* synthesis lut_function=(A (B+(C))+!A !(B+!(C))) */ ;
    defparam n953_bdd_3_lut_25076.init = 16'hb8b8;
    LUT4 index_i_6__bdd_4_lut_27884 (.A(index_i[6]), .B(index_i[5]), .C(index_i[1]), 
         .D(index_i[0]), .Z(n30578)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C))+!A (B (C)+!B !(C)))) */ ;
    defparam index_i_6__bdd_4_lut_27884.init = 16'h3cbc;
    LUT4 i1_3_lut_rep_440_4_lut (.A(index_i[2]), .B(index_i[3]), .C(index_i[4]), 
         .D(n29376), .Z(n29100)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_3_lut_rep_440_4_lut.init = 16'hfffe;
    LUT4 index_i_6__bdd_1_lut_28205 (.A(index_i[5]), .Z(n30577)) /* synthesis lut_function=(!(A)) */ ;
    defparam index_i_6__bdd_1_lut_28205.init = 16'h5555;
    LUT4 n29379_bdd_4_lut_28088 (.A(n29379), .B(index_i[6]), .C(index_i[2]), 
         .D(index_i[5]), .Z(n30582)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A !(B (C+(D))+!B (D)))) */ ;
    defparam n29379_bdd_4_lut_28088.init = 16'h5fe0;
    LUT4 mux_206_Mux_5_i308_3_lut_4_lut_3_lut_rep_823 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n32024)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_5_i308_3_lut_4_lut_3_lut_rep_823.init = 16'h4d4d;
    LUT4 n30583_bdd_3_lut (.A(n30583), .B(n30580), .C(index_i[4]), .Z(n30584)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n30583_bdd_3_lut.init = 16'hcaca;
    PFUMX i21872 (.BLUT(n23064), .ALUT(n763_adj_2985), .C0(index_i[5]), 
          .Z(n24373));
    LUT4 mux_206_Mux_0_i939_4_lut (.A(n931), .B(n29185), .C(index_i[3]), 
         .D(index_i[2]), .Z(n939)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i939_4_lut.init = 16'hfaca;
    LUT4 i20665_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n23147)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D))+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20665_3_lut_4_lut.init = 16'hccdb;
    LUT4 i11120_3_lut_4_lut (.A(n29334), .B(index_q[2]), .C(n29360), .D(n29392), 
         .Z(n444_adj_3066)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i11120_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_206_Mux_0_i923_3_lut (.A(n29409), .B(n32019), .C(index_i[3]), 
         .Z(n923_adj_3067)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i923_3_lut.init = 16'hcaca;
    LUT4 i20934_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n23416)) /* synthesis lut_function=(A (B (C)+!B (C (D)+!C !(D)))+!A !(B (C+!(D))+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i20934_3_lut_4_lut_4_lut.init = 16'ha593;
    LUT4 mux_207_Mux_6_i157_3_lut_4_lut (.A(n29334), .B(index_q[2]), .C(index_q[3]), 
         .D(n29336), .Z(n157)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_6_i157_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_207_Mux_4_i747_3_lut_4_lut (.A(n29334), .B(index_q[2]), .C(index_q[3]), 
         .D(n29388), .Z(n747_adj_3068)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_4_i747_3_lut_4_lut.init = 16'hf606;
    PFUMX i21873 (.BLUT(n23070), .ALUT(n828_adj_3069), .C0(index_i[5]), 
          .Z(n24374));
    LUT4 mux_207_Mux_6_i251_3_lut_4_lut (.A(n29334), .B(index_q[2]), .C(index_q[3]), 
         .D(n29392), .Z(n251_adj_3070)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_6_i251_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_207_Mux_6_i891_3_lut (.A(n301_adj_3071), .B(n890_adj_3072), 
         .C(index_q[4]), .Z(n891_adj_3073)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_6_i891_3_lut.init = 16'hcaca;
    LUT4 n773_bdd_3_lut_24994_4_lut (.A(n29351), .B(index_q[2]), .C(n29396), 
         .D(index_q[3]), .Z(n26639)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam n773_bdd_3_lut_24994_4_lut.init = 16'hf066;
    LUT4 mux_207_Mux_6_i828_4_lut (.A(n812_adj_3074), .B(n15114), .C(index_q[4]), 
         .D(index_q[2]), .Z(n828_adj_3075)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_6_i828_4_lut.init = 16'hfaca;
    LUT4 mux_207_Mux_6_i797_3_lut (.A(n781), .B(n29039), .C(index_q[4]), 
         .Z(n797_adj_3076)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_6_i797_3_lut.init = 16'hcaca;
    LUT4 n285_bdd_3_lut_adj_179 (.A(n29403), .B(n32020), .C(index_i[3]), 
         .Z(n26728)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n285_bdd_3_lut_adj_179.init = 16'hacac;
    LUT4 i22308_3_lut_3_lut (.A(n29467), .B(index_q[3]), .C(n32055), .Z(n24809)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam i22308_3_lut_3_lut.init = 16'h7474;
    PFUMX i21874 (.BLUT(n860_adj_3077), .ALUT(n23076), .C0(index_i[5]), 
          .Z(n24375));
    LUT4 mux_206_Mux_9_i62_3_lut_3_lut_4_lut_else_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[1]), .D(index_i[4]), .Z(n29533)) /* synthesis lut_function=(A+(B (C+!(D))+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_9_i62_3_lut_3_lut_4_lut_else_4_lut.init = 16'heaff;
    LUT4 n262_bdd_3_lut_25967 (.A(n29471), .B(n32055), .C(index_q[3]), 
         .Z(n27747)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n262_bdd_3_lut_25967.init = 16'hcaca;
    LUT4 index_q_5__bdd_3_lut_28763 (.A(index_q[5]), .B(n30637), .C(index_q[3]), 
         .Z(n30638)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam index_q_5__bdd_3_lut_28763.init = 16'hcaca;
    LUT4 index_q_6__bdd_4_lut_27929 (.A(index_q[6]), .B(index_q[5]), .C(index_q[1]), 
         .D(index_q[0]), .Z(n30636)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C))+!A (B (C)+!B !(C)))) */ ;
    defparam index_q_6__bdd_4_lut_27929.init = 16'h3cbc;
    LUT4 index_q_6__bdd_1_lut_28564 (.A(index_q[5]), .Z(n30635)) /* synthesis lut_function=(!(A)) */ ;
    defparam index_q_6__bdd_1_lut_28564.init = 16'h5555;
    LUT4 mux_207_Mux_6_i669_3_lut (.A(n653_adj_3078), .B(n668_adj_3079), 
         .C(index_q[4]), .Z(n669_adj_3080)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_6_i669_3_lut.init = 16'hcaca;
    LUT4 n29459_bdd_3_lut_28327 (.A(n29165), .B(index_q[6]), .C(index_q[5]), 
         .Z(n30639)) /* synthesis lut_function=(!(A (B)+!A (C))) */ ;
    defparam n29459_bdd_3_lut_28327.init = 16'h2727;
    LUT4 n29459_bdd_4_lut_28224 (.A(n29459), .B(index_q[6]), .C(index_q[2]), 
         .D(index_q[5]), .Z(n30640)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A !(B (C+(D))+!B (D)))) */ ;
    defparam n29459_bdd_4_lut_28224.init = 16'h5fe0;
    LUT4 n30641_bdd_3_lut (.A(n30641), .B(n30638), .C(index_q[4]), .Z(n30642)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n30641_bdd_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_3_i668_3_lut_4_lut (.A(n29351), .B(index_q[2]), .C(index_q[3]), 
         .D(n29335), .Z(n668_adj_3081)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_3_i668_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_207_Mux_4_i763_3_lut_4_lut (.A(n29351), .B(index_q[2]), .C(index_q[4]), 
         .D(n747_adj_3068), .Z(n763_adj_3082)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_4_i763_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_206_Mux_0_i716_3_lut (.A(n29430), .B(n29445), .C(index_i[3]), 
         .Z(n716_adj_3083)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i716_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_6_i542_3_lut (.A(n526_adj_2957), .B(n541_adj_3084), 
         .C(index_q[4]), .Z(n542_adj_3085)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_6_i542_3_lut.init = 16'hcaca;
    LUT4 n23269_bdd_3_lut_26845 (.A(n29036), .B(n701), .C(index_q[6]), 
         .Z(n27756)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n23269_bdd_3_lut_26845.init = 16'hacac;
    LUT4 mux_207_Mux_6_i252_4_lut (.A(index_q[2]), .B(n251_adj_3070), .C(index_q[4]), 
         .D(n12338), .Z(n252_adj_3086)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_6_i252_4_lut.init = 16'hc5ca;
    L6MUX21 i22306 (.D0(n24805), .D1(n24806), .SD(index_q[5]), .Z(n24807));
    LUT4 i24073_3_lut (.A(n28803), .B(n252_adj_3086), .C(index_q[5]), 
         .Z(n25194)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24073_3_lut.init = 16'hcaca;
    LUT4 mux_206_Mux_0_i653_3_lut (.A(n645), .B(n32028), .C(index_i[3]), 
         .Z(n653_adj_3087)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i653_3_lut.init = 16'hcaca;
    LUT4 n27759_bdd_3_lut (.A(n31750), .B(n25243), .C(index_q[8]), .Z(n27760)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n27759_bdd_3_lut.init = 16'hcaca;
    LUT4 i7126_2_lut (.A(phase_i[0]), .B(phase_i[10]), .Z(index_i_9__N_1748[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(60[14] 63[8])
    defparam i7126_2_lut.init = 16'h6666;
    LUT4 i24488_2_lut (.A(phase_i[0]), .B(phase_i[10]), .Z(index_q_9__N_1758[0])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(60[14] 63[8])
    defparam i24488_2_lut.init = 16'h9999;
    PFUMX i21893 (.BLUT(n94), .ALUT(n125_adj_3088), .C0(index_i[5]), .Z(n24394));
    LUT4 mux_206_Mux_0_i620_3_lut (.A(n32018), .B(n29442), .C(index_i[3]), 
         .Z(n620_adj_3089)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i620_3_lut.init = 16'hcaca;
    LUT4 i21477_3_lut_3_lut_4_lut (.A(n29465), .B(index_q[2]), .C(n29181), 
         .D(index_q[3]), .Z(n23959)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (B (C (D))+!B (C+!(D)))) */ ;
    defparam i21477_3_lut_3_lut_4_lut.init = 16'hf099;
    LUT4 mux_206_Mux_0_i589_3_lut (.A(n32019), .B(n931), .C(index_i[3]), 
         .Z(n589_adj_3090)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i589_3_lut.init = 16'hcaca;
    LUT4 i20715_3_lut_3_lut_4_lut (.A(n29465), .B(index_q[2]), .C(n29460), 
         .D(index_q[3]), .Z(n23197)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (B (C (D))+!B (C+!(D)))) */ ;
    defparam i20715_3_lut_3_lut_4_lut.init = 16'hf099;
    LUT4 i20608_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n23090)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A (B (C (D)+!C !(D))+!B (D))) */ ;
    defparam i20608_3_lut_4_lut.init = 16'hd926;
    LUT4 i14133_2_lut (.A(index_i[1]), .B(index_i[3]), .Z(n541_adj_3091)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i14133_2_lut.init = 16'h1111;
    LUT4 mux_206_Mux_0_i526_3_lut (.A(n29441), .B(n29429), .C(index_i[3]), 
         .Z(n526_adj_3092)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i526_3_lut.init = 16'hcaca;
    PFUMX i21894 (.BLUT(n158_adj_3093), .ALUT(n189_adj_3094), .C0(index_i[5]), 
          .Z(n24395));
    LUT4 n23287_bdd_3_lut_26832 (.A(n29038), .B(n701_adj_3095), .C(index_i[6]), 
         .Z(n27781)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n23287_bdd_3_lut_26832.init = 16'hacac;
    LUT4 mux_207_Mux_4_i507_3_lut_3_lut_4_lut (.A(n29465), .B(index_q[2]), 
         .C(n491_adj_3096), .D(index_q[4]), .Z(n507_adj_3097)) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))+!A !(B ((D)+!C)+!B !(C+(D)))) */ ;
    defparam mux_207_Mux_4_i507_3_lut_3_lut_4_lut.init = 16'h99f0;
    LUT4 mux_207_Mux_3_i860_3_lut_4_lut (.A(n29465), .B(index_q[2]), .C(index_q[4]), 
         .D(n859), .Z(n860_adj_3098)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam mux_207_Mux_3_i860_3_lut_4_lut.init = 16'hf606;
    LUT4 n27784_bdd_3_lut (.A(n31713), .B(n25169), .C(index_i[8]), .Z(n27785)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n27784_bdd_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_7_i443_3_lut_4_lut (.A(n29465), .B(index_q[2]), .C(index_q[3]), 
         .D(n29460), .Z(n443_adj_3099)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;
    defparam mux_207_Mux_7_i443_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_207_Mux_2_i700_3_lut_4_lut (.A(index_q[1]), .B(n29361), .C(index_q[4]), 
         .D(n684_adj_3100), .Z(n700_adj_3101)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_2_i700_3_lut_4_lut.init = 16'hefe0;
    PFUMX i21895 (.BLUT(n221_adj_3102), .ALUT(n252_adj_3103), .C0(index_i[5]), 
          .Z(n24396));
    LUT4 n254_bdd_4_lut_26824 (.A(index_i[5]), .B(index_i[3]), .C(index_i[6]), 
         .D(index_i[4]), .Z(n27805)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;
    defparam n254_bdd_4_lut_26824.init = 16'hf8f0;
    LUT4 mux_207_Mux_3_i1018_3_lut_4_lut (.A(index_q[1]), .B(n29361), .C(index_q[4]), 
         .D(n21714), .Z(n1018)) /* synthesis lut_function=(A (C+!(D))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_3_i1018_3_lut_4_lut.init = 16'he0ef;
    LUT4 mux_206_Mux_3_i653_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n653_adj_3104)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A !(B (D)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_3_i653_3_lut_4_lut_4_lut.init = 16'h4d99;
    LUT4 i12808_2_lut_3_lut_4_lut (.A(n29176), .B(n29374), .C(index_i[6]), 
         .D(index_i[5]), .Z(n254_adj_3105)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i12808_2_lut_3_lut_4_lut.init = 16'hfef0;
    PFUMX i21896 (.BLUT(n286_adj_3106), .ALUT(n23088), .C0(index_i[5]), 
          .Z(n24397));
    LUT4 n27810_bdd_3_lut (.A(n29559), .B(n27806), .C(index_i[7]), .Z(n27811)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n27810_bdd_3_lut.init = 16'hcaca;
    LUT4 i24093_3_lut (.A(n286_adj_3107), .B(n317), .C(index_i[5]), .Z(n25163)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24093_3_lut.init = 16'hcaca;
    PFUMX i21897 (.BLUT(n349_adj_3108), .ALUT(n23097), .C0(index_i[5]), 
          .Z(n24398));
    PFUMX i21898 (.BLUT(n413_adj_3109), .ALUT(n444_adj_3110), .C0(index_i[5]), 
          .Z(n24399));
    LUT4 mux_207_Mux_10_i637_3_lut_4_lut_4_lut (.A(n29166), .B(index_q[4]), 
         .C(index_q[5]), .D(n29079), .Z(n637)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_10_i637_3_lut_4_lut_4_lut.init = 16'h1f1c;
    L6MUX21 i22313 (.D0(n24812), .D1(n24813), .SD(index_q[5]), .Z(n24814));
    PFUMX i21899 (.BLUT(n476_adj_3111), .ALUT(n507_adj_3112), .C0(index_i[5]), 
          .Z(n24400));
    LUT4 index_i_7__bdd_4_lut_28182 (.A(index_i[7]), .B(n16828), .C(n28143), 
         .D(index_i[5]), .Z(n29029)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(B (C+(D))+!B !((D)+!C)))) */ ;
    defparam index_i_7__bdd_4_lut_28182.init = 16'h66f0;
    PFUMX i21900 (.BLUT(n23106), .ALUT(n573_adj_3046), .C0(index_i[5]), 
          .Z(n24401));
    LUT4 mux_207_Mux_5_i15_3_lut_3_lut (.A(n29373), .B(index_q[3]), .C(n29315), 
         .Z(n15_adj_3113)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam mux_207_Mux_5_i15_3_lut_3_lut.init = 16'h7474;
    LUT4 i22322_3_lut_3_lut (.A(n29373), .B(index_q[3]), .C(n29467), .Z(n24823)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;
    defparam i22322_3_lut_3_lut.init = 16'hd1d1;
    LUT4 i20643_3_lut_3_lut (.A(n29373), .B(index_q[3]), .C(n32055), .Z(n23125)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam i20643_3_lut_3_lut.init = 16'h7474;
    LUT4 n254_bdd_4_lut_26802 (.A(index_q[5]), .B(index_q[3]), .C(index_q[6]), 
         .D(index_q[4]), .Z(n27836)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;
    defparam n254_bdd_4_lut_26802.init = 16'hf8f0;
    LUT4 mux_207_Mux_0_i348_3_lut_4_lut_4_lut (.A(n29373), .B(index_q[3]), 
         .C(index_q[2]), .D(n29346), .Z(n348_adj_3114)) /* synthesis lut_function=(!(A ((C (D)+!C !(D))+!B)+!A (B (C (D)+!C !(D))))) */ ;
    defparam mux_207_Mux_0_i348_3_lut_4_lut_4_lut.init = 16'h1dd1;
    LUT4 mux_207_Mux_2_i684_3_lut_4_lut_4_lut (.A(n29373), .B(index_q[3]), 
         .C(index_q[2]), .D(n29459), .Z(n684_adj_3100)) /* synthesis lut_function=(!(A ((C (D)+!C !(D))+!B)+!A (B (C (D)+!C !(D))))) */ ;
    defparam mux_207_Mux_2_i684_3_lut_4_lut_4_lut.init = 16'h1dd1;
    PFUMX i21901 (.BLUT(n13369), .ALUT(n23112), .C0(index_i[5]), .Z(n24402));
    LUT4 mux_206_Mux_0_i627_3_lut_rep_824 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n32025)) /* synthesis lut_function=(A (B+!(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i627_3_lut_rep_824.init = 16'hdada;
    LUT4 n27841_bdd_3_lut (.A(n29553), .B(n27837), .C(index_q[7]), .Z(n27842)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n27841_bdd_3_lut.init = 16'hcaca;
    PFUMX i22325 (.BLUT(n24822), .ALUT(n24823), .C0(index_q[4]), .Z(n24826));
    LUT4 i22316_3_lut_3_lut (.A(n29373), .B(index_q[3]), .C(n108), .Z(n24817)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;
    defparam i22316_3_lut_3_lut.init = 16'hd1d1;
    LUT4 mux_206_Mux_0_i173_3_lut_4_lut (.A(n29375), .B(index_i[1]), .C(index_i[3]), 
         .D(n29441), .Z(n173_adj_3115)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i173_3_lut_4_lut.init = 16'hdfd0;
    LUT4 mux_206_Mux_1_i620_3_lut_4_lut (.A(n29375), .B(index_i[1]), .C(index_i[3]), 
         .D(n29442), .Z(n620_adj_3116)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_1_i620_3_lut_4_lut.init = 16'hdfd0;
    PFUMX i21902 (.BLUT(n669_adj_3117), .ALUT(n700_adj_3118), .C0(index_i[5]), 
          .Z(n24403));
    LUT4 n638_bdd_3_lut_26772 (.A(n638), .B(n23316), .C(index_i[7]), .Z(n27860)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n638_bdd_3_lut_26772.init = 16'hcaca;
    L6MUX21 i21903 (.D0(n23115), .D1(n763_adj_3119), .SD(index_i[5]), 
            .Z(n24404));
    LUT4 i21502_3_lut_4_lut (.A(n29375), .B(index_i[1]), .C(index_i[3]), 
         .D(n498), .Z(n23984)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21502_3_lut_4_lut.init = 16'hdfd0;
    PFUMX i21905 (.BLUT(n860_adj_3120), .ALUT(n891_adj_3121), .C0(index_i[5]), 
          .Z(n24406));
    LUT4 i20617_3_lut (.A(n29396), .B(n29336), .C(index_q[3]), .Z(n23099)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20617_3_lut.init = 16'hcaca;
    PFUMX i22326 (.BLUT(n24824), .ALUT(n24825), .C0(index_q[4]), .Z(n24827));
    LUT4 n23310_bdd_3_lut_26055 (.A(n382), .B(n509), .C(index_i[7]), .Z(n27862)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n23310_bdd_3_lut_26055.init = 16'hcaca;
    LUT4 i23776_3_lut (.A(n23098), .B(n23099), .C(index_q[4]), .Z(n23100)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23776_3_lut.init = 16'hcaca;
    LUT4 n23945_bdd_3_lut_26539 (.A(n32022), .B(n32021), .C(index_i[3]), 
         .Z(n26741)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n23945_bdd_3_lut_26539.init = 16'hcaca;
    PFUMX i21906 (.BLUT(n924), .ALUT(n23118), .C0(index_i[5]), .Z(n24407));
    PFUMX i21907 (.BLUT(n23121), .ALUT(n1018_adj_3122), .C0(index_i[5]), 
          .Z(n24408));
    LUT4 mux_207_Mux_7_i890_3_lut_4_lut (.A(index_q[0]), .B(n29367), .C(index_q[3]), 
         .D(n29168), .Z(n890_adj_3123)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A !(C+(D))) */ ;
    defparam mux_207_Mux_7_i890_3_lut_4_lut.init = 16'h808f;
    LUT4 i17712_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), .C(index_i[4]), 
         .D(n29379), .Z(n286_adj_3107)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i17712_3_lut_4_lut.init = 16'hf0e0;
    LUT4 mux_207_Mux_7_i262_3_lut_rep_853 (.A(index_q[1]), .B(index_q[0]), 
         .C(index_q[2]), .Z(n32054)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_7_i262_3_lut_rep_853.init = 16'h5858;
    LUT4 i20592_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n23074)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20592_3_lut_4_lut_4_lut.init = 16'hda5a;
    LUT4 n459_bdd_3_lut_26542 (.A(n32024), .B(n29436), .C(index_i[3]), 
         .Z(n26744)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n459_bdd_3_lut_26542.init = 16'hacac;
    LUT4 index_q_4__bdd_3_lut_26239_4_lut (.A(n29167), .B(index_q[3]), .C(index_q[5]), 
         .D(index_q[4]), .Z(n28082)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam index_q_4__bdd_3_lut_26239_4_lut.init = 16'hf080;
    LUT4 i12821_2_lut_rep_372_3_lut_4_lut (.A(n29086), .B(index_i[4]), .C(index_i[6]), 
         .D(index_i[5]), .Z(n29032)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12821_2_lut_rep_372_3_lut_4_lut.init = 16'hf080;
    L6MUX21 i22320 (.D0(n24819), .D1(n24820), .SD(index_q[5]), .Z(n24821));
    LUT4 mux_206_Mux_4_i62_4_lut (.A(n29127), .B(n61), .C(index_i[4]), 
         .D(index_i[3]), .Z(n62_adj_3124)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_4_i62_4_lut.init = 16'hc5ca;
    LUT4 mux_206_Mux_4_i31_4_lut (.A(n15_adj_3125), .B(n29190), .C(index_i[4]), 
         .D(index_i[3]), .Z(n31_adj_3126)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_4_i31_4_lut.init = 16'h3aca;
    PFUMX i21925 (.BLUT(n158_adj_3127), .ALUT(n189_adj_3036), .C0(index_i[5]), 
          .Z(n24426));
    LUT4 mux_207_Mux_2_i142_3_lut_4_lut_4_lut_4_lut_4_lut (.A(index_q[0]), 
         .B(index_q[1]), .C(index_q[3]), .D(index_q[2]), .Z(n142)) /* synthesis lut_function=(!(A (B (D)+!B (C (D)+!C !(D)))+!A (B (D)+!B (C+!(D))))) */ ;
    defparam mux_207_Mux_2_i142_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'h03ec;
    PFUMX i21926 (.BLUT(n221_adj_3128), .ALUT(n23136), .C0(index_i[5]), 
          .Z(n24427));
    LUT4 n23310_bdd_3_lut (.A(n23310), .B(n30584), .C(index_i[7]), .Z(n27863)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n23310_bdd_3_lut.init = 16'hcaca;
    LUT4 i11252_3_lut_then_4_lut (.A(index_q[4]), .B(index_q[1]), .C(index_q[0]), 
         .D(index_q[2]), .Z(n29537)) /* synthesis lut_function=(A (B (C (D))+!B !(D))+!A (B (C+(D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i11252_3_lut_then_4_lut.init = 16'hd562;
    LUT4 i12584_3_lut_4_lut (.A(index_q[0]), .B(n29367), .C(n29369), .D(index_q[5]), 
         .Z(n318_adj_2938)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (C (D))) */ ;
    defparam i12584_3_lut_4_lut.init = 16'hf800;
    LUT4 i20916_3_lut_3_lut_4_lut (.A(index_q[0]), .B(n29367), .C(index_q[3]), 
         .D(n29167), .Z(n23398)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A !(C+(D))) */ ;
    defparam i20916_3_lut_3_lut_4_lut.init = 16'h808f;
    LUT4 n24380_bdd_3_lut_26070 (.A(n24380), .B(n24381), .C(index_i[7]), 
         .Z(n27878)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n24380_bdd_3_lut_26070.init = 16'hcaca;
    PFUMX i21927 (.BLUT(n286_adj_3129), .ALUT(n317_adj_3130), .C0(index_i[5]), 
          .Z(n24428));
    LUT4 mux_207_Mux_5_i987_4_lut_4_lut_4_lut (.A(index_q[0]), .B(n29367), 
         .C(index_q[4]), .D(index_q[3]), .Z(n21712)) /* synthesis lut_function=(A (B (C+!(D))+!B (D))+!A (B (C (D)+!C !(D))+!B (D))) */ ;
    defparam mux_207_Mux_5_i987_4_lut_4_lut_4_lut.init = 16'hf38c;
    LUT4 mux_207_Mux_8_i653_3_lut_rep_380_3_lut_4_lut (.A(index_q[0]), .B(n29367), 
         .C(n29204), .D(index_q[3]), .Z(n29040)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(C+(D)))) */ ;
    defparam mux_207_Mux_8_i653_3_lut_rep_380_3_lut_4_lut.init = 16'h77f0;
    LUT4 n24382_bdd_3_lut (.A(n24382), .B(n24383), .C(index_i[7]), .Z(n27876)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n24382_bdd_3_lut.init = 16'hcaca;
    LUT4 i20874_3_lut_3_lut_4_lut (.A(index_q[0]), .B(n29367), .C(n29167), 
         .D(index_q[3]), .Z(n23356)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(C+(D)))) */ ;
    defparam i20874_3_lut_3_lut_4_lut.init = 16'h77f0;
    LUT4 mux_207_Mux_0_i397_3_lut (.A(n29470), .B(n29388), .C(index_q[3]), 
         .Z(n397)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_0_i397_3_lut.init = 16'hcaca;
    LUT4 n24380_bdd_3_lut_28642 (.A(n24379), .B(n24378), .C(index_i[7]), 
         .Z(n27879)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n24380_bdd_3_lut_28642.init = 16'hacac;
    LUT4 n557_bdd_3_lut_4_lut_4_lut (.A(n29370), .B(index_q[3]), .C(index_q[4]), 
         .D(n29168), .Z(n28285)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C))+!A !(B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam n557_bdd_3_lut_4_lut_4_lut.init = 16'h838f;
    PFUMX i21928 (.BLUT(n349_adj_3131), .ALUT(n23139), .C0(index_i[5]), 
          .Z(n24429));
    LUT4 n638_bdd_3_lut_26766 (.A(n638_adj_3132), .B(n23298), .C(index_q[7]), 
         .Z(n27897)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n638_bdd_3_lut_26766.init = 16'hcaca;
    LUT4 i22239_3_lut_3_lut_4_lut_4_lut (.A(n29370), .B(index_q[3]), .C(index_q[4]), 
         .D(n29204), .Z(n24740)) /* synthesis lut_function=(!(A (B (C)+!B ((D)+!C))+!A (B+((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i22239_3_lut_3_lut_4_lut_4_lut.init = 16'h0838;
    PFUMX i21929 (.BLUT(n413_adj_3133), .ALUT(n23142), .C0(index_i[5]), 
          .Z(n24430));
    LUT4 n62_bdd_3_lut_4_lut (.A(n29370), .B(index_q[3]), .C(index_q[4]), 
         .D(n30), .Z(n28491)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam n62_bdd_3_lut_4_lut.init = 16'hf808;
    LUT4 n23292_bdd_3_lut_26088 (.A(n382_adj_3134), .B(n509_adj_3135), .C(index_q[7]), 
         .Z(n27899)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n23292_bdd_3_lut_26088.init = 16'hcaca;
    LUT4 i11090_3_lut_4_lut_4_lut (.A(n29370), .B(index_q[3]), .C(index_q[5]), 
         .D(n29165), .Z(n13386)) /* synthesis lut_function=(A (B+(C (D)))+!A (B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i11090_3_lut_4_lut_4_lut.init = 16'hf8c8;
    LUT4 n29468_bdd_2_lut_4_lut (.A(index_q[1]), .B(index_q[0]), .C(index_q[2]), 
         .D(index_q[4]), .Z(n29904)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam n29468_bdd_2_lut_4_lut.init = 16'h5800;
    LUT4 mux_206_Mux_3_i31_3_lut (.A(n653_adj_3039), .B(n30_adj_3136), .C(index_i[4]), 
         .Z(n31_adj_3137)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_3_i31_3_lut.init = 16'hcaca;
    PFUMX i21930 (.BLUT(n23145), .ALUT(n507_adj_3138), .C0(index_i[5]), 
          .Z(n24431));
    PFUMX i22825 (.BLUT(n939_adj_3139), .ALUT(n954_adj_3140), .C0(index_q[4]), 
          .Z(n25326));
    LUT4 mux_207_Mux_3_i252_3_lut_4_lut (.A(n29167), .B(index_q[3]), .C(index_q[4]), 
         .D(n16860), .Z(n252_adj_3141)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_3_i252_3_lut_4_lut.init = 16'h08f8;
    LUT4 i11108_3_lut (.A(n13403), .B(n29442), .C(index_i[3]), .Z(n13404)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11108_3_lut.init = 16'hcaca;
    LUT4 i11149_3_lut (.A(n13444), .B(n32034), .C(index_q[3]), .Z(n13445)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i11149_3_lut.init = 16'hcaca;
    PFUMX i21329 (.BLUT(n23809), .ALUT(n23810), .C0(index_q[5]), .Z(n23811));
    LUT4 mux_207_Mux_8_i475_3_lut_3_lut_4_lut (.A(n29371), .B(index_q[1]), 
         .C(index_q[3]), .D(n29168), .Z(n475_adj_3142)) /* synthesis lut_function=(A (C+!(D))+!A (B (C+!(D))+!B !(C+(D)))) */ ;
    defparam mux_207_Mux_8_i475_3_lut_3_lut_4_lut.init = 16'he0ef;
    PFUMX i22346 (.BLUT(n221_adj_2990), .ALUT(n252_adj_2949), .C0(index_q[5]), 
          .Z(n24847));
    LUT4 mux_207_Mux_9_i124_3_lut_3_lut_4_lut (.A(n29371), .B(index_q[1]), 
         .C(index_q[3]), .D(n29168), .Z(n124)) /* synthesis lut_function=(!(A (C (D))+!A (B (C (D))+!B ((D)+!C)))) */ ;
    defparam mux_207_Mux_9_i124_3_lut_3_lut_4_lut.init = 16'h0efe;
    PFUMX i21931 (.BLUT(n23148), .ALUT(n573_adj_3045), .C0(index_i[5]), 
          .Z(n24432));
    LUT4 n23292_bdd_3_lut (.A(n23292), .B(n30642), .C(index_q[7]), .Z(n27900)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n23292_bdd_3_lut.init = 16'hcaca;
    LUT4 n557_bdd_3_lut_26377_3_lut_4_lut (.A(n29371), .B(index_q[1]), .C(index_q[4]), 
         .D(index_q[3]), .Z(n28284)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B ((D)+!C))) */ ;
    defparam n557_bdd_3_lut_26377_3_lut_4_lut.init = 16'hf10f;
    LUT4 mux_207_Mux_0_i572_3_lut_4_lut (.A(n29371), .B(index_q[1]), .C(index_q[3]), 
         .D(n29387), .Z(n572_adj_3143)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam mux_207_Mux_0_i572_3_lut_4_lut.init = 16'hefe0;
    PFUMX i27137 (.BLUT(n29579), .ALUT(n29580), .C0(index_q[1]), .Z(n29581));
    LUT4 mux_206_Mux_0_i262_3_lut_3_lut_rep_818 (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[2]), .Z(n32019)) /* synthesis lut_function=(A ((C)+!B)+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i262_3_lut_3_lut_rep_818.init = 16'ha7a7;
    LUT4 mux_207_Mux_9_i364_3_lut_3_lut_4_lut (.A(n29371), .B(index_q[1]), 
         .C(index_q[3]), .D(n29204), .Z(n364_adj_3144)) /* synthesis lut_function=(!(A (C (D))+!A (B (C (D))+!B ((D)+!C)))) */ ;
    defparam mux_207_Mux_9_i364_3_lut_3_lut_4_lut.init = 16'h0efe;
    PFUMX i21932 (.BLUT(n605_adj_3145), .ALUT(n23151), .C0(index_i[5]), 
          .Z(n24433));
    LUT4 n24892_bdd_3_lut_26111 (.A(n24894), .B(n24893), .C(index_q[7]), 
         .Z(n27924)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n24892_bdd_3_lut_26111.init = 16'hacac;
    LUT4 n24892_bdd_3_lut_26762 (.A(n24892), .B(n24891), .C(index_q[7]), 
         .Z(n27925)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n24892_bdd_3_lut_26762.init = 16'hacac;
    LUT4 mux_207_Mux_10_i62_3_lut_3_lut_4_lut (.A(n29167), .B(index_q[3]), 
         .C(n29133), .D(index_q[4]), .Z(n62_adj_3146)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_10_i62_3_lut_3_lut_4_lut.init = 16'hf077;
    LUT4 i11089_4_lut_4_lut (.A(n29371), .B(index_q[1]), .C(index_q[3]), 
         .D(n22572), .Z(n13385)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A (B (C)+!B ((D)+!C)))) */ ;
    defparam i11089_4_lut_4_lut.init = 16'h0e3e;
    LUT4 n24902_bdd_3_lut (.A(n24895), .B(n24896), .C(index_q[7]), .Z(n27922)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n24902_bdd_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_3_i251_3_lut_4_lut (.A(n29371), .B(index_q[1]), .C(index_q[3]), 
         .D(n29204), .Z(n16860)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam mux_207_Mux_3_i251_3_lut_4_lut.init = 16'hfe0e;
    LUT4 i20853_4_lut_4_lut_3_lut_4_lut (.A(n29371), .B(index_q[1]), .C(index_q[4]), 
         .D(index_q[3]), .Z(n23335)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B !((D)+!C)))) */ ;
    defparam i20853_4_lut_4_lut_3_lut_4_lut.init = 16'h11ef;
    LUT4 i20661_3_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[0]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n23143)) /* synthesis lut_function=(A (B (C+(D))+!B !(D))+!A !(B (C+(D))+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20661_3_lut_4_lut_4_lut.init = 16'h99a7;
    LUT4 mux_207_Mux_6_i955_3_lut_4_lut (.A(n29167), .B(index_q[3]), .C(index_q[4]), 
         .D(n29040), .Z(n955)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_6_i955_3_lut_4_lut.init = 16'h8f80;
    LUT4 i14157_3_lut_rep_854 (.A(index_q[2]), .B(index_q[1]), .C(index_q[0]), 
         .Z(n32055)) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i14157_3_lut_rep_854.init = 16'hc4c4;
    PFUMX i21933 (.BLUT(n669_adj_3147), .ALUT(n700_adj_3148), .C0(index_i[5]), 
          .Z(n24434));
    LUT4 i20614_3_lut (.A(n29424), .B(n32028), .C(index_i[3]), .Z(n23096)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20614_3_lut.init = 16'hcaca;
    LUT4 i14249_2_lut_3_lut_4_lut (.A(n29088), .B(index_i[4]), .C(index_i[6]), 
         .D(index_i[5]), .Z(n16668)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i14249_2_lut_3_lut_4_lut.init = 16'hfef0;
    LUT4 i20613_3_lut (.A(n32021), .B(n29447), .C(index_i[3]), .Z(n23095)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20613_3_lut.init = 16'hcaca;
    LUT4 i23924_3_lut (.A(n23095), .B(n23096), .C(index_i[4]), .Z(n23097)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23924_3_lut.init = 16'hcaca;
    LUT4 i11104_3_lut_4_lut_4_lut (.A(index_q[2]), .B(index_q[1]), .C(index_q[0]), 
         .D(n29369), .Z(n605_adj_3149)) /* synthesis lut_function=(A (B (C)+!B !(C+!(D)))+!A (B (C+!(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i11104_3_lut_4_lut_4_lut.init = 16'hc3c4;
    LUT4 mux_206_Mux_10_i574_4_lut_4_lut (.A(n29088), .B(index_i[4]), .C(index_i[5]), 
         .D(n29089), .Z(n574_adj_3150)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_10_i574_4_lut_4_lut.init = 16'h1f1c;
    L6MUX21 i22327 (.D0(n24826), .D1(n24827), .SD(index_q[5]), .Z(n24828));
    PFUMX i21934 (.BLUT(n732_adj_3151), .ALUT(n763_adj_3152), .C0(index_i[5]), 
          .Z(n24435));
    LUT4 i12546_2_lut_rep_389_3_lut_4_lut (.A(n29371), .B(index_q[1]), .C(index_q[4]), 
         .D(index_q[3]), .Z(n29049)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i12546_2_lut_rep_389_3_lut_4_lut.init = 16'hfef0;
    LUT4 i11252_3_lut_else_4_lut (.A(index_q[4]), .B(index_q[1]), .C(index_q[0]), 
         .D(index_q[2]), .Z(n29536)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A !(B (D)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i11252_3_lut_else_4_lut.init = 16'ha955;
    LUT4 mux_206_Mux_4_i269_3_lut_4_lut_3_lut_rep_827 (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .Z(n32028)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_4_i269_3_lut_4_lut_3_lut_rep_827.init = 16'h1c1c;
    LUT4 i22776_4_lut_4_lut (.A(n29095), .B(n29166), .C(index_q[5]), .D(index_q[4]), 
         .Z(n25277)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C+(D))+!B !(C (D)+!C !(D)))) */ ;
    defparam i22776_4_lut_4_lut.init = 16'hcf50;
    LUT4 i21435_3_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[0]), 
         .D(index_i[3]), .Z(n23917)) /* synthesis lut_function=(!(A (B (C)+!B !(C (D)))+!A (B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21435_3_lut_4_lut_4_lut.init = 16'h3c1c;
    LUT4 mux_207_Mux_8_i860_3_lut_4_lut (.A(n29167), .B(index_q[3]), .C(index_q[4]), 
         .D(n29133), .Z(n860_adj_3153)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_8_i860_3_lut_4_lut.init = 16'h08f8;
    LUT4 i21478_3_lut_4_lut_4_lut (.A(index_q[2]), .B(index_q[1]), .C(index_q[0]), 
         .D(index_q[3]), .Z(n23960)) /* synthesis lut_function=(A (B (C)+!B !(C+!(D)))+!A (B (C+!(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i21478_3_lut_4_lut_4_lut.init = 16'hc3c4;
    LUT4 i22240_3_lut_4_lut (.A(n29167), .B(index_q[3]), .C(index_q[4]), 
         .D(n364_adj_3144), .Z(n24741)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i22240_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_207_Mux_0_i363_3_lut_4_lut_3_lut_rep_828 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n32029)) /* synthesis lut_function=(A (B+!(C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_0_i363_3_lut_4_lut_3_lut_rep_828.init = 16'hdbdb;
    LUT4 i11258_3_lut_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n13557)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A !(B (C+(D))+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i11258_3_lut_3_lut_4_lut_4_lut.init = 16'h44db;
    LUT4 i12676_3_lut_rep_855 (.A(index_i[2]), .B(index_i[1]), .C(index_i[0]), 
         .Z(n32056)) /* synthesis lut_function=(!(A (B)+!A (B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12676_3_lut_rep_855.init = 16'h2323;
    LUT4 mux_207_Mux_3_i189_3_lut_3_lut_4_lut (.A(n29167), .B(index_q[3]), 
         .C(index_q[4]), .D(n29130), .Z(n189_adj_3154)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_3_i189_3_lut_3_lut_4_lut.init = 16'h08f8;
    LUT4 i22643_3_lut (.A(n851), .B(n29406), .C(index_i[3]), .Z(n25144)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22643_3_lut.init = 16'hcaca;
    LUT4 n26651_bdd_3_lut_26728 (.A(n26651), .B(n25196), .C(index_q[6]), 
         .Z(n27977)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n26651_bdd_3_lut_26728.init = 16'hcaca;
    PFUMX i22826 (.BLUT(n971_adj_3155), .ALUT(n986_adj_3156), .C0(index_q[4]), 
          .Z(n25327));
    LUT4 mux_207_Mux_0_i1002_3_lut_3_lut_4_lut (.A(n29465), .B(index_q[2]), 
         .C(n29373), .D(index_q[3]), .Z(n1002)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_0_i1002_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 n26651_bdd_3_lut_26159 (.A(n25197), .B(n26657), .C(index_q[6]), 
         .Z(n27976)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n26651_bdd_3_lut_26159.init = 16'hcaca;
    LUT4 n26645_bdd_3_lut_26732 (.A(n26645), .B(n25192), .C(index_q[6]), 
         .Z(n27979)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n26645_bdd_3_lut_26732.init = 16'hcaca;
    LUT4 mux_207_Mux_5_i828_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[4]), .D(n29361), .Z(n828_adj_3157)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_5_i828_4_lut_4_lut.init = 16'hc66c;
    LUT4 mux_207_Mux_6_i890_3_lut_3_lut_4_lut (.A(n29465), .B(index_q[2]), 
         .C(n29471), .D(index_q[3]), .Z(n890_adj_3072)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_6_i890_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 mux_207_Mux_3_i93_3_lut_4_lut (.A(n29465), .B(index_q[2]), .C(index_q[3]), 
         .D(n29475), .Z(n93_adj_3158)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_3_i93_3_lut_4_lut.init = 16'hefe0;
    LUT4 i26521_then_3_lut (.A(index_i[0]), .B(index_i[4]), .C(index_i[3]), 
         .Z(n29540)) /* synthesis lut_function=(A (B)+!A (B (C)+!B !(C))) */ ;
    defparam i26521_then_3_lut.init = 16'hc9c9;
    LUT4 mux_206_Mux_4_i491_3_lut_4_lut (.A(n29376), .B(index_i[2]), .C(index_i[3]), 
         .D(n32018), .Z(n491_adj_3159)) /* synthesis lut_function=(A (C+(D))+!A !(B (C+!(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_4_i491_3_lut_4_lut.init = 16'hbfb0;
    LUT4 i20754_3_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[1]), .C(index_i[0]), 
         .D(index_i[3]), .Z(n23236)) /* synthesis lut_function=(!(A (B (D)+!B !(D))+!A (B+(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20754_3_lut_4_lut_4_lut.init = 16'h2388;
    LUT4 i22642_3_lut (.A(n619), .B(n32018), .C(index_i[3]), .Z(n25143)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22642_3_lut.init = 16'hcaca;
    LUT4 mux_206_Mux_2_i908_3_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[1]), 
         .C(index_i[0]), .D(index_i[3]), .Z(n908_adj_3160)) /* synthesis lut_function=(!(A (B)+!A !(B (D)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_2_i908_3_lut_4_lut_4_lut.init = 16'h6623;
    LUT4 i23613_3_lut (.A(n716_adj_3161), .B(n731_adj_3003), .C(index_q[4]), 
         .Z(n732_adj_3162)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23613_3_lut.init = 16'hcaca;
    LUT4 n61_bdd_3_lut_25979_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n27575)) /* synthesis lut_function=(!(A (B)+!A !(B (C+(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam n61_bdd_3_lut_25979_3_lut_4_lut_4_lut.init = 16'h6663;
    LUT4 index_q_7__bdd_4_lut_28247 (.A(index_q[7]), .B(n16798), .C(n28079), 
         .D(index_q[5]), .Z(n29031)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(B (C+(D))+!B !((D)+!C)))) */ ;
    defparam index_q_7__bdd_4_lut_28247.init = 16'h66f0;
    LUT4 mux_207_Mux_11_i638_4_lut_4_lut (.A(n29049), .B(index_q[5]), .C(index_q[6]), 
         .D(n29078), .Z(n638_adj_3163)) /* synthesis lut_function=(A (B (C (D))+!B !(C))+!A (B ((D)+!C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_11_i638_4_lut_4_lut.init = 16'hc707;
    LUT4 i22636_3_lut (.A(n29407), .B(n32019), .C(index_i[3]), .Z(n25137)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22636_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_2_i669_3_lut (.A(n653_adj_3164), .B(n475_adj_3165), 
         .C(index_q[4]), .Z(n669_adj_3166)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_2_i669_3_lut.init = 16'hcaca;
    PFUMX i22827 (.BLUT(n1002), .ALUT(n1017_adj_3167), .C0(index_q[4]), 
          .Z(n25328));
    LUT4 i22635_3_lut (.A(n32056), .B(n660), .C(index_i[3]), .Z(n25136)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22635_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_2_i605_3_lut (.A(n142_adj_3168), .B(n604_adj_3013), 
         .C(index_q[4]), .Z(n605_adj_3169)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_2_i605_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_3_i221_3_lut_4_lut (.A(n29168), .B(index_q[3]), .C(index_q[4]), 
         .D(n29134), .Z(n221_adj_3170)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_3_i221_3_lut_4_lut.init = 16'h08f8;
    LUT4 i20923_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n23405)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)+!C !(D)))+!A (B (C+!(D))+!B ((D)+!C)))) */ ;
    defparam i20923_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h0e30;
    PFUMX i21437 (.BLUT(n23917), .ALUT(n23918), .C0(index_i[4]), .Z(n23919));
    LUT4 i22634_3_lut (.A(n619), .B(n29385), .C(index_i[3]), .Z(n25135)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22634_3_lut.init = 16'hcaca;
    LUT4 i23619_3_lut (.A(n29518), .B(n23372), .C(index_q[4]), .Z(n23373)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23619_3_lut.init = 16'hcaca;
    LUT4 i22633_3_lut (.A(n645), .B(n29443), .C(index_i[3]), .Z(n25134)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22633_3_lut.init = 16'hcaca;
    LUT4 i23621_3_lut (.A(n23368), .B(n23369), .C(index_q[4]), .Z(n23370)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23621_3_lut.init = 16'hcaca;
    LUT4 mux_206_Mux_4_i507_3_lut_4_lut (.A(n29376), .B(index_i[2]), .C(index_i[4]), 
         .D(n491_adj_3159), .Z(n507_adj_3171)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_4_i507_3_lut_4_lut.init = 16'h9f90;
    LUT4 i21471_3_lut_3_lut_4_lut (.A(n29376), .B(index_i[2]), .C(n29409), 
         .D(index_i[3]), .Z(n23953)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21471_3_lut_3_lut_4_lut.init = 16'hf099;
    LUT4 n811_bdd_3_lut_25637_4_lut (.A(n29376), .B(index_i[2]), .C(index_i[3]), 
         .D(n29408), .Z(n27386)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n811_bdd_3_lut_25637_4_lut.init = 16'h9f90;
    LUT4 i20628_3_lut_3_lut_4_lut (.A(n29376), .B(index_i[2]), .C(n645), 
         .D(index_i[3]), .Z(n23110)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20628_3_lut_3_lut_4_lut.init = 16'hf099;
    LUT4 mux_206_Mux_3_i860_3_lut_4_lut (.A(n29376), .B(index_i[2]), .C(index_i[4]), 
         .D(n859_adj_3172), .Z(n860_adj_3120)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_3_i860_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_206_Mux_7_i443_3_lut_4_lut (.A(n29376), .B(index_i[2]), .C(index_i[3]), 
         .D(n29409), .Z(n443_adj_3173)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_7_i443_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_206_Mux_2_i700_3_lut_4_lut (.A(index_i[1]), .B(n29372), .C(index_i[4]), 
         .D(n684_adj_3010), .Z(n700_adj_3148)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_2_i700_3_lut_4_lut.init = 16'hefe0;
    LUT4 mux_206_Mux_3_i1018_3_lut_4_lut (.A(index_i[1]), .B(n29372), .C(index_i[4]), 
         .D(n21706), .Z(n1018_adj_3122)) /* synthesis lut_function=(A (C+!(D))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_3_i1018_3_lut_4_lut.init = 16'he0ef;
    LUT4 n954_bdd_3_lut_26227 (.A(n21704), .B(n29100), .C(index_i[5]), 
         .Z(n28073)) /* synthesis lut_function=(A (B (C))+!A (B+!(C))) */ ;
    defparam n954_bdd_3_lut_26227.init = 16'hc5c5;
    LUT4 mux_207_Mux_3_i157_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n157_adj_3174)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B !(C+(D))))) */ ;
    defparam mux_207_Mux_3_i157_3_lut_3_lut_4_lut.init = 16'h1ff0;
    LUT4 i24172_3_lut (.A(n30467), .B(n29571), .C(index_q[5]), .Z(n24889)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24172_3_lut.init = 16'hcaca;
    LUT4 i24176_3_lut (.A(n542_adj_3175), .B(n573_adj_3020), .C(index_q[5]), 
         .Z(n24883)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24176_3_lut.init = 16'hcaca;
    L6MUX21 i21936 (.D0(n860_adj_3176), .D1(n891_adj_3177), .SD(index_i[5]), 
            .Z(n24437));
    LUT4 i24179_3_lut (.A(n29574), .B(n444), .C(index_q[5]), .Z(n24881)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24179_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_1_i732_3_lut (.A(n716_adj_2945), .B(n491_adj_3178), 
         .C(index_q[4]), .Z(n732_adj_3179)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_1_i732_3_lut.init = 16'hcaca;
    LUT4 i26521_else_3_lut (.A(index_i[2]), .B(index_i[0]), .C(index_i[4]), 
         .D(index_i[3]), .Z(n29539)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)+!C !(D)))+!A (B (C+!(D))+!B !(C)))) */ ;
    defparam i26521_else_3_lut.init = 16'h1e38;
    LUT4 n924_bdd_3_lut_26617 (.A(n924_adj_3180), .B(n28075), .C(index_i[5]), 
         .Z(n28076)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n924_bdd_3_lut_26617.init = 16'hcaca;
    LUT4 i12554_3_lut_4_lut (.A(n29034), .B(index_q[7]), .C(index_q[8]), 
         .D(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_1783[14])) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (D))) */ ;
    defparam i12554_3_lut_4_lut.init = 16'hffe0;
    LUT4 index_q_4__bdd_4_lut_27750 (.A(index_q[4]), .B(n29161), .C(index_q[7]), 
         .D(n29134), .Z(n28079)) /* synthesis lut_function=(A ((C)+!B)+!A ((D)+!C)) */ ;
    defparam index_q_4__bdd_4_lut_27750.init = 16'hf7a7;
    LUT4 i20757_3_lut_3_lut_4_lut (.A(n29379), .B(index_i[2]), .C(n1001), 
         .D(index_i[3]), .Z(n23239)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20757_3_lut_3_lut_4_lut.init = 16'hf077;
    LUT4 mux_206_Mux_6_i939_3_lut_rep_382_3_lut_4_lut (.A(n29379), .B(index_i[2]), 
         .C(index_i[3]), .D(n29177), .Z(n29042)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_6_i939_3_lut_rep_382_3_lut_4_lut.init = 16'h08f8;
    LUT4 n316_bdd_3_lut (.A(n316_adj_3181), .B(n285_adj_3182), .C(index_i[5]), 
         .Z(n28100)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n316_bdd_3_lut.init = 16'hacac;
    LUT4 n28103_bdd_3_lut (.A(n28103), .B(n28102), .C(index_i[5]), .Z(n28104)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n28103_bdd_3_lut.init = 16'hcaca;
    LUT4 mux_206_Mux_7_i173_3_lut (.A(n29443), .B(n645), .C(index_i[3]), 
         .Z(n173_adj_2958)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_7_i173_3_lut.init = 16'hcaca;
    LUT4 mux_206_Mux_1_i317_3_lut (.A(n301), .B(n908_adj_3160), .C(index_i[4]), 
         .Z(n317_adj_3183)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_1_i317_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_2_i413_3_lut (.A(n397_adj_3184), .B(n954), .C(index_q[4]), 
         .Z(n413_adj_3185)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_2_i413_3_lut.init = 16'hcaca;
    LUT4 mux_206_Mux_6_i732_3_lut_4_lut (.A(n29385), .B(index_i[3]), .C(index_i[4]), 
         .D(n731_adj_3186), .Z(n732_adj_3187)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_6_i732_3_lut_4_lut.init = 16'hf909;
    LUT4 mux_206_Mux_6_i700_3_lut_4_lut (.A(n29385), .B(index_i[3]), .C(index_i[4]), 
         .D(n684_adj_3188), .Z(n700_adj_3189)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_6_i700_3_lut_4_lut.init = 16'h9f90;
    LUT4 i22475_3_lut_4_lut (.A(n29168), .B(index_q[3]), .C(index_q[4]), 
         .D(n46), .Z(n24976)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i22475_3_lut_4_lut.init = 16'h8f80;
    LUT4 i22476_3_lut_3_lut_4_lut (.A(n29168), .B(index_q[3]), .C(n93_adj_3190), 
         .D(index_q[4]), .Z(n24977)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i22476_3_lut_3_lut_4_lut.init = 16'hf077;
    PFUMX i20785 (.BLUT(n445_adj_2978), .ALUT(n508), .C0(index_q[6]), 
          .Z(n23267));
    LUT4 i24406_3_lut_rep_378_4_lut (.A(n29100), .B(index_i[5]), .C(index_i[8]), 
         .D(n1021), .Z(n29038)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i24406_3_lut_rep_378_4_lut.init = 16'hf808;
    LUT4 mux_206_Mux_6_i875_3_lut_4_lut (.A(n29379), .B(index_i[2]), .C(index_i[3]), 
         .D(n29377), .Z(n875_adj_3033)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_6_i875_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_207_Mux_2_i317_3_lut (.A(n668_adj_3081), .B(n316_adj_3191), 
         .C(index_q[4]), .Z(n317_adj_3192)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_2_i317_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_2_i286_3_lut (.A(n270), .B(n653_adj_3193), .C(index_q[4]), 
         .Z(n286_adj_3194)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_2_i286_3_lut.init = 16'hcaca;
    LUT4 n24437_bdd_3_lut (.A(n24437), .B(index_i[7]), .C(n27418), .Z(n28106)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n24437_bdd_3_lut.init = 16'he2e2;
    PFUMX i21440 (.BLUT(n23920), .ALUT(n23921), .C0(index_i[4]), .Z(n23922));
    LUT4 index_i_7__bdd_4_lut_26293 (.A(index_i[4]), .B(index_i[5]), .C(n908_adj_3160), 
         .D(n29522), .Z(n28107)) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C))) */ ;
    defparam index_i_7__bdd_4_lut_26293.init = 16'hdc10;
    LUT4 mux_206_Mux_1_i732_3_lut (.A(n716_adj_2982), .B(n491_adj_3195), 
         .C(index_i[4]), .Z(n732_adj_3196)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_1_i732_3_lut.init = 16'hcaca;
    LUT4 mux_206_Mux_8_i15_3_lut_4_lut (.A(n29379), .B(index_i[2]), .C(index_i[3]), 
         .D(n29408), .Z(n188)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_8_i15_3_lut_4_lut.init = 16'hf808;
    PFUMX i20591 (.BLUT(n23071), .ALUT(n23072), .C0(index_q[4]), .Z(n23073));
    LUT4 mux_206_Mux_3_i251_3_lut_4_lut (.A(n29379), .B(index_i[2]), .C(index_i[3]), 
         .D(n29179), .Z(n16610)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_3_i251_3_lut_4_lut.init = 16'h8f80;
    LUT4 n811_bdd_3_lut_4_lut (.A(n29379), .B(index_i[2]), .C(index_i[3]), 
         .D(n29177), .Z(n27387)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A !(C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n811_bdd_3_lut_4_lut.init = 16'h808f;
    LUT4 mux_206_Mux_6_i844_3_lut_4_lut (.A(n29379), .B(index_i[2]), .C(index_i[3]), 
         .D(n29380), .Z(n844_adj_2999)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_6_i844_3_lut_4_lut.init = 16'hf808;
    LUT4 i24214_3_lut (.A(n27391), .B(n23816), .C(index_q[5]), .Z(n23817)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24214_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut (.A(index_q[6]), .B(n29133), .C(index_q[5]), .D(index_q[4]), 
         .Z(n22201)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i1_4_lut.init = 16'hfffe;
    LUT4 i19370_4_lut (.A(n29360), .B(n892), .C(index_q[6]), .D(index_q[5]), 
         .Z(n21709)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D))))) */ ;
    defparam i19370_4_lut.init = 16'h3a35;
    LUT4 i24408_3_lut (.A(n21709), .B(n22201), .C(index_q[7]), .Z(n24458)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24408_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_6_i732_3_lut_4_lut (.A(n29467), .B(index_q[3]), .C(index_q[4]), 
         .D(n731), .Z(n732_adj_3197)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_6_i732_3_lut_4_lut.init = 16'hf909;
    LUT4 n28108_bdd_3_lut_26535 (.A(n28108), .B(n29587), .C(index_i[4]), 
         .Z(n28109)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n28108_bdd_3_lut_26535.init = 16'hcaca;
    LUT4 i12548_2_lut_rep_544_3_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .Z(n29204)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i12548_2_lut_rep_544_3_lut.init = 16'he0e0;
    LUT4 n28110_bdd_3_lut (.A(n28110), .B(n28106), .C(index_i[6]), .Z(n28111)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n28110_bdd_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_14_i511_4_lut_4_lut (.A(n29034), .B(index_q[7]), .C(index_q[8]), 
         .D(n254), .Z(n511)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (B (C+!(D))+!B !(C)))) */ ;
    defparam mux_207_Mux_14_i511_4_lut_4_lut.init = 16'h1c10;
    LUT4 mux_206_Mux_9_i364_3_lut_3_lut_4_lut (.A(n29379), .B(index_i[2]), 
         .C(n29179), .D(index_i[3]), .Z(n364_adj_3198)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_9_i364_3_lut_3_lut_4_lut.init = 16'h77f0;
    LUT4 n954_bdd_3_lut_26613_3_lut_4_lut (.A(n29379), .B(index_i[2]), .C(n29377), 
         .D(index_i[3]), .Z(n28074)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n954_bdd_3_lut_26613_3_lut_4_lut.init = 16'hf077;
    LUT4 index_i_4__bdd_4_lut_27751 (.A(index_i[4]), .B(n29173), .C(index_i[7]), 
         .D(n29143), .Z(n28143)) /* synthesis lut_function=(A ((C)+!B)+!A ((D)+!C)) */ ;
    defparam index_i_4__bdd_4_lut_27751.init = 16'hf7a7;
    LUT4 i24640_2_lut_rep_387_3_lut_4_lut (.A(n29379), .B(index_i[2]), .C(index_i[5]), 
         .D(n29374), .Z(n29047)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i24640_2_lut_rep_387_3_lut_4_lut.init = 16'h0f7f;
    LUT4 i24245_3_lut (.A(n30204), .B(n27467), .C(index_i[5]), .Z(n24376)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24245_3_lut.init = 16'hcaca;
    PFUMX i21446 (.BLUT(n23926), .ALUT(n23927), .C0(index_i[4]), .Z(n23928));
    LUT4 i24249_3_lut (.A(n542_adj_3199), .B(n573_adj_3050), .C(index_i[5]), 
         .Z(n24370)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24249_3_lut.init = 16'hcaca;
    LUT4 i24251_3_lut (.A(n27073), .B(n444_adj_3200), .C(index_i[5]), 
         .Z(n24368)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24251_3_lut.init = 16'hcaca;
    PFUMX i22443 (.BLUT(n31_adj_3201), .ALUT(n62_adj_3202), .C0(index_q[5]), 
          .Z(n24944));
    LUT4 mux_206_Mux_2_i142_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n142_adj_3203)) /* synthesis lut_function=(!(A (B)+!A (B (C)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_2_i142_3_lut_4_lut_4_lut_4_lut.init = 16'h3626;
    LUT4 n557_bdd_2_lut_3_lut_4_lut (.A(n29379), .B(index_i[2]), .C(index_i[6]), 
         .D(index_i[3]), .Z(n28344)) /* synthesis lut_function=(A (B (C)+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n557_bdd_2_lut_3_lut_4_lut.init = 16'hf087;
    LUT4 mux_207_Mux_0_i795_3_lut_3_lut_rep_830 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n32031)) /* synthesis lut_function=(A (B+(C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_0_i795_3_lut_3_lut_rep_830.init = 16'hadad;
    LUT4 mux_207_Mux_0_i796_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n796_adj_3204)) /* synthesis lut_function=(A (B (C+(D))+!B (C (D)))+!A !(B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_0_i796_3_lut_4_lut_4_lut.init = 16'hadc0;
    PFUMX i21449 (.BLUT(n23929), .ALUT(n23930), .C0(index_i[4]), .Z(n23931));
    LUT4 n954_bdd_3_lut_26304 (.A(n21712), .B(n29099), .C(index_q[5]), 
         .Z(n28170)) /* synthesis lut_function=(A (B (C))+!A (B+!(C))) */ ;
    defparam n954_bdd_3_lut_26304.init = 16'hc5c5;
    LUT4 mux_206_Mux_7_i890_3_lut_3_lut_4_lut (.A(index_i[0]), .B(n29400), 
         .C(index_i[3]), .D(n29180), .Z(n890_adj_3205)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A !(C+(D))) */ ;
    defparam mux_206_Mux_7_i890_3_lut_3_lut_4_lut.init = 16'h808f;
    LUT4 i12837_3_lut_4_lut (.A(index_i[0]), .B(n29400), .C(n29374), .D(index_i[5]), 
         .Z(n318)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (C (D))) */ ;
    defparam i12837_3_lut_4_lut.init = 16'hf800;
    LUT4 n924_bdd_3_lut_26404 (.A(n924_adj_3206), .B(n28172), .C(index_q[5]), 
         .Z(n28173)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n924_bdd_3_lut_26404.init = 16'hcaca;
    LUT4 i20739_3_lut_3_lut_4_lut (.A(index_i[0]), .B(n29400), .C(index_i[3]), 
         .D(n29179), .Z(n23221)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A !(C+(D))) */ ;
    defparam i20739_3_lut_3_lut_4_lut.init = 16'h808f;
    LUT4 mux_206_Mux_5_i987_4_lut_4_lut_4_lut (.A(index_i[0]), .B(n29400), 
         .C(index_i[4]), .D(index_i[3]), .Z(n21704)) /* synthesis lut_function=(A (B (C+!(D))+!B (D))+!A (B (C (D)+!C !(D))+!B (D))) */ ;
    defparam mux_206_Mux_5_i987_4_lut_4_lut_4_lut.init = 16'hf38c;
    LUT4 i20658_3_lut_3_lut_4_lut (.A(index_i[0]), .B(n29400), .C(n29179), 
         .D(index_i[3]), .Z(n23140)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(C+(D)))) */ ;
    defparam i20658_3_lut_3_lut_4_lut.init = 16'h77f0;
    LUT4 mux_207_Mux_6_i700_3_lut_4_lut (.A(n29467), .B(index_q[3]), .C(index_q[4]), 
         .D(n684_adj_3207), .Z(n700_adj_3208)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_6_i700_3_lut_4_lut.init = 16'h9f90;
    LUT4 i23786_3_lut (.A(n23092), .B(n23093), .C(index_q[4]), .Z(n23094)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23786_3_lut.init = 16'hcaca;
    LUT4 i23631_3_lut (.A(n142), .B(n15165), .C(index_q[4]), .Z(n158_adj_3209)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23631_3_lut.init = 16'hcaca;
    LUT4 n62_bdd_3_lut_4_lut_adj_180 (.A(n29418), .B(index_i[3]), .C(index_i[4]), 
         .D(n30_adj_3210), .Z(n28537)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n62_bdd_3_lut_4_lut_adj_180.init = 16'hf808;
    LUT4 i24272_3_lut (.A(n27539), .B(n23912), .C(index_i[5]), .Z(n23913)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24272_3_lut.init = 16'hcaca;
    LUT4 i19392_4_lut (.A(n29365), .B(n16898), .C(index_i[6]), .D(index_i[5]), 
         .Z(n21737)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D))))) */ ;
    defparam i19392_4_lut.init = 16'h3a35;
    LUT4 i24420_3_lut (.A(n21737), .B(n22131), .C(index_i[7]), .Z(n24719)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24420_3_lut.init = 16'hcaca;
    LUT4 i24297_3_lut (.A(n13387), .B(n892_adj_3211), .C(index_q[6]), 
         .Z(n25228)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24297_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_4_lut_adj_181 (.A(n29049), .B(index_q[5]), .C(index_q[8]), 
         .D(n29250), .Z(n22031)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i1_3_lut_4_lut_adj_181.init = 16'hfff8;
    LUT4 n236_bdd_3_lut_26520_4_lut_4_lut (.A(n29418), .B(index_i[3]), .C(index_i[4]), 
         .D(n29180), .Z(n28364)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C))+!A !(B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n236_bdd_3_lut_26520_4_lut_4_lut.init = 16'h838f;
    LUT4 i22281_3_lut_3_lut_4_lut_4_lut (.A(n29418), .B(index_i[3]), .C(index_i[4]), 
         .D(n29176), .Z(n24782)) /* synthesis lut_function=(!(A (B (C)+!B ((D)+!C))+!A (B+((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i22281_3_lut_3_lut_4_lut_4_lut.init = 16'h0838;
    LUT4 i11232_3_lut_4_lut_4_lut (.A(n29418), .B(index_i[3]), .C(index_i[5]), 
         .D(n29177), .Z(n13529)) /* synthesis lut_function=(A (B+(C (D)))+!A (B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11232_3_lut_4_lut_4_lut.init = 16'hf8c8;
    LUT4 mux_206_Mux_9_i124_3_lut_3_lut_4_lut (.A(n29375), .B(index_i[1]), 
         .C(index_i[3]), .D(n29180), .Z(n124_adj_3044)) /* synthesis lut_function=(!(A (C (D))+!A (B (C (D))+!B ((D)+!C)))) */ ;
    defparam mux_206_Mux_9_i124_3_lut_3_lut_4_lut.init = 16'h0efe;
    LUT4 mux_206_Mux_8_i475_3_lut_3_lut_4_lut (.A(n29375), .B(index_i[1]), 
         .C(index_i[3]), .D(n29180), .Z(n475_adj_3212)) /* synthesis lut_function=(A (C+!(D))+!A (B (C+!(D))+!B !(C+(D)))) */ ;
    defparam mux_206_Mux_8_i475_3_lut_3_lut_4_lut.init = 16'he0ef;
    LUT4 mux_206_Mux_0_i572_3_lut_4_lut (.A(n29375), .B(index_i[1]), .C(index_i[3]), 
         .D(n32021), .Z(n572_adj_3213)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam mux_206_Mux_0_i572_3_lut_4_lut.init = 16'hefe0;
    LUT4 i11231_4_lut_4_lut (.A(n29375), .B(index_i[1]), .C(index_i[3]), 
         .D(n22576), .Z(n13528)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A (B (C)+!B ((D)+!C)))) */ ;
    defparam i11231_4_lut_4_lut.init = 16'h0e3e;
    LUT4 n236_bdd_3_lut_26449_3_lut_4_lut (.A(n29375), .B(index_i[1]), .C(index_i[4]), 
         .D(index_i[3]), .Z(n28363)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B ((D)+!C))) */ ;
    defparam n236_bdd_3_lut_26449_3_lut_4_lut.init = 16'hf10f;
    LUT4 i21402_4_lut_4_lut_3_lut_4_lut (.A(n29375), .B(index_i[1]), .C(index_i[4]), 
         .D(index_i[3]), .Z(n23884)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B !((D)+!C)))) */ ;
    defparam i21402_4_lut_4_lut_3_lut_4_lut.init = 16'h11ef;
    LUT4 i12817_2_lut_rep_393_3_lut_4_lut (.A(n29375), .B(index_i[1]), .C(index_i[4]), 
         .D(index_i[3]), .Z(n29053)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i12817_2_lut_rep_393_3_lut_4_lut.init = 16'hfef0;
    PFUMX i21452 (.BLUT(n23932), .ALUT(n23933), .C0(index_i[4]), .Z(n23934));
    LUT4 i21480_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n23962)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A !(B (D)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i21480_3_lut_3_lut_4_lut.init = 16'ha955;
    LUT4 i22579_3_lut (.A(n28664), .B(n25071), .C(index_q[6]), .Z(n25080)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22579_3_lut.init = 16'hcaca;
    LUT4 mux_206_Mux_6_i890_3_lut_3_lut_4_lut (.A(n29376), .B(index_i[2]), 
         .C(n29382), .D(index_i[3]), .Z(n890_adj_3034)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_6_i890_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 i12869_4_lut (.A(n29101), .B(index_i[7]), .C(n16898), .D(index_i[6]), 
         .Z(n1021)) /* synthesis lut_function=(A (B+(C (D)))+!A (B+(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12869_4_lut.init = 16'hfcdd;
    LUT4 mux_206_Mux_3_i93_3_lut_4_lut (.A(n29376), .B(index_i[2]), .C(index_i[3]), 
         .D(n29377), .Z(n93)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_3_i93_3_lut_4_lut.init = 16'hefe0;
    LUT4 mux_206_Mux_8_i124_3_lut_3_lut_4_lut (.A(n29376), .B(index_i[2]), 
         .C(n29380), .D(index_i[3]), .Z(n124_adj_3214)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_8_i124_3_lut_3_lut_4_lut.init = 16'h11f0;
    PFUMX i21455 (.BLUT(n23935), .ALUT(n23936), .C0(index_i[4]), .Z(n23937));
    LUT4 mux_206_Mux_0_i1002_3_lut_3_lut_4_lut (.A(n29376), .B(index_i[2]), 
         .C(n1001), .D(index_i[3]), .Z(n1002_adj_3215)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i1002_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 mux_207_Mux_9_i62_3_lut_3_lut_4_lut_then_4_lut (.A(index_q[2]), .B(index_q[1]), 
         .C(index_q[0]), .D(index_q[4]), .Z(n29549)) /* synthesis lut_function=(!(A (B+(C+!(D)))+!A !(B (D)+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_9_i62_3_lut_3_lut_4_lut_then_4_lut.init = 16'h5701;
    LUT4 mux_206_Mux_11_i638_4_lut_4_lut (.A(n29053), .B(index_i[5]), .C(index_i[6]), 
         .D(n29087), .Z(n638_adj_3216)) /* synthesis lut_function=(A (B (C (D))+!B !(C))+!A (B ((D)+!C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_11_i638_4_lut_4_lut.init = 16'hc707;
    LUT4 i20946_3_lut (.A(n29336), .B(n29393), .C(index_q[3]), .Z(n23428)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20946_3_lut.init = 16'hcaca;
    LUT4 i23737_3_lut (.A(n23428), .B(n23429), .C(index_q[4]), .Z(n23430)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23737_3_lut.init = 16'hcaca;
    LUT4 i20724_3_lut_4_lut (.A(n29379), .B(index_i[2]), .C(index_i[3]), 
         .D(n29409), .Z(n23206)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20724_3_lut_4_lut.init = 16'hdfd0;
    LUT4 i22558_3_lut (.A(n94_adj_3052), .B(n476), .C(index_q[5]), .Z(n25059)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22558_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_7_i572_3_lut_rep_379_3_lut_3_lut_4_lut (.A(index_q[0]), 
         .B(index_q[1]), .C(index_q[3]), .D(index_q[2]), .Z(n29039)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)+!C !(D)))) */ ;
    defparam mux_207_Mux_7_i572_3_lut_rep_379_3_lut_3_lut_4_lut.init = 16'hfe01;
    LUT4 i22598_3_lut (.A(n32019), .B(n29384), .C(index_i[3]), .Z(n25099)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22598_3_lut.init = 16'hcaca;
    LUT4 i22597_3_lut (.A(n1001), .B(n29407), .C(index_i[3]), .Z(n25098)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22597_3_lut.init = 16'hcaca;
    PFUMX i20803 (.BLUT(n445), .ALUT(n508_adj_3037), .C0(index_i[6]), 
          .Z(n23285));
    LUT4 n698_bdd_3_lut_25716_4_lut (.A(n29379), .B(index_i[2]), .C(index_i[3]), 
         .D(n29385), .Z(n27465)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n698_bdd_3_lut_25716_4_lut.init = 16'hdfd0;
    LUT4 i21451_3_lut_4_lut (.A(n29379), .B(index_i[2]), .C(index_i[3]), 
         .D(n29446), .Z(n23933)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21451_3_lut_4_lut.init = 16'hdfd0;
    LUT4 mux_207_Mux_0_i915_3_lut_rep_800 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29460)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C)+!B !(C))) */ ;
    defparam mux_207_Mux_0_i915_3_lut_rep_800.init = 16'he3e3;
    LUT4 i22595_3_lut (.A(n29384), .B(n645), .C(index_i[3]), .Z(n25096)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22595_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_0_i333_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n333)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B (D))) */ ;
    defparam mux_207_Mux_0_i333_3_lut_3_lut_4_lut.init = 16'hf10e;
    LUT4 i24346_3_lut (.A(n13530), .B(n892_adj_3217), .C(index_i[6]), 
         .Z(n24835)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24346_3_lut.init = 16'hcaca;
    LUT4 n922_bdd_3_lut_26608 (.A(n32019), .B(index_i[3]), .C(n32018), 
         .Z(n27185)) /* synthesis lut_function=(A (B+(C))+!A !(B+!(C))) */ ;
    defparam n922_bdd_3_lut_26608.init = 16'hb8b8;
    LUT4 i20943_3_lut (.A(n29373), .B(n588), .C(index_q[3]), .Z(n23425)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20943_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_9_i62_3_lut_3_lut_4_lut_else_4_lut (.A(index_q[2]), .B(index_q[1]), 
         .C(index_q[0]), .D(index_q[4]), .Z(n29548)) /* synthesis lut_function=(A+(B (C+!(D))+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_9_i62_3_lut_3_lut_4_lut_else_4_lut.init = 16'heaff;
    LUT4 i23739_3_lut (.A(n23425), .B(n23426), .C(index_q[4]), .Z(n23427)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23739_3_lut.init = 16'hcaca;
    LUT4 i12824_3_lut_4_lut (.A(n29032), .B(index_i[7]), .C(index_i[8]), 
         .D(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_1768[14])) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (D))) */ ;
    defparam i12824_3_lut_4_lut.init = 16'hffe0;
    LUT4 i22512_3_lut (.A(n236), .B(n251), .C(index_i[4]), .Z(n25013)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22512_3_lut.init = 16'hcaca;
    LUT4 i12670_4_lut (.A(n29102), .B(index_q[7]), .C(n892), .D(index_q[6]), 
         .Z(n1021_adj_3218)) /* synthesis lut_function=(A (B+(C (D)))+!A (B+(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i12670_4_lut.init = 16'hfcdd;
    LUT4 i22841_3_lut (.A(n25339), .B(n25340), .C(index_q[7]), .Z(n25342)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22841_3_lut.init = 16'hcaca;
    LUT4 i22840_3_lut (.A(n25337), .B(n25338), .C(index_q[7]), .Z(n25341)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22840_3_lut.init = 16'hcaca;
    LUT4 i22808_3_lut (.A(n25304), .B(n25305), .C(index_i[7]), .Z(n25309)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22808_3_lut.init = 16'hcaca;
    LUT4 i22800_3_lut (.A(n25288), .B(n26746), .C(index_i[6]), .Z(n25301)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22800_3_lut.init = 16'hcaca;
    LUT4 i22799_3_lut (.A(n26730), .B(n25287), .C(index_i[6]), .Z(n25300)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22799_3_lut.init = 16'hcaca;
    LUT4 i22797_3_lut (.A(n26724), .B(n25283), .C(index_i[6]), .Z(n25298)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22797_3_lut.init = 16'hcaca;
    LUT4 i22772_3_lut (.A(n25270), .B(n25271), .C(index_i[7]), .Z(n25273)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22772_3_lut.init = 16'hcaca;
    LUT4 mux_206_Mux_3_i30_3_lut_3_lut_4_lut_3_lut_4_lut (.A(index_i[1]), 
         .B(index_i[0]), .C(index_i[3]), .D(index_i[2]), .Z(n30_adj_3136)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_3_i30_3_lut_3_lut_4_lut_3_lut_4_lut.init = 16'hfe11;
    LUT4 i22771_3_lut (.A(n25268), .B(n25269), .C(index_i[7]), .Z(n25272)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22771_3_lut.init = 16'hcaca;
    LUT4 i22730_3_lut (.A(n25224), .B(n25225), .C(index_q[7]), .Z(n25231)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22730_3_lut.init = 16'hcaca;
    LUT4 i22729_3_lut (.A(n25222), .B(n25223), .C(index_q[7]), .Z(n25230)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22729_3_lut.init = 16'hcaca;
    PFUMX i22376 (.BLUT(n158_adj_3219), .ALUT(n189_adj_3220), .C0(index_q[5]), 
          .Z(n24877));
    PFUMX i22344 (.BLUT(n94_adj_3221), .ALUT(n125_adj_3222), .C0(index_q[5]), 
          .Z(n24845));
    LUT4 i22734_3_lut (.A(n25232), .B(n25233), .C(index_q[8]), .Z(n25235)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22734_3_lut.init = 16'hcaca;
    LUT4 i22717_3_lut (.A(n25213), .B(n25214), .C(index_q[7]), .Z(n25218)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22717_3_lut.init = 16'hcaca;
    PFUMX i22345 (.BLUT(n20006), .ALUT(n16248), .C0(index_q[5]), .Z(n24846));
    LUT4 index_q_8__bdd_3_lut_26186_then_4_lut (.A(index_q[4]), .B(index_q[6]), 
         .C(index_q[5]), .D(n29095), .Z(n29552)) /* synthesis lut_function=(!(A (B (C+(D)))+!A (B (C)))) */ ;
    defparam index_q_8__bdd_3_lut_26186_then_4_lut.init = 16'h373f;
    LUT4 n27757_bdd_3_lut_3_lut (.A(n1021_adj_3218), .B(index_q[8]), .C(n27757), 
         .Z(n27758)) /* synthesis lut_function=(A (B+(C))+!A !(B+!(C))) */ ;
    defparam n27757_bdd_3_lut_3_lut.init = 16'hb8b8;
    LUT4 index_q_8__bdd_3_lut_26186_else_4_lut (.A(n29161), .B(index_q[4]), 
         .C(index_q[6]), .D(index_q[5]), .Z(n29551)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;
    defparam index_q_8__bdd_3_lut_26186_else_4_lut.init = 16'hf080;
    LUT4 i22534_3_lut (.A(n25032), .B(n25033), .C(index_i[7]), .Z(n25035)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22534_3_lut.init = 16'hcaca;
    LUT4 i22533_3_lut (.A(n25030), .B(n25031), .C(index_i[7]), .Z(n25034)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22533_3_lut.init = 16'hcaca;
    LUT4 i22503_3_lut (.A(n25001), .B(n25002), .C(index_q[7]), .Z(n25004)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22503_3_lut.init = 16'hcaca;
    LUT4 i22502_3_lut (.A(n24999), .B(n25000), .C(index_q[7]), .Z(n25003)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22502_3_lut.init = 16'hcaca;
    LUT4 i22401_3_lut (.A(n24897), .B(n24898), .C(index_q[7]), .Z(n24902)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22401_3_lut.init = 16'hcaca;
    LUT4 i21970_3_lut (.A(n24464), .B(n24465), .C(index_q[7]), .Z(n24471)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21970_3_lut.init = 16'hcaca;
    PFUMX i22374 (.BLUT(n31_adj_3223), .ALUT(n62_adj_3224), .C0(index_q[5]), 
          .Z(n24875));
    LUT4 i21969_3_lut (.A(n24462), .B(n24463), .C(index_q[7]), .Z(n24470)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21969_3_lut.init = 16'hcaca;
    LUT4 n26753_bdd_3_lut (.A(n26753), .B(n157_adj_3225), .C(index_i[4]), 
         .Z(n26754)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n26753_bdd_3_lut.init = 16'hcaca;
    LUT4 i22337_3_lut (.A(n24831), .B(n24832), .C(index_i[7]), .Z(n24838)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22337_3_lut.init = 16'hcaca;
    LUT4 i14123_3_lut (.A(index_i[2]), .B(index_i[1]), .C(index_i[0]), 
         .Z(n1001)) /* synthesis lut_function=(A (B)+!A (B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i14123_3_lut.init = 16'hdcdc;
    LUT4 i22336_3_lut (.A(n24829), .B(n24830), .C(index_i[7]), .Z(n24837)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22336_3_lut.init = 16'hcaca;
    LUT4 i22341_3_lut (.A(n24839), .B(n24840), .C(index_i[8]), .Z(n24842)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22341_3_lut.init = 16'hcaca;
    LUT4 i12908_2_lut_rep_513_3_lut (.A(index_i[2]), .B(index_i[3]), .C(index_i[1]), 
         .Z(n29173)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12908_2_lut_rep_513_3_lut.init = 16'hfefe;
    LUT4 i1_3_lut_4_lut_adj_182 (.A(n29053), .B(index_i[5]), .C(index_i[8]), 
         .D(n29251), .Z(n22033)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_3_lut_4_lut_adj_182.init = 16'hfff8;
    LUT4 i21888_3_lut (.A(n24384), .B(n24385), .C(index_i[7]), .Z(n24389)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21888_3_lut.init = 16'hcaca;
    LUT4 mux_206_Mux_14_i511_4_lut_4_lut (.A(n29032), .B(index_i[7]), .C(index_i[8]), 
         .D(n254_adj_3105), .Z(n511_adj_3226)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (B (C+!(D))+!B !(C)))) */ ;
    defparam mux_206_Mux_14_i511_4_lut_4_lut.init = 16'h1c10;
    LUT4 mux_206_Mux_11_i766_3_lut (.A(n638_adj_3216), .B(n16882), .C(index_i[7]), 
         .Z(n766)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_11_i766_3_lut.init = 16'h3a3a;
    LUT4 i22231_3_lut (.A(n27195), .B(n24726), .C(index_i[7]), .Z(n24732)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22231_3_lut.init = 16'hcaca;
    LUT4 i22230_3_lut (.A(n24723), .B(n24724), .C(index_i[7]), .Z(n24731)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22230_3_lut.init = 16'hcaca;
    PFUMX i21386 (.BLUT(n23866), .ALUT(n23867), .C0(index_i[5]), .Z(n23868));
    LUT4 n62_bdd_4_lut (.A(n29372), .B(n29173), .C(index_i[6]), .D(index_i[4]), 
         .Z(n31711)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C+(D)))+!A (B ((D)+!C)+!B !(C)))) */ ;
    defparam n62_bdd_4_lut.init = 16'h3af0;
    LUT4 n25172_bdd_4_lut (.A(n252_adj_3227), .B(n29143), .C(index_i[4]), 
         .D(index_i[5]), .Z(n31708)) /* synthesis lut_function=(A (B (D)+!B ((D)+!C))+!A !(B+(C+(D)))) */ ;
    defparam n25172_bdd_4_lut.init = 16'haa03;
    LUT4 n62_bdd_3_lut (.A(n62_adj_3228), .B(n125_adj_3049), .C(index_i[6]), 
         .Z(n31710)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n62_bdd_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_11_i766_3_lut (.A(n638_adj_3163), .B(n16930), .C(index_q[7]), 
         .Z(n766_adj_3229)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_11_i766_3_lut.init = 16'h3a3a;
    LUT4 i24426_3_lut (.A(n25230), .B(n25231), .C(index_q[8]), .Z(n25234)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24426_3_lut.init = 16'hcaca;
    PFUMX i21968 (.BLUT(n956_adj_3230), .ALUT(n22170), .C0(index_q[6]), 
          .Z(n24469));
    LUT4 i22505_3_lut (.A(n15_adj_3231), .B(n30_adj_3232), .C(index_i[4]), 
         .Z(n25006)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22505_3_lut.init = 16'hcaca;
    LUT4 i20935_3_lut (.A(n29395), .B(n32036), .C(index_q[3]), .Z(n23417)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20935_3_lut.init = 16'hcaca;
    LUT4 i22586_3_lut (.A(n25084), .B(n25085), .C(index_q[8]), .Z(n25087)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22586_3_lut.init = 16'hcaca;
    LUT4 i22585_3_lut (.A(n25082), .B(n25083), .C(index_q[8]), .Z(n25086)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22585_3_lut.init = 16'hcaca;
    LUT4 n62_bdd_3_lut_adj_183 (.A(n62_adj_3146), .B(n125_adj_3016), .C(index_q[6]), 
         .Z(n31747)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n62_bdd_3_lut_adj_183.init = 16'hcaca;
    LUT4 i22370_3_lut (.A(n24866), .B(n28174), .C(index_q[7]), .Z(n24871)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22370_3_lut.init = 16'hcaca;
    LUT4 i22369_3_lut (.A(n24864), .B(n24865), .C(index_q[7]), .Z(n24870)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22369_3_lut.init = 16'hcaca;
    LUT4 i24475_3_lut (.A(n24870), .B(n24871), .C(index_q[8]), .Z(n24873)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24475_3_lut.init = 16'hcaca;
    LUT4 n25277_bdd_4_lut (.A(n252_adj_3233), .B(n29134), .C(index_q[4]), 
         .D(index_q[5]), .Z(n31745)) /* synthesis lut_function=(A (B (D)+!B ((D)+!C))+!A !(B+(C+(D)))) */ ;
    defparam n25277_bdd_4_lut.init = 16'haa03;
    LUT4 n62_bdd_4_lut_adj_184 (.A(n29361), .B(n29161), .C(index_q[6]), 
         .D(index_q[4]), .Z(n31748)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C+(D)))+!A (B ((D)+!C)+!B !(C)))) */ ;
    defparam n62_bdd_4_lut_adj_184.init = 16'h3af0;
    LUT4 i24448_3_lut (.A(n24837), .B(n24838), .C(index_i[8]), .Z(n24841)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24448_3_lut.init = 16'hcaca;
    L6MUX21 i22347 (.D0(n23967), .D1(n23970), .SD(index_q[5]), .Z(n24848));
    LUT4 i21952_3_lut (.A(n24450), .B(n28111), .C(index_i[8]), .Z(n24453)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21952_3_lut.init = 16'hcaca;
    LUT4 i21951_3_lut (.A(n24448), .B(n24449), .C(index_i[8]), .Z(n24452)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21951_3_lut.init = 16'hcaca;
    PFUMX i21389 (.BLUT(n23869), .ALUT(n23870), .C0(index_i[5]), .Z(n23871));
    LUT4 i12835_4_lut (.A(n16668), .B(index_i[8]), .C(n16882), .D(index_i[7]), 
         .Z(n1022)) /* synthesis lut_function=(A (B+(C (D)))+!A (B+(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12835_4_lut.init = 16'hfcdd;
    LUT4 i12570_4_lut (.A(n16844), .B(index_q[8]), .C(n16930), .D(index_q[7]), 
         .Z(n1022_adj_3234)) /* synthesis lut_function=(A (B+(C (D)))+!A (B+(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i12570_4_lut.init = 16'hfcdd;
    LUT4 i20766_3_lut (.A(n28148), .B(n23286), .C(index_i[8]), .Z(n23248)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20766_3_lut.init = 16'hcaca;
    LUT4 i21513_3_lut_4_lut (.A(index_i[0]), .B(n29400), .C(index_i[3]), 
         .D(n29429), .Z(n23995)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A ((D)+!C)) */ ;
    defparam i21513_3_lut_4_lut.init = 16'hfd0d;
    LUT4 i21857_3_lut (.A(n24353), .B(n28077), .C(index_i[7]), .Z(n24358)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21857_3_lut.init = 16'hcaca;
    LUT4 i21856_3_lut (.A(n24351), .B(n24352), .C(index_i[7]), .Z(n24357)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21856_3_lut.init = 16'hcaca;
    LUT4 i24483_3_lut (.A(n24357), .B(n24358), .C(index_i[8]), .Z(n24360)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24483_3_lut.init = 16'hcaca;
    LUT4 index_i_8__bdd_3_lut_then_4_lut (.A(index_i[4]), .B(index_i[6]), 
         .C(index_i[5]), .D(n29086), .Z(n29558)) /* synthesis lut_function=(!(A (B (C+(D)))+!A (B (C)))) */ ;
    defparam index_i_8__bdd_3_lut_then_4_lut.init = 16'h373f;
    LUT4 mux_206_Mux_5_i731_3_lut (.A(n29424), .B(n32020), .C(index_i[3]), 
         .Z(n731_adj_3235)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_5_i731_3_lut.init = 16'hcaca;
    LUT4 n922_bdd_3_lut_25476 (.A(n32019), .B(n29385), .C(index_i[3]), 
         .Z(n27184)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;
    defparam n922_bdd_3_lut_25476.init = 16'h3a3a;
    LUT4 i20727_3_lut (.A(n28084), .B(n23268), .C(index_q[8]), .Z(n23209)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20727_3_lut.init = 16'hcaca;
    LUT4 i11250_3_lut_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n13549)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A !(B (C+(D))+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11250_3_lut_3_lut_4_lut_4_lut.init = 16'h44db;
    LUT4 i22472_3_lut (.A(n24970), .B(n24971), .C(index_q[8]), .Z(n24973)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22472_3_lut.init = 16'hcaca;
    LUT4 i22471_3_lut (.A(n24968), .B(n24969), .C(index_q[8]), .Z(n24972)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22471_3_lut.init = 16'hcaca;
    LUT4 i22036_3_lut (.A(n24534), .B(n24535), .C(index_q[8]), .Z(n24537)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22036_3_lut.init = 16'hcaca;
    LUT4 i22035_3_lut (.A(n24532), .B(n24533), .C(index_q[8]), .Z(n24536)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22035_3_lut.init = 16'hcaca;
    LUT4 i22371_3_lut (.A(n24868), .B(n24869), .C(index_q[8]), .Z(n24872)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22371_3_lut.init = 16'hcaca;
    LUT4 i22005_3_lut (.A(n24503), .B(n24504), .C(index_i[8]), .Z(n24506)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22005_3_lut.init = 16'hcaca;
    LUT4 i22004_3_lut (.A(n24501), .B(n24502), .C(index_i[8]), .Z(n24505)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22004_3_lut.init = 16'hcaca;
    LUT4 i21921_3_lut (.A(n24419), .B(n24420), .C(index_i[8]), .Z(n24422)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21921_3_lut.init = 16'hcaca;
    LUT4 i21920_3_lut (.A(n24417), .B(n24418), .C(index_i[8]), .Z(n24421)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21920_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_6_i325_3_lut_4_lut_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n325)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_6_i325_3_lut_4_lut_3_lut.init = 16'h6d6d;
    PFUMX i27135 (.BLUT(n29575), .ALUT(n29576), .C0(index_i[1]), .Z(n29577));
    LUT4 i24479_3_lut (.A(n574_adj_3150), .B(n637_adj_3236), .C(index_i[6]), 
         .Z(n23287)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24479_3_lut.init = 16'hcaca;
    LUT4 i20731_3_lut_4_lut (.A(index_i[0]), .B(n29418), .C(index_i[3]), 
         .D(n29433), .Z(n23213)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20731_3_lut_4_lut.init = 16'hfb0b;
    LUT4 i21858_3_lut (.A(n24355), .B(n24356), .C(index_i[8]), .Z(n24359)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21858_3_lut.init = 16'hcaca;
    L6MUX21 i22348 (.D0(n23973), .D1(n23073), .SD(index_q[5]), .Z(n24849));
    LUT4 i24485_3_lut (.A(n574_adj_3056), .B(n637), .C(index_q[6]), .Z(n23269)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24485_3_lut.init = 16'hcaca;
    LUT4 index_i_8__bdd_3_lut_else_4_lut (.A(n29173), .B(index_i[4]), .C(index_i[6]), 
         .D(index_i[5]), .Z(n29557)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;
    defparam index_i_8__bdd_3_lut_else_4_lut.init = 16'hf080;
    PFUMX i22349 (.BLUT(n413_adj_3237), .ALUT(n444_adj_3066), .C0(index_q[5]), 
          .Z(n24850));
    LUT4 mux_207_Mux_8_i285_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n285_adj_3238)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C (D)+!C !(D))+!B (C)))) */ ;
    defparam mux_207_Mux_8_i285_3_lut_3_lut_4_lut.init = 16'h0fc1;
    PFUMX i21482 (.BLUT(n23962), .ALUT(n23963), .C0(index_q[4]), .Z(n23964));
    LUT4 mux_207_Mux_0_i557_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n557_adj_3239)) /* synthesis lut_function=(A ((D)+!C)+!A !((D)+!B)) */ ;
    defparam mux_207_Mux_0_i557_3_lut_4_lut.init = 16'haa4e;
    LUT4 mux_207_Mux_0_i699_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n699_adj_3240)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (D))+!A (B (C+!(D))+!B !(C+!(D))))) */ ;
    defparam mux_207_Mux_0_i699_3_lut_3_lut_4_lut.init = 16'h1c33;
    LUT4 i20937_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n23419)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C (D)))+!A (B (C+(D))+!B !(C)))) */ ;
    defparam i20937_4_lut_4_lut_4_lut.init = 16'h301c;
    LUT4 i21475_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n23957)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B (C (D)+!C !(D))))) */ ;
    defparam i21475_3_lut_3_lut_4_lut.init = 16'h0f1c;
    LUT4 mux_207_Mux_0_i15_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n15_adj_3053)) /* synthesis lut_function=(A (B (C)+!B ((D)+!C))+!A (B (C)+!B !(C))) */ ;
    defparam mux_207_Mux_0_i15_3_lut_4_lut_4_lut.init = 16'he3c3;
    LUT4 i1_2_lut_rep_805 (.A(index_q[1]), .B(index_q[0]), .Z(n29465)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i1_2_lut_rep_805.init = 16'h8888;
    LUT4 mux_207_Mux_6_i781_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), 
         .B(index_q[0]), .C(index_q[3]), .D(index_q[2]), .Z(n781)) /* synthesis lut_function=(A (B (D)+!B (C (D)+!C !(D)))+!A !(D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_6_i781_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'ha857;
    LUT4 mux_206_Mux_10_i413_3_lut_4_lut (.A(n29176), .B(index_i[3]), .C(index_i[4]), 
         .D(n29146), .Z(n413_adj_3241)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_10_i413_3_lut_4_lut.init = 16'hf101;
    LUT4 mux_207_Mux_1_i348_3_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[0]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n348_adj_3242)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_1_i348_3_lut_4_lut_4_lut.init = 16'h5f80;
    L6MUX21 i25232 (.D0(n26901), .D1(n26899), .SD(index_i[5]), .Z(n26902));
    LUT4 i20917_3_lut_4_lut_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[0]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n23399)) /* synthesis lut_function=(!(A (B (C)+!B (C+(D)))+!A !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i20917_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'h585f;
    LUT4 i12706_2_lut_2_lut_3_lut (.A(index_q[1]), .B(index_q[0]), .C(index_q[3]), 
         .Z(n15114)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i12706_2_lut_2_lut_3_lut.init = 16'h0808;
    LUT4 n27398_bdd_3_lut_26538_4_lut (.A(n29176), .B(index_i[3]), .C(index_i[5]), 
         .D(n27400), .Z(n28108)) /* synthesis lut_function=(!(A (C+!(D))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n27398_bdd_3_lut_26538_4_lut.init = 16'h1f10;
    LUT4 mux_207_Mux_7_i491_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[0]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n491_adj_3243)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C+!(D)))+!A !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_7_i491_3_lut_4_lut_4_lut_4_lut.init = 16'h5780;
    LUT4 i24735_2_lut_rep_472_3_lut_4_lut (.A(index_q[1]), .B(index_q[0]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n29132)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i24735_2_lut_rep_472_3_lut_4_lut.init = 16'h0007;
    LUT4 n28442_bdd_3_lut (.A(n28442), .B(n476_adj_3244), .C(index_i[5]), 
         .Z(n28443)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n28442_bdd_3_lut.init = 16'hcaca;
    PFUMX i21398 (.BLUT(n23878), .ALUT(n23879), .C0(index_i[5]), .Z(n23880));
    PFUMX i21485 (.BLUT(n23965), .ALUT(n23966), .C0(index_q[4]), .Z(n23967));
    PFUMX i21977 (.BLUT(n94_adj_3245), .ALUT(n23202), .C0(index_i[5]), 
          .Z(n24478));
    LUT4 mux_207_Mux_9_i316_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[0]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n316_adj_3246)) /* synthesis lut_function=(!(A (B (C (D))+!B (C (D)+!C !(D)))+!A !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_9_i316_3_lut_4_lut_4_lut_4_lut.init = 16'h5ff8;
    LUT4 n285_bdd_3_lut_4_lut_4_lut_4_lut_adj_185 (.A(index_q[1]), .B(index_q[0]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n27559)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)+!C !(D)))+!A ((D)+!C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam n285_bdd_3_lut_4_lut_4_lut_4_lut_adj_185.init = 16'hf58f;
    L6MUX21 i21978 (.D0(n23205), .D1(n23208), .SD(index_i[5]), .Z(n24479));
    LUT4 i11254_3_lut_4_lut_3_lut (.A(index_q[1]), .B(index_q[0]), .C(index_q[4]), 
         .Z(n13553)) /* synthesis lut_function=(A (B)+!A !(B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i11254_3_lut_4_lut_3_lut.init = 16'h9898;
    LUT4 mux_207_Mux_8_i526_3_lut_3_lut_3_lut_4_lut (.A(index_q[1]), .B(index_q[0]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n526_adj_3247)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_8_i526_3_lut_3_lut_3_lut_4_lut.init = 16'h0f70;
    LUT4 mux_206_Mux_3_i828_3_lut_3_lut_4_lut (.A(n29176), .B(index_i[3]), 
         .C(n157_adj_3248), .D(index_i[4]), .Z(n828_adj_3249)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_3_i828_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 mux_207_Mux_4_i1002_3_lut_3_lut_3_lut_4_lut (.A(index_q[1]), .B(index_q[0]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n1002_adj_3250)) /* synthesis lut_function=(A (B (C (D))+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_4_i1002_3_lut_3_lut_3_lut_4_lut.init = 16'hf007;
    LUT4 n28446_bdd_3_lut (.A(n29541), .B(n28444), .C(index_i[5]), .Z(n28447)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n28446_bdd_3_lut.init = 16'hcaca;
    LUT4 i22300_3_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[0]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n24801)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A !(C (D)+!C !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i22300_3_lut_4_lut_4_lut.init = 16'h8f50;
    PFUMX i25230 (.BLUT(n26900), .ALUT(n645), .C0(index_i[3]), .Z(n26901));
    LUT4 mux_207_Mux_8_i732_3_lut (.A(index_q[3]), .B(n16858), .C(index_q[5]), 
         .Z(n732_adj_3251)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_8_i732_3_lut.init = 16'h3a3a;
    LUT4 i12511_2_lut_rep_420_3_lut_4_lut (.A(index_q[1]), .B(index_q[0]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n29080)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i12511_2_lut_rep_420_3_lut_4_lut.init = 16'hf080;
    LUT4 mux_207_Mux_7_i526_3_lut_3_lut_4_lut_4_lut_3_lut_4_lut (.A(index_q[1]), 
         .B(index_q[0]), .C(index_q[3]), .D(index_q[2]), .Z(n526_adj_3252)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(D))+!A !(D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_7_i526_3_lut_3_lut_4_lut_4_lut_3_lut_4_lut.init = 16'h887f;
    LUT4 n172_bdd_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[0]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n27390)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam n172_bdd_3_lut_4_lut_4_lut_4_lut.init = 16'h0f58;
    LUT4 i12514_2_lut_rep_508_3_lut (.A(index_q[1]), .B(index_q[0]), .C(index_q[2]), 
         .Z(n29168)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i12514_2_lut_rep_508_3_lut.init = 16'hf8f8;
    PFUMX i21488 (.BLUT(n23968), .ALUT(n23969), .C0(index_q[4]), .Z(n23970));
    LUT4 i20607_3_lut (.A(n29389), .B(n32029), .C(index_q[3]), .Z(n23089)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20607_3_lut.init = 16'hcaca;
    PFUMX i22350 (.BLUT(n476_adj_3253), .ALUT(n507_adj_3254), .C0(index_q[5]), 
          .Z(n24851));
    LUT4 index_q_6__bdd_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[0]), 
         .C(index_q[6]), .D(n29361), .Z(n28502)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam index_q_6__bdd_4_lut_4_lut_4_lut.init = 16'h0f7a;
    LUT4 mux_207_Mux_6_i812_3_lut_4_lut_3_lut_4_lut (.A(index_q[1]), .B(index_q[0]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n812_adj_3074)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(D))+!A !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_6_i812_3_lut_4_lut_3_lut_4_lut.init = 16'h7780;
    LUT4 mux_207_Mux_3_i1002_3_lut_3_lut_4_lut (.A(index_q[1]), .B(index_q[0]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n21714)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (D))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_3_i1002_3_lut_3_lut_4_lut.init = 16'hf708;
    LUT4 mux_207_Mux_8_i635_3_lut_4_lut_3_lut_4_lut (.A(index_q[1]), .B(index_q[0]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n635_adj_3255)) /* synthesis lut_function=(!(A (B (C (D))+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_8_i635_3_lut_4_lut_3_lut_4_lut.init = 16'h0ff8;
    PFUMX i21491 (.BLUT(n23971), .ALUT(n23972), .C0(index_q[4]), .Z(n23973));
    LUT4 i21810_2_lut (.A(index_q[3]), .B(index_q[5]), .Z(n24311)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i21810_2_lut.init = 16'h8888;
    LUT4 n77_bdd_3_lut_26950_3_lut_4_lut_4_lut_3_lut_4_lut (.A(index_q[1]), 
         .B(index_q[0]), .C(index_q[3]), .D(index_q[2]), .Z(n27573)) /* synthesis lut_function=(A (B (C)+!B !(D))+!A !(D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam n77_bdd_3_lut_26950_3_lut_4_lut_4_lut_3_lut_4_lut.init = 16'h80f7;
    LUT4 i20648_then_4_lut (.A(index_q[2]), .B(index_q[1]), .C(index_q[4]), 
         .D(index_q[3]), .Z(n29479)) /* synthesis lut_function=(A (B (C+(D))+!B !(C))+!A !(B (C+(D))+!B !(C+!(D)))) */ ;
    defparam i20648_then_4_lut.init = 16'h9a97;
    LUT4 n301_bdd_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[0]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n27557)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (D))+!A !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam n301_bdd_3_lut_4_lut_4_lut_4_lut.init = 16'h50f7;
    PFUMX i21401 (.BLUT(n23881), .ALUT(n23882), .C0(index_i[5]), .Z(n23883));
    LUT4 i12775_2_lut_rep_397_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[0]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n29057)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i12775_2_lut_rep_397_4_lut_4_lut_4_lut.init = 16'h0058;
    LUT4 mux_207_Mux_7_i747_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[0]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n747_adj_3256)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))+!A (C (D)+!C !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_7_i747_3_lut_4_lut_4_lut_4_lut.init = 16'hf0a7;
    LUT4 i20922_3_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[0]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n23404)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i20922_3_lut_4_lut_4_lut.init = 16'h5a8a;
    PFUMX i25228 (.BLUT(n26898), .ALUT(n23615), .C0(index_i[4]), .Z(n26899));
    LUT4 i12702_3_lut_3_lut_3_lut_4_lut (.A(index_q[1]), .B(index_q[0]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n15110)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (D))+!A (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i12702_3_lut_3_lut_3_lut_4_lut.init = 16'h00f7;
    LUT4 mux_207_Mux_7_i141_3_lut_4_lut_3_lut (.A(index_q[1]), .B(index_q[0]), 
         .C(index_q[2]), .Z(n141)) /* synthesis lut_function=(A ((C)+!B)+!A (B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_7_i141_3_lut_4_lut_3_lut.init = 16'he7e7;
    LUT4 i1_2_lut_rep_474_3_lut_4_lut (.A(index_q[1]), .B(index_q[0]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n29134)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i1_2_lut_rep_474_3_lut_4_lut.init = 16'h8000;
    LUT4 mux_207_Mux_7_i92_3_lut_rep_807 (.A(index_q[1]), .B(index_q[0]), 
         .C(index_q[2]), .Z(n29467)) /* synthesis lut_function=(A (B+!(C))+!A !((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_7_i92_3_lut_rep_807.init = 16'h8e8e;
    LUT4 mux_207_Mux_8_i124_3_lut_3_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[0]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n124_adj_3257)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (B (C+!(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_8_i124_3_lut_3_lut_4_lut_4_lut.init = 16'h07a1;
    LUT4 mux_207_Mux_0_i581_3_lut_3_lut_rep_810 (.A(index_q[1]), .B(index_q[0]), 
         .C(index_q[2]), .Z(n29470)) /* synthesis lut_function=(A ((C)+!B)+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_0_i581_3_lut_3_lut_rep_810.init = 16'ha7a7;
    LUT4 i23655_3_lut (.A(n23155), .B(n23156), .C(index_q[4]), .Z(n23157)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i23655_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_8_i29_3_lut_rep_811 (.A(index_q[1]), .B(index_q[0]), 
         .C(index_q[2]), .Z(n29471)) /* synthesis lut_function=(!(A (B (C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_8_i29_3_lut_rep_811.init = 16'h7e7e;
    LUT4 mux_207_Mux_7_i7_3_lut_4_lut_3_lut_rep_812 (.A(index_q[1]), .B(index_q[0]), 
         .C(index_q[2]), .Z(n29472)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_7_i7_3_lut_4_lut_3_lut_rep_812.init = 16'h1818;
    LUT4 i20648_else_4_lut (.A(index_q[2]), .B(index_q[1]), .C(index_q[4]), 
         .D(index_q[3]), .Z(n29478)) /* synthesis lut_function=(!(A (B (C)+!B (C+(D)))+!A !(B (C (D)+!C !(D))+!B (C+!(D))))) */ ;
    defparam i20648_else_4_lut.init = 16'h581f;
    LUT4 mux_207_Mux_8_i172_3_lut_3_lut_rep_815 (.A(index_q[1]), .B(index_q[0]), 
         .C(index_q[2]), .Z(n29475)) /* synthesis lut_function=(!(A (B (C))+!A !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_8_i172_3_lut_3_lut_rep_815.init = 16'h7a7a;
    LUT4 mux_207_Mux_7_i716_3_lut_3_lut_4_lut (.A(index_q[1]), .B(index_q[0]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n716_adj_3258)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C+!(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_7_i716_3_lut_3_lut_4_lut.init = 16'h0f81;
    PFUMX i21404 (.BLUT(n23884), .ALUT(n23885), .C0(index_i[5]), .Z(n23886));
    LUT4 mux_207_Mux_5_i30_3_lut_4_lut (.A(index_q[1]), .B(index_q[0]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n30_adj_3259)) /* synthesis lut_function=(A ((D)+!B)+!A !(B (D)+!B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_5_i30_3_lut_4_lut.init = 16'haa67;
    LUT4 mux_207_Mux_2_i557_3_lut_3_lut_4_lut (.A(index_q[1]), .B(index_q[0]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n557_adj_3014)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C+!(D))+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_2_i557_3_lut_3_lut_4_lut.init = 16'h0f18;
    LUT4 i20902_3_lut_4_lut (.A(index_q[1]), .B(index_q[0]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n23384)) /* synthesis lut_function=(!(A (B (C (D))+!B (D))+!A (B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i20902_3_lut_4_lut.init = 16'h18aa;
    LUT4 mux_207_Mux_4_i526_3_lut_3_lut_4_lut (.A(index_q[1]), .B(index_q[0]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n526_adj_3260)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A !(B ((D)+!C)+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_4_i526_3_lut_3_lut_4_lut.init = 16'h7e0f;
    LUT4 i20886_3_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[0]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n23368)) /* synthesis lut_function=(A (B (C+(D))+!B !(D))+!A !(B (C+(D))+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i20886_3_lut_4_lut_4_lut.init = 16'h99a7;
    LUT4 n262_bdd_3_lut_26871_3_lut_4_lut (.A(index_q[1]), .B(index_q[0]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n27748)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C (D)))+!A (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam n262_bdd_3_lut_26871_3_lut_4_lut.init = 16'h0fa7;
    LUT4 mux_207_Mux_7_i620_3_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[0]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n620_adj_3261)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_7_i620_3_lut_4_lut_4_lut.init = 16'h85a5;
    LUT4 mux_207_Mux_8_i93_3_lut_3_lut_4_lut (.A(index_q[1]), .B(index_q[0]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n93_adj_3262)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_8_i93_3_lut_3_lut_4_lut.init = 16'h0f85;
    LUT4 i20691_3_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[0]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n23173)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i20691_3_lut_4_lut_4_lut.init = 16'h5a58;
    LUT4 i21474_3_lut_3_lut_4_lut (.A(index_q[1]), .B(index_q[0]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n23956)) /* synthesis lut_function=(!(A (B (D)+!B !(C+!(D)))+!A !(B (C (D))+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i21474_3_lut_3_lut_4_lut.init = 16'h71aa;
    LUT4 mux_207_Mux_0_i762_3_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[0]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n762_adj_3263)) /* synthesis lut_function=(A (B+!(D))+!A !(B ((D)+!C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_0_i762_3_lut_4_lut_4_lut.init = 16'h98fa;
    LUT4 i24617_2_lut_rep_816 (.A(index_q[4]), .B(index_q[3]), .Z(n29476)) /* synthesis lut_function=((B)+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i24617_2_lut_rep_816.init = 16'hdddd;
    LUT4 mux_207_Mux_3_i797_3_lut_4_lut (.A(index_q[4]), .B(index_q[3]), 
         .C(n796), .D(n29475), .Z(n797)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_3_i797_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_206_Mux_2_i716_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), 
         .B(index_i[2]), .C(index_i[3]), .D(index_i[0]), .Z(n716_adj_3264)) /* synthesis lut_function=(!(A (B)+!A !(B (C+!(D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_2_i716_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h6367;
    LUT4 n699_bdd_4_lut (.A(n29068), .B(index_q[6]), .C(n29133), .D(index_q[5]), 
         .Z(n28501)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C+!(D))+!B (D))) */ ;
    defparam n699_bdd_4_lut.init = 16'hd1cc;
    LUT4 n28504_bdd_3_lut (.A(n28504), .B(n28501), .C(index_q[4]), .Z(n23298)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n28504_bdd_3_lut.init = 16'hcaca;
    LUT4 i22280_3_lut_3_lut_4_lut (.A(n29177), .B(index_i[3]), .C(n316), 
         .D(index_i[4]), .Z(n24781)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i22280_3_lut_3_lut_4_lut.init = 16'hf011;
    PFUMX i21980 (.BLUT(n23214), .ALUT(n317_adj_3183), .C0(index_i[5]), 
          .Z(n24481));
    PFUMX i21503 (.BLUT(n23983), .ALUT(n23984), .C0(index_i[4]), .Z(n23985));
    LUT4 i20931_3_lut_3_lut_4_lut (.A(n29459), .B(index_q[2]), .C(n29373), 
         .D(index_q[3]), .Z(n23413)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i20931_3_lut_3_lut_4_lut.init = 16'hf077;
    LUT4 i5071_2_lut_rep_657 (.A(index_q[0]), .B(index_q[2]), .Z(n29317)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i5071_2_lut_rep_657.init = 16'h6666;
    LUT4 mux_207_Mux_8_i301_3_lut_4_lut (.A(n29459), .B(index_q[2]), .C(index_q[3]), 
         .D(n29475), .Z(n301_adj_3071)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_8_i301_3_lut_4_lut.init = 16'h8f80;
    LUT4 i11126_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n13422)) /* synthesis lut_function=(!(A (B (D)+!B (C+!(D)))+!A !(B (D)+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i11126_3_lut_4_lut_4_lut.init = 16'h4699;
    LUT4 i14391_1_lut_2_lut_3_lut_4_lut (.A(n29176), .B(index_i[3]), .C(index_i[5]), 
         .D(index_i[4]), .Z(n381)) /* synthesis lut_function=(!(A (C+(D))+!A (B (C+(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i14391_1_lut_2_lut_3_lut_4_lut.init = 16'h010f;
    LUT4 n954_bdd_3_lut_26400_3_lut_4_lut (.A(n29459), .B(index_q[2]), .C(n29475), 
         .D(index_q[3]), .Z(n28171)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam n954_bdd_3_lut_26400_3_lut_4_lut.init = 16'hf077;
    LUT4 i24628_2_lut_rep_385_3_lut_4_lut (.A(n29459), .B(index_q[2]), .C(index_q[5]), 
         .D(n29369), .Z(n29045)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i24628_2_lut_rep_385_3_lut_4_lut.init = 16'h0f7f;
    LUT4 mux_206_Mux_10_i637_3_lut_4_lut_4_lut (.A(n29178), .B(index_i[4]), 
         .C(index_i[5]), .D(n29088), .Z(n637_adj_3236)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_10_i637_3_lut_4_lut_4_lut.init = 16'h1f1c;
    PFUMX i22351 (.BLUT(n19977), .ALUT(n573_adj_3265), .C0(index_q[5]), 
          .Z(n24852));
    LUT4 mux_206_Mux_8_i860_3_lut_4_lut (.A(n29179), .B(index_i[3]), .C(index_i[4]), 
         .D(n29147), .Z(n860_adj_3266)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_8_i860_3_lut_4_lut.init = 16'h08f8;
    LUT4 n986_bdd_4_lut (.A(n29064), .B(index_i[6]), .C(n29147), .D(index_i[5]), 
         .Z(n28575)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C+!(D))+!B (D))) */ ;
    defparam n986_bdd_4_lut.init = 16'hd1cc;
    PFUMX i21407 (.BLUT(n23887), .ALUT(n23888), .C0(index_i[5]), .Z(n23889));
    LUT4 n28578_bdd_3_lut (.A(n28578), .B(n28575), .C(index_i[4]), .Z(n23316)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n28578_bdd_3_lut.init = 16'hcaca;
    LUT4 index_i_4__bdd_3_lut_26288_4_lut (.A(n29179), .B(index_i[3]), .C(index_i[5]), 
         .D(index_i[4]), .Z(n28146)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam index_i_4__bdd_3_lut_26288_4_lut.init = 16'hf080;
    LUT4 mux_206_Mux_3_i252_3_lut_4_lut (.A(n29179), .B(index_i[3]), .C(index_i[4]), 
         .D(n16610), .Z(n252_adj_3103)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_3_i252_3_lut_4_lut.init = 16'h08f8;
    LUT4 mux_206_Mux_10_i62_3_lut_3_lut_4_lut (.A(n29179), .B(index_i[3]), 
         .C(n29147), .D(index_i[4]), .Z(n62_adj_3228)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_10_i62_3_lut_3_lut_4_lut.init = 16'hf077;
    LUT4 mux_206_Mux_6_i955_3_lut_4_lut (.A(n29179), .B(index_i[3]), .C(index_i[4]), 
         .D(n29042), .Z(n955_adj_3267)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_6_i955_3_lut_4_lut.init = 16'h8f80;
    LUT4 i20598_3_lut_4_lut_4_lut (.A(index_q[0]), .B(n29395), .C(index_q[3]), 
         .D(n29367), .Z(n23080)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i20598_3_lut_4_lut_4_lut.init = 16'hcfc5;
    LUT4 mux_207_Mux_3_i62_3_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[4]), .D(n812_adj_3074), .Z(n62_adj_3202)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_3_i62_3_lut_4_lut.init = 16'h6f60;
    LUT4 i22282_3_lut_4_lut (.A(n29179), .B(index_i[3]), .C(index_i[4]), 
         .D(n364_adj_3198), .Z(n24783)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i22282_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_206_Mux_3_i189_3_lut_3_lut_4_lut (.A(n29179), .B(index_i[3]), 
         .C(index_i[4]), .D(n29146), .Z(n189_adj_3094)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_3_i189_3_lut_3_lut_4_lut.init = 16'h08f8;
    LUT4 i22507_3_lut_3_lut_4_lut (.A(n29180), .B(index_i[3]), .C(n93_adj_3268), 
         .D(index_i[4]), .Z(n25008)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i22507_3_lut_3_lut_4_lut.init = 16'hf077;
    PFUMX mux_207_Mux_1_i636 (.BLUT(n620), .ALUT(n635), .C0(index_q[4]), 
          .Z(n636_adj_3269)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 i12689_3_lut_3_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n15097)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12689_3_lut_3_lut_3_lut_4_lut.init = 16'h10ff;
    LUT4 mux_206_Mux_10_i252_3_lut_4_lut_4_lut (.A(n29180), .B(index_i[3]), 
         .C(index_i[4]), .D(n29176), .Z(n252_adj_3227)) /* synthesis lut_function=(!(A (B (C)+!B !(C+(D)))+!A !(B+(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_10_i252_3_lut_4_lut_4_lut.init = 16'h7f7c;
    PFUMX i21413 (.BLUT(n23893), .ALUT(n23894), .C0(index_i[5]), .Z(n23895));
    LUT4 i22506_3_lut_4_lut (.A(n29180), .B(index_i[3]), .C(index_i[4]), 
         .D(n46_adj_3270), .Z(n25007)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i22506_3_lut_4_lut.init = 16'h8f80;
    LUT4 i22511_3_lut_4_lut (.A(n29180), .B(index_i[3]), .C(index_i[4]), 
         .D(n220), .Z(n25012)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i22511_3_lut_4_lut.init = 16'hf808;
    PFUMX i21416 (.BLUT(n23896), .ALUT(n23897), .C0(index_i[5]), .Z(n23898));
    LUT4 mux_206_Mux_3_i221_3_lut_4_lut (.A(n29180), .B(index_i[3]), .C(index_i[4]), 
         .D(n29143), .Z(n221_adj_3102)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_3_i221_3_lut_4_lut.init = 16'h08f8;
    LUT4 i12705_3_lut (.A(index_q[2]), .B(index_q[1]), .C(index_q[0]), 
         .Z(n85)) /* synthesis lut_function=(!(A (B (C))+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i12705_3_lut.init = 16'h3b3b;
    PFUMX i21419 (.BLUT(n23899), .ALUT(n23900), .C0(index_i[5]), .Z(n23901));
    LUT4 i23668_3_lut (.A(n23980), .B(n29502), .C(index_q[4]), .Z(n23982)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23668_3_lut.init = 16'hcaca;
    LUT4 n557_bdd_3_lut_3_lut_4_lut (.A(n29180), .B(index_i[3]), .C(index_i[6]), 
         .D(n29146), .Z(n28343)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n557_bdd_3_lut_3_lut_4_lut.init = 16'h08f8;
    LUT4 i24695_2_lut (.A(index_i[5]), .B(index_i[4]), .Z(n24303)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i24695_2_lut.init = 16'heeee;
    LUT4 mux_206_Mux_3_i747_3_lut (.A(n29432), .B(n498), .C(index_i[3]), 
         .Z(n747_adj_3271)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_3_i747_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut (.A(index_i[0]), .B(index_i[4]), .C(index_i[2]), .Z(n22576)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_3_lut.init = 16'hfefe;
    LUT4 n627_bdd_3_lut_26738 (.A(n29333), .B(n29387), .C(index_q[3]), 
         .Z(n28662)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n627_bdd_3_lut_26738.init = 16'hcaca;
    LUT4 mux_207_Mux_3_i924_3_lut (.A(n908_adj_2960), .B(index_q[0]), .C(index_q[4]), 
         .Z(n924_adj_3272)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_3_i924_3_lut.init = 16'hcaca;
    LUT4 n27782_bdd_3_lut_3_lut (.A(n1021), .B(index_i[8]), .C(n27782), 
         .Z(n27783)) /* synthesis lut_function=(A (B+(C))+!A !(B+!(C))) */ ;
    defparam n27782_bdd_3_lut_3_lut.init = 16'hb8b8;
    LUT4 mux_207_Mux_3_i891_3_lut (.A(n541_adj_3084), .B(n890_adj_3273), 
         .C(index_q[4]), .Z(n891_adj_3274)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_3_i891_3_lut.init = 16'hcaca;
    PFUMX i21422 (.BLUT(n23902), .ALUT(n23903), .C0(index_i[5]), .Z(n23904));
    PFUMX i21506 (.BLUT(n23986), .ALUT(n23987), .C0(index_i[4]), .Z(n23988));
    LUT4 i20920_3_lut (.A(n32031), .B(n29392), .C(index_q[3]), .Z(n23402)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20920_3_lut.init = 16'hcaca;
    PFUMX i21981 (.BLUT(n349_adj_3275), .ALUT(n23217), .C0(index_i[5]), 
          .Z(n24482));
    L6MUX21 i21982 (.D0(n23220), .D1(n23223), .SD(index_i[5]), .Z(n24483));
    L6MUX21 i21983 (.D0(n23229), .D1(n23232), .SD(index_i[5]), .Z(n24484));
    PFUMX i22352 (.BLUT(n605_adj_3276), .ALUT(n636_adj_3277), .C0(index_q[5]), 
          .Z(n24853));
    LUT4 i21406_3_lut_3_lut_4_lut (.A(n29177), .B(index_i[3]), .C(n93_adj_3278), 
         .D(index_i[4]), .Z(n23888)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21406_3_lut_3_lut_4_lut.init = 16'h11f0;
    LUT4 mux_206_Mux_5_i15_3_lut (.A(n29443), .B(n32056), .C(index_i[3]), 
         .Z(n15_adj_3279)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_5_i15_3_lut.init = 16'hcaca;
    LUT4 mux_206_Mux_6_i653_3_lut (.A(n29435), .B(n619), .C(index_i[3]), 
         .Z(n653_adj_3047)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_6_i653_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_3_i669_3_lut (.A(n653_adj_3193), .B(n668_adj_3081), 
         .C(index_q[4]), .Z(n669_adj_3280)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_3_i669_3_lut.init = 16'hcaca;
    LUT4 mux_206_Mux_5_i124_3_lut (.A(n645), .B(n29427), .C(index_i[3]), 
         .Z(n124_adj_3281)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_5_i124_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_0_i986_3_lut (.A(n29391), .B(n985_adj_3282), .C(index_q[3]), 
         .Z(n986_adj_3156)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_0_i986_3_lut.init = 16'hcaca;
    PFUMX i22353 (.BLUT(n23082), .ALUT(n700_adj_3283), .C0(index_q[5]), 
          .Z(n24854));
    PFUMX mux_207_Mux_2_i891 (.BLUT(n875_adj_3284), .ALUT(n890_adj_3285), 
          .C0(index_q[4]), .Z(n891_adj_3286)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    L6MUX21 i22354 (.D0(n732_adj_3287), .D1(n23091), .SD(index_q[5]), 
            .Z(n24855));
    LUT4 mux_206_Mux_5_i397_3_lut (.A(n29447), .B(n204), .C(index_i[3]), 
         .Z(n397_adj_3288)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_5_i397_3_lut.init = 16'hcaca;
    PFUMX i22355 (.BLUT(n797_adj_3289), .ALUT(n828_adj_3157), .C0(index_q[5]), 
          .Z(n24856));
    LUT4 i11136_4_lut (.A(n29367), .B(n29168), .C(index_q[3]), .D(index_q[4]), 
         .Z(n13432)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B ((D)+!C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i11136_4_lut.init = 16'h3afa;
    LUT4 n262_bdd_3_lut_26744 (.A(n29389), .B(n32055), .C(index_q[3]), 
         .Z(n28676)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n262_bdd_3_lut_26744.init = 16'hcaca;
    PFUMX i21425 (.BLUT(n23905), .ALUT(n23906), .C0(index_i[5]), .Z(n23907));
    PFUMX mux_207_Mux_2_i860 (.BLUT(n844_adj_2953), .ALUT(n859_adj_3290), 
          .C0(index_q[4]), .Z(n860_adj_3291)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    PFUMX i21428 (.BLUT(n23908), .ALUT(n23909), .C0(index_i[5]), .Z(n23910));
    LUT4 n627_bdd_3_lut (.A(n29333), .B(n588), .C(index_q[3]), .Z(n28678)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n627_bdd_3_lut.init = 16'hacac;
    LUT4 mux_206_Mux_5_i506_3_lut (.A(n32028), .B(n32023), .C(index_i[3]), 
         .Z(n506_adj_3292)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_5_i506_3_lut.init = 16'hcaca;
    L6MUX21 i21985 (.D0(n23238), .D1(n636_adj_3293), .SD(index_i[5]), 
            .Z(n24486));
    LUT4 mux_207_Mux_0_i188_3_lut (.A(n29472), .B(n101), .C(index_q[3]), 
         .Z(n188_adj_3294)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_0_i188_3_lut.init = 16'hcaca;
    PFUMX i21986 (.BLUT(n23241), .ALUT(n700_adj_3029), .C0(index_i[5]), 
          .Z(n24487));
    PFUMX i20678 (.BLUT(n23158), .ALUT(n23159), .C0(index_q[4]), .Z(n23160));
    LUT4 index_i_5__bdd_3_lut_25646 (.A(index_i[5]), .B(n645), .C(n32018), 
         .Z(n27187)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam index_i_5__bdd_3_lut_25646.init = 16'he4e4;
    LUT4 i23686_3_lut (.A(n23956), .B(n23957), .C(index_q[4]), .Z(n23958)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23686_3_lut.init = 16'hcaca;
    PFUMX i22356 (.BLUT(n860_adj_3295), .ALUT(n891_adj_3296), .C0(index_q[5]), 
          .Z(n24857));
    LUT4 mux_207_Mux_3_i476_3_lut (.A(n460_adj_3024), .B(n285_adj_3025), 
         .C(index_q[4]), .Z(n476_adj_3297)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_3_i476_3_lut.init = 16'hcaca;
    LUT4 i20913_3_lut (.A(n29395), .B(n32029), .C(index_q[3]), .Z(n23395)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20913_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_3_i413_3_lut (.A(n397_adj_3298), .B(n29281), .C(index_q[4]), 
         .Z(n413_adj_3299)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_3_i413_3_lut.init = 16'hcaca;
    LUT4 index_i_0__bdd_4_lut_27100 (.A(index_i[0]), .B(index_i[3]), .C(index_i[1]), 
         .D(index_i[2]), .Z(n29481)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C (D)))+!A !(B (C+!(D))+!B !(C+(D))))) */ ;
    defparam index_i_0__bdd_4_lut_27100.init = 16'h4ae7;
    LUT4 mux_207_Mux_3_i286_4_lut (.A(n93_adj_3158), .B(index_q[2]), .C(index_q[4]), 
         .D(n16645), .Z(n286_adj_3300)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_3_i286_4_lut.init = 16'h3aca;
    L6MUX21 i21988 (.D0(n23244), .D1(n23931), .SD(index_i[5]), .Z(n24489));
    PFUMX i21990 (.BLUT(n924_adj_3301), .ALUT(n23940), .C0(index_i[5]), 
          .Z(n24491));
    LUT4 mux_207_Mux_3_i158_3_lut (.A(n142_adj_3168), .B(n157_adj_3174), 
         .C(index_q[4]), .Z(n158_adj_3302)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_3_i158_3_lut.init = 16'hcaca;
    PFUMX i27133 (.BLUT(n29572), .ALUT(n29573), .C0(index_q[0]), .Z(n29574));
    LUT4 mux_207_Mux_3_i125_3_lut (.A(n46_adj_2991), .B(n526_adj_3260), 
         .C(index_q[4]), .Z(n125_adj_3303)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_3_i125_3_lut.init = 16'hcaca;
    LUT4 mux_206_Mux_0_i397_3_lut (.A(n32019), .B(n32020), .C(index_i[3]), 
         .Z(n397_adj_3304)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i397_3_lut.init = 16'hcaca;
    LUT4 i23765_3_lut (.A(n23392), .B(n23393), .C(index_q[4]), .Z(n23394)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23765_3_lut.init = 16'hcaca;
    LUT4 mux_206_Mux_5_i859_3_lut (.A(n851), .B(n29443), .C(index_i[3]), 
         .Z(n859_adj_3305)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_5_i859_3_lut.init = 16'hcaca;
    PFUMX i21991 (.BLUT(n987), .ALUT(n23943), .C0(index_i[5]), .Z(n24492));
    LUT4 mux_206_Mux_5_i875_3_lut (.A(n645), .B(n32018), .C(index_i[3]), 
         .Z(n875_adj_3306)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_5_i875_3_lut.init = 16'hcaca;
    LUT4 mux_206_Mux_0_i285_3_lut (.A(n29382), .B(n32039), .C(index_i[3]), 
         .Z(n285_adj_3182)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i285_3_lut.init = 16'hcaca;
    LUT4 mux_206_Mux_5_i781_3_lut_4_lut_4_lut_then_4_lut (.A(index_i[3]), 
         .B(index_i[0]), .C(index_i[4]), .D(index_i[2]), .Z(n29483)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_5_i781_3_lut_4_lut_4_lut_then_4_lut.init = 16'hece0;
    LUT4 mux_207_Mux_1_i301_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n301_adj_3307)) /* synthesis lut_function=(A (B (C+(D))+!B !(D))+!A !(B (C+(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_1_i301_3_lut_4_lut_4_lut.init = 16'h99b6;
    LUT4 mux_207_Mux_5_i31_3_lut (.A(n15_adj_3113), .B(n30_adj_3259), .C(index_q[4]), 
         .Z(n31_adj_3308)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_5_i31_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_1_i317_3_lut (.A(n301_adj_3307), .B(n908_adj_3309), 
         .C(index_q[4]), .Z(n317_adj_3310)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_1_i317_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_3_i30_3_lut_4_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n30_adj_3311)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C+!(D)))) */ ;
    defparam mux_207_Mux_3_i30_3_lut_4_lut_3_lut_4_lut.init = 16'hfe11;
    LUT4 i20603_then_4_lut (.A(index_i[0]), .B(index_i[4]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n29516)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C))+!A (B (C)+!B !(C+!(D)))) */ ;
    defparam i20603_then_4_lut.init = 16'hc34a;
    LUT4 i11257_3_lut_4_lut_3_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[4]), 
         .Z(n13556)) /* synthesis lut_function=(!(A (B)+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i11257_3_lut_4_lut_3_lut.init = 16'h6262;
    LUT4 mux_207_Mux_6_i7_3_lut_4_lut_3_lut_rep_736 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29396)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_6_i7_3_lut_4_lut_3_lut_rep_736.init = 16'hd6d6;
    PFUMX i20837 (.BLUT(n23317), .ALUT(n23318), .C0(index_q[5]), .Z(n23319));
    LUT4 mux_206_Mux_5_i781_3_lut_4_lut_4_lut_else_4_lut (.A(index_i[3]), 
         .B(index_i[0]), .C(index_i[4]), .Z(n29482)) /* synthesis lut_function=(!(A (C)+!A (B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_5_i781_3_lut_4_lut_4_lut_else_4_lut.init = 16'h1f1f;
    LUT4 mux_206_Mux_4_i61_3_lut (.A(n29429), .B(n29445), .C(index_i[3]), 
         .Z(n61)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_4_i61_3_lut.init = 16'hcaca;
    PFUMX i22375 (.BLUT(n94_adj_3312), .ALUT(n23094), .C0(index_q[5]), 
          .Z(n24876));
    LUT4 mux_206_Mux_0_i188_3_lut (.A(n29384), .B(n187), .C(index_i[3]), 
         .Z(n188_adj_3313)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i188_3_lut.init = 16'hcaca;
    PFUMX i22008 (.BLUT(n94_adj_3314), .ALUT(n23382), .C0(index_q[5]), 
          .Z(n24509));
    LUT4 mux_206_Mux_4_i270_3_lut (.A(n29442), .B(n32028), .C(index_i[3]), 
         .Z(n270_adj_3315)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_4_i270_3_lut.init = 16'hcaca;
    LUT4 mux_206_Mux_4_i15_3_lut (.A(n32023), .B(n931), .C(index_i[3]), 
         .Z(n15_adj_3125)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_4_i15_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_0_i908_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n908_adj_3031)) /* synthesis lut_function=(!(A (B (C (D))+!B !(D))+!A (B+((D)+!C)))) */ ;
    defparam mux_207_Mux_0_i908_3_lut_4_lut_4_lut.init = 16'h2a98;
    LUT4 mux_207_Mux_7_i762_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), 
         .B(index_q[1]), .C(index_q[3]), .D(index_q[2]), .Z(n762_adj_3316)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A (B (C (D)+!C !(D))+!B !(C)))) */ ;
    defparam mux_207_Mux_7_i762_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h1cf0;
    PFUMX i20840 (.BLUT(n23320), .ALUT(n23321), .C0(index_q[5]), .Z(n23322));
    LUT4 i23645_3_lut (.A(n29523), .B(n124_adj_3032), .C(index_i[4]), 
         .Z(n25009)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23645_3_lut.init = 16'hcaca;
    PFUMX mux_207_Mux_3_i763 (.BLUT(n747_adj_3317), .ALUT(n762_adj_3062), 
          .C0(index_q[4]), .Z(n763_adj_3318)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 i3906_2_lut_rep_766 (.A(index_i[0]), .B(index_i[1]), .Z(n29426)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i3906_2_lut_rep_766.init = 16'h6666;
    LUT4 i20901_3_lut (.A(n900_adj_3319), .B(n32036), .C(index_q[3]), 
         .Z(n23383)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20901_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_2_i716_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), 
         .B(index_q[1]), .C(index_q[3]), .D(index_q[2]), .Z(n716_adj_3161)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)+!C !(D)))+!A (B (D)+!B !((D)+!C)))) */ ;
    defparam mux_207_Mux_2_i716_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h31cf;
    LUT4 mux_206_Mux_4_i348_3_lut (.A(n32025), .B(n29441), .C(index_i[3]), 
         .Z(n348)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_4_i348_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_0_i219_3_lut_3_lut_rep_832 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n32033)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_0_i219_3_lut_3_lut_rep_832.init = 16'h9393;
    PFUMX i22377 (.BLUT(n221_adj_3320), .ALUT(n252_adj_3321), .C0(index_q[5]), 
          .Z(n24878));
    LUT4 mux_206_Mux_4_i668_3_lut (.A(n29385), .B(n32039), .C(index_i[3]), 
         .Z(n668_adj_3322)) /* synthesis lut_function=(A (B (C))+!A (B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_4_i668_3_lut.init = 16'hc5c5;
    PFUMX i21509 (.BLUT(n23989), .ALUT(n23990), .C0(index_i[4]), .Z(n23991));
    LUT4 mux_206_Mux_4_i684_3_lut (.A(n619), .B(n660), .C(index_i[3]), 
         .Z(n684_adj_3323)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_4_i684_3_lut.init = 16'hcaca;
    PFUMX i21512 (.BLUT(n23992), .ALUT(n23993), .C0(index_i[4]), .Z(n23994));
    PFUMX i22378 (.BLUT(n286_adj_3324), .ALUT(n23100), .C0(index_q[5]), 
          .Z(n24879));
    LUT4 i23784_3_lut (.A(n29519), .B(n23381), .C(index_q[4]), .Z(n23382)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23784_3_lut.init = 16'hcaca;
    PFUMX i22379 (.BLUT(n349_adj_3325), .ALUT(n23103), .C0(index_q[5]), 
          .Z(n24880));
    LUT4 mux_207_Mux_7_i108_3_lut_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n108)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_7_i108_3_lut_3_lut.init = 16'hc6c6;
    L6MUX21 i22009 (.D0(n23385), .D1(n23388), .SD(index_q[5]), .Z(n24510));
    LUT4 i13094_2_lut_rep_473_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n29133)) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;
    defparam i13094_2_lut_rep_473_3_lut_4_lut.init = 16'he000;
    PFUMX i21518 (.BLUT(n23998), .ALUT(n23999), .C0(index_i[4]), .Z(n24000));
    PFUMX i22011 (.BLUT(n23391), .ALUT(n317_adj_3310), .C0(index_q[5]), 
          .Z(n24512));
    LUT4 i23505_3_lut (.A(n27620), .B(n124_adj_3326), .C(index_q[4]), 
         .Z(n24978)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23505_3_lut.init = 16'hcaca;
    LUT4 i20605_3_lut (.A(n32039), .B(n29435), .C(index_i[3]), .Z(n23087)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20605_3_lut.init = 16'hcaca;
    LUT4 i20604_3_lut (.A(n29385), .B(n619), .C(index_i[3]), .Z(n23086)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20604_3_lut.init = 16'hcaca;
    LUT4 i20868_3_lut (.A(n526_adj_3252), .B(n15_adj_3053), .C(index_q[4]), 
         .Z(n23350)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20868_3_lut.init = 16'hcaca;
    PFUMX i22012 (.BLUT(n349_adj_3327), .ALUT(n23394), .C0(index_q[5]), 
          .Z(n24513));
    LUT4 mux_207_Mux_0_i963_3_lut_3_lut_rep_727 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29387)) /* synthesis lut_function=(!(A (B)+!A (B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_0_i963_3_lut_3_lut_rep_727.init = 16'h3636;
    LUT4 i23926_3_lut (.A(n23086), .B(n23087), .C(index_i[4]), .Z(n23088)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23926_3_lut.init = 16'hcaca;
    L6MUX21 i22013 (.D0(n23397), .D1(n23400), .SD(index_q[5]), .Z(n24514));
    LUT4 i20865_3_lut (.A(n397_adj_3328), .B(n475_adj_2987), .C(index_q[4]), 
         .Z(n23347)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20865_3_lut.init = 16'hcaca;
    LUT4 i20892_3_lut (.A(n404), .B(n29357), .C(index_q[3]), .Z(n23374)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20892_3_lut.init = 16'hcaca;
    L6MUX21 i22014 (.D0(n23403), .D1(n23406), .SD(index_q[5]), .Z(n24515));
    LUT4 i23617_3_lut (.A(n23374), .B(n23375), .C(index_q[4]), .Z(n23376)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23617_3_lut.init = 16'hcaca;
    LUT4 i20863_3_lut (.A(n348_adj_3329), .B(n443_adj_3099), .C(index_q[4]), 
         .Z(n23345)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20863_3_lut.init = 16'hcaca;
    LUT4 i20862_3_lut (.A(n397_adj_3328), .B(n731), .C(index_q[4]), .Z(n23344)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20862_3_lut.init = 16'hcaca;
    LUT4 i20860_3_lut (.A(n364_adj_3055), .B(n379_adj_3063), .C(index_q[4]), 
         .Z(n23342)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20860_3_lut.init = 16'hcaca;
    LUT4 i20859_3_lut (.A(n333_adj_3330), .B(n348_adj_3329), .C(index_q[4]), 
         .Z(n23341)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20859_3_lut.init = 16'hcaca;
    LUT4 i20686_3_lut (.A(n29388), .B(n325), .C(index_q[3]), .Z(n23168)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20686_3_lut.init = 16'hcaca;
    PFUMX i20849 (.BLUT(n23329), .ALUT(n23330), .C0(index_q[5]), .Z(n23331));
    LUT4 i23744_3_lut (.A(n23167), .B(n23168), .C(index_q[4]), .Z(n23169)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23744_3_lut.init = 16'hcaca;
    PFUMX i27131 (.BLUT(n29569), .ALUT(n29570), .C0(index_q[1]), .Z(n29571));
    LUT4 i12684_3_lut (.A(index_i[3]), .B(index_i[1]), .C(index_i[0]), 
         .Z(n15092)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12684_3_lut.init = 16'hc8c8;
    LUT4 mux_206_Mux_3_i348_3_lut (.A(n29436), .B(n29446), .C(index_i[3]), 
         .Z(n348_adj_3331)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_3_i348_3_lut.init = 16'hcaca;
    PFUMX i22384 (.BLUT(n669_adj_3332), .ALUT(n700_adj_3333), .C0(index_q[5]), 
          .Z(n24885));
    LUT4 i20682_3_lut (.A(n588), .B(n29395), .C(index_q[3]), .Z(n23164)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20682_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_1_i924_3_lut (.A(n316_adj_3334), .B(n412_adj_3335), 
         .C(index_q[4]), .Z(n924_adj_3336)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_1_i924_3_lut.init = 16'hcaca;
    LUT4 i25856_then_4_lut (.A(index_q[0]), .B(index_q[4]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n29570)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)+!C !(D))+!B (C (D)))) */ ;
    defparam i25856_then_4_lut.init = 16'hda0e;
    LUT4 i22389_4_lut (.A(n23175), .B(n1002_adj_3250), .C(index_q[5]), 
         .D(index_q[4]), .Z(n24890)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;
    defparam i22389_4_lut.init = 16'hfaca;
    LUT4 mux_206_Mux_3_i908_3_lut (.A(n29431), .B(n29445), .C(index_i[3]), 
         .Z(n908_adj_3337)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_3_i908_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_4_i860_3_lut (.A(n506_adj_3338), .B(n15_adj_3339), 
         .C(index_q[4]), .Z(n860_adj_3340)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_4_i860_3_lut.init = 16'hcaca;
    PFUMX i22385 (.BLUT(n23133), .ALUT(n763_adj_3082), .C0(index_q[5]), 
          .Z(n24886));
    LUT4 mux_207_Mux_5_i731_3_lut (.A(n32029), .B(n29388), .C(index_q[3]), 
         .Z(n731_adj_3341)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_5_i731_3_lut.init = 16'hcaca;
    LUT4 i23746_3_lut (.A(n23164), .B(n23165), .C(index_q[4]), .Z(n23166)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23746_3_lut.init = 16'hcaca;
    LUT4 i12756_3_lut_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n15165)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B !(C+!(D))))) */ ;
    defparam i12756_3_lut_3_lut_3_lut_4_lut.init = 16'h10ff;
    L6MUX21 i22016 (.D0(n23412), .D1(n636_adj_3269), .SD(index_q[5]), 
            .Z(n24517));
    PFUMX i22017 (.BLUT(n23415), .ALUT(n700_adj_3342), .C0(index_q[5]), 
          .Z(n24518));
    LUT4 mux_206_Mux_2_i270_3_lut (.A(n29443), .B(n29407), .C(index_i[3]), 
         .Z(n270_adj_3343)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_2_i270_3_lut.init = 16'hcaca;
    LUT4 mux_206_Mux_2_i316_3_lut (.A(n29444), .B(n29429), .C(index_i[3]), 
         .Z(n316_adj_3344)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_2_i316_3_lut.init = 16'hcaca;
    PFUMX i20852 (.BLUT(n23332), .ALUT(n23333), .C0(index_q[5]), .Z(n23334));
    LUT4 i20851_3_lut (.A(n491_adj_3345), .B(n506_adj_3346), .C(index_q[4]), 
         .Z(n23333)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20851_3_lut.init = 16'hcaca;
    LUT4 i20850_3_lut (.A(n460), .B(n475_adj_3142), .C(index_q[4]), .Z(n23332)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20850_3_lut.init = 16'hcaca;
    LUT4 mux_206_Mux_2_i397_3_lut (.A(n32039), .B(n29409), .C(index_i[3]), 
         .Z(n397_adj_3347)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_2_i397_3_lut.init = 16'hcaca;
    LUT4 i23753_3_lut (.A(n23413), .B(n23414), .C(index_q[4]), .Z(n23415)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23753_3_lut.init = 16'hcaca;
    LUT4 i25856_else_4_lut (.A(index_q[0]), .B(index_q[4]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n29569)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C))+!A (B (C)+!B (C+(D)))) */ ;
    defparam i25856_else_4_lut.init = 16'hf178;
    LUT4 i23756_3_lut (.A(n23131), .B(n23132), .C(index_q[4]), .Z(n23133)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23756_3_lut.init = 16'hcaca;
    L6MUX21 i22019 (.D0(n23418), .D1(n23421), .SD(index_q[5]), .Z(n24520));
    LUT4 mux_207_Mux_4_i700_3_lut (.A(n684_adj_3348), .B(index_q[1]), .C(index_q[4]), 
         .Z(n700_adj_3333)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_4_i700_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_4_i669_3_lut (.A(n781), .B(n668_adj_3054), .C(index_q[4]), 
         .Z(n669_adj_3332)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_4_i669_3_lut.init = 16'hcaca;
    PFUMX i22386 (.BLUT(n23166), .ALUT(n828_adj_3349), .C0(index_q[5]), 
          .Z(n24887));
    LUT4 i20848_3_lut (.A(n251_adj_2952), .B(n443_adj_2969), .C(index_q[4]), 
         .Z(n23330)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20848_3_lut.init = 16'hcaca;
    LUT4 i20847_3_lut (.A(n460), .B(n16626), .C(index_q[4]), .Z(n23329)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;
    defparam i20847_3_lut.init = 16'h3a3a;
    PFUMX mux_207_Mux_5_i732 (.BLUT(n13422), .ALUT(n731_adj_3341), .C0(index_q[4]), 
          .Z(n732_adj_3287)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 mux_207_Mux_4_i542_3_lut (.A(n526_adj_3260), .B(n506_adj_3346), 
         .C(index_q[4]), .Z(n542_adj_3175)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_4_i542_3_lut.init = 16'hcaca;
    LUT4 i22383_4_lut (.A(n29136), .B(n29480), .C(index_q[5]), .D(index_q[4]), 
         .Z(n24884)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam i22383_4_lut.init = 16'hc5ca;
    PFUMX i22387 (.BLUT(n860_adj_3340), .ALUT(n23169), .C0(index_q[5]), 
          .Z(n24888));
    LUT4 i21526_3_lut (.A(n29441), .B(n29432), .C(index_i[3]), .Z(n24008)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21526_3_lut.init = 16'hcaca;
    LUT4 i21525_3_lut (.A(n29403), .B(n325_adj_2972), .C(index_i[3]), 
         .Z(n24007)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21525_3_lut.init = 16'hcaca;
    LUT4 i25816_then_4_lut (.A(index_q[2]), .B(index_q[3]), .C(index_q[1]), 
         .D(index_q[4]), .Z(n29573)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B (C)))) */ ;
    defparam i25816_then_4_lut.init = 16'h0fe1;
    LUT4 i23949_3_lut (.A(n24007), .B(n24008), .C(index_i[4]), .Z(n24009)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23949_3_lut.init = 16'hcaca;
    PFUMX mux_206_Mux_1_i636 (.BLUT(n620_adj_3116), .ALUT(n635_adj_3350), 
          .C0(index_i[4]), .Z(n636_adj_3293)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    PFUMX i20855 (.BLUT(n23335), .ALUT(n23336), .C0(index_q[5]), .Z(n23337));
    LUT4 i21523_3_lut (.A(n29433), .B(n32028), .C(index_i[3]), .Z(n24005)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21523_3_lut.init = 16'hcaca;
    LUT4 i23951_3_lut (.A(n24004), .B(n24005), .C(index_i[4]), .Z(n24006)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23951_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_1_i349_3_lut (.A(n506_adj_3346), .B(n348_adj_3242), 
         .C(index_q[4]), .Z(n349_adj_3327)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_1_i349_3_lut.init = 16'hcaca;
    PFUMX i22021 (.BLUT(n924_adj_3336), .ALUT(n23427), .C0(index_q[5]), 
          .Z(n24522));
    PFUMX i22022 (.BLUT(n987_adj_3351), .ALUT(n23430), .C0(index_q[5]), 
          .Z(n24523));
    LUT4 i23767_3_lut (.A(n23389), .B(n23390), .C(index_q[4]), .Z(n23391)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23767_3_lut.init = 16'hcaca;
    LUT4 index_q_0__bdd_4_lut_27096 (.A(index_q[0]), .B(index_q[1]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n29486)) /* synthesis lut_function=(A (B (D)+!B !((D)+!C))+!A !(B (C+!(D))+!B (D))) */ ;
    defparam index_q_0__bdd_4_lut_27096.init = 16'h8c31;
    PFUMX i20858 (.BLUT(n23338), .ALUT(n23339), .C0(index_q[5]), .Z(n23340));
    LUT4 i23954_3_lut (.A(n24001), .B(n24002), .C(index_i[4]), .Z(n24003)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23954_3_lut.init = 16'hcaca;
    LUT4 i25816_else_4_lut (.A(index_q[2]), .B(index_q[3]), .C(index_q[1]), 
         .D(index_q[4]), .Z(n29572)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A (B (D)+!B !(C (D)+!C !(D))))) */ ;
    defparam i25816_else_4_lut.init = 16'h38c7;
    LUT4 i21516_3_lut (.A(n29432), .B(n29424), .C(index_i[3]), .Z(n23998)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21516_3_lut.init = 16'hcaca;
    PFUMX i20861 (.BLUT(n23341), .ALUT(n23342), .C0(index_q[5]), .Z(n23343));
    PFUMX i20864 (.BLUT(n23344), .ALUT(n23345), .C0(index_q[5]), .Z(n23346));
    PFUMX i20867 (.BLUT(n23347), .ALUT(n23348), .C0(index_q[5]), .Z(n23349));
    PFUMX i11093 (.BLUT(n13553), .ALUT(n13554), .C0(n24093), .Z(n13389));
    PFUMX mux_207_Mux_1_i891 (.BLUT(n882), .ALUT(n890_adj_3352), .C0(n29476), 
          .Z(n891_adj_3353)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 i22381_3_lut (.A(n476), .B(n507_adj_3097), .C(index_q[5]), .Z(n24882)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22381_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_3_i94_3_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[4]), .D(n93_adj_3158), .Z(n94_adj_3354)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_3_i94_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_206_Mux_5_i700_3_lut (.A(n460_adj_3355), .B(n29437), .C(index_i[4]), 
         .Z(n700)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_5_i700_3_lut.init = 16'hcaca;
    PFUMX i20870 (.BLUT(n23350), .ALUT(n23351), .C0(index_q[5]), .Z(n23352));
    LUT4 mux_207_Mux_4_i286_3_lut (.A(n270_adj_3356), .B(n15_adj_3357), 
         .C(index_q[4]), .Z(n286_adj_3324)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_4_i286_3_lut.init = 16'hcaca;
    PFUMX i20873 (.BLUT(n23353), .ALUT(n23354), .C0(index_q[5]), .Z(n23355));
    LUT4 i21510_3_lut (.A(n325_adj_2972), .B(n29424), .C(index_i[3]), 
         .Z(n23992)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21510_3_lut.init = 16'hcaca;
    PFUMX i20693 (.BLUT(n23173), .ALUT(n23174), .C0(index_q[4]), .Z(n23175));
    LUT4 i21508_3_lut (.A(n29447), .B(n32020), .C(index_i[3]), .Z(n23990)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21508_3_lut.init = 16'hcaca;
    LUT4 i21507_3_lut (.A(n29446), .B(n32021), .C(index_i[3]), .Z(n23989)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21507_3_lut.init = 16'hcaca;
    LUT4 i20887_3_lut (.A(n404), .B(n29355), .C(index_q[3]), .Z(n23369)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20887_3_lut.init = 16'hcaca;
    PFUMX i26895 (.BLUT(n28839), .ALUT(n29422), .C0(index_i[4]), .Z(n28840));
    LUT4 mux_207_Mux_3_i747_3_lut (.A(n29389), .B(n404), .C(index_q[3]), 
         .Z(n747_adj_3317)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_3_i747_3_lut.init = 16'hcaca;
    LUT4 i24064_3_lut (.A(n29511), .B(n29514), .C(index_q[5]), .Z(n23325)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24064_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_0_i971_3_lut (.A(n29387), .B(n29471), .C(index_q[3]), 
         .Z(n971_adj_3155)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_0_i971_3_lut.init = 16'hcaca;
    LUT4 i20838_3_lut (.A(n301_adj_3071), .B(n93_adj_3262), .C(index_q[4]), 
         .Z(n23320)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20838_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_0_i396_3_lut_4_lut_3_lut_rep_728 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29388)) /* synthesis lut_function=(A ((C)+!B)+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_0_i396_3_lut_4_lut_3_lut_rep_728.init = 16'hb6b6;
    LUT4 i14216_3_lut_rep_713 (.A(index_q[2]), .B(index_q[1]), .C(index_q[0]), 
         .Z(n29373)) /* synthesis lut_function=(A (B)+!A (B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i14216_3_lut_rep_713.init = 16'hdcdc;
    LUT4 mux_207_Mux_6_i442_rep_729 (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .Z(n29389)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_6_i442_rep_729.init = 16'h6464;
    LUT4 mux_207_Mux_1_i94_3_lut (.A(index_q[0]), .B(n93_adj_3358), .C(index_q[4]), 
         .Z(n94_adj_3314)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_1_i94_3_lut.init = 16'hcaca;
    PFUMX i20903 (.BLUT(n23383), .ALUT(n23384), .C0(index_q[4]), .Z(n23385));
    PFUMX mux_206_Mux_2_i891 (.BLUT(n875), .ALUT(n890), .C0(index_i[4]), 
          .Z(n891_adj_3177)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 mux_207_Mux_2_i763_4_lut_4_lut (.A(index_q[0]), .B(n13436), .C(index_q[4]), 
         .D(n157), .Z(n763_adj_3359)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_2_i763_4_lut_4_lut.init = 16'hdfd0;
    PFUMX mux_206_Mux_2_i860 (.BLUT(n844), .ALUT(n859_adj_3360), .C0(index_i[4]), 
          .Z(n860_adj_3176)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 mux_207_Mux_4_i94_3_lut (.A(n61_adj_3361), .B(n29283), .C(index_q[4]), 
         .Z(n94_adj_3312)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_4_i94_3_lut.init = 16'hcaca;
    LUT4 i23628_3_lut (.A(n23362), .B(n23363), .C(index_q[4]), .Z(n23364)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23628_3_lut.init = 16'hcaca;
    LUT4 i20878_3_lut (.A(n29355), .B(n29463), .C(index_q[3]), .Z(n23360)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20878_3_lut.init = 16'hcaca;
    PFUMX i22509 (.BLUT(n142_adj_3362), .ALUT(n157_adj_3363), .C0(index_i[4]), 
          .Z(n25010));
    LUT4 i20835_3_lut (.A(n15), .B(n526_adj_3260), .C(index_q[4]), .Z(n23317)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20835_3_lut.init = 16'hcaca;
    PFUMX i27074 (.BLUT(n29482), .ALUT(n29483), .C0(index_i[1]), .Z(n29484));
    LUT4 mux_207_Mux_0_i134_3_lut_4_lut_3_lut_rep_730 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29390)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_0_i134_3_lut_4_lut_3_lut_rep_730.init = 16'h6969;
    PFUMX i26856 (.BLUT(n28802), .ALUT(n29317), .C0(index_q[4]), .Z(n28803));
    LUT4 mux_207_Mux_0_i123_3_lut_3_lut_rep_731 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29391)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_0_i123_3_lut_3_lut_rep_731.init = 16'h6c6c;
    LUT4 i23625_3_lut (.A(n23359), .B(n23360), .C(index_q[4]), .Z(n23361)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23625_3_lut.init = 16'hcaca;
    PFUMX i20906 (.BLUT(n23386), .ALUT(n23387), .C0(index_q[4]), .Z(n23388));
    PFUMX i22510 (.BLUT(n173_adj_3115), .ALUT(n188_adj_3313), .C0(index_i[4]), 
          .Z(n25011));
    LUT4 mux_207_Mux_2_i908_3_lut_4_lut_4_lut (.A(index_q[2]), .B(index_q[1]), 
         .C(index_q[0]), .D(index_q[3]), .Z(n908_adj_3309)) /* synthesis lut_function=(!(A (B)+!A !(B (D)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_2_i908_3_lut_4_lut_4_lut.init = 16'h6623;
    LUT4 i23623_3_lut (.A(n23356), .B(n23357), .C(index_q[4]), .Z(n23358)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23623_3_lut.init = 16'hcaca;
    LUT4 i23725_3_lut (.A(n620_adj_3261), .B(n15110), .C(index_q[4]), 
         .Z(n23354)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23725_3_lut.init = 16'hcaca;
    LUT4 i22596_3_lut_3_lut (.A(n29385), .B(index_i[3]), .C(n32039), .Z(n25097)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam i22596_3_lut_3_lut.init = 16'h7474;
    LUT4 mux_207_Mux_5_i573_3_lut_3_lut (.A(index_q[0]), .B(index_q[4]), 
         .C(n572), .Z(n573_adj_3265)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_5_i573_3_lut_3_lut.init = 16'hd1d1;
    PFUMX i22478 (.BLUT(n142_adj_3364), .ALUT(n157_adj_3365), .C0(index_q[4]), 
          .Z(n24979));
    LUT4 mux_206_Mux_1_i924_3_lut (.A(n316_adj_3181), .B(n29419), .C(index_i[4]), 
         .Z(n924_adj_3301)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_1_i924_3_lut.init = 16'hcaca;
    LUT4 n811_bdd_4_lut_then_4_lut (.A(index_i[3]), .B(index_i[4]), .C(index_i[0]), 
         .D(index_i[2]), .Z(n29576)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B+(C (D)+!C !(D)))) */ ;
    defparam n811_bdd_4_lut_then_4_lut.init = 16'hf44f;
    LUT4 mux_207_Mux_4_i221_3_lut_3_lut (.A(index_q[0]), .B(index_q[4]), 
         .C(n205), .Z(n221_adj_3320)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_4_i221_3_lut_3_lut.init = 16'h7474;
    LUT4 mux_206_Mux_7_i892_3_lut (.A(n62_adj_3366), .B(n891_adj_3367), 
         .C(index_i[5]), .Z(n892_adj_3368)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_7_i892_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_5_i891_3_lut (.A(n875_adj_3369), .B(n379_adj_3063), 
         .C(index_q[4]), .Z(n891_adj_3296)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_5_i891_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_5_i860_3_lut (.A(n15_adj_3113), .B(n859_adj_3370), 
         .C(index_q[4]), .Z(n860_adj_3295)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_5_i860_3_lut.init = 16'hcaca;
    LUT4 i20677_3_lut (.A(n29461), .B(n141), .C(index_q[3]), .Z(n23159)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20677_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_2_i507_3_lut_3_lut (.A(index_q[0]), .B(index_q[4]), 
         .C(n491_adj_3371), .Z(n507_adj_3372)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_2_i507_3_lut_3_lut.init = 16'h7474;
    LUT4 i20928_3_lut_3_lut_4_lut_4_lut (.A(index_q[2]), .B(index_q[1]), 
         .C(index_q[0]), .D(index_q[3]), .Z(n23410)) /* synthesis lut_function=(!(A (B (D)+!B !(D))+!A (B+(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i20928_3_lut_3_lut_4_lut_4_lut.init = 16'h2388;
    LUT4 i20676_3_lut (.A(n29315), .B(n29460), .C(index_q[3]), .Z(n23158)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20676_3_lut.init = 16'hcaca;
    LUT4 i23798_3_lut (.A(n23239), .B(n23240), .C(index_i[4]), .Z(n23241)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23798_3_lut.init = 16'hcaca;
    LUT4 i21495_3_lut_4_lut_4_lut (.A(index_q[0]), .B(n29393), .C(index_q[3]), 
         .D(n29370), .Z(n23977)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i21495_3_lut_4_lut_4_lut.init = 16'hc5c0;
    LUT4 i21427_3_lut (.A(n747), .B(n908), .C(index_i[4]), .Z(n23909)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21427_3_lut.init = 16'hcaca;
    LUT4 i21426_3_lut (.A(n716), .B(n16744), .C(index_i[4]), .Z(n23908)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21426_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_6_i653_3_lut (.A(n29464), .B(n85), .C(index_q[3]), 
         .Z(n653_adj_3078)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_6_i653_3_lut.init = 16'hcaca;
    LUT4 i21424_3_lut (.A(n93_adj_3373), .B(n699), .C(index_i[4]), .Z(n23906)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21424_3_lut.init = 16'hcaca;
    LUT4 i21423_3_lut (.A(n653_adj_3012), .B(n29058), .C(index_i[4]), 
         .Z(n23905)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21423_3_lut.init = 16'hcaca;
    LUT4 i20674_3_lut (.A(n29461), .B(n29181), .C(index_q[3]), .Z(n23156)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20674_3_lut.init = 16'hcaca;
    LUT4 i20673_3_lut (.A(n29472), .B(n141), .C(index_q[3]), .Z(n23155)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20673_3_lut.init = 16'hcaca;
    LUT4 i11148_3_lut_4_lut_4_lut (.A(index_q[0]), .B(n588), .C(index_q[4]), 
         .D(n29370), .Z(n13444)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B ((D)+!C)+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i11148_3_lut_4_lut_4_lut.init = 16'h5c0c;
    LUT4 mux_207_Mux_7_i173_3_lut (.A(n29315), .B(n29181), .C(index_q[3]), 
         .Z(n173_adj_3374)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_7_i173_3_lut.init = 16'hcaca;
    PFUMX i22343 (.BLUT(n31_adj_3308), .ALUT(n23952), .C0(index_q[5]), 
          .Z(n24844));
    LUT4 mux_207_Mux_2_i859_3_lut_4_lut_4_lut (.A(index_q[0]), .B(n29357), 
         .C(index_q[3]), .D(n29370), .Z(n859_adj_3290)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B ((D)+!C)+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_2_i859_3_lut_4_lut_4_lut.init = 16'h5c0c;
    LUT4 i23806_3_lut (.A(n23080), .B(n23081), .C(index_q[4]), .Z(n23082)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23806_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_4_i15_3_lut (.A(n32031), .B(n588), .C(index_q[3]), 
         .Z(n15_adj_3357)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_4_i15_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_4_i61_3_lut (.A(n29395), .B(n32035), .C(index_q[3]), 
         .Z(n61_adj_3361)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_4_i61_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_1_i890_4_lut_4_lut_4_lut_4_lut (.A(index_q[4]), .B(index_q[0]), 
         .C(n29181), .D(index_q[3]), .Z(n890_adj_3352)) /* synthesis lut_function=(!(A (B)+!A !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam mux_207_Mux_1_i890_4_lut_4_lut_4_lut_4_lut.init = 16'h7277;
    PFUMX i22515 (.BLUT(n333_adj_3375), .ALUT(n348_adj_2975), .C0(index_i[4]), 
          .Z(n25016));
    LUT4 mux_207_Mux_0_i698_3_lut_rep_801 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29461)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B (C)+!B !(C)))) */ ;
    defparam mux_207_Mux_0_i698_3_lut_rep_801.init = 16'h1c1c;
    LUT4 mux_207_Mux_5_i636_4_lut (.A(n157_adj_3376), .B(n29112), .C(index_q[4]), 
         .D(index_q[3]), .Z(n636_adj_3277)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_5_i636_4_lut.init = 16'h3aca;
    LUT4 mux_207_Mux_3_i444_3_lut_4_lut (.A(index_q[0]), .B(index_q[3]), 
         .C(n29367), .D(index_q[4]), .Z(n444_adj_3377)) /* synthesis lut_function=(!(A (B (D)+!B (C (D)))+!A !(B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_3_i444_3_lut_4_lut.init = 16'h46aa;
    PFUMX i22516 (.BLUT(n364), .ALUT(n379), .C0(index_i[4]), .Z(n25017));
    LUT4 i21505_3_lut (.A(n32024), .B(n32021), .C(index_i[3]), .Z(n23987)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21505_3_lut.init = 16'hcaca;
    PFUMX mux_206_Mux_1_i891 (.BLUT(n882_adj_3378), .ALUT(n890_adj_3379), 
          .C0(n29311), .Z(n891_adj_3380)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 mux_207_Mux_4_i252_4_lut_4_lut (.A(index_q[0]), .B(index_q[3]), 
         .C(n29370), .D(index_q[4]), .Z(n252_adj_3321)) /* synthesis lut_function=(!(A (B (D)+!B !(D))+!A !(B ((D)+!C)+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_4_i252_4_lut_4_lut.init = 16'h669d;
    LUT4 i24500_2_lut_rep_625 (.A(index_q[1]), .B(index_q[2]), .Z(n29285)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i24500_2_lut_rep_625.init = 16'h9999;
    PFUMX i22444 (.BLUT(n94_adj_3354), .ALUT(n125_adj_3303), .C0(index_q[5]), 
          .Z(n24945));
    LUT4 mux_207_Mux_0_i93_3_lut_3_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .Z(n93_adj_3190)) /* synthesis lut_function=(A (B)+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_0_i93_3_lut_3_lut.init = 16'h9c9c;
    PFUMX i22517 (.BLUT(n397_adj_3304), .ALUT(n412), .C0(index_i[4]), 
          .Z(n25018));
    LUT4 mux_206_Mux_1_i349_3_lut (.A(n541_adj_3381), .B(n348_adj_2944), 
         .C(index_i[4]), .Z(n349_adj_3275)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_1_i349_3_lut.init = 16'hcaca;
    PFUMX i22518 (.BLUT(n428_adj_2964), .ALUT(n443), .C0(index_i[4]), 
          .Z(n25019));
    PFUMX i22445 (.BLUT(n158_adj_3302), .ALUT(n189_adj_3154), .C0(index_q[5]), 
          .Z(n24946));
    LUT4 n262_bdd_2_lut_26743_3_lut (.A(index_q[1]), .B(index_q[2]), .C(index_q[3]), 
         .Z(n28675)) /* synthesis lut_function=(A (B+(C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam n262_bdd_2_lut_26743_3_lut.init = 16'hf9f9;
    LUT4 i21417_3_lut (.A(n526_adj_3382), .B(n15_adj_3231), .C(index_i[4]), 
         .Z(n23899)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21417_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_5_i397_3_lut (.A(n29353), .B(n332), .C(index_q[3]), 
         .Z(n397_adj_3383)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_5_i397_3_lut.init = 16'hcaca;
    PFUMX i22446 (.BLUT(n221_adj_3170), .ALUT(n252_adj_3141), .C0(index_q[5]), 
          .Z(n24947));
    LUT4 mux_207_Mux_5_i506_3_lut (.A(n29336), .B(n32031), .C(index_q[3]), 
         .Z(n506_adj_3338)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_5_i506_3_lut.init = 16'hcaca;
    PFUMX i22519 (.BLUT(n460_adj_2956), .ALUT(n475), .C0(index_i[4]), 
          .Z(n25020));
    LUT4 i21414_3_lut (.A(n397_adj_3384), .B(n475_adj_3011), .C(index_i[4]), 
         .Z(n23896)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21414_3_lut.init = 16'hcaca;
    LUT4 i21412_3_lut (.A(n348_adj_3385), .B(n443_adj_3173), .C(index_i[4]), 
         .Z(n23894)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21412_3_lut.init = 16'hcaca;
    LUT4 n811_bdd_4_lut_else_4_lut (.A(index_i[3]), .B(index_i[4]), .C(index_i[0]), 
         .D(index_i[2]), .Z(n29575)) /* synthesis lut_function=(!(A (B (D)+!B ((D)+!C))+!A !(B+!((D)+!C)))) */ ;
    defparam n811_bdd_4_lut_else_4_lut.init = 16'h44fc;
    PFUMX i22447 (.BLUT(n286_adj_3300), .ALUT(n23190), .C0(index_q[5]), 
          .Z(n24948));
    LUT4 i21411_3_lut (.A(n397_adj_3384), .B(n731_adj_3186), .C(index_i[4]), 
         .Z(n23893)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21411_3_lut.init = 16'hcaca;
    LUT4 i20599_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n23081)) /* synthesis lut_function=(A (B (C)+!B !(C (D)+!C !(D)))+!A (B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i20599_3_lut_4_lut_4_lut.init = 16'hd6a5;
    PFUMX i22520 (.BLUT(n491_adj_3386), .ALUT(n12581), .C0(index_i[4]), 
          .Z(n25021));
    PFUMX i22448 (.BLUT(n349_adj_3387), .ALUT(n23949), .C0(index_q[5]), 
          .Z(n24949));
    LUT4 mux_207_Mux_2_i62_3_lut_3_lut (.A(index_q[1]), .B(index_q[4]), 
         .C(n526_adj_2957), .Z(n62)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_2_i62_3_lut_3_lut.init = 16'h7474;
    LUT4 mux_207_Mux_10_i252_3_lut_4_lut_4_lut (.A(n29204), .B(index_q[3]), 
         .C(index_q[4]), .D(n29168), .Z(n252_adj_3233)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B (C (D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_10_i252_3_lut_4_lut_4_lut.init = 16'h3efe;
    LUT4 mux_207_Mux_6_i636_4_lut_4_lut (.A(index_q[1]), .B(index_q[4]), 
         .C(n635_adj_3388), .D(n16249), .Z(n636_adj_3389)) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_6_i636_4_lut_4_lut.init = 16'hf3d1;
    LUT4 mux_206_Mux_7_i348_3_lut (.A(n32018), .B(n32019), .C(index_i[3]), 
         .Z(n348_adj_3385)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_7_i348_3_lut.init = 16'hcaca;
    LUT4 mux_206_Mux_7_i397_3_lut (.A(n32018), .B(n29385), .C(index_i[3]), 
         .Z(n397_adj_3384)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_7_i397_3_lut.init = 16'hcaca;
    LUT4 mux_206_Mux_6_i731_3_lut (.A(n29409), .B(n29406), .C(index_i[3]), 
         .Z(n731_adj_3186)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_6_i731_3_lut.init = 16'hcaca;
    LUT4 i23825_3_lut (.A(n19975), .B(n19976), .C(index_q[4]), .Z(n19977)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23825_3_lut.init = 16'hcaca;
    LUT4 i13839_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[4]), 
         .C(n29326), .D(index_q[0]), .Z(n16248)) /* synthesis lut_function=(!(A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i13839_3_lut_4_lut_4_lut_4_lut.init = 16'h55d5;
    LUT4 mux_207_Mux_3_i349_3_lut_3_lut (.A(index_q[1]), .B(index_q[4]), 
         .C(n348_adj_3390), .Z(n349_adj_3387)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_3_i349_3_lut_3_lut.init = 16'hd1d1;
    PFUMX i22449 (.BLUT(n413_adj_3299), .ALUT(n444_adj_3377), .C0(index_q[5]), 
          .Z(n24950));
    PFUMX i20915 (.BLUT(n23395), .ALUT(n23396), .C0(index_q[4]), .Z(n23397));
    LUT4 mux_207_Mux_6_i475_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n475_adj_3165)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A !(B (C+(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_6_i475_3_lut_4_lut_4_lut.init = 16'h9936;
    PFUMX i22450 (.BLUT(n476_adj_3297), .ALUT(n507), .C0(index_q[5]), 
          .Z(n24951));
    PFUMX i22479 (.BLUT(n173_adj_2942), .ALUT(n188_adj_3294), .C0(index_q[4]), 
          .Z(n24980));
    PFUMX i22451 (.BLUT(n23958), .ALUT(n573_adj_3021), .C0(index_q[5]), 
          .Z(n24952));
    LUT4 i21501_3_lut (.A(n29432), .B(n32021), .C(index_i[3]), .Z(n23983)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21501_3_lut.init = 16'hcaca;
    LUT4 i23827_3_lut (.A(n23212), .B(n23213), .C(index_i[4]), .Z(n23214)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23827_3_lut.init = 16'hcaca;
    PFUMX i20918 (.BLUT(n23398), .ALUT(n23399), .C0(index_q[4]), .Z(n23400));
    L6MUX21 i26741 (.D0(n28679), .D1(n28677), .SD(index_q[5]), .Z(n28680));
    LUT4 i21496_3_lut (.A(n325), .B(n32036), .C(index_q[3]), .Z(n23978)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21496_3_lut.init = 16'hcaca;
    LUT4 i23674_3_lut (.A(n23977), .B(n23978), .C(index_q[4]), .Z(n23979)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23674_3_lut.init = 16'hcaca;
    PFUMX i26739 (.BLUT(n572), .ALUT(n28678), .C0(index_q[4]), .Z(n28679));
    LUT4 i21400_3_lut (.A(n491_adj_3391), .B(n541_adj_3381), .C(index_i[4]), 
         .Z(n23882)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21400_3_lut.init = 16'hcaca;
    LUT4 i21493_3_lut (.A(n29427), .B(n32039), .C(index_i[3]), .Z(n23975)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21493_3_lut.init = 16'hcaca;
    LUT4 n23615_bdd_3_lut (.A(n29443), .B(n29409), .C(index_i[3]), .Z(n26898)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n23615_bdd_3_lut.init = 16'hcaca;
    PFUMX i26736 (.BLUT(n28676), .ALUT(n28675), .C0(index_q[4]), .Z(n28677));
    LUT4 i21399_3_lut (.A(n557), .B(n475_adj_3212), .C(index_i[4]), .Z(n23881)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21399_3_lut.init = 16'hcaca;
    LUT4 i23976_3_lut (.A(n23974), .B(n23975), .C(index_i[4]), .Z(n23976)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23976_3_lut.init = 16'hcaca;
    LUT4 i21490_3_lut (.A(n29353), .B(n29388), .C(index_q[3]), .Z(n23972)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21490_3_lut.init = 16'hcaca;
    LUT4 i21489_3_lut (.A(n32036), .B(n29387), .C(index_q[3]), .Z(n23971)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21489_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_5_i507_3_lut (.A(n491_adj_3178), .B(n506_adj_3338), 
         .C(index_q[4]), .Z(n507_adj_3254)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_5_i507_3_lut.init = 16'hcaca;
    LUT4 i20581_3_lut (.A(n900), .B(n325_adj_2972), .C(index_i[3]), .Z(n23063)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20581_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_5_i476_3_lut (.A(n460_adj_3392), .B(n475_adj_3393), 
         .C(index_q[4]), .Z(n476_adj_3253)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_5_i476_3_lut.init = 16'hcaca;
    LUT4 i21487_3_lut (.A(n29355), .B(n29387), .C(index_q[3]), .Z(n23969)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21487_3_lut.init = 16'hcaca;
    PFUMX i22452 (.BLUT(n13432), .ALUT(n23961), .C0(index_q[5]), .Z(n24953));
    LUT4 mux_207_Mux_5_i859_3_lut (.A(n141), .B(n29315), .C(index_q[3]), 
         .Z(n859_adj_3370)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_5_i859_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_5_i875_3_lut (.A(n29181), .B(n29461), .C(index_q[3]), 
         .Z(n875_adj_3369)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_5_i875_3_lut.init = 16'hcaca;
    PFUMX i27071 (.BLUT(n29478), .ALUT(n29479), .C0(index_q[0]), .Z(n29480));
    LUT4 i23730_3_lut (.A(n491_adj_3243), .B(n506_adj_3394), .C(index_q[4]), 
         .Z(n23348)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23730_3_lut.init = 16'hcaca;
    LUT4 mux_206_Mux_1_i94_3_lut (.A(index_i[0]), .B(n93_adj_3395), .C(index_i[4]), 
         .Z(n94_adj_3245)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_1_i94_3_lut.init = 16'hcaca;
    L6MUX21 i26720 (.D0(n28663), .D1(n28660), .SD(index_q[5]), .Z(n28664));
    LUT4 i21483_3_lut (.A(n29389), .B(n29387), .C(index_q[3]), .Z(n23965)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21483_3_lut.init = 16'hcaca;
    LUT4 i21397_3_lut (.A(n251_adj_2955), .B(n443_adj_2962), .C(index_i[4]), 
         .Z(n23879)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21397_3_lut.init = 16'hcaca;
    LUT4 i21396_3_lut (.A(n557), .B(n16744), .C(index_i[4]), .Z(n23878)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;
    defparam i21396_3_lut.init = 16'h3a3a;
    LUT4 mux_207_Mux_5_i700_3_lut (.A(n460_adj_3392), .B(n29390), .C(index_q[4]), 
         .Z(n700_adj_3283)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_5_i700_3_lut.init = 16'hcaca;
    PFUMX i22453 (.BLUT(n669_adj_3280), .ALUT(n700_adj_3396), .C0(index_q[5]), 
          .Z(n24954));
    LUT4 mux_207_Mux_5_i413_3_lut (.A(n397_adj_3383), .B(n251_adj_3070), 
         .C(index_q[4]), .Z(n413_adj_3237)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_5_i413_3_lut.init = 16'hcaca;
    LUT4 i21481_3_lut (.A(n29352), .B(n29388), .C(index_q[3]), .Z(n23963)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21481_3_lut.init = 16'hcaca;
    PFUMX i26718 (.BLUT(n28662), .ALUT(n28661), .C0(index_q[4]), .Z(n28663));
    LUT4 i22246_3_lut_4_lut (.A(n29204), .B(index_q[3]), .C(index_q[4]), 
         .D(n29132), .Z(n24747)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i22246_3_lut_4_lut.init = 16'hfe0e;
    LUT4 mux_206_Mux_1_i986_3_lut (.A(n32018), .B(n29436), .C(index_i[3]), 
         .Z(n986_adj_3397)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_1_i986_3_lut.init = 16'hcaca;
    PFUMX i26715 (.BLUT(n29054), .ALUT(n28659), .C0(index_q[4]), .Z(n28660));
    L6MUX21 i22454 (.D0(n23964), .D1(n763_adj_3318), .SD(index_q[5]), 
            .Z(n24955));
    LUT4 i14198_2_lut_rep_641 (.A(index_i[2]), .B(index_i[0]), .Z(n29301)) /* synthesis lut_function=(A (B)) */ ;
    defparam i14198_2_lut_rep_641.init = 16'h8888;
    PFUMX i20921 (.BLUT(n23401), .ALUT(n23402), .C0(index_q[4]), .Z(n23403));
    LUT4 mux_206_Mux_4_i828_3_lut_4_lut (.A(index_i[4]), .B(index_i[3]), 
         .C(n812_adj_2950), .D(n29404), .Z(n828_adj_3069)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_4_i828_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_206_Mux_5_i797_3_lut_4_lut (.A(index_i[4]), .B(index_i[3]), 
         .C(n29484), .D(n29432), .Z(n797_adj_3018)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_5_i797_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i22456 (.BLUT(n860_adj_3098), .ALUT(n891_adj_3274), .C0(index_q[5]), 
          .Z(n24957));
    PFUMX i20924 (.BLUT(n23404), .ALUT(n23405), .C0(index_q[4]), .Z(n23406));
    LUT4 mux_206_Mux_1_i763_3_lut_4_lut (.A(index_i[4]), .B(index_i[3]), 
         .C(n29577), .D(n29432), .Z(n763_adj_3398)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_1_i763_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i14407_1_lut_2_lut_3_lut_4_lut (.A(n29204), .B(index_q[3]), .C(index_q[5]), 
         .D(index_q[4]), .Z(n381_adj_2939)) /* synthesis lut_function=(!(A (C+(D))+!A (B (C+(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i14407_1_lut_2_lut_3_lut_4_lut.init = 16'h010f;
    PFUMX i22457 (.BLUT(n924_adj_3272), .ALUT(n23979), .C0(index_q[5]), 
          .Z(n24958));
    PFUMX mux_206_Mux_3_i763 (.BLUT(n747_adj_3271), .ALUT(n762), .C0(index_i[4]), 
          .Z(n763_adj_3119)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 i21390_3_lut (.A(n205_adj_3399), .B(n188), .C(index_i[4]), .Z(n23872)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21390_3_lut.init = 16'hcaca;
    LUT4 i24234_3_lut (.A(n23872), .B(n29501), .C(index_i[5]), .Z(n23874)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24234_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_4_i270_3_lut (.A(n32034), .B(n29336), .C(index_q[3]), 
         .Z(n270_adj_3356)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_4_i270_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_4_i348_3_lut (.A(n29333), .B(n29335), .C(index_q[3]), 
         .Z(n348_adj_3400)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_4_i348_3_lut.init = 16'hcaca;
    LUT4 i21387_3_lut (.A(n875_adj_3033), .B(n93_adj_3373), .C(index_i[4]), 
         .Z(n23869)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21387_3_lut.init = 16'hcaca;
    LUT4 index_i_1__bdd_4_lut_27597 (.A(index_i[1]), .B(index_i[0]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n29578)) /* synthesis lut_function=(!(A (B (D)+!B (C+!(D)))+!A !(B (C (D)+!C !(D))+!B !((D)+!C)))) */ ;
    defparam index_i_1__bdd_4_lut_27597.init = 16'h429c;
    LUT4 i20881_3_lut_4_lut_4_lut (.A(index_q[2]), .B(n141), .C(index_q[3]), 
         .D(n29459), .Z(n23363)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i20881_3_lut_4_lut_4_lut.init = 16'hc5c0;
    LUT4 n627_bdd_3_lut_26717_4_lut_4_lut (.A(index_q[2]), .B(n85), .C(index_q[3]), 
         .D(n29459), .Z(n28661)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B ((D)+!C)+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam n627_bdd_3_lut_26717_4_lut_4_lut.init = 16'h5c0c;
    LUT4 i23684_3_lut (.A(n23959), .B(n23960), .C(index_q[4]), .Z(n23961)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23684_3_lut.init = 16'hcaca;
    PFUMX i22458 (.BLUT(n23982), .ALUT(n1018), .C0(index_q[5]), .Z(n24959));
    LUT4 mux_207_Mux_4_i684_3_lut (.A(n85), .B(n108), .C(index_q[3]), 
         .Z(n684_adj_3348)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_4_i684_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_7_i506_3_lut_4_lut_4_lut (.A(index_q[2]), .B(n29461), 
         .C(index_q[3]), .D(n29459), .Z(n506_adj_3394)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B ((D)+!C)+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_7_i506_3_lut_4_lut_4_lut.init = 16'h5c0c;
    LUT4 mux_207_Mux_4_i491_3_lut_4_lut_4_lut (.A(index_q[2]), .B(n29461), 
         .C(index_q[3]), .D(n29465), .Z(n491_adj_3096)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_4_i491_3_lut_4_lut_4_lut.init = 16'hfc5c;
    LUT4 i21384_3_lut (.A(n188), .B(n526), .C(index_i[4]), .Z(n23866)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21384_3_lut.init = 16'hcaca;
    LUT4 i23517_3_lut (.A(n23953), .B(n23954), .C(index_i[4]), .Z(n23955)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23517_3_lut.init = 16'hcaca;
    LUT4 i21469_3_lut (.A(n29463), .B(n32055), .C(index_q[3]), .Z(n23951)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21469_3_lut.init = 16'hcaca;
    LUT4 i23704_3_lut (.A(n23950), .B(n23951), .C(index_q[4]), .Z(n23952)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23704_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_5_i924_4_lut_3_lut (.A(index_q[2]), .B(n16637), .C(index_q[4]), 
         .Z(n924_adj_3206)) /* synthesis lut_function=(!(A (B+(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_5_i924_4_lut_3_lut.init = 16'h5656;
    LUT4 i21466_3_lut (.A(n32029), .B(n29336), .C(index_q[3]), .Z(n23948)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21466_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_1_i986_3_lut (.A(n29461), .B(n32033), .C(index_q[3]), 
         .Z(n986_adj_3401)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_1_i986_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_4_i62_4_lut (.A(n29368), .B(n61_adj_3361), .C(index_q[4]), 
         .D(index_q[3]), .Z(n62_adj_3224)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_4_i62_4_lut.init = 16'hc5ca;
    LUT4 i12677_2_lut_rep_426_3_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n29086)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12677_2_lut_rep_426_3_lut_4_lut.init = 16'hfef0;
    LUT4 n20177_bdd_4_lut_then_4_lut (.A(index_q[3]), .B(index_q[4]), .C(index_q[0]), 
         .D(index_q[2]), .Z(n29580)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B+(C (D)+!C !(D)))) */ ;
    defparam n20177_bdd_4_lut_then_4_lut.init = 16'hf44f;
    LUT4 mux_207_Mux_4_i31_4_lut (.A(n15_adj_3357), .B(n29059), .C(index_q[4]), 
         .D(index_q[3]), .Z(n31_adj_3223)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_4_i31_4_lut.init = 16'h3aca;
    LUT4 i21465_3_lut (.A(n29387), .B(n29353), .C(index_q[3]), .Z(n23947)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21465_3_lut.init = 16'hcaca;
    LUT4 i23690_3_lut (.A(n23947), .B(n23948), .C(index_q[4]), .Z(n23949)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23690_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_6_i15_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n15_adj_3339)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C))+!A !(B (C+!(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_6_i15_3_lut_4_lut_4_lut.init = 16'h5ad6;
    LUT4 i21463_3_lut (.A(n498), .B(n29446), .C(index_i[3]), .Z(n23945)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21463_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_649 (.A(index_i[4]), .B(index_i[5]), .Z(n29309)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_2_lut_rep_649.init = 16'heeee;
    LUT4 i1_3_lut_4_lut_adj_186 (.A(index_i[4]), .B(index_i[5]), .C(index_i[3]), 
         .D(n29400), .Z(n22180)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_3_lut_4_lut_adj_186.init = 16'hfffe;
    LUT4 mux_207_Mux_10_i413_3_lut_3_lut_4_lut (.A(n29204), .B(index_q[3]), 
         .C(n29130), .D(index_q[4]), .Z(n413_adj_3402)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_10_i413_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 mux_207_Mux_7_i333_3_lut (.A(n29467), .B(n29181), .C(index_q[3]), 
         .Z(n333_adj_3330)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_7_i333_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_7_i348_3_lut (.A(n29461), .B(n29470), .C(index_q[3]), 
         .Z(n348_adj_3329)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_7_i348_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_7_i397_3_lut (.A(n29461), .B(n29467), .C(index_q[3]), 
         .Z(n397_adj_3328)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_7_i397_3_lut.init = 16'hcaca;
    LUT4 i24623_2_lut (.A(index_q[3]), .B(index_q[2]), .Z(n24093)) /* synthesis lut_function=(A+!(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i24623_2_lut.init = 16'hbbbb;
    LUT4 mux_207_Mux_4_i142_3_lut_3_lut (.A(index_q[0]), .B(index_q[2]), 
         .C(index_q[3]), .Z(n142_adj_3403)) /* synthesis lut_function=(A (B (C))+!A !(B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_4_i142_3_lut_3_lut.init = 16'h9595;
    LUT4 i17692_3_lut (.A(n20004), .B(n20005), .C(index_q[4]), .Z(n20006)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17692_3_lut.init = 16'hcaca;
    LUT4 i21459_3_lut (.A(n32028), .B(n29431), .C(index_i[3]), .Z(n23941)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21459_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_5_i125_3_lut (.A(n109), .B(n124_adj_3051), .C(index_q[4]), 
         .Z(n125_adj_3222)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_5_i125_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_1_i62_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[2]), 
         .C(index_q[4]), .D(index_q[3]), .Z(n62_adj_3404)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))+!A !(B (C)+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_1_i62_3_lut_4_lut_4_lut.init = 16'ha5a6;
    LUT4 i23790_3_lut (.A(n23941), .B(n23942), .C(index_i[4]), .Z(n23943)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23790_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_5_i94_3_lut (.A(n653_adj_3078), .B(n635_adj_3388), 
         .C(index_q[4]), .Z(n94_adj_3221)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_5_i94_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_4_i158_3_lut (.A(n142_adj_3403), .B(n157_adj_3376), 
         .C(index_q[4]), .Z(n158_adj_3219)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_4_i158_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_3_i828_3_lut_3_lut_4_lut (.A(n29204), .B(index_q[3]), 
         .C(n157_adj_3174), .D(index_q[4]), .Z(n828)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_3_i828_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 mux_207_Mux_4_i812_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[2]), 
         .C(index_q[3]), .D(index_q[4]), .Z(n812_adj_3405)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A !(B (D)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_4_i812_3_lut_3_lut_4_lut.init = 16'ha955;
    LUT4 mux_206_Mux_3_i700_3_lut_4_lut (.A(index_i[4]), .B(index_i[3]), 
         .C(n684_adj_3406), .D(n29404), .Z(n700_adj_3118)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_3_i700_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i24630_2_lut_rep_651 (.A(index_i[4]), .B(index_i[3]), .Z(n29311)) /* synthesis lut_function=((B)+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i24630_2_lut_rep_651.init = 16'hdddd;
    PFUMX i26639 (.BLUT(n28577), .ALUT(n28576), .C0(index_i[5]), .Z(n28578));
    LUT4 i22571_4_lut_4_lut (.A(index_q[4]), .B(index_q[5]), .C(n29508), 
         .D(n908_adj_3309), .Z(n25072)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam i22571_4_lut_4_lut.init = 16'hd1c0;
    LUT4 mux_206_Mux_7_i250_3_lut_4_lut_3_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[2]), .Z(n851)) /* synthesis lut_function=(A ((C)+!B)+!A (B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_7_i250_3_lut_4_lut_3_lut.init = 16'he7e7;
    LUT4 mux_206_Mux_3_i797_3_lut_4_lut (.A(index_i[4]), .B(index_i[3]), 
         .C(n796_adj_3407), .D(n29377), .Z(n797_adj_3408)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_3_i797_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_206_Mux_5_i924_4_lut_3_lut (.A(index_i[2]), .B(n16591), .C(index_i[4]), 
         .Z(n924_adj_3180)) /* synthesis lut_function=(!(A (B+(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_5_i924_4_lut_3_lut.init = 16'h5656;
    LUT4 i23782_3_lut (.A(n109_adj_2967), .B(n124_adj_3257), .C(index_q[4]), 
         .Z(n23321)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23782_3_lut.init = 16'hcaca;
    LUT4 i20737_3_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[0]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n23219)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20737_3_lut_4_lut_4_lut.init = 16'hfa1a;
    LUT4 i21456_3_lut (.A(n1001), .B(n931), .C(index_i[3]), .Z(n23938)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21456_3_lut.init = 16'hcaca;
    LUT4 i23792_3_lut (.A(n23938), .B(n23939), .C(index_i[4]), .Z(n23940)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23792_3_lut.init = 16'hcaca;
    LUT4 i21454_3_lut (.A(n498), .B(n29405), .C(index_i[3]), .Z(n23936)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21454_3_lut.init = 16'hcaca;
    LUT4 i11224_4_lut_4_lut (.A(index_i[4]), .B(n24296), .C(n13566), .D(n29377), 
         .Z(n13520)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam i11224_4_lut_4_lut.init = 16'hf4b0;
    L6MUX21 i26603 (.D0(n28538), .D1(n28536), .SD(index_i[6]), .Z(n23310));
    PFUMX i26601 (.BLUT(n28537), .ALUT(n62_adj_3366), .C0(index_i[5]), 
          .Z(n28538));
    LUT4 i21453_3_lut (.A(n29441), .B(n325_adj_2972), .C(index_i[3]), 
         .Z(n23935)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21453_3_lut.init = 16'hcaca;
    PFUMX i26599 (.BLUT(n28535), .ALUT(n28534), .C0(index_i[5]), .Z(n28536));
    LUT4 i21486_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n23968)) /* synthesis lut_function=(A (B (C (D))+!B !(C (D)))+!A !(B (D)+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i21486_3_lut_4_lut_4_lut.init = 16'h9366;
    LUT4 mux_207_Mux_3_i700_3_lut_4_lut (.A(index_q[4]), .B(index_q[3]), 
         .C(n684_adj_3409), .D(n29354), .Z(n700_adj_3396)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_3_i700_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i14226_3_lut (.A(index_q[3]), .B(index_q[1]), .C(index_q[0]), 
         .Z(n16645)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i14226_3_lut.init = 16'hc8c8;
    LUT4 mux_207_Mux_3_i348_3_lut (.A(n32033), .B(n32036), .C(index_q[3]), 
         .Z(n348_adj_3390)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_3_i348_3_lut.init = 16'hcaca;
    LUT4 i12531_2_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n844_adj_3410)) /* synthesis lut_function=(A (B+!(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i12531_2_lut_3_lut_4_lut.init = 16'h9ff9;
    LUT4 i20593_3_lut (.A(n32020), .B(n325_adj_2972), .C(index_i[3]), 
         .Z(n23075)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20593_3_lut.init = 16'hcaca;
    PFUMX i20930 (.BLUT(n23410), .ALUT(n23411), .C0(index_q[4]), .Z(n23412));
    LUT4 i11086_4_lut_4_lut (.A(index_q[4]), .B(n24311), .C(n29538), .D(n29475), 
         .Z(n13382)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam i11086_4_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_207_Mux_3_i31_3_lut (.A(n781), .B(n30_adj_3311), .C(index_q[4]), 
         .Z(n31_adj_3201)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_3_i31_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_4_i349_3_lut_4_lut (.A(index_q[0]), .B(index_q[2]), 
         .C(index_q[4]), .D(n348_adj_3400), .Z(n349_adj_3325)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_4_i349_3_lut_4_lut.init = 16'hf606;
    LUT4 i23936_3_lut (.A(n23074), .B(n23075), .C(index_i[4]), .Z(n23076)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23936_3_lut.init = 16'hcaca;
    L6MUX21 mux_207_Mux_7_i253 (.D0(n13389), .D1(n23160), .SD(index_q[5]), 
            .Z(n253)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 i21445_3_lut (.A(n29441), .B(n29405), .C(index_i[3]), .Z(n23927)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21445_3_lut.init = 16'hcaca;
    LUT4 mux_206_Mux_4_i541_3_lut_4_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n541_adj_3381)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_4_i541_3_lut_4_lut_3_lut_4_lut.init = 16'h0ef0;
    LUT4 mux_206_Mux_5_i828_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[4]), .D(n29372), .Z(n828_adj_3019)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_5_i828_4_lut_4_lut.init = 16'hc66c;
    LUT4 i21444_3_lut (.A(n325_adj_2972), .B(n204), .C(index_i[3]), .Z(n23926)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21444_3_lut.init = 16'hcaca;
    PFUMX i26573 (.BLUT(n28503), .ALUT(n28502), .C0(index_q[5]), .Z(n28504));
    LUT4 mux_206_Mux_6_i660_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n660)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_6_i660_3_lut_3_lut.init = 16'hc6c6;
    LUT4 i11063_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n812_adj_3057)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+(D)))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11063_3_lut_4_lut_4_lut.init = 16'h666c;
    LUT4 i22244_3_lut_3_lut_4_lut (.A(n29204), .B(index_q[3]), .C(n412_adj_3335), 
         .D(index_q[4]), .Z(n24745)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i22244_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 i8865_2_lut_rep_714 (.A(index_i[3]), .B(index_i[4]), .Z(n29374)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i8865_2_lut_rep_714.init = 16'heeee;
    PFUMX mux_207_Mux_7_i190 (.BLUT(n23157), .ALUT(n173_adj_3374), .C0(index_q[5]), 
          .Z(n190_adj_3411)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 n124_bdd_3_lut_4_lut (.A(n29177), .B(index_i[3]), .C(index_i[4]), 
         .D(n93_adj_3278), .Z(n28535)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n124_bdd_3_lut_4_lut.init = 16'hfe0e;
    L6MUX21 i26563 (.D0(n28492), .D1(n28490), .SD(index_q[6]), .Z(n23292));
    LUT4 i17662_3_lut_3_lut (.A(index_q[0]), .B(index_q[2]), .C(index_q[3]), 
         .Z(n19976)) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i17662_3_lut_3_lut.init = 16'h6a6a;
    PFUMX i26561 (.BLUT(n28491), .ALUT(n62_adj_3412), .C0(index_q[5]), 
          .Z(n28492));
    LUT4 mux_207_Mux_6_i573_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[4]), .D(n572_adj_3413), .Z(n573_adj_3414)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_6_i573_3_lut_4_lut.init = 16'hf909;
    LUT4 i11132_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[4]), .D(n29326), .Z(n189_adj_3220)) /* synthesis lut_function=(A (B (C (D)))+!A !(B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i11132_3_lut_4_lut_4_lut_4_lut.init = 16'h9555;
    PFUMX i26559 (.BLUT(n28489), .ALUT(n28488), .C0(index_q[5]), .Z(n28490));
    LUT4 i11043_3_lut_4_lut (.A(index_i[3]), .B(index_i[4]), .C(n29434), 
         .D(n32039), .Z(n605_adj_3415)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11043_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_206_Mux_0_i236_3_lut_3_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[3]), .Z(n236)) /* synthesis lut_function=(A (B+(C))+!A !(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i236_3_lut_3_lut.init = 16'ha9a9;
    LUT4 i23816_3_lut (.A(n620_adj_3416), .B(n16308), .C(index_i[4]), 
         .Z(n23903)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23816_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_6_i924_3_lut_4_lut (.A(index_q[2]), .B(index_q[3]), 
         .C(index_q[4]), .D(n762_adj_3316), .Z(n924_adj_3417)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_6_i924_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_206_Mux_7_i891_3_lut_4_lut (.A(n29177), .B(index_i[3]), .C(index_i[4]), 
         .D(n890_adj_3205), .Z(n891_adj_3367)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_7_i891_3_lut_4_lut.init = 16'hfe0e;
    LUT4 i23819_3_lut (.A(n491), .B(n506), .C(index_i[4]), .Z(n23897)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23819_3_lut.init = 16'hcaca;
    LUT4 n61_bdd_3_lut_25998_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n27486)) /* synthesis lut_function=(!(A (B)+!A !(B (C+(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n61_bdd_3_lut_25998_4_lut_4_lut_4_lut.init = 16'h6663;
    LUT4 mux_207_Mux_7_i892_3_lut (.A(n62_adj_3412), .B(n891_adj_3418), 
         .C(index_q[5]), .Z(n892_adj_3419)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_7_i892_3_lut.init = 16'hcaca;
    LUT4 i11057_3_lut_3_lut_4_lut (.A(index_i[3]), .B(index_i[4]), .C(n29429), 
         .D(index_i[0]), .Z(n605)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11057_3_lut_3_lut_4_lut.init = 16'h10fe;
    LUT4 i20746_3_lut (.A(n32023), .B(n29440), .C(index_i[3]), .Z(n23228)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20746_3_lut.init = 16'hcaca;
    LUT4 i14158_2_lut_rep_616 (.A(index_q[2]), .B(index_q[0]), .Z(n29276)) /* synthesis lut_function=(A (B)) */ ;
    defparam i14158_2_lut_rep_616.init = 16'h8888;
    LUT4 mux_206_Mux_5_i116_3_lut_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n645)) /* synthesis lut_function=(!(A (B)+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_5_i116_3_lut_3_lut_3_lut.init = 16'h6363;
    LUT4 i23884_3_lut (.A(n716_adj_3264), .B(n731_adj_3420), .C(index_i[4]), 
         .Z(n732_adj_3151)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23884_3_lut.init = 16'hcaca;
    PFUMX i20609 (.BLUT(n23089), .ALUT(n23090), .C0(index_q[4]), .Z(n23091));
    PFUMX mux_207_Mux_8_i764 (.BLUT(n716_adj_2946), .ALUT(n732_adj_3251), 
          .C0(n24091), .Z(n764)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 i3220_1_lut_rep_658 (.A(index_i[0]), .Z(n29318)) /* synthesis lut_function=(!(A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i3220_1_lut_rep_658.init = 16'h5555;
    LUT4 mux_206_Mux_2_i349_3_lut_3_lut (.A(index_i[0]), .B(index_i[4]), 
         .C(n348_adj_3421), .Z(n349_adj_3131)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_2_i349_3_lut_3_lut.init = 16'hd1d1;
    PFUMX i26523 (.BLUT(n28447), .ALUT(n28443), .C0(index_i[6]), .Z(n28448));
    PFUMX i27123 (.BLUT(n29557), .ALUT(n29558), .C0(index_i[8]), .Z(n29559));
    LUT4 i14150_2_lut_rep_715 (.A(index_i[2]), .B(index_i[0]), .Z(n29375)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i14150_2_lut_rep_715.init = 16'heeee;
    LUT4 i11107_3_lut_4_lut_4_lut (.A(index_i[0]), .B(n931), .C(index_i[4]), 
         .D(n29418), .Z(n13403)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B ((D)+!C)+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11107_3_lut_4_lut_4_lut.init = 16'h5c0c;
    PFUMX mux_207_Mux_8_i574 (.BLUT(n542_adj_3422), .ALUT(n13385), .C0(index_q[5]), 
          .Z(n574)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 n20177_bdd_4_lut_else_4_lut (.A(index_q[3]), .B(index_q[4]), .C(index_q[0]), 
         .D(index_q[2]), .Z(n29579)) /* synthesis lut_function=(!(A (B (D)+!B ((D)+!C))+!A !(B+!((D)+!C)))) */ ;
    defparam n20177_bdd_4_lut_else_4_lut.init = 16'h44fc;
    LUT4 mux_206_Mux_2_i507_3_lut_3_lut (.A(index_i[0]), .B(index_i[4]), 
         .C(n491_adj_3423), .Z(n507_adj_3138)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_2_i507_3_lut_3_lut.init = 16'h7474;
    PFUMX mux_206_Mux_5_i732 (.BLUT(n13357), .ALUT(n731_adj_3235), .C0(index_i[4]), 
          .Z(n732_adj_3017)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 mux_206_Mux_8_i45_3_lut_rep_720 (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[2]), .Z(n29380)) /* synthesis lut_function=(A (C)+!A !(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_8_i45_3_lut_rep_720.init = 16'ha1a1;
    LUT4 mux_206_Mux_2_i669_3_lut (.A(n653_adj_3424), .B(n475_adj_3009), 
         .C(index_i[4]), .Z(n669_adj_3147)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_2_i669_3_lut.init = 16'hcaca;
    LUT4 i14451_3_lut_4_lut (.A(n29177), .B(index_i[3]), .C(n11112), .D(index_i[6]), 
         .Z(n16882)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i14451_3_lut_4_lut.init = 16'hffe0;
    LUT4 mux_206_Mux_2_i763_4_lut_4_lut (.A(index_i[0]), .B(n13373), .C(index_i[4]), 
         .D(n157_adj_3225), .Z(n763_adj_3152)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_2_i763_4_lut_4_lut.init = 16'hdfd0;
    LUT4 mux_206_Mux_0_i684_3_lut_4_lut_4_lut (.A(index_i[0]), .B(n29439), 
         .C(index_i[3]), .D(n29418), .Z(n684_adj_3425)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B ((D)+!C)+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i684_3_lut_4_lut_4_lut.init = 16'h5c0c;
    LUT4 mux_206_Mux_4_i221_3_lut_3_lut (.A(index_i[0]), .B(index_i[4]), 
         .C(n205_adj_3426), .Z(n221_adj_3041)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_4_i221_3_lut_3_lut.init = 16'h7474;
    LUT4 mux_206_Mux_2_i605_3_lut (.A(n142_adj_3427), .B(n604_adj_3428), 
         .C(index_i[4]), .Z(n605_adj_3145)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_2_i605_3_lut.init = 16'hcaca;
    PFUMX i21860 (.BLUT(n24359), .ALUT(n24360), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_1768[5]));
    PFUMX i21922 (.BLUT(n24421), .ALUT(n24422), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_1768[3]));
    PFUMX i22006 (.BLUT(n24505), .ALUT(n24506), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_1768[1]));
    PFUMX i22373 (.BLUT(n24872), .ALUT(n24873), .C0(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_1783[5]));
    PFUMX i22037 (.BLUT(n24536), .ALUT(n24537), .C0(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_1783[1]));
    PFUMX i22473 (.BLUT(n24972), .ALUT(n24973), .C0(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_1783[3]));
    PFUMX i20729 (.BLUT(n23209), .ALUT(n23210), .C0(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_1783[11]));
    LUT4 mux_206_Mux_2_i859_3_lut_4_lut_4_lut (.A(index_i[0]), .B(n29403), 
         .C(index_i[3]), .D(n29418), .Z(n859_adj_3360)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B ((D)+!C)+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_2_i859_3_lut_4_lut_4_lut.init = 16'h5c0c;
    LUT4 i23844_3_lut (.A(n109_adj_2954), .B(n124_adj_3214), .C(index_i[4]), 
         .Z(n23870)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23844_3_lut.init = 16'hcaca;
    LUT4 mux_206_Mux_4_i142_3_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[3]), 
         .C(index_i[2]), .Z(n142_adj_3429)) /* synthesis lut_function=(A (B (C))+!A !(B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_4_i142_3_lut_4_lut_3_lut.init = 16'h9595;
    LUT4 i23893_3_lut (.A(n29481), .B(n23147), .C(index_i[4]), .Z(n23148)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23893_3_lut.init = 16'hcaca;
    LUT4 mux_206_Mux_5_i573_3_lut_3_lut (.A(index_i[0]), .B(index_i[4]), 
         .C(n572_adj_3430), .Z(n573)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_5_i573_3_lut_3_lut.init = 16'hd1d1;
    PFUMX i20768 (.BLUT(n23248), .ALUT(n23249), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_1768[11]));
    LUT4 mux_207_Mux_0_i939_4_lut (.A(n588), .B(n29334), .C(index_q[3]), 
         .D(index_q[2]), .Z(n939_adj_3139)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_0_i939_4_lut.init = 16'hfaca;
    LUT4 i21328_3_lut (.A(n747_adj_3256), .B(n762_adj_3316), .C(index_q[4]), 
         .Z(n23810)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21328_3_lut.init = 16'hcaca;
    LUT4 i21327_3_lut (.A(n716_adj_3258), .B(n16626), .C(index_q[4]), 
         .Z(n23809)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21327_3_lut.init = 16'hcaca;
    PFUMX i20936 (.BLUT(n23416), .ALUT(n23417), .C0(index_q[4]), .Z(n23418));
    LUT4 i20841_3_lut_then_4_lut (.A(index_q[4]), .B(index_q[0]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n29510)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A !(B (C)+!B !((D)+!C))) */ ;
    defparam i20841_3_lut_then_4_lut.init = 16'h95a5;
    LUT4 mux_206_Mux_6_i157_3_lut_4_lut (.A(n29185), .B(index_i[2]), .C(index_i[3]), 
         .D(n32028), .Z(n157_adj_3225)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_6_i157_3_lut_4_lut.init = 16'hf606;
    LUT4 i11249_3_lut_4_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[4]), .Z(n13548)) /* synthesis lut_function=(!(A (B)+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11249_3_lut_4_lut_4_lut_3_lut.init = 16'h6262;
    LUT4 i20634_3_lut_4_lut_4_lut (.A(index_i[0]), .B(n29431), .C(index_i[3]), 
         .D(n29418), .Z(n23116)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20634_3_lut_4_lut_4_lut.init = 16'hc5c0;
    LUT4 i23896_3_lut (.A(n23143), .B(n23144), .C(index_i[4]), .Z(n23145)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23896_3_lut.init = 16'hcaca;
    L6MUX21 i14989394_i1 (.D0(n25036), .D1(n25274), .SD(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_1768[0]));
    L6MUX21 i14983391_i1 (.D0(n25005), .D1(n25343), .SD(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_1783[0]));
    L6MUX21 i28747 (.D0(n31749), .D1(n31746), .SD(index_q[7]), .Z(n31750));
    PFUMX i21953 (.BLUT(n24452), .ALUT(n24453), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_1768[2]));
    PFUMX i28745 (.BLUT(n31748), .ALUT(n31747), .C0(index_q[5]), .Z(n31749));
    PFUMX i22342 (.BLUT(n24841), .ALUT(n24842), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_1768[8]));
    LUT4 mux_206_Mux_6_i251_3_lut_4_lut (.A(n29185), .B(index_i[2]), .C(index_i[3]), 
         .D(n29440), .Z(n251_adj_3064)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_6_i251_3_lut_4_lut.init = 16'hf606;
    PFUMX mux_206_Mux_14_i1023 (.BLUT(n511_adj_3226), .ALUT(n22033), .C0(index_i[9]), 
          .Z(quarter_wave_sample_register_i_15__N_1768[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    PFUMX i28743 (.BLUT(n25277), .ALUT(n31745), .C0(index_q[6]), .Z(n31746));
    PFUMX i22587 (.BLUT(n25086), .ALUT(n25087), .C0(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_1783[2]));
    L6MUX21 i22495 (.D0(n24985), .D1(n24986), .SD(index_q[5]), .Z(n24996));
    L6MUX21 i22496 (.D0(n24987), .D1(n24988), .SD(index_q[5]), .Z(n24997));
    LUT4 i11055_3_lut_4_lut (.A(n29185), .B(index_i[2]), .C(n29365), .D(n29440), 
         .Z(n444_adj_3002)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11055_3_lut_4_lut.init = 16'h6f60;
    PFUMX mux_207_Mux_14_i1023 (.BLUT(n511), .ALUT(n22031), .C0(index_q[9]), 
          .Z(quarter_wave_sample_register_q_15__N_1783[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 mux_206_Mux_2_i413_3_lut (.A(n397_adj_3347), .B(n954_adj_3431), 
         .C(index_i[4]), .Z(n413_adj_3133)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_2_i413_3_lut.init = 16'hcaca;
    PFUMX i22592 (.BLUT(n25089), .ALUT(n25090), .C0(index_i[4]), .Z(n25093));
    L6MUX21 i22497 (.D0(n24989), .D1(n24990), .SD(index_q[5]), .Z(n24998));
    PFUMX i22521 (.BLUT(n25006), .ALUT(n25007), .C0(index_i[5]), .Z(n25022));
    LUT4 mux_206_Mux_4_i747_3_lut_4_lut (.A(n29185), .B(index_i[2]), .C(index_i[3]), 
         .D(n32020), .Z(n747_adj_2984)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_4_i747_3_lut_4_lut.init = 16'hf606;
    PFUMX i22735 (.BLUT(n25234), .ALUT(n25235), .C0(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_1783[8]));
    LUT4 mux_206_Mux_2_i317_3_lut (.A(n668), .B(n316_adj_3344), .C(index_i[4]), 
         .Z(n317_adj_3130)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_2_i317_3_lut.init = 16'hcaca;
    L6MUX21 i28715 (.D0(n31712), .D1(n31709), .SD(index_i[7]), .Z(n31713));
    PFUMX i28713 (.BLUT(n31711), .ALUT(n31710), .C0(index_i[5]), .Z(n31712));
    L6MUX21 i22809 (.D0(n25306), .D1(n25307), .SD(index_i[8]), .Z(n25310));
    PFUMX i22593 (.BLUT(n25091), .ALUT(n25092), .C0(index_i[4]), .Z(n25094));
    PFUMX i28711 (.BLUT(n25172), .ALUT(n31708), .C0(index_i[6]), .Z(n31709));
    LUT4 mux_206_Mux_2_i286_3_lut (.A(n270_adj_3343), .B(n653_adj_3104), 
         .C(index_i[4]), .Z(n286_adj_3129)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_2_i286_3_lut.init = 16'hcaca;
    PFUMX i22522 (.BLUT(n25008), .ALUT(n25009), .C0(index_i[5]), .Z(n25023));
    LUT4 mux_206_Mux_4_i252_4_lut_4_lut (.A(index_i[0]), .B(index_i[3]), 
         .C(n29418), .D(index_i[4]), .Z(n252_adj_3042)) /* synthesis lut_function=(!(A (B (D)+!B !(D))+!A !(B ((D)+!C)+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_4_i252_4_lut_4_lut.init = 16'h669d;
    PFUMX i25104 (.BLUT(n26754), .ALUT(n29422), .C0(index_i[5]), .Z(n26755));
    LUT4 i23905_3_lut (.A(n142_adj_3203), .B(n15097), .C(index_i[4]), 
         .Z(n158_adj_3127)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23905_3_lut.init = 16'hcaca;
    L6MUX21 i26452 (.D0(n28365), .D1(n29026), .SD(index_i[6]), .Z(n638));
    PFUMX i26450 (.BLUT(n28364), .ALUT(n28363), .C0(index_i[5]), .Z(n28365));
    PFUMX i22234 (.BLUT(n24731), .ALUT(n24732), .C0(index_i[8]), .Z(n24735));
    LUT4 mux_206_Mux_3_i444_3_lut_4_lut (.A(index_i[0]), .B(index_i[3]), 
         .C(n29400), .D(index_i[4]), .Z(n444_adj_3110)) /* synthesis lut_function=(!(A (B (D)+!B (C (D)))+!A !(B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_3_i444_3_lut_4_lut.init = 16'h46aa;
    LUT4 i23909_3_lut (.A(n23119), .B(n29477), .C(index_i[4]), .Z(n23121)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23909_3_lut.init = 16'hcaca;
    LUT4 i24624_2_lut (.A(index_q[5]), .B(index_q[4]), .Z(n24091)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i24624_2_lut.init = 16'heeee;
    L6MUX21 i22235 (.D0(n24733), .D1(n24734), .SD(index_i[8]), .Z(n24736));
    LUT4 mux_206_Mux_3_i796_3_lut_3_lut (.A(index_i[4]), .B(n731_adj_3186), 
         .C(index_i[2]), .Z(n796_adj_3407)) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam mux_206_Mux_3_i796_3_lut_3_lut.init = 16'he4e4;
    PFUMX i20939 (.BLUT(n23419), .ALUT(n23420), .C0(index_q[4]), .Z(n23421));
    LUT4 i1_3_lut_adj_187 (.A(index_q[0]), .B(index_q[4]), .C(index_q[2]), 
         .Z(n22572)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_3_lut_adj_187.init = 16'hfefe;
    LUT4 mux_206_Mux_3_i924_3_lut (.A(n908_adj_3337), .B(index_i[0]), .C(index_i[4]), 
         .Z(n924)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_3_i924_3_lut.init = 16'hcaca;
    LUT4 i24494_2_lut_rep_664 (.A(index_i[1]), .B(index_i[2]), .Z(n29324)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i24494_2_lut_rep_664.init = 16'h9999;
    LUT4 mux_206_Mux_3_i891_3_lut (.A(n541_adj_3058), .B(n890_adj_2973), 
         .C(index_i[4]), .Z(n891_adj_3121)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_3_i891_3_lut.init = 16'hcaca;
    L6MUX21 i21919 (.D0(n24415), .D1(n24416), .SD(index_i[7]), .Z(n24420));
    LUT4 mux_206_Mux_2_i731_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n731_adj_3420)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_2_i731_3_lut_4_lut_4_lut.init = 16'h6cc6;
    LUT4 i22324_3_lut (.A(n141), .B(n32054), .C(index_q[3]), .Z(n24825)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22324_3_lut.init = 16'hcaca;
    LUT4 i22323_3_lut (.A(n85), .B(n29461), .C(index_q[3]), .Z(n24824)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22323_3_lut.init = 16'hcaca;
    L6MUX21 i26433 (.D0(n28345), .D1(n28342), .SD(index_i[4]), .Z(n509));
    LUT4 n442_bdd_2_lut_25675_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[3]), 
         .Z(n27413)) /* synthesis lut_function=(A (B+(C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n442_bdd_2_lut_25675_3_lut.init = 16'hf9f9;
    LUT4 mux_206_Mux_0_i93_3_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .Z(n93_adj_3268)) /* synthesis lut_function=(A (B)+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i93_3_lut_3_lut.init = 16'h9c9c;
    LUT4 i22321_3_lut (.A(n32054), .B(n29470), .C(index_q[3]), .Z(n24822)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22321_3_lut.init = 16'hcaca;
    LUT4 mux_206_Mux_3_i669_3_lut (.A(n653_adj_3104), .B(n668), .C(index_i[4]), 
         .Z(n669_adj_3117)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_3_i669_3_lut.init = 16'hcaca;
    PFUMX i26431 (.BLUT(n28344), .ALUT(n28343), .C0(index_i[5]), .Z(n28345));
    LUT4 i11073_4_lut (.A(n29400), .B(n29180), .C(index_i[3]), .D(index_i[4]), 
         .Z(n13369)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B ((D)+!C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11073_4_lut.init = 16'h3afa;
    LUT4 i20667_3_lut (.A(n498), .B(n29403), .C(index_i[3]), .Z(n23149)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20667_3_lut.init = 16'hcaca;
    LUT4 i23891_3_lut (.A(n23149), .B(n23150), .C(index_i[4]), .Z(n23151)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23891_3_lut.init = 16'hcaca;
    LUT4 i21918_3_lut (.A(n24413), .B(n24414), .C(index_i[7]), .Z(n24419)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21918_3_lut.init = 16'hcaca;
    PFUMX i21973 (.BLUT(n24470), .ALUT(n24471), .C0(index_q[8]), .Z(n24474));
    L6MUX21 i21974 (.D0(n24472), .D1(n24473), .SD(index_q[8]), .Z(n24475));
    L6MUX21 i22003 (.D0(n24499), .D1(n24500), .SD(index_i[7]), .Z(n24504));
    LUT4 i21913_3_lut (.A(n24403), .B(n24404), .C(index_i[6]), .Z(n24414)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21913_3_lut.init = 16'hcaca;
    L6MUX21 i22034 (.D0(n24530), .D1(n24531), .SD(index_q[7]), .Z(n24535));
    LUT4 i20841_3_lut_else_4_lut (.A(index_q[4]), .B(index_q[0]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n29509)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A !(C (D)+!C !(D)))) */ ;
    defparam i20841_3_lut_else_4_lut.init = 16'h5a85;
    LUT4 i22000_3_lut (.A(n24493), .B(n24494), .C(index_i[7]), .Z(n24501)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22000_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_2_i491_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n491_adj_3371)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A !(B (C)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_2_i491_3_lut_4_lut_4_lut.init = 16'h6a5a;
    LUT4 i21993_3_lut (.A(n24479), .B(n27488), .C(index_i[6]), .Z(n24494)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21993_3_lut.init = 16'hcaca;
    LUT4 i22002_3_lut (.A(n24497), .B(n24498), .C(index_i[7]), .Z(n24503)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22002_3_lut.init = 16'hcaca;
    LUT4 i21996_3_lut (.A(n27513), .B(n24486), .C(index_i[6]), .Z(n24497)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21996_3_lut.init = 16'hcaca;
    L6MUX21 i22470 (.D0(n24966), .D1(n24967), .SD(index_q[7]), .Z(n24971));
    PFUMX i22504 (.BLUT(n25003), .ALUT(n25004), .C0(index_q[8]), .Z(n25005));
    PFUMX i22535 (.BLUT(n25034), .ALUT(n25035), .C0(index_i[8]), .Z(n25036));
    LUT4 i22031_3_lut (.A(n24524), .B(n24525), .C(index_q[7]), .Z(n24532)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22031_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_519_3_lut (.A(index_i[2]), .B(index_i[0]), .C(index_i[1]), 
         .Z(n29179)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_2_lut_rep_519_3_lut.init = 16'hfefe;
    LUT4 i22024_3_lut (.A(n24510), .B(n27577), .C(index_q[6]), .Z(n24525)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22024_3_lut.init = 16'hcaca;
    L6MUX21 i22523 (.D0(n25010), .D1(n25011), .SD(index_i[5]), .Z(n25024));
    PFUMX i22524 (.BLUT(n25012), .ALUT(n25013), .C0(index_i[5]), .Z(n25025));
    LUT4 i22033_3_lut (.A(n24528), .B(n24529), .C(index_q[7]), .Z(n24534)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22033_3_lut.init = 16'hcaca;
    LUT4 i22027_3_lut (.A(n27588), .B(n24517), .C(index_q[6]), .Z(n24528)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22027_3_lut.init = 16'hcaca;
    LUT4 mux_206_Mux_0_i739_3_lut_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n931)) /* synthesis lut_function=(!(A (B+(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i739_3_lut_3_lut_3_lut.init = 16'h5656;
    PFUMX i25102 (.BLUT(n29426), .ALUT(n26752), .C0(index_i[2]), .Z(n26753));
    PFUMX i22820 (.BLUT(n781_adj_3432), .ALUT(n796_adj_3204), .C0(index_q[4]), 
          .Z(n25321));
    LUT4 i23919_3_lut (.A(n23104), .B(n23105), .C(index_i[4]), .Z(n23106)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23919_3_lut.init = 16'hcaca;
    PFUMX i26428 (.BLUT(n28341), .ALUT(n28340), .C0(index_i[6]), .Z(n28342));
    PFUMX i27119 (.BLUT(n29551), .ALUT(n29552), .C0(index_q[8]), .Z(n29553));
    LUT4 i11071_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[4]), .Z(n444_adj_3200)) /* synthesis lut_function=(!(A (B)+!A !(B (C (D))+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11071_3_lut_4_lut_4_lut_4_lut.init = 16'h6333;
    LUT4 i22469_3_lut (.A(n24964), .B(n24965), .C(index_q[7]), .Z(n24970)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22469_3_lut.init = 16'hcaca;
    LUT4 i22464_3_lut (.A(n24954), .B(n24955), .C(index_q[6]), .Z(n24965)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22464_3_lut.init = 16'hcaca;
    LUT4 mux_206_Mux_1_i882_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n882_adj_3378)) /* synthesis lut_function=(A ((C)+!B)+!A !((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_1_i882_3_lut_3_lut.init = 16'ha6a6;
    LUT4 mux_206_Mux_3_i476_3_lut (.A(n460_adj_3028), .B(n285_adj_3027), 
         .C(index_i[4]), .Z(n476_adj_3111)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_3_i476_3_lut.init = 16'hcaca;
    LUT4 mux_206_Mux_8_i716_3_lut_4_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[1]), .D(index_i[3]), .Z(n716_adj_2965)) /* synthesis lut_function=(!(A (D)+!A !(B+(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_8_i716_3_lut_4_lut_4_lut_4_lut.init = 16'h55fe;
    LUT4 mux_207_Mux_5_i53_3_lut_4_lut_3_lut_rep_803 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29463)) /* synthesis lut_function=(A ((C)+!B)+!A (B)) */ ;
    defparam mux_207_Mux_5_i53_3_lut_4_lut_3_lut_rep_803.init = 16'he6e6;
    PFUMX i20942 (.BLUT(n23422), .ALUT(n23423), .C0(index_q[4]), .Z(n23424));
    LUT4 i11053_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(n29329), .D(index_i[4]), .Z(n221)) /* synthesis lut_function=(!(A (B)+!A (B (C+(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11053_3_lut_4_lut_4_lut_4_lut.init = 16'h3336;
    LUT4 mux_206_Mux_3_i413_3_lut (.A(n397_adj_3433), .B(n29322), .C(index_i[4]), 
         .Z(n413_adj_3109)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_3_i413_3_lut.init = 16'hcaca;
    PFUMX i22773 (.BLUT(n25272), .ALUT(n25273), .C0(index_i[8]), .Z(n25274));
    PFUMX i22805 (.BLUT(n25298), .ALUT(n25299), .C0(index_i[7]), .Z(n25306));
    LUT4 mux_206_Mux_5_i954_3_lut_3_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[1]), .Z(n954_adj_3431)) /* synthesis lut_function=(!(A (C)+!A (B+((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_5_i954_3_lut_3_lut_4_lut_4_lut.init = 16'h0a1a;
    PFUMX i22806 (.BLUT(n25300), .ALUT(n25301), .C0(index_i[7]), .Z(n25307));
    LUT4 i21851_3_lut (.A(n24341), .B(n24342), .C(index_i[6]), .Z(n24352)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21851_3_lut.init = 16'hcaca;
    PFUMX i22842 (.BLUT(n25341), .ALUT(n25342), .C0(index_q[8]), .Z(n25343));
    PFUMX i27117 (.BLUT(n29548), .ALUT(n29549), .C0(index_q[3]), .Z(n62_adj_3412));
    LUT4 mux_206_Mux_3_i286_4_lut (.A(n93), .B(index_i[2]), .C(index_i[4]), 
         .D(n15092), .Z(n286_adj_3106)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_3_i286_4_lut.init = 16'h3aca;
    LUT4 mux_207_Mux_0_i923_3_lut (.A(n29460), .B(n29470), .C(index_q[3]), 
         .Z(n923)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_0_i923_3_lut.init = 16'hcaca;
    LUT4 i7619_2_lut (.A(index_q[4]), .B(index_q[5]), .Z(n9850)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i7619_2_lut.init = 16'h8888;
    L6MUX21 i22232 (.D0(n24727), .D1(n24728), .SD(index_i[7]), .Z(n24733));
    L6MUX21 i22233 (.D0(n24729), .D1(n24730), .SD(index_i[7]), .Z(n24734));
    LUT4 mux_206_Mux_3_i507_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[4]), .D(n491_adj_2976), .Z(n507_adj_3112)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_3_i507_3_lut_4_lut.init = 16'h6f60;
    L6MUX21 i21854 (.D0(n24347), .D1(n24348), .SD(index_i[7]), .Z(n24355));
    L6MUX21 i21855 (.D0(n24349), .D1(n24350), .SD(index_i[7]), .Z(n24356));
    LUT4 mux_206_Mux_4_i363_3_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n325_adj_2972)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_4_i363_3_lut_4_lut_3_lut.init = 16'h6d6d;
    L6MUX21 i21914 (.D0(n24405), .D1(n24406), .SD(index_i[6]), .Z(n24415));
    L6MUX21 i21916 (.D0(n24409), .D1(n24410), .SD(index_i[7]), .Z(n24417));
    L6MUX21 i21917 (.D0(n24411), .D1(n24412), .SD(index_i[7]), .Z(n24418));
    LUT4 i12682_2_lut_rep_428_3_lut_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[1]), .Z(n29088)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12682_2_lut_rep_428_3_lut_4_lut.init = 16'hf0e0;
    LUT4 mux_206_Mux_0_i747_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n747_adj_3434)) /* synthesis lut_function=(!(A (B+!(C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i747_3_lut_4_lut_4_lut_4_lut.init = 16'h6556;
    L6MUX21 i20786 (.D0(n23266), .D1(n23267), .SD(index_q[7]), .Z(n23268));
    LUT4 mux_206_Mux_3_i158_3_lut (.A(n142_adj_3427), .B(n157_adj_3248), 
         .C(index_i[4]), .Z(n158_adj_3093)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_3_i158_3_lut.init = 16'hcaca;
    LUT4 i8881_2_lut (.A(index_i[4]), .B(index_i[5]), .Z(n11112)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i8881_2_lut.init = 16'h8888;
    L6MUX21 i22338 (.D0(n24833), .D1(n24834), .SD(index_i[7]), .Z(n24839));
    LUT4 i17716_4_lut (.A(index_q[0]), .B(index_q[4]), .C(index_q[1]), 
         .D(n29361), .Z(n286_adj_3435)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i17716_4_lut.init = 16'hccc8;
    L6MUX21 i21948 (.D0(n24442), .D1(n24443), .SD(index_i[7]), .Z(n24449));
    LUT4 i21947_3_lut (.A(n28448), .B(n24441), .C(index_i[7]), .Z(n24448)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21947_3_lut.init = 16'hcaca;
    L6MUX21 i21949 (.D0(n24444), .D1(n24445), .SD(index_i[7]), .Z(n24450));
    LUT4 i22739_3_lut_4_lut_4_lut (.A(n29132), .B(index_q[4]), .C(index_q[5]), 
         .D(n29130), .Z(n25240)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C)+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i22739_3_lut_4_lut_4_lut.init = 16'h0434;
    LUT4 i22364_3_lut (.A(n24854), .B(n24855), .C(index_q[6]), .Z(n24865)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22364_3_lut.init = 16'hcaca;
    LUT4 i12703_2_lut_rep_666 (.A(index_q[2]), .B(index_q[3]), .Z(n29326)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i12703_2_lut_rep_666.init = 16'h8888;
    L6MUX21 i22526 (.D0(n25016), .D1(n25017), .SD(index_i[5]), .Z(n25027));
    LUT4 mux_206_Mux_5_i53_3_lut_4_lut_3_lut_rep_767 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29427)) /* synthesis lut_function=(A ((C)+!B)+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_5_i53_3_lut_4_lut_3_lut_rep_767.init = 16'he6e6;
    PFUMX i22339 (.BLUT(n24835), .ALUT(n24836), .C0(index_i[7]), .Z(n24840));
    LUT4 i13840_2_lut_2_lut_3_lut (.A(index_q[2]), .B(index_q[3]), .C(index_q[0]), 
         .Z(n16249)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i13840_2_lut_2_lut_3_lut.init = 16'h0808;
    LUT4 mux_206_Mux_3_i125_3_lut (.A(n109_adj_2961), .B(n526), .C(index_i[4]), 
         .Z(n125_adj_3088)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_3_i125_3_lut.init = 16'hcaca;
    LUT4 mux_206_Mux_5_i581_3_lut_3_lut_rep_769 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29429)) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_5_i581_3_lut_3_lut_rep_769.init = 16'h6a6a;
    LUT4 mux_207_Mux_8_i892_3_lut_4_lut (.A(n29132), .B(index_q[4]), .C(index_q[5]), 
         .D(n860_adj_3153), .Z(n892_adj_3211)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_8_i892_3_lut_4_lut.init = 16'h4f40;
    PFUMX i22599 (.BLUT(n25096), .ALUT(n25097), .C0(index_i[4]), .Z(n25100));
    LUT4 i13955_2_lut_rep_470_3_lut (.A(index_q[2]), .B(index_q[3]), .C(index_q[1]), 
         .Z(n29130)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i13955_2_lut_rep_470_3_lut.init = 16'h8080;
    L6MUX21 i22527 (.D0(n25018), .D1(n25019), .SD(index_i[5]), .Z(n25028));
    L6MUX21 i26380 (.D0(n28286), .D1(n29028), .SD(index_q[6]), .Z(n638_adj_3132));
    LUT4 i21809_1_lut_2_lut (.A(index_q[2]), .B(index_q[3]), .Z(n24310)) /* synthesis lut_function=(!(A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i21809_1_lut_2_lut.init = 16'h7777;
    LUT4 mux_206_Mux_0_i708_3_lut_4_lut_4_lut_3_lut_rep_770 (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[2]), .Z(n29430)) /* synthesis lut_function=(!(A (B)+!A ((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i708_3_lut_4_lut_4_lut_3_lut_rep_770.init = 16'h2626;
    LUT4 i22247_3_lut_3_lut_3_lut_4_lut (.A(index_q[2]), .B(index_q[3]), 
         .C(index_q[4]), .D(index_q[1]), .Z(n24748)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i22247_3_lut_3_lut_3_lut_4_lut.init = 16'h878f;
    LUT4 i17691_3_lut_3_lut_3_lut_4_lut (.A(index_q[2]), .B(index_q[3]), 
         .C(index_q[1]), .D(index_q[0]), .Z(n20005)) /* synthesis lut_function=(!(A (B (C)+!B !(C (D)+!C !(D)))+!A !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i17691_3_lut_3_lut_3_lut_4_lut.init = 16'h780f;
    PFUMX i26378 (.BLUT(n28285), .ALUT(n28284), .C0(index_q[5]), .Z(n28286));
    PFUMX i22600 (.BLUT(n25098), .ALUT(n25099), .C0(index_i[4]), .Z(n25101));
    LUT4 index_q_6__bdd_3_lut_4_lut (.A(index_q[2]), .B(index_q[3]), .C(n29465), 
         .D(index_q[6]), .Z(n28503)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(D))+!A !(D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam index_q_6__bdd_3_lut_4_lut.init = 16'h887f;
    LUT4 i22581_3_lut (.A(n25074), .B(n25075), .C(index_q[7]), .Z(n25082)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22581_3_lut.init = 16'hcaca;
    L6MUX21 i22528 (.D0(n25020), .D1(n25021), .SD(index_i[5]), .Z(n25029));
    LUT4 i11102_3_lut_3_lut_3_lut_4_lut (.A(index_q[2]), .B(index_q[3]), 
         .C(index_q[1]), .D(index_q[0]), .Z(n541_adj_3084)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i11102_3_lut_3_lut_3_lut_4_lut.init = 16'h870f;
    LUT4 i21876_4_lut (.A(n29517), .B(n1002_adj_3436), .C(index_i[5]), 
         .D(index_i[4]), .Z(n24377)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;
    defparam i21876_4_lut.init = 16'hfaca;
    LUT4 i17690_3_lut_3_lut_4_lut (.A(index_q[2]), .B(index_q[3]), .C(index_q[1]), 
         .D(index_q[0]), .Z(n20004)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i17690_3_lut_3_lut_4_lut.init = 16'hf078;
    LUT4 i12659_2_lut_rep_407_3_lut_4_lut (.A(index_q[2]), .B(index_q[3]), 
         .C(index_q[4]), .D(n29459), .Z(n29067)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i12659_2_lut_rep_407_3_lut_4_lut.init = 16'hf8f0;
    LUT4 mux_206_Mux_4_i860_3_lut (.A(n506_adj_3292), .B(n26722), .C(index_i[4]), 
         .Z(n860_adj_3077)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_4_i860_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_7_i924_3_lut_3_lut_4_lut (.A(index_q[2]), .B(index_q[3]), 
         .C(index_q[4]), .D(n29459), .Z(n924_adj_3437)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_7_i924_3_lut_3_lut_4_lut.init = 16'h878f;
    LUT4 mux_206_Mux_5_i459_3_lut_4_lut_3_lut_rep_771 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29431)) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_5_i459_3_lut_4_lut_3_lut_rep_771.init = 16'h6b6b;
    LUT4 mux_206_Mux_0_i30_3_lut (.A(n29380), .B(n29408), .C(index_i[3]), 
         .Z(n30_adj_3232)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i30_3_lut.init = 16'hcaca;
    LUT4 i12583_2_lut_rep_406_3_lut_4_lut (.A(index_q[2]), .B(index_q[3]), 
         .C(index_q[4]), .D(n29465), .Z(n29066)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i12583_2_lut_rep_406_3_lut_4_lut.init = 16'hf8f0;
    PFUMX i22559 (.BLUT(n158_adj_3209), .ALUT(n189_adj_3006), .C0(index_q[5]), 
          .Z(n25060));
    LUT4 mux_206_Mux_9_i285_3_lut_3_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[1]), .Z(n285_adj_3043)) /* synthesis lut_function=(A (C)+!A !(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_9_i285_3_lut_3_lut_4_lut_4_lut.init = 16'ha0a1;
    LUT4 mux_206_Mux_6_i889_3_lut_rep_722 (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[2]), .Z(n29382)) /* synthesis lut_function=(!(A (B (C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_6_i889_3_lut_rep_722.init = 16'h7e7e;
    LUT4 i22223_3_lut (.A(n190), .B(n26902), .C(index_i[6]), .Z(n24724)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22223_3_lut.init = 16'hcaca;
    LUT4 i22245_3_lut_4_lut_3_lut (.A(index_q[3]), .B(index_q[4]), .C(n29168), 
         .Z(n24746)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i22245_3_lut_4_lut_3_lut.init = 16'h6464;
    LUT4 mux_206_Mux_5_i262_3_lut_4_lut_3_lut_rep_772 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29432)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_5_i262_3_lut_4_lut_3_lut_rep_772.init = 16'h6464;
    LUT4 i21405_3_lut_4_lut_4_lut (.A(n29177), .B(index_i[4]), .C(index_i[3]), 
         .D(n29176), .Z(n23887)) /* synthesis lut_function=(A (B (C)+!B !(C+!(D)))+!A (B (C)+!B (C+(D)))) */ ;
    defparam i21405_3_lut_4_lut_4_lut.init = 16'hd3d0;
    L6MUX21 i20804 (.D0(n23284), .D1(n23285), .SD(index_i[7]), .Z(n23286));
    LUT4 i1_2_lut_rep_590 (.A(index_q[6]), .B(index_q[7]), .Z(n29250)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i1_2_lut_rep_590.init = 16'heeee;
    LUT4 mux_207_Mux_2_i221_4_lut_4_lut (.A(index_q[3]), .B(index_q[4]), 
         .C(n29165), .D(n29080), .Z(n221_adj_3438)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (B+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_2_i221_4_lut_4_lut.init = 16'hf7c4;
    LUT4 mux_206_Mux_6_i7_3_lut_4_lut_3_lut_rep_773 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29433)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_6_i7_3_lut_4_lut_3_lut_rep_773.init = 16'hd6d6;
    LUT4 i10024_4_lut_4_lut (.A(index_q[3]), .B(index_q[0]), .C(index_q[1]), 
         .D(index_q[2]), .Z(n12256)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (D)+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i10024_4_lut_4_lut.init = 16'h0bf4;
    LUT4 i23939_3_lut (.A(n23068), .B(n23069), .C(index_i[4]), .Z(n23070)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23939_3_lut.init = 16'hcaca;
    LUT4 i12532_4_lut_4_lut (.A(index_q[3]), .B(index_q[2]), .C(index_q[0]), 
         .D(index_q[1]), .Z(n875_adj_3026)) /* synthesis lut_function=((B (C)+!B (D))+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i12532_4_lut_4_lut.init = 16'hf7d5;
    LUT4 mux_207_Mux_1_i987_3_lut_4_lut_4_lut (.A(index_q[3]), .B(n986_adj_3401), 
         .C(index_q[4]), .D(n32054), .Z(n987_adj_3351)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_1_i987_3_lut_4_lut_4_lut.init = 16'hc5c0;
    LUT4 i22330_3_lut (.A(n27464), .B(n25095), .C(index_i[6]), .Z(n24831)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22330_3_lut.init = 16'hcaca;
    L6MUX21 i21971 (.D0(n24466), .D1(n24467), .SD(index_q[7]), .Z(n24472));
    L6MUX21 i21972 (.D0(n24468), .D1(n24469), .SD(index_q[7]), .Z(n24473));
    LUT4 i22335_3_lut_4_lut (.A(n29074), .B(n29069), .C(index_i[5]), .D(index_i[6]), 
         .Z(n24836)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (B+((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i22335_3_lut_4_lut.init = 16'hffc5;
    LUT4 i12527_2_lut_4_lut_4_lut_4_lut (.A(index_q[3]), .B(index_q[2]), 
         .C(index_q[1]), .D(index_q[0]), .Z(n668_adj_3439)) /* synthesis lut_function=(!(A+!(B (C)+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i12527_2_lut_4_lut_4_lut_4_lut.init = 16'h5041;
    LUT4 i21962_3_lut (.A(n190_adj_3411), .B(n253), .C(index_q[6]), .Z(n24463)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21962_3_lut.init = 16'hcaca;
    L6MUX21 i21997 (.D0(n24487), .D1(n24488), .SD(index_i[6]), .Z(n24498));
    L6MUX21 i21998 (.D0(n24489), .D1(n24490), .SD(index_i[6]), .Z(n24499));
    LUT4 i21334_4_lut_3_lut (.A(index_q[3]), .B(index_q[4]), .C(n29165), 
         .Z(n23816)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i21334_4_lut_3_lut.init = 16'h6565;
    L6MUX21 i22367 (.D0(n24860), .D1(n24861), .SD(index_q[7]), .Z(n24868));
    L6MUX21 i22368 (.D0(n24862), .D1(n24863), .SD(index_q[7]), .Z(n24869));
    L6MUX21 i22001 (.D0(n24495), .D1(n24496), .SD(index_i[7]), .Z(n24502));
    L6MUX21 i22028 (.D0(n24518), .D1(n24519), .SD(index_q[6]), .Z(n24529));
    LUT4 n45_bdd_2_lut_3_lut_3_lut_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[1]), .D(index_i[3]), .Z(n27537)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n45_bdd_2_lut_3_lut_3_lut_4_lut.init = 16'h00fe;
    LUT4 i11091_3_lut_3_lut (.A(index_q[3]), .B(index_q[4]), .C(n13386), 
         .Z(n13387)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i11091_3_lut_3_lut.init = 16'h7474;
    L6MUX21 i22029 (.D0(n24520), .D1(n24521), .SD(index_q[6]), .Z(n24530));
    L6MUX21 i22032 (.D0(n24526), .D1(n24527), .SD(index_q[7]), .Z(n24533));
    LUT4 i21963_3_lut (.A(n24828), .B(n23343), .C(index_q[6]), .Z(n24464)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21963_3_lut.init = 16'hcaca;
    L6MUX21 i22465 (.D0(n24956), .D1(n24957), .SD(index_q[6]), .Z(n24966));
    L6MUX21 i22467 (.D0(n24960), .D1(n24961), .SD(index_q[7]), .Z(n24968));
    L6MUX21 i22468 (.D0(n24962), .D1(n24963), .SD(index_q[7]), .Z(n24969));
    L6MUX21 i22582 (.D0(n25076), .D1(n25077), .SD(index_q[7]), .Z(n25083));
    L6MUX21 i22583 (.D0(n25078), .D1(n25079), .SD(index_q[7]), .Z(n25084));
    PFUMX i22584 (.BLUT(n25080), .ALUT(n25081), .C0(index_q[7]), .Z(n25085));
    LUT4 n22_bdd_3_lut_25601_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n26722)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C))+!A !(B (C+!(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n22_bdd_3_lut_25601_4_lut_4_lut.init = 16'h5ad6;
    LUT4 mux_206_Mux_0_i46_3_lut_4_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[1]), .D(index_i[3]), .Z(n46_adj_3270)) /* synthesis lut_function=(A (D)+!A (B+(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i46_3_lut_4_lut_4_lut_4_lut.init = 16'hfe55;
    LUT4 i21514_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n23996)) /* synthesis lut_function=(A (B (C)+!B !(C (D)+!C !(D)))+!A (B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21514_3_lut_4_lut_4_lut.init = 16'hd6a5;
    L6MUX21 i22668 (.D0(n25167), .D1(n25168), .SD(index_i[7]), .Z(n25169));
    LUT4 i22499_3_lut (.A(n24993), .B(n29906), .C(index_q[6]), .Z(n25000)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22499_3_lut.init = 16'hcaca;
    LUT4 i22500_3_lut (.A(n27750), .B(n24996), .C(index_q[6]), .Z(n25001)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22500_3_lut.init = 16'hcaca;
    LUT4 i22530_3_lut (.A(n25024), .B(n25025), .C(index_i[6]), .Z(n25031)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22530_3_lut.init = 16'hcaca;
    LUT4 i22531_3_lut (.A(n28105), .B(n25027), .C(index_i[6]), .Z(n25032)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22531_3_lut.init = 16'hcaca;
    LUT4 mux_206_Mux_0_i220_3_lut (.A(n29406), .B(n29436), .C(index_i[3]), 
         .Z(n220)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i220_3_lut.init = 16'hcaca;
    LUT4 i23941_3_lut (.A(n23062), .B(n23063), .C(index_i[4]), .Z(n23064)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23941_3_lut.init = 16'hcaca;
    LUT4 i22723_3_lut (.A(n27561), .B(n24807), .C(index_q[6]), .Z(n25224)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22723_3_lut.init = 16'hcaca;
    L6MUX21 i22716 (.D0(n25211), .D1(n25212), .SD(index_q[7]), .Z(n25217));
    L6MUX21 i22731 (.D0(n25226), .D1(n25227), .SD(index_q[7]), .Z(n25232));
    PFUMX i22732 (.BLUT(n25228), .ALUT(n25229), .C0(index_q[7]), .Z(n25233));
    LUT4 mux_207_Mux_10_i701_4_lut_4_lut (.A(n29134), .B(index_q[4]), .C(index_q[5]), 
         .D(n29068), .Z(n701)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B (C (D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_10_i701_4_lut_4_lut.init = 16'h3efe;
    L6MUX21 i22742 (.D0(n25241), .D1(n25242), .SD(index_q[7]), .Z(n25243));
    LUT4 i20580_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n23062)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20580_3_lut_4_lut.init = 16'h64cc;
    LUT4 mux_207_Mux_7_i956_3_lut_3_lut_4_lut (.A(n29134), .B(index_q[4]), 
         .C(n924_adj_3437), .D(index_q[5]), .Z(n956_adj_3230)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_7_i956_3_lut_3_lut_4_lut.init = 16'h11f0;
    L6MUX21 i22807 (.D0(n25302), .D1(n25303), .SD(index_i[7]), .Z(n25308));
    LUT4 mux_206_Mux_5_i460_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n460_adj_3355)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A !(B (C)+!B !(C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_5_i460_3_lut_4_lut_4_lut.init = 16'h6b5a;
    LUT4 i1_2_lut_rep_591 (.A(index_i[6]), .B(index_i[7]), .Z(n29251)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_2_lut_rep_591.init = 16'heeee;
    L6MUX21 i22222 (.D0(n25102), .D1(n25140), .SD(index_i[6]), .Z(n24723));
    L6MUX21 i22225 (.D0(n23895), .D1(n23898), .SD(index_i[6]), .Z(n24726));
    L6MUX21 i22226 (.D0(n23901), .D1(n23904), .SD(index_i[6]), .Z(n24727));
    L6MUX21 i22227 (.D0(n23907), .D1(n23910), .SD(index_i[6]), .Z(n24728));
    PFUMX i22228 (.BLUT(n23913), .ALUT(n892_adj_3368), .C0(index_i[6]), 
          .Z(n24729));
    LUT4 i20637_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n23119)) /* synthesis lut_function=(!(A (B)+!A (B (C+(D))+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20637_3_lut_3_lut_4_lut.init = 16'h3326;
    L6MUX21 i22243 (.D0(n24742), .D1(n24743), .SD(index_q[6]), .Z(n382_adj_3134));
    L6MUX21 i22250 (.D0(n24749), .D1(n24750), .SD(index_q[6]), .Z(n509_adj_3135));
    LUT4 mux_206_Mux_4_i700_3_lut (.A(n684_adj_3323), .B(index_i[1]), .C(index_i[4]), 
         .Z(n700_adj_3061)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_4_i700_3_lut.init = 16'hcaca;
    LUT4 mux_206_Mux_6_i667_3_lut_rep_724 (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[2]), .Z(n29384)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_6_i667_3_lut_rep_724.init = 16'h1818;
    LUT4 mux_206_Mux_2_i491_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n491_adj_3423)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A !(B (C)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_2_i491_3_lut_4_lut_4_lut.init = 16'h6a5a;
    LUT4 i11040_2_lut_rep_669 (.A(index_i[2]), .B(index_i[3]), .Z(n29329)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11040_2_lut_rep_669.init = 16'h8888;
    LUT4 i1_2_lut_rep_716 (.A(index_i[1]), .B(index_i[0]), .Z(n29376)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_2_lut_rep_716.init = 16'h8888;
    LUT4 mux_206_Mux_4_i669_3_lut (.A(n653_adj_3039), .B(n668_adj_3322), 
         .C(index_i[4]), .Z(n669_adj_3060)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_4_i669_3_lut.init = 16'hcaca;
    LUT4 i14178_3_lut (.A(index_i[3]), .B(index_i[1]), .C(index_i[0]), 
         .Z(n16591)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i14178_3_lut.init = 16'hecec;
    PFUMX i22560 (.BLUT(n221_adj_3438), .ALUT(n23364), .C0(index_q[5]), 
          .Z(n25061));
    LUT4 i11267_3_lut (.A(n13565), .B(n188), .C(index_i[4]), .Z(n13566)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11267_3_lut.init = 16'hcaca;
    LUT4 i21795_2_lut (.A(index_i[3]), .B(index_i[5]), .Z(n24296)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21795_2_lut.init = 16'h8888;
    PFUMX i26307 (.BLUT(n28173), .ALUT(n28170), .C0(index_q[6]), .Z(n28174));
    LUT4 mux_206_Mux_5_i30_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n30_adj_3440)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A (B+!(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_5_i30_3_lut_4_lut.init = 16'hcc67;
    PFUMX i26305 (.BLUT(n28171), .ALUT(n954), .C0(index_q[4]), .Z(n28172));
    L6MUX21 i21846 (.D0(n24331), .D1(n24332), .SD(index_i[6]), .Z(n24347));
    LUT4 i21247_3_lut (.A(n93_adj_3262), .B(n699_adj_2981), .C(index_q[4]), 
         .Z(n23729)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21247_3_lut.init = 16'hcaca;
    LUT4 i22737_3_lut_4_lut_4_lut (.A(n29133), .B(index_q[4]), .C(index_q[5]), 
         .D(n29095), .Z(n25238)) /* synthesis lut_function=(A ((C+!(D))+!B)+!A (B (C+!(D))+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i22737_3_lut_4_lut_4_lut.init = 16'he3ef;
    LUT4 i21246_3_lut (.A(n653), .B(n29063), .C(index_q[4]), .Z(n23728)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21246_3_lut.init = 16'hcaca;
    LUT4 i22238_3_lut_3_lut_4_lut (.A(n29165), .B(index_q[3]), .C(n316_adj_3246), 
         .D(index_q[4]), .Z(n24739)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i22238_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 mux_207_Mux_2_i270_3_lut (.A(n29315), .B(n29316), .C(index_q[3]), 
         .Z(n270)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_2_i270_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_2_i316_3_lut (.A(n29352), .B(n29395), .C(index_q[3]), 
         .Z(n316_adj_3191)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_2_i316_3_lut.init = 16'hcaca;
    LUT4 index_i_6__bdd_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[6]), .D(n29372), .Z(n28576)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam index_i_6__bdd_4_lut_4_lut_4_lut.init = 16'h0f7a;
    L6MUX21 i26286 (.D0(n28147), .D1(n29029), .SD(index_i[6]), .Z(n28148));
    L6MUX21 i21847 (.D0(n24333), .D1(n24334), .SD(index_i[6]), .Z(n24348));
    L6MUX21 i21848 (.D0(n24335), .D1(n24336), .SD(index_i[6]), .Z(n24349));
    PFUMX i26284 (.BLUT(n28146), .ALUT(n29047), .C0(index_i[7]), .Z(n28147));
    PFUMX i27111 (.BLUT(n29539), .ALUT(n29540), .C0(index_i[1]), .Z(n29541));
    L6MUX21 i21849 (.D0(n24337), .D1(n24338), .SD(index_i[6]), .Z(n24350));
    LUT4 mux_206_Mux_6_i635_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n635_adj_3441)) /* synthesis lut_function=(A (B (C+(D))+!B !(D))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_6_i635_3_lut_4_lut.init = 16'hcce6;
    LUT4 mux_207_Mux_10_i317_3_lut_3_lut_4_lut (.A(n29165), .B(index_q[3]), 
         .C(n29130), .D(index_q[4]), .Z(n317_adj_3442)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_10_i317_3_lut_3_lut_4_lut.init = 16'hf011;
    L6MUX21 i21850 (.D0(n24339), .D1(n24340), .SD(index_i[6]), .Z(n24351));
    L6MUX21 i22285 (.D0(n24784), .D1(n24785), .SD(index_i[6]), .Z(n382));
    LUT4 mux_206_Mux_4_i653_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n653_adj_3039)) /* synthesis lut_function=(A (B (D)+!B (C (D)+!C !(D)))+!A !(D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_4_i653_3_lut_4_lut_4_lut_4_lut.init = 16'ha857;
    LUT4 i20857_3_lut_3_lut_4_lut (.A(n29165), .B(index_q[3]), .C(n93_adj_3443), 
         .D(index_q[4]), .Z(n23339)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i20857_3_lut_3_lut_4_lut.init = 16'h11f0;
    LUT4 mux_206_Mux_4_i542_3_lut (.A(n526), .B(n541_adj_3381), .C(index_i[4]), 
         .Z(n542_adj_3199)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_4_i542_3_lut.init = 16'hcaca;
    L6MUX21 i21852 (.D0(n24343), .D1(n24344), .SD(index_i[6]), .Z(n24353));
    L6MUX21 i21877 (.D0(n24362), .D1(n24363), .SD(index_i[6]), .Z(n24378));
    L6MUX21 i21878 (.D0(n24364), .D1(n24365), .SD(index_i[6]), .Z(n24379));
    LUT4 i24496_2_lut_rep_774 (.A(index_i[0]), .B(index_i[1]), .Z(n29434)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i24496_2_lut_rep_774.init = 16'h9999;
    L6MUX21 i21879 (.D0(n24366), .D1(n24367), .SD(index_i[6]), .Z(n24380));
    PFUMX i21880 (.BLUT(n24368), .ALUT(n24369), .C0(index_i[6]), .Z(n24381));
    LUT4 i14218_3_lut (.A(index_q[3]), .B(index_q[1]), .C(index_q[0]), 
         .Z(n16637)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i14218_3_lut.init = 16'hecec;
    PFUMX i21881 (.BLUT(n24370), .ALUT(n24371), .C0(index_i[6]), .Z(n24382));
    L6MUX21 i21882 (.D0(n24372), .D1(n24373), .SD(index_i[6]), .Z(n24383));
    L6MUX21 i21883 (.D0(n24374), .D1(n24375), .SD(index_i[6]), .Z(n24384));
    PFUMX i21884 (.BLUT(n24376), .ALUT(n24377), .C0(index_i[6]), .Z(n24385));
    LUT4 mux_206_Mux_5_i889_3_lut_rep_725 (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[2]), .Z(n29385)) /* synthesis lut_function=(A (B+!(C))+!A !((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_5_i889_3_lut_rep_725.init = 16'h8e8e;
    LUT4 i20622_3_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[0]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n23104)) /* synthesis lut_function=(!(A (B (D)+!B !(C+!(D)))+!A !(B (C (D))+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20622_3_lut_3_lut_4_lut.init = 16'h71aa;
    L6MUX21 i22721 (.D0(n23319), .D1(n23322), .SD(index_q[6]), .Z(n25222));
    PFUMX i21904 (.BLUT(n797_adj_3408), .ALUT(n828_adj_3249), .C0(index_i[5]), 
          .Z(n24405));
    LUT4 i13012_2_lut_rep_486_3_lut (.A(index_i[2]), .B(index_i[3]), .C(index_i[1]), 
         .Z(n29146)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i13012_2_lut_rep_486_3_lut.init = 16'h8080;
    LUT4 i21870_4_lut (.A(n29148), .B(n27388), .C(index_i[5]), .D(index_i[4]), 
         .Z(n24371)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam i21870_4_lut.init = 16'hc5ca;
    LUT4 mux_207_Mux_2_i397_3_lut (.A(n32055), .B(n29460), .C(index_q[3]), 
         .Z(n397_adj_3184)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_2_i397_3_lut.init = 16'hcaca;
    L6MUX21 i21908 (.D0(n24393), .D1(n24394), .SD(index_i[6]), .Z(n24409));
    L6MUX21 i21909 (.D0(n24395), .D1(n24396), .SD(index_i[6]), .Z(n24410));
    L6MUX21 i21910 (.D0(n24397), .D1(n24398), .SD(index_i[6]), .Z(n24411));
    L6MUX21 i21911 (.D0(n24399), .D1(n24400), .SD(index_i[6]), .Z(n24412));
    L6MUX21 i21912 (.D0(n24401), .D1(n24402), .SD(index_i[6]), .Z(n24413));
    L6MUX21 i21915 (.D0(n24407), .D1(n24408), .SD(index_i[6]), .Z(n24416));
    L6MUX21 i22328 (.D0(n23868), .D1(n23871), .SD(index_i[6]), .Z(n24829));
    PFUMX i22329 (.BLUT(n13520), .ALUT(n23874), .C0(index_i[6]), .Z(n24830));
    LUT4 i12518_2_lut_rep_429_3_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n29089)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12518_2_lut_rep_429_3_lut_4_lut.init = 16'hf080;
    LUT4 n124_bdd_3_lut_4_lut_adj_188 (.A(n29165), .B(index_q[3]), .C(index_q[4]), 
         .D(n93_adj_3443), .Z(n28489)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam n124_bdd_3_lut_4_lut_adj_188.init = 16'hfe0e;
    L6MUX21 i22331 (.D0(n23880), .D1(n23883), .SD(index_i[6]), .Z(n24832));
    L6MUX21 i22332 (.D0(n574_adj_2971), .D1(n23886), .SD(index_i[6]), 
            .Z(n24833));
    L6MUX21 i22333 (.D0(n23889), .D1(n764_adj_2966), .SD(index_i[6]), 
            .Z(n24834));
    LUT4 i11041_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n541_adj_3058)) /* synthesis lut_function=(A (B (C (D))+!B !(C (D)))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11041_3_lut_4_lut_4_lut_4_lut.init = 16'h9333;
    LUT4 mux_207_Mux_4_i828_3_lut_4_lut (.A(index_q[4]), .B(index_q[3]), 
         .C(n812_adj_3405), .D(n29354), .Z(n828_adj_3349)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_4_i828_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i21868_3_lut (.A(n476_adj_3244), .B(n507_adj_3171), .C(index_i[5]), 
         .Z(n24369)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21868_3_lut.init = 16'hcaca;
    L6MUX21 i21940 (.D0(n24426), .D1(n24427), .SD(index_i[6]), .Z(n24441));
    L6MUX21 i21941 (.D0(n24428), .D1(n24429), .SD(index_i[6]), .Z(n24442));
    LUT4 index_i_6__bdd_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), .C(n29376), 
         .D(index_i[6]), .Z(n28577)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(D))+!A !(D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam index_i_6__bdd_3_lut_4_lut.init = 16'h887f;
    PFUMX i26279 (.BLUT(n28140), .ALUT(n28139), .C0(index_q[3]), .Z(n28141));
    LUT4 i13850_2_lut_2_lut_3_lut (.A(index_i[2]), .B(index_i[3]), .C(index_i[0]), 
         .Z(n16259)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i13850_2_lut_2_lut_3_lut.init = 16'h0808;
    L6MUX21 i21942 (.D0(n24430), .D1(n24431), .SD(index_i[6]), .Z(n24443));
    LUT4 i21498_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n23980)) /* synthesis lut_function=(!(A (B)+!A (B (C+(D))+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i21498_3_lut_3_lut_4_lut.init = 16'h3326;
    LUT4 i12864_2_lut_rep_409_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[4]), .D(n29376), .Z(n29069)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12864_2_lut_rep_409_3_lut_4_lut.init = 16'hf8f0;
    L6MUX21 i21943 (.D0(n24432), .D1(n24433), .SD(index_i[6]), .Z(n24444));
    L6MUX21 i21944 (.D0(n24434), .D1(n24435), .SD(index_i[6]), .Z(n24445));
    LUT4 mux_207_Mux_7_i891_3_lut_4_lut (.A(n29165), .B(index_q[3]), .C(index_q[4]), 
         .D(n890_adj_3123), .Z(n891_adj_3418)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_7_i891_3_lut_4_lut.init = 16'hfe0e;
    LUT4 i14494_3_lut_4_lut (.A(n29165), .B(index_q[3]), .C(n9850), .D(index_q[6]), 
         .Z(n16930)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i14494_3_lut_4_lut.init = 16'hffe0;
    LUT4 i21817_1_lut_2_lut (.A(index_i[2]), .B(index_i[3]), .Z(n24318)) /* synthesis lut_function=(!(A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21817_1_lut_2_lut.init = 16'h7777;
    LUT4 mux_206_Mux_4_i286_3_lut (.A(n270_adj_3315), .B(n15_adj_3125), 
         .C(index_i[4]), .Z(n286)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_4_i286_3_lut.init = 16'hcaca;
    LUT4 mux_206_Mux_0_i698_3_lut_rep_817 (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[2]), .Z(n32018)) /* synthesis lut_function=(!(A (C)+!A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i698_3_lut_rep_817.init = 16'h1a1a;
    PFUMX i26255 (.BLUT(n28109), .ALUT(n28107), .C0(index_i[7]), .Z(n28110));
    LUT4 i20736_3_lut (.A(n29429), .B(n29424), .C(index_i[3]), .Z(n23218)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20736_3_lut.init = 16'hcaca;
    L6MUX21 i25096 (.D0(n26745), .D1(n26742), .SD(index_i[5]), .Z(n26746));
    L6MUX21 i21961 (.D0(n24814), .D1(n24821), .SD(index_q[6]), .Z(n24462));
    L6MUX21 i21964 (.D0(n23346), .D1(n23349), .SD(index_q[6]), .Z(n24465));
    L6MUX21 i21965 (.D0(n23352), .D1(n23355), .SD(index_q[6]), .Z(n24466));
    L6MUX21 i21966 (.D0(n23730), .D1(n23811), .SD(index_q[6]), .Z(n24467));
    PFUMX i21967 (.BLUT(n23817), .ALUT(n892_adj_3419), .C0(index_q[6]), 
          .Z(n24468));
    LUT4 i17688_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n20002)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i17688_3_lut_4_lut_4_lut_4_lut.init = 16'h3999;
    LUT4 i14466_2_lut_rep_414_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[4]), .D(n29379), .Z(n29074)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i14466_2_lut_rep_414_3_lut_4_lut.init = 16'hf8f0;
    LUT4 mux_206_Mux_7_i924_3_lut_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[4]), .D(n29379), .Z(n924_adj_3444)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_7_i924_3_lut_3_lut_4_lut.init = 16'h878f;
    LUT4 mux_206_Mux_2_i604_3_lut_4_lut_4_lut_4_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n604_adj_3428)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)+!C !(D)))+!A (B (C)+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_2_i604_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'h3c9f;
    LUT4 mux_206_Mux_1_i890_4_lut_4_lut_4_lut_4_lut (.A(index_i[3]), .B(index_i[4]), 
         .C(n645), .D(index_i[0]), .Z(n890_adj_3379)) /* synthesis lut_function=(!(A (B (D)+!B !(C))+!A (B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_1_i890_4_lut_4_lut_4_lut_4_lut.init = 16'h31fd;
    LUT4 i13899_3_lut_3_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n16308)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (D))+!A (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i13899_3_lut_3_lut_3_lut_4_lut.init = 16'h00f7;
    PFUMX i22561 (.BLUT(n286_adj_3194), .ALUT(n317_adj_3192), .C0(index_q[5]), 
          .Z(n25062));
    LUT4 i25647_then_4_lut (.A(index_i[1]), .B(index_i[5]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n29586)) /* synthesis lut_function=(A (B (C)+!B !(C+!(D)))+!A (B (C+(D))+!B !(C (D)))) */ ;
    defparam i25647_then_4_lut.init = 16'hc7d1;
    LUT4 mux_206_Mux_6_i924_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[4]), .D(n908), .Z(n924_adj_3445)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_6_i924_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_206_Mux_4_i94_3_lut (.A(n61), .B(n29319), .C(index_i[4]), 
         .Z(n94_adj_3030)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_4_i94_3_lut.init = 16'hcaca;
    PFUMX i21987 (.BLUT(n732_adj_3196), .ALUT(n763_adj_3398), .C0(index_i[5]), 
          .Z(n24488));
    L6MUX21 i22359 (.D0(n24844), .D1(n24845), .SD(index_q[6]), .Z(n24860));
    L6MUX21 i21989 (.D0(n23934), .D1(n891_adj_3380), .SD(index_i[5]), 
            .Z(n24490));
    L6MUX21 i21992 (.D0(n24477), .D1(n24478), .SD(index_i[6]), .Z(n24493));
    LUT4 mux_206_Mux_0_i699_3_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n699_adj_3446)) /* synthesis lut_function=(!(A (C+!(D))+!A (B (D)+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i699_3_lut_3_lut_4_lut.init = 16'h1a55;
    L6MUX21 i22360 (.D0(n24846), .D1(n24847), .SD(index_q[6]), .Z(n24861));
    PFUMX i22562 (.BLUT(n349_adj_2994), .ALUT(n23361), .C0(index_q[5]), 
          .Z(n25063));
    LUT4 i12884_3_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[3]), 
         .Z(n12338)) /* synthesis lut_function=(!((B (C))+!A)) */ ;
    defparam i12884_3_lut.init = 16'h2a2a;
    LUT4 mux_206_Mux_5_i109_3_lut_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .Z(n109_adj_3447)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_5_i109_3_lut_3_lut_3_lut.init = 16'h3939;
    PFUMX i22563 (.BLUT(n413_adj_3185), .ALUT(n23358), .C0(index_q[5]), 
          .Z(n25064));
    PFUMX i26253 (.BLUT(n28104), .ALUT(n28100), .C0(index_i[4]), .Z(n28105));
    LUT4 mux_207_Mux_5_i797_3_lut_4_lut (.A(index_q[4]), .B(index_q[3]), 
         .C(n29505), .D(n29389), .Z(n797_adj_3289)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_5_i797_3_lut_4_lut.init = 16'hf1e0;
    L6MUX21 i21994 (.D0(n24481), .D1(n24482), .SD(index_i[6]), .Z(n24495));
    L6MUX21 i21995 (.D0(n24483), .D1(n24484), .SD(index_i[6]), .Z(n24496));
    LUT4 mux_206_Mux_1_i987_3_lut_4_lut_4_lut (.A(index_i[3]), .B(n986_adj_3397), 
         .C(index_i[4]), .D(n29406), .Z(n987)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_1_i987_3_lut_4_lut_4_lut.init = 16'hc5c0;
    LUT4 i10323_4_lut_4_lut (.A(index_i[3]), .B(index_i[0]), .C(index_i[1]), 
         .D(index_i[2]), .Z(n12581)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (D)+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i10323_4_lut_4_lut.init = 16'h0bf4;
    LUT4 i12455_4_lut_4_lut (.A(index_i[3]), .B(index_i[2]), .C(index_i[0]), 
         .D(index_i[1]), .Z(n875_adj_3448)) /* synthesis lut_function=((B (C)+!B (D))+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12455_4_lut_4_lut.init = 16'hf7d5;
    L6MUX21 i22361 (.D0(n24848), .D1(n24849), .SD(index_q[6]), .Z(n24862));
    L6MUX21 i22362 (.D0(n24850), .D1(n24851), .SD(index_q[6]), .Z(n24863));
    PFUMX i26250 (.BLUT(n28101), .ALUT(n29318), .C0(index_i[3]), .Z(n28102));
    L6MUX21 i26237 (.D0(n28083), .D1(n29031), .SD(index_q[6]), .Z(n28084));
    PFUMX i26235 (.BLUT(n28082), .ALUT(n29045), .C0(index_q[7]), .Z(n28083));
    LUT4 i21430_4_lut_3_lut (.A(index_i[3]), .B(index_i[4]), .C(n29177), 
         .Z(n23912)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21430_4_lut_3_lut.init = 16'h6565;
    PFUMX i26230 (.BLUT(n28076), .ALUT(n28073), .C0(index_i[6]), .Z(n28077));
    LUT4 mux_206_Mux_2_i221_4_lut_4_lut (.A(index_i[3]), .B(index_i[4]), 
         .C(n29177), .D(n29089), .Z(n221_adj_3128)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (B+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_2_i221_4_lut_4_lut.init = 16'hf7c4;
    L6MUX21 i22363 (.D0(n24852), .D1(n24853), .SD(index_q[6]), .Z(n24864));
    L6MUX21 i22365 (.D0(n24856), .D1(n24857), .SD(index_q[6]), .Z(n24866));
    L6MUX21 i21999 (.D0(n24491), .D1(n24492), .SD(index_i[6]), .Z(n24500));
    PFUMX i22018 (.BLUT(n732_adj_3179), .ALUT(n763), .C0(index_q[5]), 
          .Z(n24519));
    L6MUX21 i22020 (.D0(n23424), .D1(n891_adj_3353), .SD(index_q[5]), 
            .Z(n24521));
    L6MUX21 i22390 (.D0(n24875), .D1(n24876), .SD(index_q[6]), .Z(n24891));
    L6MUX21 i22391 (.D0(n24877), .D1(n24878), .SD(index_q[6]), .Z(n24892));
    L6MUX21 i22023 (.D0(n24508), .D1(n24509), .SD(index_q[6]), .Z(n24524));
    L6MUX21 i22025 (.D0(n24512), .D1(n24513), .SD(index_q[6]), .Z(n24526));
    L6MUX21 i22026 (.D0(n24514), .D1(n24515), .SD(index_q[6]), .Z(n24527));
    L6MUX21 i22392 (.D0(n24879), .D1(n24880), .SD(index_q[6]), .Z(n24893));
    PFUMX i26228 (.BLUT(n28074), .ALUT(n954_adj_3431), .C0(index_i[4]), 
          .Z(n28075));
    PFUMX i22393 (.BLUT(n24881), .ALUT(n24882), .C0(index_q[6]), .Z(n24894));
    L6MUX21 i22030 (.D0(n24522), .D1(n24523), .SD(index_q[6]), .Z(n24531));
    PFUMX i22394 (.BLUT(n24883), .ALUT(n24884), .C0(index_q[6]), .Z(n24895));
    LUT4 i20745_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n23227)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !(B (C+!(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20745_3_lut_4_lut_4_lut.init = 16'ha5a9;
    L6MUX21 i22395 (.D0(n24885), .D1(n24886), .SD(index_q[6]), .Z(n24896));
    LUT4 i11233_3_lut_3_lut (.A(index_i[3]), .B(index_i[4]), .C(n13529), 
         .Z(n13530)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11233_3_lut_3_lut.init = 16'h7474;
    L6MUX21 i22396 (.D0(n24887), .D1(n24888), .SD(index_q[6]), .Z(n24897));
    PFUMX i22397 (.BLUT(n24889), .ALUT(n24890), .C0(index_q[6]), .Z(n24898));
    LUT4 i12575_2_lut_2_lut_3_lut (.A(index_i[1]), .B(index_i[0]), .C(index_i[3]), 
         .Z(n14983)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12575_2_lut_2_lut_3_lut.init = 16'h0808;
    LUT4 i12444_2_lut_rep_670 (.A(index_q[0]), .B(index_q[1]), .Z(n29330)) /* synthesis lut_function=((B)+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i12444_2_lut_rep_670.init = 16'hdddd;
    PFUMX i22564 (.BLUT(n23370), .ALUT(n507_adj_3372), .C0(index_q[5]), 
          .Z(n25065));
    LUT4 mux_207_Mux_6_i668_3_lut (.A(n108), .B(n29472), .C(index_q[3]), 
         .Z(n668_adj_3079)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_6_i668_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_6_i684_3_lut (.A(n29181), .B(n32055), .C(index_q[3]), 
         .Z(n684_adj_3207)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_6_i684_3_lut.init = 16'hcaca;
    LUT4 i25647_else_4_lut (.A(index_i[1]), .B(index_i[5]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n29585)) /* synthesis lut_function=(A (B (C)+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B (D))) */ ;
    defparam i25647_else_4_lut.init = 16'h86f1;
    LUT4 n122_bdd_3_lut_25962_4_lut_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .Z(n26658)) /* synthesis lut_function=(A (B)+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam n122_bdd_3_lut_25962_4_lut_3_lut.init = 16'hd9d9;
    LUT4 i20697_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n23179)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (D))+!A !(D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i20697_3_lut_4_lut_4_lut_4_lut.init = 16'ha25d;
    PFUMX i22637 (.BLUT(n25134), .ALUT(n25135), .C0(index_i[4]), .Z(n25138));
    LUT4 mux_207_Mux_0_i635_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n635_adj_3449)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_0_i635_3_lut_4_lut_4_lut.init = 16'hfd0a;
    PFUMX i22565 (.BLUT(n23373), .ALUT(n573_adj_3015), .C0(index_q[5]), 
          .Z(n25066));
    LUT4 mux_207_Mux_0_i316_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n316_adj_3334)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+(D)))+!A (B (C+(D))+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_0_i316_3_lut_4_lut_4_lut_4_lut.init = 16'h332d;
    PFUMX i22638 (.BLUT(n25136), .ALUT(n25137), .C0(index_i[4]), .Z(n25139));
    LUT4 mux_207_Mux_6_i564_3_lut_4_lut_3_lut_rep_671 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29331)) /* synthesis lut_function=(A (B)+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_6_i564_3_lut_4_lut_3_lut_rep_671.init = 16'hd9d9;
    PFUMX i22566 (.BLUT(n605_adj_3169), .ALUT(n23376), .C0(index_q[5]), 
          .Z(n25067));
    LUT4 mux_207_Mux_0_i627_3_lut_rep_673 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29333)) /* synthesis lut_function=(A (B+!(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_0_i627_3_lut_rep_673.init = 16'hdada;
    LUT4 mux_206_Mux_5_i891_3_lut (.A(n875_adj_3306), .B(n27184), .C(index_i[4]), 
         .Z(n891)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_5_i891_3_lut.init = 16'hcaca;
    LUT4 i20685_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n23167)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i20685_3_lut_4_lut_4_lut.init = 16'hda5a;
    PFUMX i22567 (.BLUT(n669_adj_3166), .ALUT(n700_adj_3101), .C0(index_q[5]), 
          .Z(n25068));
    LUT4 i12466_2_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n668_adj_3450)) /* synthesis lut_function=(!(A ((D)+!B)+!A (B ((D)+!C)+!B (C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12466_2_lut_4_lut_4_lut_4_lut.init = 16'h00c9;
    LUT4 mux_206_Mux_5_i860_3_lut (.A(n15_adj_3279), .B(n859_adj_3305), 
         .C(index_i[4]), .Z(n860_adj_3022)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_5_i860_3_lut.init = 16'hcaca;
    LUT4 i20929_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n23411)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C))+!A !(B (C)+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i20929_3_lut_4_lut_4_lut.init = 16'h5ad3;
    LUT4 i17687_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n20001)) /* synthesis lut_function=(A (B)+!A !(B (C (D))+!B !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i17687_3_lut_4_lut_4_lut.init = 16'h9ccc;
    LUT4 i12890_3_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .Z(n12265)) /* synthesis lut_function=(!((B (C))+!A)) */ ;
    defparam i12890_3_lut.init = 16'h2a2a;
    LUT4 i20907_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n23389)) /* synthesis lut_function=(!(A (B (C (D))+!B (C (D)+!C !(D)))+!A !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i20907_3_lut_4_lut_4_lut.init = 16'h5aad;
    PFUMX i22568 (.BLUT(n732_adj_3162), .ALUT(n763_adj_3359), .C0(index_q[5]), 
          .Z(n25069));
    LUT4 i1_2_lut_rep_483_3_lut_4_lut (.A(index_i[1]), .B(index_i[0]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n29143)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_2_lut_rep_483_3_lut_4_lut.init = 16'h8000;
    LUT4 n773_bdd_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n26640)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam n773_bdd_3_lut_4_lut_4_lut.init = 16'ha5ad;
    LUT4 mux_206_Mux_6_i573_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[4]), .D(n572_adj_3451), .Z(n573_adj_3452)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_6_i573_3_lut_4_lut.init = 16'hf909;
    PFUMX i22645 (.BLUT(n25143), .ALUT(n25144), .C0(index_i[4]), .Z(n25146));
    LUT4 mux_207_Mux_6_i645_3_lut_4_lut_3_lut_rep_804 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29464)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B))) */ ;
    defparam mux_207_Mux_6_i645_3_lut_4_lut_3_lut_rep_804.init = 16'h1919;
    PFUMX i25094 (.BLUT(n26744), .ALUT(n475_adj_3009), .C0(index_i[4]), 
          .Z(n26745));
    LUT4 mux_207_Mux_6_i572_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n572_adj_3413)) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_6_i572_3_lut_4_lut.init = 16'hccd9;
    LUT4 i12783_2_lut_rep_674 (.A(index_q[0]), .B(index_q[1]), .Z(n29334)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i12783_2_lut_rep_674.init = 16'h2222;
    L6MUX21 i22570 (.D0(n860_adj_3291), .D1(n891_adj_3286), .SD(index_q[5]), 
            .Z(n25071));
    LUT4 mux_207_Mux_0_i985_3_lut_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n985_adj_3282)) /* synthesis lut_function=(!(A (B+!(C))+!A (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_0_i985_3_lut_3_lut.init = 16'h2525;
    L6MUX21 i26164 (.D0(n27980), .D1(n27978), .SD(index_q[8]), .Z(n27981));
    PFUMX i26162 (.BLUT(n27979), .ALUT(n25208), .C0(index_q[7]), .Z(n27980));
    PFUMX i27109 (.BLUT(n29536), .ALUT(n29537), .C0(index_q[3]), .Z(n29538));
    LUT4 i23963_3_lut (.A(n23995), .B(n23996), .C(index_i[4]), .Z(n23997)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23963_3_lut.init = 16'hcaca;
    PFUMX i20696 (.BLUT(n23176), .ALUT(n23177), .C0(index_q[4]), .Z(n23178));
    L6MUX21 i22594 (.D0(n25093), .D1(n25094), .SD(index_i[5]), .Z(n25095));
    LUT4 i24742_2_lut_rep_485_3_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n29145)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i24742_2_lut_rep_485_3_lut_4_lut.init = 16'h0007;
    LUT4 mux_206_Mux_5_i636_4_lut (.A(n157_adj_3453), .B(n29186), .C(index_i[4]), 
         .D(index_i[3]), .Z(n636)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_5_i636_4_lut.init = 16'h3aca;
    PFUMX i26160 (.BLUT(n27977), .ALUT(n27976), .C0(index_q[7]), .Z(n27978));
    LUT4 i23966_3_lut (.A(n20015), .B(n20016), .C(index_i[4]), .Z(n20017)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23966_3_lut.init = 16'hcaca;
    LUT4 mux_206_Mux_8_i526_3_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n526_adj_3005)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_8_i526_3_lut_3_lut_4_lut.init = 16'h0f70;
    LUT4 i12456_2_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n844_adj_3454)) /* synthesis lut_function=(A (B+!(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12456_2_lut_3_lut_4_lut.init = 16'h9ff9;
    LUT4 mux_207_Mux_4_i205_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n205)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_4_i205_3_lut_4_lut_4_lut.init = 16'h5a2a;
    LUT4 mux_207_Mux_0_i165_3_lut_4_lut_3_lut_rep_675 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29335)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_0_i165_3_lut_4_lut_3_lut_rep_675.init = 16'h9292;
    PFUMX i22007 (.BLUT(n13445), .ALUT(n62_adj_3404), .C0(index_q[5]), 
          .Z(n24508));
    LUT4 mux_207_Mux_6_i70_3_lut_rep_676 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29336)) /* synthesis lut_function=(!(A (B+(C))+!A !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_6_i70_3_lut_rep_676.init = 16'h5252;
    LUT4 mux_207_Mux_2_i348_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n348_adj_2993)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_2_i348_3_lut_4_lut_4_lut.init = 16'h52a5;
    L6MUX21 i26114 (.D0(n27926), .D1(n27923), .SD(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_1783[4]));
    PFUMX i26112 (.BLUT(n27925), .ALUT(n27924), .C0(index_q[8]), .Z(n27926));
    LUT4 i20694_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n23176)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C))+!A !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i20694_3_lut_4_lut_4_lut.init = 16'h5a52;
    LUT4 n316_bdd_3_lut_26868_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n27745)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A !(B ((D)+!C)+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam n316_bdd_3_lut_26868_3_lut_4_lut.init = 16'h552c;
    PFUMX i26109 (.BLUT(n27922), .ALUT(n24902), .C0(index_q[8]), .Z(n27923));
    LUT4 mux_206_Mux_6_i668_3_lut (.A(n660), .B(n29384), .C(index_i[3]), 
         .Z(n668_adj_3048)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_6_i668_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_0_i812_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n812_adj_3023)) /* synthesis lut_function=(A (B (C+(D))+!B !(C))+!A (B (D)+!B !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_0_i812_3_lut_4_lut_4_lut_4_lut.init = 16'hcf92;
    L6MUX21 i26091 (.D0(n27901), .D1(n27898), .SD(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_1783[9]));
    PFUMX i26089 (.BLUT(n27900), .ALUT(n27899), .C0(index_q[8]), .Z(n27901));
    LUT4 i20877_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n23359)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C))+!A !(B ((D)+!C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i20877_3_lut_4_lut_4_lut.init = 16'h925a;
    LUT4 mux_206_Mux_6_i684_3_lut (.A(n645), .B(n32039), .C(index_i[3]), 
         .Z(n684_adj_3188)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_6_i684_3_lut.init = 16'hcaca;
    PFUMX i21976 (.BLUT(n13404), .ALUT(n62_adj_3455), .C0(index_i[5]), 
          .Z(n24477));
    LUT4 mux_206_Mux_5_i507_3_lut (.A(n491_adj_3195), .B(n506_adj_3292), 
         .C(index_i[4]), .Z(n507_adj_3008)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_5_i507_3_lut.init = 16'hcaca;
    PFUMX i22484 (.BLUT(n333), .ALUT(n348_adj_3114), .C0(index_q[4]), 
          .Z(n24985));
    LUT4 mux_206_Mux_5_i476_3_lut (.A(n460_adj_3355), .B(n475_adj_3456), 
         .C(index_i[4]), .Z(n476_adj_3007)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_5_i476_3_lut.init = 16'hcaca;
    PFUMX i21892 (.BLUT(n31_adj_3137), .ALUT(n62_adj_2947), .C0(index_i[5]), 
          .Z(n24393));
    PFUMX i22485 (.BLUT(n364_adj_3457), .ALUT(n379_adj_2970), .C0(index_q[4]), 
          .Z(n24986));
    PFUMX i26086 (.BLUT(n27897), .ALUT(n24458), .C0(index_q[8]), .Z(n27898));
    L6MUX21 i26073 (.D0(n27880), .D1(n27877), .SD(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_1768[4]));
    PFUMX i22486 (.BLUT(n397), .ALUT(n412_adj_2986), .C0(index_q[4]), 
          .Z(n24987));
    PFUMX i26071 (.BLUT(n27879), .ALUT(n27878), .C0(index_i[8]), .Z(n27880));
    LUT4 mux_207_Mux_5_i460_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n460_adj_3392)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A !(B (C)+!B !(C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_5_i460_3_lut_4_lut_4_lut.init = 16'h6b5a;
    LUT4 i24465_3_lut_4_lut (.A(n29102), .B(n29250), .C(index_q[8]), .D(n766_adj_3229), 
         .Z(n23210)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i24465_3_lut_4_lut.init = 16'hefe0;
    PFUMX i26068 (.BLUT(n27876), .ALUT(n24389), .C0(index_i[8]), .Z(n27877));
    PFUMX i21861 (.BLUT(n31_adj_3126), .ALUT(n62_adj_3124), .C0(index_i[5]), 
          .Z(n24362));
    L6MUX21 i26058 (.D0(n27864), .D1(n27861), .SD(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_1768[9]));
    PFUMX i26056 (.BLUT(n27863), .ALUT(n27862), .C0(index_i[8]), .Z(n27864));
    PFUMX i27107 (.BLUT(n29533), .ALUT(n29534), .C0(index_i[3]), .Z(n62_adj_3366));
    PFUMX i20699 (.BLUT(n23179), .ALUT(n23180), .C0(index_q[4]), .Z(n23181));
    L6MUX21 i22601 (.D0(n25100), .D1(n25101), .SD(index_i[5]), .Z(n25102));
    LUT4 mux_206_Mux_5_i413_3_lut (.A(n397_adj_3288), .B(n251_adj_3064), 
         .C(index_i[4]), .Z(n413)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_5_i413_3_lut.init = 16'hcaca;
    LUT4 n133_bdd_3_lut_25946_4_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .Z(n26752)) /* synthesis lut_function=(A (B)+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n133_bdd_3_lut_25946_4_lut_3_lut.init = 16'hd9d9;
    PFUMX i22487 (.BLUT(n428), .ALUT(n443_adj_2951), .C0(index_q[4]), 
          .Z(n24988));
    PFUMX i25091 (.BLUT(n26741), .ALUT(n23945), .C0(index_i[4]), .Z(n26742));
    LUT4 mux_206_Mux_6_i498_3_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n498)) /* synthesis lut_function=(A (B+!(C))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_6_i498_3_lut_4_lut_3_lut.init = 16'h9b9b;
    LUT4 mux_206_Mux_8_i635_3_lut_4_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n635_adj_3004)) /* synthesis lut_function=(!(A (B (C (D))+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_8_i635_3_lut_4_lut_3_lut_4_lut.init = 16'h0ff8;
    LUT4 i22317_3_lut (.A(n29316), .B(n29470), .C(index_q[3]), .Z(n24818)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22317_3_lut.init = 16'hcaca;
    LUT4 i17689_3_lut (.A(n20001), .B(n20002), .C(index_i[4]), .Z(n20003)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17689_3_lut.init = 16'hcaca;
    LUT4 i11069_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(n29329), .D(index_i[4]), .Z(n189)) /* synthesis lut_function=(A (B (C (D)))+!A !(B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11069_3_lut_4_lut_4_lut_4_lut.init = 16'h9555;
    PFUMX i26053 (.BLUT(n27860), .ALUT(n24719), .C0(index_i[8]), .Z(n27861));
    LUT4 mux_206_Mux_5_i572_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n572_adj_3430)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A !(B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_5_i572_3_lut_4_lut_4_lut.init = 16'ha9a5;
    LUT4 mux_206_Mux_5_i125_3_lut (.A(n109_adj_3447), .B(n124_adj_3281), 
         .C(index_i[4]), .Z(n125)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_5_i125_3_lut.init = 16'hcaca;
    LUT4 mux_206_Mux_5_i94_3_lut (.A(n653_adj_3047), .B(n635_adj_3441), 
         .C(index_i[4]), .Z(n94_adj_2996)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_5_i94_3_lut.init = 16'hcaca;
    LUT4 i22236_3_lut (.A(n24735), .B(n24736), .C(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_1768[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22236_3_lut.init = 16'hcaca;
    PFUMX i26039 (.BLUT(n27842), .ALUT(n1022_adj_3234), .C0(index_q[9]), 
          .Z(quarter_wave_sample_register_q_15__N_1783[12]));
    LUT4 i22811_3_lut (.A(n25310), .B(n25311), .C(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_1768[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22811_3_lut.init = 16'hcaca;
    LUT4 i22810_3_lut (.A(n25308), .B(n25309), .C(index_i[8]), .Z(n25311)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22810_3_lut.init = 16'hcaca;
    LUT4 mux_206_Mux_6_i812_3_lut_4_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n812)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(D))+!A !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_6_i812_3_lut_4_lut_3_lut_4_lut.init = 16'h7780;
    LUT4 mux_160_i16_3_lut (.A(\quarter_wave_sample_register_i[15] ), .B(o_val_pipeline_i_0__15__N_1799[15]), 
         .C(phase_negation_i[1]), .Z(n670[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam mux_160_i16_3_lut.init = 16'hcaca;
    LUT4 i20650_3_lut (.A(n900_adj_3319), .B(n325), .C(index_q[3]), .Z(n23132)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20650_3_lut.init = 16'hcaca;
    LUT4 mux_160_i15_3_lut (.A(quarter_wave_sample_register_i[14]), .B(o_val_pipeline_i_0__15__N_1799[14]), 
         .C(phase_negation_i[1]), .Z(n670[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam mux_160_i15_3_lut.init = 16'hcaca;
    PFUMX i26035 (.BLUT(n254_adj_3458), .ALUT(n27836), .C0(index_q[8]), 
          .Z(n27837));
    LUT4 mux_160_i14_3_lut (.A(quarter_wave_sample_register_i[13]), .B(o_val_pipeline_i_0__15__N_1799[13]), 
         .C(phase_negation_i[1]), .Z(n670[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam mux_160_i14_3_lut.init = 16'hcaca;
    LUT4 mux_206_Mux_5_i31_3_lut (.A(n15_adj_3279), .B(n30_adj_3440), .C(index_i[4]), 
         .Z(n31)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_5_i31_3_lut.init = 16'hcaca;
    LUT4 mux_160_i13_3_lut (.A(quarter_wave_sample_register_i[12]), .B(o_val_pipeline_i_0__15__N_1799[12]), 
         .C(phase_negation_i[1]), .Z(n670[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam mux_160_i13_3_lut.init = 16'hcaca;
    LUT4 mux_160_i12_3_lut (.A(quarter_wave_sample_register_i[11]), .B(o_val_pipeline_i_0__15__N_1799[11]), 
         .C(phase_negation_i[1]), .Z(n670[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam mux_160_i12_3_lut.init = 16'hcaca;
    LUT4 mux_160_i11_3_lut (.A(quarter_wave_sample_register_i[10]), .B(o_val_pipeline_i_0__15__N_1799[10]), 
         .C(phase_negation_i[1]), .Z(n670[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam mux_160_i11_3_lut.init = 16'hcaca;
    LUT4 mux_160_i10_3_lut (.A(quarter_wave_sample_register_i[9]), .B(o_val_pipeline_i_0__15__N_1799[9]), 
         .C(phase_negation_i[1]), .Z(n670[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam mux_160_i10_3_lut.init = 16'hcaca;
    LUT4 mux_206_Mux_2_i269_3_lut_3_lut_rep_747_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29407)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_2_i269_3_lut_3_lut_rep_747_3_lut.init = 16'h3939;
    LUT4 mux_160_i9_3_lut (.A(quarter_wave_sample_register_i[8]), .B(o_val_pipeline_i_0__15__N_1799[8]), 
         .C(phase_negation_i[1]), .Z(n670[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam mux_160_i9_3_lut.init = 16'hcaca;
    LUT4 mux_160_i8_3_lut (.A(quarter_wave_sample_register_i[7]), .B(o_val_pipeline_i_0__15__N_1799[7]), 
         .C(phase_negation_i[1]), .Z(n670[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam mux_160_i8_3_lut.init = 16'hcaca;
    LUT4 i20603_else_4_lut (.A(index_i[0]), .B(index_i[4]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n29515)) /* synthesis lut_function=(A (C)+!A !(B ((D)+!C)+!B !(C))) */ ;
    defparam i20603_else_4_lut.init = 16'hb0f0;
    LUT4 mux_160_i7_3_lut (.A(quarter_wave_sample_register_i[6]), .B(o_val_pipeline_i_0__15__N_1799[6]), 
         .C(phase_negation_i[1]), .Z(n670[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam mux_160_i7_3_lut.init = 16'hcaca;
    LUT4 mux_160_i6_3_lut (.A(quarter_wave_sample_register_i[5]), .B(o_val_pipeline_i_0__15__N_1799[5]), 
         .C(phase_negation_i[1]), .Z(n670[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam mux_160_i6_3_lut.init = 16'hcaca;
    LUT4 mux_160_i5_3_lut (.A(quarter_wave_sample_register_i[4]), .B(o_val_pipeline_i_0__15__N_1799[4]), 
         .C(phase_negation_i[1]), .Z(n670[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam mux_160_i5_3_lut.init = 16'hcaca;
    LUT4 mux_160_i4_3_lut (.A(quarter_wave_sample_register_i[3]), .B(o_val_pipeline_i_0__15__N_1799[3]), 
         .C(phase_negation_i[1]), .Z(n670[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam mux_160_i4_3_lut.init = 16'hcaca;
    LUT4 mux_160_i3_3_lut (.A(quarter_wave_sample_register_i[2]), .B(o_val_pipeline_i_0__15__N_1799[2]), 
         .C(phase_negation_i[1]), .Z(n670[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam mux_160_i3_3_lut.init = 16'hcaca;
    LUT4 mux_160_i2_3_lut (.A(quarter_wave_sample_register_i[1]), .B(o_val_pipeline_i_0__15__N_1799[1]), 
         .C(phase_negation_i[1]), .Z(n670[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam mux_160_i2_3_lut.init = 16'hcaca;
    LUT4 mux_160_i1_3_lut (.A(quarter_wave_sample_register_i[0]), .B(o_val_pipeline_i_0__15__N_1799[0]), 
         .C(phase_negation_i[1]), .Z(n670[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[29:60])
    defparam mux_160_i1_3_lut.init = 16'hcaca;
    PFUMX i22488 (.BLUT(n460_adj_2968), .ALUT(n475_adj_3459), .C0(index_q[4]), 
          .Z(n24989));
    LUT4 i12784_2_lut_rep_686 (.A(index_q[0]), .B(index_q[1]), .Z(n29346)) /* synthesis lut_function=(A+!(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i12784_2_lut_rep_686.init = 16'hbbbb;
    PFUMX i26016 (.BLUT(n27811), .ALUT(n1022), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_1768[12]));
    LUT4 i21975_3_lut (.A(n24474), .B(n24475), .C(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_1783[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21975_3_lut.init = 16'hcaca;
    LUT4 i22720_3_lut (.A(n27981), .B(n25220), .C(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_1783[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22720_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_6_i498_3_lut_4_lut_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n404)) /* synthesis lut_function=(A (B+!(C))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_6_i498_3_lut_4_lut_3_lut.init = 16'h9b9b;
    LUT4 i20893_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n23375)) /* synthesis lut_function=(A (C+(D))+!A !(B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i20893_3_lut_4_lut_4_lut.init = 16'haba5;
    LUT4 i22719_3_lut (.A(n25217), .B(n25218), .C(index_q[8]), .Z(n25220)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22719_3_lut.init = 16'hcaca;
    LUT4 i24514_2_lut (.A(phase_i[9]), .B(phase_i[10]), .Z(index_q_9__N_1758[9])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(60[14] 63[8])
    defparam i24514_2_lut.init = 16'h9999;
    LUT4 i24516_2_lut (.A(phase_i[8]), .B(phase_i[10]), .Z(index_q_9__N_1758[8])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(60[14] 63[8])
    defparam i24516_2_lut.init = 16'h9999;
    LUT4 n166_bdd_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n28802)) /* synthesis lut_function=(!(A (D)+!A !(B (D)+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam n166_bdd_4_lut_4_lut_4_lut.init = 16'h54bb;
    LUT4 i24518_2_lut (.A(phase_i[7]), .B(phase_i[10]), .Z(index_q_9__N_1758[7])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(60[14] 63[8])
    defparam i24518_2_lut.init = 16'h9999;
    LUT4 mux_207_Mux_6_i332_3_lut_3_lut_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n332)) /* synthesis lut_function=(!(A (C)+!A !((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_6_i332_3_lut_3_lut_3_lut.init = 16'h5b5b;
    LUT4 i24520_2_lut (.A(phase_i[6]), .B(phase_i[10]), .Z(index_q_9__N_1758[6])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(60[14] 63[8])
    defparam i24520_2_lut.init = 16'h9999;
    LUT4 mux_207_Mux_4_i900_3_lut_4_lut_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n900_adj_3319)) /* synthesis lut_function=(A ((C)+!B)+!A !(B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_4_i900_3_lut_4_lut_3_lut.init = 16'hb2b2;
    LUT4 i24522_2_lut (.A(phase_i[5]), .B(phase_i[10]), .Z(index_q_9__N_1758[5])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(60[14] 63[8])
    defparam i24522_2_lut.init = 16'h9999;
    PFUMX i26011 (.BLUT(n254_adj_3460), .ALUT(n27805), .C0(index_i[8]), 
          .Z(n27806));
    LUT4 i11145_3_lut_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n875_adj_3284)) /* synthesis lut_function=(A (C (D))+!A !(B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i11145_3_lut_3_lut_4_lut_4_lut.init = 16'hb555;
    LUT4 i20616_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n23098)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A !(B (C+!(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i20616_3_lut_4_lut_4_lut.init = 16'ha52b;
    PFUMX i25996 (.BLUT(n27785), .ALUT(n27783), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_1768[10]));
    LUT4 i24524_2_lut (.A(phase_i[4]), .B(phase_i[10]), .Z(index_q_9__N_1758[4])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(60[14] 63[8])
    defparam i24524_2_lut.init = 16'h9999;
    LUT4 mux_207_Mux_0_i364_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n364_adj_3457)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A ((C+!(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_0_i364_3_lut_3_lut_4_lut.init = 16'hdb55;
    LUT4 i20890_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n23372)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D))+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i20890_3_lut_4_lut.init = 16'hccdb;
    L6MUX21 i22639 (.D0(n25138), .D1(n25139), .SD(index_i[5]), .Z(n25140));
    LUT4 i24526_2_lut (.A(phase_i[3]), .B(phase_i[10]), .Z(index_q_9__N_1758[3])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(60[14] 63[8])
    defparam i24526_2_lut.init = 16'h9999;
    LUT4 i24528_2_lut (.A(phase_i[2]), .B(phase_i[10]), .Z(index_q_9__N_1758[2])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(60[14] 63[8])
    defparam i24528_2_lut.init = 16'h9999;
    LUT4 i24530_2_lut (.A(phase_i[1]), .B(phase_i[10]), .Z(index_q_9__N_1758[1])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(60[14] 63[8])
    defparam i24530_2_lut.init = 16'h9999;
    LUT4 i7149_2_lut (.A(phase_i[9]), .B(phase_i[10]), .Z(index_i_9__N_1748[9])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(60[14] 63[8])
    defparam i7149_2_lut.init = 16'h6666;
    LUT4 i7150_2_lut (.A(phase_i[8]), .B(phase_i[10]), .Z(index_i_9__N_1748[8])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(60[14] 63[8])
    defparam i7150_2_lut.init = 16'h6666;
    PFUMX i22743 (.BLUT(n526_adj_3092), .ALUT(n541_adj_3091), .C0(index_i[4]), 
          .Z(n25244));
    LUT4 i7151_2_lut (.A(phase_i[7]), .B(phase_i[10]), .Z(index_i_9__N_1748[7])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(60[14] 63[8])
    defparam i7151_2_lut.init = 16'h6666;
    LUT4 i7152_2_lut (.A(phase_i[6]), .B(phase_i[10]), .Z(index_i_9__N_1748[6])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(60[14] 63[8])
    defparam i7152_2_lut.init = 16'h6666;
    LUT4 i7153_2_lut (.A(phase_i[5]), .B(phase_i[10]), .Z(index_i_9__N_1748[5])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(60[14] 63[8])
    defparam i7153_2_lut.init = 16'h6666;
    PFUMX i25994 (.BLUT(n23287), .ALUT(n27781), .C0(index_i[7]), .Z(n27782));
    LUT4 mux_207_Mux_4_i262_3_lut_3_lut_rep_833 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n32034)) /* synthesis lut_function=(A (B+(C))+!A !(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_4_i262_3_lut_3_lut_rep_833.init = 16'ha9a9;
    LUT4 i7154_2_lut (.A(phase_i[4]), .B(phase_i[10]), .Z(index_i_9__N_1748[4])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(60[14] 63[8])
    defparam i7154_2_lut.init = 16'h6666;
    LUT4 mux_207_Mux_3_i397_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n397_adj_3298)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !(B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_3_i397_3_lut_4_lut_4_lut.init = 16'ha95a;
    PFUMX i22744 (.BLUT(n557_adj_3461), .ALUT(n572_adj_3213), .C0(index_i[4]), 
          .Z(n25245));
    LUT4 i7155_2_lut (.A(phase_i[3]), .B(phase_i[10]), .Z(index_i_9__N_1748[3])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(60[14] 63[8])
    defparam i7155_2_lut.init = 16'h6666;
    LUT4 i7156_2_lut (.A(phase_i[2]), .B(phase_i[10]), .Z(index_i_9__N_1748[2])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(60[14] 63[8])
    defparam i7156_2_lut.init = 16'h6666;
    LUT4 i7157_2_lut (.A(phase_i[1]), .B(phase_i[10]), .Z(index_i_9__N_1748[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(60[14] 63[8])
    defparam i7157_2_lut.init = 16'h6666;
    LUT4 mux_161_i16_3_lut (.A(\quarter_wave_sample_register_i[15] ), .B(o_val_pipeline_q_0__15__N_1831[15]), 
         .C(phase_negation_q[1]), .Z(n671[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(81[29:60])
    defparam mux_161_i16_3_lut.init = 16'hcaca;
    LUT4 mux_161_i15_3_lut (.A(quarter_wave_sample_register_q[14]), .B(o_val_pipeline_q_0__15__N_1831[14]), 
         .C(phase_negation_q[1]), .Z(n671[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(81[29:60])
    defparam mux_161_i15_3_lut.init = 16'hcaca;
    LUT4 mux_161_i14_3_lut (.A(quarter_wave_sample_register_q[13]), .B(o_val_pipeline_q_0__15__N_1831[13]), 
         .C(phase_negation_q[1]), .Z(n671[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(81[29:60])
    defparam mux_161_i14_3_lut.init = 16'hcaca;
    PFUMX i22745 (.BLUT(n589_adj_3090), .ALUT(n604_adj_2977), .C0(index_i[4]), 
          .Z(n25246));
    LUT4 mux_161_i13_3_lut (.A(quarter_wave_sample_register_q[12]), .B(o_val_pipeline_q_0__15__N_1831[12]), 
         .C(phase_negation_q[1]), .Z(n671[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(81[29:60])
    defparam mux_161_i13_3_lut.init = 16'hcaca;
    LUT4 i12452_2_lut_rep_691 (.A(index_q[0]), .B(index_q[1]), .Z(n29351)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i12452_2_lut_rep_691.init = 16'h4444;
    LUT4 i8307_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n157_adj_3376)) /* synthesis lut_function=(!(A (C (D))+!A !(B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i8307_3_lut_4_lut_4_lut.init = 16'h4aaa;
    LUT4 mux_161_i12_3_lut (.A(quarter_wave_sample_register_q[11]), .B(o_val_pipeline_q_0__15__N_1831[11]), 
         .C(phase_negation_q[1]), .Z(n671[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(81[29:60])
    defparam mux_161_i12_3_lut.init = 16'hcaca;
    LUT4 mux_161_i11_3_lut (.A(quarter_wave_sample_register_q[10]), .B(o_val_pipeline_q_0__15__N_1831[10]), 
         .C(phase_negation_q[1]), .Z(n671[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(81[29:60])
    defparam mux_161_i11_3_lut.init = 16'hcaca;
    LUT4 mux_161_i10_3_lut (.A(quarter_wave_sample_register_q[9]), .B(o_val_pipeline_q_0__15__N_1831[9]), 
         .C(phase_negation_q[1]), .Z(n671[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(81[29:60])
    defparam mux_161_i10_3_lut.init = 16'hcaca;
    PFUMX i22746 (.BLUT(n620_adj_3089), .ALUT(n635_adj_3462), .C0(index_i[4]), 
          .Z(n25247));
    LUT4 mux_207_Mux_0_i954_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n954_adj_3140)) /* synthesis lut_function=(A (D)+!A !(B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_0_i954_3_lut_4_lut_4_lut.init = 16'haf40;
    LUT4 mux_161_i9_3_lut (.A(quarter_wave_sample_register_q[8]), .B(o_val_pipeline_q_0__15__N_1831[8]), 
         .C(phase_negation_q[1]), .Z(n671[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(81[29:60])
    defparam mux_161_i9_3_lut.init = 16'hcaca;
    LUT4 n994_bdd_3_lut_25780_3_lut_4_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n27484)) /* synthesis lut_function=(A (B (C)+!B !(D))+!A !(D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n994_bdd_3_lut_25780_3_lut_4_lut_3_lut_4_lut.init = 16'h80f7;
    LUT4 mux_161_i8_3_lut (.A(quarter_wave_sample_register_q[7]), .B(o_val_pipeline_q_0__15__N_1831[7]), 
         .C(phase_negation_q[1]), .Z(n671[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(81[29:60])
    defparam mux_161_i8_3_lut.init = 16'hcaca;
    LUT4 mux_161_i7_3_lut (.A(quarter_wave_sample_register_q[6]), .B(o_val_pipeline_q_0__15__N_1831[6]), 
         .C(phase_negation_q[1]), .Z(n671[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(81[29:60])
    defparam mux_161_i7_3_lut.init = 16'hcaca;
    LUT4 mux_161_i6_3_lut (.A(quarter_wave_sample_register_q[5]), .B(o_val_pipeline_q_0__15__N_1831[5]), 
         .C(phase_negation_q[1]), .Z(n671[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(81[29:60])
    defparam mux_161_i6_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_3_i676_3_lut_4_lut_3_lut_rep_692 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29352)) /* synthesis lut_function=(A (B (C))+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_3_i676_3_lut_4_lut_3_lut_rep_692.init = 16'h9494;
    LUT4 mux_161_i5_3_lut (.A(quarter_wave_sample_register_q[4]), .B(o_val_pipeline_q_0__15__N_1831[4]), 
         .C(phase_negation_q[1]), .Z(n671[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(81[29:60])
    defparam mux_161_i5_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_6_i356_3_lut_4_lut_3_lut_rep_693 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29353)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_6_i356_3_lut_4_lut_3_lut_rep_693.init = 16'h4949;
    LUT4 mux_161_i4_3_lut (.A(quarter_wave_sample_register_q[3]), .B(o_val_pipeline_q_0__15__N_1831[3]), 
         .C(phase_negation_q[1]), .Z(n671[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(81[29:60])
    defparam mux_161_i4_3_lut.init = 16'hcaca;
    PFUMX i25977 (.BLUT(n27760), .ALUT(n27758), .C0(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_1783[10]));
    LUT4 mux_161_i3_3_lut (.A(quarter_wave_sample_register_q[2]), .B(o_val_pipeline_q_0__15__N_1831[2]), 
         .C(phase_negation_q[1]), .Z(n671[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(81[29:60])
    defparam mux_161_i3_3_lut.init = 16'hcaca;
    LUT4 mux_206_Mux_7_i526_3_lut_3_lut_4_lut_3_lut_4_lut (.A(index_i[1]), 
         .B(index_i[0]), .C(index_i[3]), .D(index_i[2]), .Z(n526_adj_3382)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(D))+!A !(D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_7_i526_3_lut_3_lut_4_lut_3_lut_4_lut.init = 16'h887f;
    LUT4 mux_161_i2_3_lut (.A(quarter_wave_sample_register_q[1]), .B(o_val_pipeline_q_0__15__N_1831[1]), 
         .C(phase_negation_q[1]), .Z(n671[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(81[29:60])
    defparam mux_161_i2_3_lut.init = 16'hcaca;
    LUT4 mux_207_Mux_6_i22_rep_694 (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .Z(n29354)) /* synthesis lut_function=(!(A (C)+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_6_i22_rep_694.init = 16'h4a4a;
    LUT4 mux_206_Mux_5_i38_3_lut_4_lut_3_lut_rep_775 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29435)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_5_i38_3_lut_4_lut_3_lut_rep_775.init = 16'h1919;
    LUT4 mux_207_Mux_2_i284_rep_695 (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .Z(n29355)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_2_i284_rep_695.init = 16'h4d4d;
    LUT4 mux_207_Mux_0_i490_3_lut_4_lut_3_lut_rep_696 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29356)) /* synthesis lut_function=(!(A (B+!(C))+!A ((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_0_i490_3_lut_4_lut_3_lut_rep_696.init = 16'h2424;
    PFUMX i22747 (.BLUT(n653_adj_3087), .ALUT(n668_adj_3450), .C0(index_i[4]), 
          .Z(n25248));
    LUT4 mux_207_Mux_0_i953_3_lut_rep_697 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29357)) /* synthesis lut_function=(A (C)+!A !((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_0_i953_3_lut_rep_697.init = 16'ha4a4;
    L6MUX21 i22691 (.D0(n23178), .D1(n23181), .SD(index_q[5]), .Z(n25192));
    LUT4 mux_161_i1_3_lut (.A(quarter_wave_sample_register_q[0]), .B(o_val_pipeline_q_0__15__N_1831[0]), 
         .C(phase_negation_q[1]), .Z(n671[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(81[29:60])
    defparam mux_161_i1_3_lut.init = 16'hcaca;
    LUT4 i20932_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n23414)) /* synthesis lut_function=(!(A ((D)+!C)+!A !(B ((D)+!C)+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i20932_3_lut_3_lut_4_lut.init = 16'h55a4;
    LUT4 mux_207_Mux_0_i491_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n491_adj_3463)) /* synthesis lut_function=(!(A (B (D)+!B !(C+!(D)))+!A ((C+!(D))+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_0_i491_3_lut_4_lut.init = 16'h24aa;
    LUT4 i1_2_lut (.A(o_phase[11]), .B(o_phase[10]), .Z(phase_q_11__N_1874[11])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i1_2_lut.init = 16'h9999;
    LUT4 mux_207_Mux_2_i890_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n890_adj_3285)) /* synthesis lut_function=(A (B (D)+!B !((D)+!C))+!A !(B (C+(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_2_i890_3_lut_4_lut_4_lut.init = 16'h9934;
    L6MUX21 i22695 (.D0(n23187), .D1(n19983), .SD(index_q[5]), .Z(n25196));
    LUT4 mux_207_Mux_3_i653_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n653_adj_3193)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A !(B (D)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_3_i653_3_lut_4_lut_4_lut.init = 16'h4d99;
    PFUMX i22748 (.BLUT(n684_adj_3425), .ALUT(n699_adj_3446), .C0(index_i[4]), 
          .Z(n25249));
    LUT4 mux_207_Mux_5_i475_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n475_adj_3393)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_5_i475_3_lut_4_lut_4_lut.init = 16'hd4a5;
    L6MUX21 i22696 (.D0(n23193), .D1(n13394), .SD(index_q[5]), .Z(n25197));
    LUT4 mux_207_Mux_0_i157_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n157_adj_3365)) /* synthesis lut_function=(A (B (C+!(D))+!B !(D))+!A (B (D)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_0_i157_3_lut_4_lut.init = 16'hd4aa;
    LUT4 mux_207_Mux_5_i491_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n491_adj_3178)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A !(B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_5_i491_3_lut_4_lut_4_lut.init = 16'ha54a;
    PFUMX i22698 (.BLUT(n542_adj_3085), .ALUT(n573_adj_3414), .C0(index_q[5]), 
          .Z(n25199));
    LUT4 i20910_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n23392)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (D))+!A !(B (C (D))+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i20910_3_lut_3_lut_4_lut.init = 16'h4933;
    LUT4 n572_bdd_3_lut_26943_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n27583)) /* synthesis lut_function=(A (B (C+(D)))+!A (B ((D)+!C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam n572_bdd_3_lut_26943_4_lut.init = 16'hcc94;
    LUT4 mux_207_Mux_3_i684_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[4]), .Z(n684_adj_3409)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A !(B ((D)+!C)+!B (C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_3_i684_3_lut_3_lut_4_lut.init = 16'h5594;
    PFUMX i22749 (.BLUT(n716_adj_3083), .ALUT(n731_adj_2948), .C0(index_i[4]), 
          .Z(n25250));
    LUT4 mux_207_Mux_2_i653_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n653_adj_3164)) /* synthesis lut_function=(A (B (C+!(D))+!B !(D))+!A !(B (C+!(D))+!B !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_2_i653_3_lut_4_lut.init = 16'h94aa;
    LUT4 mux_207_Mux_0_i781_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n781_adj_3432)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A (B (C)+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_0_i781_4_lut_4_lut_4_lut.init = 16'h0cb4;
    PFUMX i25975 (.BLUT(n23269), .ALUT(n27756), .C0(index_q[7]), .Z(n27757));
    LUT4 mux_206_Mux_0_i219_3_lut_3_lut_3_lut_rep_776 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29436)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i219_3_lut_3_lut_3_lut_rep_776.init = 16'h9393;
    L6MUX21 i25970 (.D0(n27749), .D1(n27746), .SD(index_q[5]), .Z(n27750));
    PFUMX i25968 (.BLUT(n27748), .ALUT(n27747), .C0(index_q[4]), .Z(n27749));
    L6MUX21 i25081 (.D0(n26729), .D1(n26727), .SD(index_i[5]), .Z(n26730));
    PFUMX i22699 (.BLUT(n605_adj_3149), .ALUT(n636_adj_3389), .C0(index_q[5]), 
          .Z(n25200));
    LUT4 mux_206_Mux_6_i284_3_lut_4_lut_3_lut_rep_777 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29437)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_6_i284_3_lut_4_lut_3_lut_rep_777.init = 16'h6969;
    PFUMX i27919 (.BLUT(n30640), .ALUT(n30639), .C0(index_q[3]), .Z(n30641));
    PFUMX i22750 (.BLUT(n747_adj_3434), .ALUT(n762_adj_3464), .C0(index_i[4]), 
          .Z(n25251));
    PFUMX i25079 (.BLUT(n26728), .ALUT(n285_adj_3027), .C0(index_i[4]), 
          .Z(n26729));
    PFUMX i22700 (.BLUT(n669_adj_3080), .ALUT(n700_adj_3208), .C0(index_q[5]), 
          .Z(n25201));
    PFUMX i22751 (.BLUT(n781_adj_3465), .ALUT(n796_adj_3466), .C0(index_i[4]), 
          .Z(n25252));
    LUT4 i14174_2_lut_rep_700 (.A(index_q[3]), .B(index_q[4]), .Z(n29360)) /* synthesis lut_function=(A (B)) */ ;
    defparam i14174_2_lut_rep_700.init = 16'h8888;
    PFUMX i22701 (.BLUT(n732_adj_3197), .ALUT(n23199), .C0(index_q[5]), 
          .Z(n25202));
    LUT4 i24459_3_lut_4_lut (.A(n29101), .B(n29251), .C(index_i[8]), .D(n766), 
         .Z(n23249)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i24459_3_lut_4_lut.init = 16'hefe0;
    PFUMX i27915 (.BLUT(n30636), .ALUT(n30635), .C0(index_q[2]), .Z(n30637));
    LUT4 i22738_3_lut_3_lut_4_lut (.A(index_q[3]), .B(index_q[4]), .C(n413_adj_3402), 
         .D(index_q[5]), .Z(n25239)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(C+(D)))) */ ;
    defparam i22738_3_lut_3_lut_4_lut.init = 16'h77f0;
    PFUMX i22752 (.BLUT(n812_adj_3467), .ALUT(n13320), .C0(index_i[4]), 
          .Z(n25253));
    LUT4 i14195_2_lut_rep_442_3_lut (.A(index_q[3]), .B(index_q[4]), .C(index_q[5]), 
         .Z(n29102)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam i14195_2_lut_rep_442_3_lut.init = 16'hf8f8;
    PFUMX i22702 (.BLUT(n797_adj_3076), .ALUT(n828_adj_3075), .C0(index_q[5]), 
          .Z(n25203));
    LUT4 i1_2_lut_3_lut (.A(index_q[3]), .B(index_q[4]), .C(index_q[5]), 
         .Z(n22328)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h8080;
    LUT4 i14371_2_lut_3_lut_4_lut (.A(index_q[3]), .B(index_q[4]), .C(index_q[2]), 
         .D(n29465), .Z(n16798)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i14371_2_lut_3_lut_4_lut.init = 16'h8880;
    LUT4 i1_2_lut_rep_701 (.A(index_q[3]), .B(index_q[2]), .Z(n29361)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i1_2_lut_rep_701.init = 16'heeee;
    PFUMX i25965 (.BLUT(n27745), .ALUT(n316_adj_3334), .C0(index_q[4]), 
          .Z(n27746));
    LUT4 i21391_3_lut_then_4_lut (.A(index_i[4]), .B(index_i[2]), .C(index_i[3]), 
         .D(index_i[0]), .Z(n29500)) /* synthesis lut_function=(!(A (B (C)+!B ((D)+!C))+!A !((C)+!B))) */ ;
    defparam i21391_3_lut_then_4_lut.init = 16'h5979;
    LUT4 i21391_3_lut_else_4_lut (.A(index_i[4]), .B(index_i[2]), .C(index_i[3]), 
         .D(index_i[0]), .Z(n29499)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A !(B (C+!(D))+!B !(C)))) */ ;
    defparam i21391_3_lut_else_4_lut.init = 16'h6965;
    PFUMX i22703 (.BLUT(n860), .ALUT(n891_adj_3073), .C0(index_q[5]), 
          .Z(n25204));
    PFUMX i22754 (.BLUT(n875_adj_3448), .ALUT(n890_adj_2983), .C0(index_i[4]), 
          .Z(n25255));
    PFUMX i25077 (.BLUT(n26726), .ALUT(n26725), .C0(index_i[4]), .Z(n26727));
    PFUMX i22755 (.BLUT(n908_adj_2992), .ALUT(n923_adj_3067), .C0(index_i[4]), 
          .Z(n25256));
    LUT4 i13059_2_lut_rep_501_3_lut (.A(index_q[3]), .B(index_q[2]), .C(index_q[1]), 
         .Z(n29161)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i13059_2_lut_rep_501_3_lut.init = 16'hfefe;
    L6MUX21 i22759 (.D0(n25244), .D1(n25245), .SD(index_i[5]), .Z(n25260));
    L6MUX21 i22760 (.D0(n25246), .D1(n25247), .SD(index_i[5]), .Z(n25261));
    L6MUX21 i22761 (.D0(n25248), .D1(n25249), .SD(index_i[5]), .Z(n25262));
    PFUMX i22756 (.BLUT(n939), .ALUT(n954_adj_3468), .C0(index_i[4]), 
          .Z(n25257));
    L6MUX21 i22762 (.D0(n25250), .D1(n25251), .SD(index_i[5]), .Z(n25263));
    PFUMX i27881 (.BLUT(n30582), .ALUT(n30581), .C0(index_i[3]), .Z(n30583));
    L6MUX21 i22763 (.D0(n25252), .D1(n25253), .SD(index_i[5]), .Z(n25264));
    PFUMX i22757 (.BLUT(n971), .ALUT(n986), .C0(index_i[4]), .Z(n25258));
    L6MUX21 i22764 (.D0(n25254), .D1(n25255), .SD(index_i[5]), .Z(n25265));
    L6MUX21 i22765 (.D0(n25256), .D1(n25257), .SD(index_i[5]), .Z(n25266));
    L6MUX21 i22766 (.D0(n25258), .D1(n25259), .SD(index_i[5]), .Z(n25267));
    L6MUX21 i22782 (.D0(n23919), .D1(n23922), .SD(index_i[5]), .Z(n25283));
    PFUMX i22758 (.BLUT(n1002_adj_3215), .ALUT(n1017), .C0(index_i[4]), 
          .Z(n25259));
    PFUMX i27877 (.BLUT(n30578), .ALUT(n30577), .C0(index_i[2]), .Z(n30579));
    PFUMX i22489 (.BLUT(n491_adj_3463), .ALUT(n12256), .C0(index_q[4]), 
          .Z(n24990));
    L6MUX21 i25074 (.D0(n26723), .D1(n26720), .SD(index_i[5]), .Z(n26724));
    L6MUX21 i22786 (.D0(n23928), .D1(n20014), .SD(index_i[5]), .Z(n25287));
    PFUMX i20705 (.BLUT(n23185), .ALUT(n23186), .C0(index_q[4]), .Z(n23187));
    PFUMX i25072 (.BLUT(n26722), .ALUT(n26721), .C0(index_i[4]), .Z(n26723));
    L6MUX21 i22787 (.D0(n23937), .D1(n13335), .SD(index_i[5]), .Z(n25288));
    PFUMX i22789 (.BLUT(n542_adj_3059), .ALUT(n573_adj_3452), .C0(index_i[5]), 
          .Z(n25290));
    LUT4 n284_bdd_3_lut_25833_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n27585)) /* synthesis lut_function=(A (B (C+(D))+!B ((D)+!C))+!A !(B (C+(D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam n284_bdd_3_lut_25833_4_lut.init = 16'haa96;
    LUT4 i21468_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n23950)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(D))+!A (B))) */ ;
    defparam i21468_3_lut_3_lut_4_lut.init = 16'h3319;
    PFUMX i25069 (.BLUT(n26719), .ALUT(n26718), .C0(index_i[4]), .Z(n26720));
    LUT4 mux_207_Mux_8_i506_3_lut_4_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n506_adj_3346)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B ((D)+!C)))) */ ;
    defparam mux_207_Mux_8_i506_3_lut_4_lut_3_lut_4_lut.init = 16'h0ef0;
    PFUMX i22790 (.BLUT(n605_adj_3415), .ALUT(n636_adj_3469), .C0(index_i[5]), 
          .Z(n25291));
    LUT4 i14251_2_lut_rep_705 (.A(index_i[3]), .B(index_i[4]), .Z(n29365)) /* synthesis lut_function=(A (B)) */ ;
    defparam i14251_2_lut_rep_705.init = 16'h8888;
    LUT4 i22664_3_lut_3_lut_4_lut (.A(index_i[3]), .B(index_i[4]), .C(n413_adj_3241), 
         .D(index_i[5]), .Z(n25165)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(C+(D)))) */ ;
    defparam i22664_3_lut_3_lut_4_lut.init = 16'h77f0;
    LUT4 i12469_2_lut_rep_520_3_lut (.A(index_i[1]), .B(index_i[0]), .C(index_i[2]), 
         .Z(n29180)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12469_2_lut_rep_520_3_lut.init = 16'hf8f8;
    LUT4 n27194_bdd_3_lut_28072 (.A(n27194), .B(n27190), .C(index_i[6]), 
         .Z(n27195)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n27194_bdd_3_lut_28072.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_adj_189 (.A(index_i[3]), .B(index_i[4]), .C(index_i[5]), 
         .Z(n22332)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_3_lut_adj_189.init = 16'h8080;
    LUT4 mux_206_Mux_5_i761_3_lut_4_lut_3_lut_rep_778 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29438)) /* synthesis lut_function=(A (B)+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_5_i761_3_lut_4_lut_3_lut_rep_778.init = 16'hd9d9;
    PFUMX i22490 (.BLUT(n24975), .ALUT(n24976), .C0(index_q[5]), .Z(n24991));
    LUT4 i14273_2_lut_rep_441_3_lut (.A(index_i[3]), .B(index_i[4]), .C(index_i[5]), 
         .Z(n29101)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam i14273_2_lut_rep_441_3_lut.init = 16'hf8f8;
    LUT4 i14400_2_lut_3_lut_4_lut (.A(index_i[3]), .B(index_i[4]), .C(index_i[2]), 
         .D(n29376), .Z(n16828)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i14400_2_lut_3_lut_4_lut.init = 16'h8880;
    LUT4 mux_206_Mux_8_i732_3_lut (.A(index_i[3]), .B(n16900), .C(index_i[5]), 
         .Z(n732)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_8_i732_3_lut.init = 16'h3a3a;
    PFUMX i25867 (.BLUT(n27619), .ALUT(n32055), .C0(index_q[3]), .Z(n27620));
    LUT4 mux_207_Mux_0_i124_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n124_adj_3326)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A !(B (D)+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_0_i124_3_lut_4_lut_4_lut.init = 16'h6c99;
    LUT4 mux_206_Mux_0_i900_3_lut_4_lut_3_lut_rep_779 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29439)) /* synthesis lut_function=(A (B)+!A !(B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i900_3_lut_4_lut_3_lut_rep_779.init = 16'h9898;
    LUT4 mux_206_Mux_4_i1002_3_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n1002_adj_3436)) /* synthesis lut_function=(A (B (C (D))+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_4_i1002_3_lut_3_lut_4_lut.init = 16'hf007;
    CCU2D unary_minus_27_add_3_17 (.A0(\quarter_wave_sample_register_i[15] ), 
          .B0(GND_net), .C0(GND_net), .D0(GND_net), .A1(GND_net), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n19713), .S0(o_val_pipeline_q_0__15__N_1831[15]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(81[29:60])
    defparam unary_minus_27_add_3_17.INIT0 = 16'hf555;
    defparam unary_minus_27_add_3_17.INIT1 = 16'h0000;
    defparam unary_minus_27_add_3_17.INJECT1_0 = "NO";
    defparam unary_minus_27_add_3_17.INJECT1_1 = "NO";
    PFUMX i22791 (.BLUT(n669), .ALUT(n700_adj_3189), .C0(index_i[5]), 
          .Z(n25292));
    PFUMX i22792 (.BLUT(n732_adj_3187), .ALUT(n23955), .C0(index_i[5]), 
          .Z(n25293));
    LUT4 i23990_3_lut (.A(n23611), .B(n23612), .C(index_i[4]), .Z(n23613)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i23990_3_lut.init = 16'hcaca;
    LUT4 i21447_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[0]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n23929)) /* synthesis lut_function=(!(A (C+(D))+!A !(B (C (D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21447_4_lut_4_lut_4_lut.init = 16'h501a;
    LUT4 i14181_2_lut_rep_740 (.A(index_i[1]), .B(index_i[2]), .Z(n29400)) /* synthesis lut_function=(A (B)) */ ;
    defparam i14181_2_lut_rep_740.init = 16'h8888;
    LUT4 mux_206_Mux_4_i93_3_lut_4_lut_3_lut_rep_659_4_lut (.A(index_i[1]), 
         .B(index_i[2]), .C(index_i[3]), .D(index_i[0]), .Z(n29319)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D)))) */ ;
    defparam mux_206_Mux_4_i93_3_lut_4_lut_3_lut_rep_659_4_lut.init = 16'h07f0;
    LUT4 mux_207_Mux_0_i715_3_lut_3_lut_rep_834 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n32035)) /* synthesis lut_function=(A (B (C))+!A !(B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_0_i715_3_lut_3_lut_rep_834.init = 16'h9595;
    LUT4 mux_206_Mux_6_i134_3_lut_4_lut_3_lut_rep_780 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29440)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_6_i134_3_lut_4_lut_3_lut_rep_780.init = 16'h9696;
    LUT4 mux_206_Mux_3_i142_3_lut_3_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .Z(n142_adj_3427)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B+!(C)))) */ ;
    defparam mux_206_Mux_3_i142_3_lut_3_lut_3_lut.init = 16'h3838;
    PFUMX i22793 (.BLUT(n797_adj_3040), .ALUT(n828_adj_3038), .C0(index_i[5]), 
          .Z(n25294));
    LUT4 i13083_2_lut_rep_467_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[0]), 
         .Z(n29127)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13083_2_lut_rep_467_3_lut.init = 16'h7070;
    LUT4 i11077_2_lut_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[3]), 
         .Z(n13373)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i11077_2_lut_3_lut.init = 16'h8080;
    LUT4 mux_206_Mux_3_i1002_3_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n21706)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (D))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_3_i1002_3_lut_3_lut_4_lut.init = 16'hf708;
    LUT4 n953_bdd_3_lut_26722_4_lut (.A(n29346), .B(index_q[2]), .C(index_q[3]), 
         .D(n29333), .Z(n26647)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam n953_bdd_3_lut_26722_4_lut.init = 16'hf606;
    LUT4 i12678_2_lut_rep_488_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[3]), 
         .Z(n29148)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam i12678_2_lut_rep_488_3_lut.init = 16'hf8f8;
    LUT4 mux_206_Mux_6_i340_3_lut_4_lut_4_lut_3_lut_rep_781 (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[2]), .Z(n29441)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_6_i340_3_lut_4_lut_4_lut_3_lut_rep_781.init = 16'h9292;
    L6MUX21 i25836 (.D0(n27587), .D1(n27584), .SD(index_q[5]), .Z(n27588));
    PFUMX i22794 (.BLUT(n860_adj_3000), .ALUT(n891_adj_3035), .C0(index_i[5]), 
          .Z(n25295));
    PFUMX i25834 (.BLUT(n27586), .ALUT(n27585), .C0(index_q[4]), .Z(n27587));
    LUT4 mux_207_Mux_3_i890_3_lut_4_lut (.A(n29346), .B(index_q[2]), .C(index_q[3]), 
         .D(n325), .Z(n890_adj_3273)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_3_i890_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_207_Mux_1_i93_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n93_adj_3358)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C+(D)))+!A !(B (C (D)+!C !(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_1_i93_3_lut_4_lut_4_lut.init = 16'h955a;
    LUT4 i13845_2_lut_rep_526_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[0]), 
         .Z(n29186)) /* synthesis lut_function=(A (B+!(C))+!A !(C)) */ ;
    defparam i13845_2_lut_rep_526_3_lut.init = 16'h8f8f;
    LUT4 mux_206_Mux_3_i396_3_lut_3_lut_rep_782 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29442)) /* synthesis lut_function=(A (B+(C))+!A !(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_3_i396_3_lut_3_lut_rep_782.init = 16'ha9a9;
    LUT4 i20695_3_lut_4_lut (.A(n29346), .B(index_q[2]), .C(index_q[3]), 
         .D(n29390), .Z(n23177)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i20695_3_lut_4_lut.init = 16'hf606;
    LUT4 i22315_3_lut (.A(n85), .B(n29467), .C(index_q[3]), .Z(n24816)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22315_3_lut.init = 16'hcaca;
    LUT4 mux_206_Mux_2_i262_3_lut_3_lut_rep_783 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29443)) /* synthesis lut_function=(A (B)+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_2_i262_3_lut_3_lut_rep_783.init = 16'h9c9c;
    LUT4 i12892_2_lut_rep_517_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[0]), 
         .Z(n29177)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i12892_2_lut_rep_517_3_lut.init = 16'h8080;
    PFUMX i20711 (.BLUT(n23191), .ALUT(n23192), .C0(index_q[4]), .Z(n23193));
    LUT4 i20659_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .D(index_i[3]), .Z(n23141)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(D))+!A (B+!(D)))) */ ;
    defparam i20659_3_lut_4_lut_4_lut_4_lut.init = 16'h3380;
    LUT4 i22314_3_lut (.A(n29181), .B(n29315), .C(index_q[3]), .Z(n24815)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22314_3_lut.init = 16'hcaca;
    LUT4 mux_206_Mux_9_i30_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .D(index_i[3]), .Z(n30_adj_3210)) /* synthesis lut_function=(A (B (C (D))+!B !(D))+!A !(B+(D))) */ ;
    defparam mux_206_Mux_9_i30_3_lut_4_lut_4_lut_4_lut.init = 16'h8033;
    LUT4 i12580_2_lut_rep_404_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n29064)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;
    defparam i12580_2_lut_rep_404_3_lut_4_lut.init = 16'hf8f0;
    LUT4 mux_206_Mux_8_i491_3_lut_3_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n491_adj_3391)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A !(C))) */ ;
    defparam mux_206_Mux_8_i491_3_lut_3_lut_3_lut_4_lut.init = 16'h7870;
    LUT4 i21520_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n24002)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C (D)+!C !(D)))+!A !(B (D)+!B (C (D)+!C !(D))))) */ ;
    defparam i21520_3_lut_4_lut_4_lut_4_lut.init = 16'h7c03;
    LUT4 i20587_3_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[3]), 
         .D(index_i[0]), .Z(n23069)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D))) */ ;
    defparam i20587_3_lut_3_lut_4_lut.init = 16'hf80f;
    LUT4 mux_207_Mux_12_i254_4_lut (.A(n29045), .B(n22328), .C(index_q[6]), 
         .D(n29168), .Z(n254_adj_3458)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_12_i254_4_lut.init = 16'hca0a;
    PFUMX i25831 (.BLUT(n27583), .ALUT(n29057), .C0(index_q[4]), .Z(n27584));
    L6MUX21 i25823 (.D0(n27576), .D1(n27574), .SD(index_q[4]), .Z(n27577));
    PFUMX i25821 (.BLUT(n29080), .ALUT(n27575), .C0(index_q[5]), .Z(n27576));
    CCU2D unary_minus_27_add_3_15 (.A0(quarter_wave_sample_register_q[13]), 
          .B0(GND_net), .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_q[14]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19712), .COUT(n19713), 
          .S0(o_val_pipeline_q_0__15__N_1831[13]), .S1(o_val_pipeline_q_0__15__N_1831[14]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(81[29:60])
    defparam unary_minus_27_add_3_15.INIT0 = 16'hf555;
    defparam unary_minus_27_add_3_15.INIT1 = 16'hf555;
    defparam unary_minus_27_add_3_15.INJECT1_0 = "NO";
    defparam unary_minus_27_add_3_15.INJECT1_1 = "NO";
    PFUMX i25819 (.BLUT(n27573), .ALUT(n27572), .C0(index_q[5]), .Z(n27574));
    LUT4 i22665_3_lut_4_lut_4_lut (.A(n29145), .B(index_i[4]), .C(index_i[5]), 
         .D(n29146), .Z(n25166)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C)+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i22665_3_lut_4_lut_4_lut.init = 16'h0434;
    CCU2D unary_minus_27_add_3_13 (.A0(quarter_wave_sample_register_q[11]), 
          .B0(GND_net), .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_q[12]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19711), .COUT(n19712), 
          .S0(o_val_pipeline_q_0__15__N_1831[11]), .S1(o_val_pipeline_q_0__15__N_1831[12]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(81[29:60])
    defparam unary_minus_27_add_3_13.INIT0 = 16'hf555;
    defparam unary_minus_27_add_3_13.INIT1 = 16'hf555;
    defparam unary_minus_27_add_3_13.INJECT1_0 = "NO";
    defparam unary_minus_27_add_3_13.INJECT1_1 = "NO";
    CCU2D unary_minus_27_add_3_11 (.A0(quarter_wave_sample_register_q[9]), 
          .B0(GND_net), .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_q[10]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19710), .COUT(n19711), 
          .S0(o_val_pipeline_q_0__15__N_1831[9]), .S1(o_val_pipeline_q_0__15__N_1831[10]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(81[29:60])
    defparam unary_minus_27_add_3_11.INIT0 = 16'hf555;
    defparam unary_minus_27_add_3_11.INIT1 = 16'hf555;
    defparam unary_minus_27_add_3_11.INJECT1_0 = "NO";
    defparam unary_minus_27_add_3_11.INJECT1_1 = "NO";
    LUT4 mux_206_Mux_3_i723_3_lut_4_lut_3_lut_rep_784 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29444)) /* synthesis lut_function=(A (B (C))+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_3_i723_3_lut_4_lut_3_lut_rep_784.init = 16'h9494;
    LUT4 mux_206_Mux_6_i867_3_lut_3_lut_rep_717 (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[2]), .Z(n29377)) /* synthesis lut_function=(!(A (B (C))+!A !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_6_i867_3_lut_3_lut_rep_717.init = 16'h7a7a;
    LUT4 mux_207_Mux_3_i491_3_lut_4_lut (.A(n29276), .B(index_q[1]), .C(index_q[3]), 
         .D(n32033), .Z(n491_adj_2959)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_3_i491_3_lut_4_lut.init = 16'h4f40;
    L6MUX21 i25808 (.D0(n27560), .D1(n27558), .SD(index_q[5]), .Z(n27561));
    PFUMX i25806 (.BLUT(n27559), .ALUT(n285_adj_3238), .C0(index_q[4]), 
          .Z(n27560));
    LUT4 mux_206_Mux_4_i77_3_lut_3_lut_rep_785 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29445)) /* synthesis lut_function=(A (B (C))+!A !(B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_4_i77_3_lut_3_lut_rep_785.init = 16'h9595;
    LUT4 mux_206_Mux_8_i892_3_lut_4_lut (.A(n29145), .B(index_i[4]), .C(index_i[5]), 
         .D(n860_adj_3266), .Z(n892_adj_3217)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_8_i892_3_lut_4_lut.init = 16'h4f40;
    PFUMX i25804 (.BLUT(n301_adj_3071), .ALUT(n27557), .C0(index_q[4]), 
          .Z(n27558));
    LUT4 index_i_5__bdd_3_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n28103)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C (D)))+!A (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam index_i_5__bdd_3_lut_3_lut_4_lut.init = 16'h0fa7;
    LUT4 i12462_2_lut_rep_742 (.A(index_i[0]), .B(index_i[1]), .Z(n29402)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12462_2_lut_rep_742.init = 16'h4444;
    LUT4 i7789_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n157_adj_3453)) /* synthesis lut_function=(!(A (C (D))+!A !(B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i7789_3_lut_4_lut_4_lut.init = 16'h4aaa;
    LUT4 mux_207_Mux_0_i475_3_lut_4_lut (.A(n29276), .B(index_q[1]), .C(index_q[3]), 
         .D(n29168), .Z(n475_adj_3459)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_0_i475_3_lut_4_lut.init = 16'h4f40;
    PFUMX i25785 (.BLUT(n27538), .ALUT(n27537), .C0(index_i[4]), .Z(n27539));
    LUT4 mux_206_Mux_0_i954_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n954_adj_3468)) /* synthesis lut_function=(A (D)+!A !(B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i954_3_lut_4_lut_4_lut.init = 16'haf40;
    LUT4 mux_206_Mux_6_i505_3_lut_rep_786 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29446)) /* synthesis lut_function=(A (B)+!A (B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_6_i505_3_lut_rep_786.init = 16'hc9c9;
    LUT4 mux_206_Mux_6_i378_3_lut_4_lut_3_lut_rep_787 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29447)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_6_i378_3_lut_4_lut_3_lut_rep_787.init = 16'h4949;
    LUT4 mux_206_Mux_8_i205_3_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n205_adj_3399)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_8_i205_3_lut_3_lut_4_lut.init = 16'h7a0f;
    LUT4 mux_206_Mux_6_i269_rep_743 (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .Z(n29403)) /* synthesis lut_function=(A (C)+!A !((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_6_i269_rep_743.init = 16'ha4a4;
    LUT4 i20733_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n23215)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (D))+!A !(B (C (D))+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20733_3_lut_3_lut_4_lut.init = 16'h4933;
    LUT4 mux_206_Mux_5_i483_rep_744 (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .Z(n29404)) /* synthesis lut_function=(!(A (C)+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_5_i483_rep_744.init = 16'h4a4a;
    LUT4 mux_206_Mux_0_i557_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n557_adj_3461)) /* synthesis lut_function=(A ((D)+!C)+!A !((D)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i557_3_lut_4_lut.init = 16'haa4e;
    LUT4 mux_206_Mux_0_i781_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n781_adj_3465)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A (B (C)+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i781_4_lut_4_lut_4_lut.init = 16'h0cb4;
    LUT4 mux_206_Mux_5_i491_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n491_adj_3195)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A !(B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_5_i491_3_lut_4_lut_4_lut.init = 16'ha54a;
    LUT4 i20758_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n23240)) /* synthesis lut_function=(!(A ((D)+!C)+!A !(B ((D)+!C)+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20758_3_lut_3_lut_4_lut.init = 16'h55a4;
    CCU2D unary_minus_27_add_3_9 (.A0(quarter_wave_sample_register_q[7]), 
          .B0(GND_net), .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_q[8]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19709), .COUT(n19710), 
          .S0(o_val_pipeline_q_0__15__N_1831[7]), .S1(o_val_pipeline_q_0__15__N_1831[8]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(81[29:60])
    defparam unary_minus_27_add_3_9.INIT0 = 16'hf555;
    defparam unary_minus_27_add_3_9.INIT1 = 16'hf555;
    defparam unary_minus_27_add_3_9.INJECT1_0 = "NO";
    defparam unary_minus_27_add_3_9.INJECT1_1 = "NO";
    FD1S3BX quarter_wave_sample_register_i_i15 (.D(n32066), .CK(dac_clk_p_c), 
            .PD(i_sw0_c), .Q(\quarter_wave_sample_register_i[15] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_i_i15.GSR = "DISABLED";
    L6MUX21 i25764 (.D0(n27512), .D1(n27509), .SD(index_i[5]), .Z(n27513));
    PFUMX i25762 (.BLUT(n27511), .ALUT(n27510), .C0(index_i[4]), .Z(n27512));
    LUT4 n476_bdd_3_lut_3_lut (.A(index_i[1]), .B(index_i[4]), .C(n124_adj_3281), 
         .Z(n28442)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n476_bdd_3_lut_3_lut.init = 16'hd1d1;
    LUT4 n23123_bdd_3_lut_3_lut (.A(index_i[1]), .B(n812_adj_3057), .C(index_i[4]), 
         .Z(n28444)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n23123_bdd_3_lut_3_lut.init = 16'h5c5c;
    LUT4 mux_206_Mux_0_i985_3_lut_4_lut_3_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .Z(n985)) /* synthesis lut_function=(!(A (B+(C))+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i985_3_lut_4_lut_3_lut_3_lut.init = 16'h4343;
    PFUMX i25758 (.BLUT(n27508), .ALUT(n29070), .C0(index_i[4]), .Z(n27509));
    FD1S3BX quarter_wave_sample_register_i_i14 (.D(quarter_wave_sample_register_i_15__N_1768[14]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_i[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_i_i14.GSR = "DISABLED";
    LUT4 i21457_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n23939)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C+(D)))+!A (B (C)+!B !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21457_3_lut_4_lut_4_lut.init = 16'hc95a;
    FD1S3BX quarter_wave_sample_register_i_i13 (.D(quarter_wave_sample_register_i_15__N_1768[13]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_i[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_i_i13.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i12 (.D(quarter_wave_sample_register_i_15__N_1768[12]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_i[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_i_i12.GSR = "DISABLED";
    LUT4 i12715_2_lut_rep_525_2_lut (.A(index_i[1]), .B(index_i[0]), .Z(n29185)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12715_2_lut_rep_525_2_lut.init = 16'h4444;
    FD1S3BX quarter_wave_sample_register_i_i11 (.D(quarter_wave_sample_register_i_15__N_1768[11]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_i[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_i_i11.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i10 (.D(quarter_wave_sample_register_i_15__N_1768[10]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_i[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_i_i10.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i9 (.D(quarter_wave_sample_register_i_15__N_1768[9]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_i[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_i_i9.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i8 (.D(quarter_wave_sample_register_i_15__N_1768[8]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_i[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_i_i8.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i7 (.D(quarter_wave_sample_register_i_15__N_1768[7]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_i[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_i_i7.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i6 (.D(quarter_wave_sample_register_i_15__N_1768[6]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_i[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_i_i6.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i5 (.D(quarter_wave_sample_register_i_15__N_1768[5]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_i[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_i_i5.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i4 (.D(quarter_wave_sample_register_i_15__N_1768[4]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_i[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_i_i4.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i3 (.D(quarter_wave_sample_register_i_15__N_1768[3]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_i[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_i_i3.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i2 (.D(quarter_wave_sample_register_i_15__N_1768[2]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_i[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_i_i2.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i1 (.D(quarter_wave_sample_register_i_15__N_1768[1]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_i[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_i_i1.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i32 (.D(n670[15]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_i[0] [15])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i32.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i31 (.D(n670[14]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_i[0] [14])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i31.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i30 (.D(n670[13]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_i[0] [13])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i30.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i29 (.D(n670[12]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_i[0] [12])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i29.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i28 (.D(n670[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_i[0] [11])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i28.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i27 (.D(n670[10]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_i[0] [10])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i27.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i26 (.D(n670[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_i[0] [9])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i26.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i25 (.D(n670[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_i[0] [8])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i25.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i24 (.D(n670[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_i[0] [7])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i24.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i23 (.D(n670[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_i[0] [6])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i23.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i22 (.D(n670[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_i[0] [5])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i22.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i21 (.D(n670[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_i[0] [4])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i21.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i20 (.D(n670[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_i[0] [3])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i20.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i19 (.D(n670[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_i[0] [2])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i19.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i18 (.D(n670[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_i[0] [1])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i18.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i17 (.D(n670[0]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_i[0] [0])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i17.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i16 (.D(\o_val_pipeline_i[0] [15]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(o_sample_i[15])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i16.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i15 (.D(\o_val_pipeline_i[0] [14]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(o_sample_i[14])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i15.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i14 (.D(\o_val_pipeline_i[0] [13]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(o_sample_i[13])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i14.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i13 (.D(\o_val_pipeline_i[0] [12]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(o_sample_i[12])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i13.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i12 (.D(\o_val_pipeline_i[0] [11]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(o_sample_i[11])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i12.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i11 (.D(\o_val_pipeline_i[0] [10]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(o_sample_i[10])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i11.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i10 (.D(\o_val_pipeline_i[0] [9]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(o_sample_i[9])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i10.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i9 (.D(\o_val_pipeline_i[0] [8]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(o_sample_i[8])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i9.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i8 (.D(\o_val_pipeline_i[0] [7]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(o_sample_i[7])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i8.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i7 (.D(\o_val_pipeline_i[0] [6]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(o_sample_i[6])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i7.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i6 (.D(\o_val_pipeline_i[0] [5]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(o_sample_i[5])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i6.GSR = "DISABLED";
    LUT4 mux_206_Mux_1_i93_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n93_adj_3395)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C+(D)))+!A !(B (C (D)+!C !(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_1_i93_3_lut_4_lut_4_lut.init = 16'h955a;
    FD1S3DX o_val_pipeline_i_1__i5 (.D(\o_val_pipeline_i[0] [4]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(o_sample_i[4])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i5.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i4 (.D(\o_val_pipeline_i[0] [3]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(o_sample_i[3])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i4.GSR = "DISABLED";
    LUT4 mux_206_Mux_7_i956_3_lut_3_lut_4_lut (.A(n29143), .B(index_i[4]), 
         .C(n924_adj_3444), .D(index_i[5]), .Z(n956)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_7_i956_3_lut_3_lut_4_lut.init = 16'h11f0;
    PFUMX i22491 (.BLUT(n24977), .ALUT(n24978), .C0(index_q[5]), .Z(n24992));
    LUT4 mux_206_Mux_10_i701_4_lut_4_lut (.A(n29143), .B(index_i[4]), .C(index_i[5]), 
         .D(n29064), .Z(n701_adj_3095)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B (C (D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_10_i701_4_lut_4_lut.init = 16'h3efe;
    FD1S3DX o_val_pipeline_i_1__i3 (.D(\o_val_pipeline_i[0] [2]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(o_sample_i[2])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i3.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i2 (.D(\o_val_pipeline_i[0] [1]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(o_sample_i[1])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_i_1__i2.GSR = "DISABLED";
    LUT4 mux_206_Mux_3_i349_3_lut_3_lut (.A(index_i[1]), .B(index_i[4]), 
         .C(n348_adj_3331), .Z(n349_adj_3108)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_3_i349_3_lut_3_lut.init = 16'hd1d1;
    FD1S3BX quarter_wave_sample_register_q_i14 (.D(quarter_wave_sample_register_q_15__N_1783[14]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_q[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_q_i14.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i13 (.D(quarter_wave_sample_register_q_15__N_1783[13]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_q[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_q_i13.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i12 (.D(quarter_wave_sample_register_q_15__N_1783[12]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_q[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_q_i12.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i11 (.D(quarter_wave_sample_register_q_15__N_1783[11]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_q[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_q_i11.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i10 (.D(quarter_wave_sample_register_q_15__N_1783[10]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_q[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_q_i10.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i9 (.D(quarter_wave_sample_register_q_15__N_1783[9]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_q[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_q_i9.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i8 (.D(quarter_wave_sample_register_q_15__N_1783[8]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_q[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_q_i8.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i7 (.D(quarter_wave_sample_register_q_15__N_1783[7]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_q[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_q_i7.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i6 (.D(quarter_wave_sample_register_q_15__N_1783[6]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_q[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_q_i6.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i5 (.D(quarter_wave_sample_register_q_15__N_1783[5]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_q[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_q_i5.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i4 (.D(quarter_wave_sample_register_q_15__N_1783[4]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_q[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_q_i4.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i3 (.D(quarter_wave_sample_register_q_15__N_1783[3]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_q[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_q_i3.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i2 (.D(quarter_wave_sample_register_q_15__N_1783[2]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_q[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_q_i2.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i1 (.D(quarter_wave_sample_register_q_15__N_1783[1]), 
            .CK(dac_clk_p_c), .PD(i_sw0_c), .Q(quarter_wave_sample_register_q[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam quarter_wave_sample_register_q_i1.GSR = "DISABLED";
    FD1S3DX index_q_i9 (.D(index_q_9__N_1758[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(index_q[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam index_q_i9.GSR = "DISABLED";
    LUT4 i13849_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(n29329), .C(index_i[4]), 
         .D(index_i[0]), .Z(n16258)) /* synthesis lut_function=(!(A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i13849_3_lut_4_lut_4_lut_4_lut.init = 16'h55d5;
    FD1S3DX index_q_i8 (.D(index_q_9__N_1758[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(index_q[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam index_q_i8.GSR = "DISABLED";
    FD1S3DX index_q_i7 (.D(index_q_9__N_1758[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(index_q[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam index_q_i7.GSR = "DISABLED";
    FD1S3DX index_q_i6 (.D(index_q_9__N_1758[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(index_q[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam index_q_i6.GSR = "DISABLED";
    FD1S3DX index_q_i5 (.D(index_q_9__N_1758[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(index_q[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam index_q_i5.GSR = "DISABLED";
    FD1S3DX index_q_i4 (.D(index_q_9__N_1758[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(index_q[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam index_q_i4.GSR = "DISABLED";
    FD1S3DX index_q_i3 (.D(index_q_9__N_1758[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(index_q[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam index_q_i3.GSR = "DISABLED";
    FD1S3DX index_q_i2 (.D(index_q_9__N_1758[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(index_q[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam index_q_i2.GSR = "DISABLED";
    LUT4 n572_bdd_3_lut_26956_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n27508)) /* synthesis lut_function=(A (B (C+(D)))+!A (B ((D)+!C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n572_bdd_3_lut_26956_4_lut.init = 16'hcc94;
    FD1S3DX index_q_i1 (.D(index_q_9__N_1758[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(index_q[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam index_q_i1.GSR = "DISABLED";
    FD1S3DX index_i_i9 (.D(index_i_9__N_1748[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(index_i[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam index_i_i9.GSR = "DISABLED";
    FD1S3DX index_i_i8 (.D(index_i_9__N_1748[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(index_i[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam index_i_i8.GSR = "DISABLED";
    FD1S3DX index_i_i7 (.D(index_i_9__N_1748[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(index_i[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam index_i_i7.GSR = "DISABLED";
    FD1S3DX index_i_i6 (.D(index_i_9__N_1748[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(index_i[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam index_i_i6.GSR = "DISABLED";
    FD1S3DX index_i_i5 (.D(index_i_9__N_1748[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(index_i[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam index_i_i5.GSR = "DISABLED";
    FD1S3DX index_i_i4 (.D(index_i_9__N_1748[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(index_i[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam index_i_i4.GSR = "DISABLED";
    FD1S3DX index_i_i3 (.D(index_i_9__N_1748[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(index_i[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam index_i_i3.GSR = "DISABLED";
    FD1S3DX index_i_i2 (.D(index_i_9__N_1748[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(index_i[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam index_i_i2.GSR = "DISABLED";
    FD1S3DX index_i_i1 (.D(index_i_9__N_1748[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(index_i[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam index_i_i1.GSR = "DISABLED";
    FD1S3DX phase_negation_q_i1 (.D(phase_negation_q[0]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(phase_negation_q[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam phase_negation_q_i1.GSR = "DISABLED";
    FD1S3DX phase_negation_i_i1 (.D(phase_negation_i[0]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(phase_negation_i[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam phase_negation_i_i1.GSR = "DISABLED";
    LUT4 mux_206_Mux_0_i187_3_lut_4_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .Z(n187)) /* synthesis lut_function=(!(A (B)+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i187_3_lut_4_lut_3_lut.init = 16'h7676;
    FD1S3DX o_val_pipeline_q_1__i32 (.D(n671[15]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_q[0] [15])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_q_1__i32.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i31 (.D(n671[14]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_q[0] [14])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_q_1__i31.GSR = "DISABLED";
    LUT4 index_q_1__bdd_4_lut_27097 (.A(index_q[1]), .B(index_q[3]), .C(index_q[0]), 
         .D(index_q[2]), .Z(n29502)) /* synthesis lut_function=(!(A (B (D)+!B (C))+!A (B (C+!(D))+!B !(C+!(D))))) */ ;
    defparam index_q_1__bdd_4_lut_27097.init = 16'h169b;
    LUT4 mux_206_Mux_3_i684_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[4]), .Z(n684_adj_3406)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A !(B ((D)+!C)+!B (C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_3_i684_3_lut_3_lut_4_lut.init = 16'h5594;
    LUT4 mux_206_Mux_4_i205_3_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[3]), 
         .C(index_i[2]), .D(index_i[0]), .Z(n205_adj_3426)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(D))+!A (B (C (D)+!C !(D))+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_4_i205_3_lut_4_lut_4_lut.init = 16'h37c0;
    FD1S3DX o_val_pipeline_q_1__i30 (.D(n671[13]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_q[0] [13])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_q_1__i30.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i29 (.D(n671[12]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_q[0] [12])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_q_1__i29.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i28 (.D(n671[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_q[0] [11])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_q_1__i28.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i27 (.D(n671[10]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_q[0] [10])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_q_1__i27.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i26 (.D(n671[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_q[0] [9])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_q_1__i26.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i25 (.D(n671[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_q[0] [8])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_q_1__i25.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i24 (.D(n671[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_q[0] [7])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_q_1__i24.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i23 (.D(n671[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_q[0] [6])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_q_1__i23.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i22 (.D(n671[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_q[0] [5])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_q_1__i22.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i21 (.D(n671[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_q[0] [4])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_q_1__i21.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i20 (.D(n671[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_q[0] [3])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_q_1__i20.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i19 (.D(n671[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_q[0] [2])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_q_1__i19.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i18 (.D(n671[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_q[0] [1])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_q_1__i18.GSR = "DISABLED";
    LUT4 mux_206_Mux_2_i653_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n653_adj_3424)) /* synthesis lut_function=(A (B (C+!(D))+!B !(D))+!A !(B (C+!(D))+!B !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_2_i653_3_lut_4_lut.init = 16'h94aa;
    FD1S3DX o_val_pipeline_q_1__i17 (.D(n671[0]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(\o_val_pipeline_q[0] [0])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_q_1__i17.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i16 (.D(\o_val_pipeline_q[0] [15]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(o_sample_q[15])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_q_1__i16.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i15 (.D(\o_val_pipeline_q[0] [14]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(o_sample_q[14])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_q_1__i15.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i14 (.D(\o_val_pipeline_q[0] [13]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(o_sample_q[13])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_q_1__i14.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i13 (.D(\o_val_pipeline_q[0] [12]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(o_sample_q[12])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_q_1__i13.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i12 (.D(\o_val_pipeline_q[0] [11]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(o_sample_q[11])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_q_1__i12.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i11 (.D(\o_val_pipeline_q[0] [10]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(o_sample_q[10])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_q_1__i11.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i10 (.D(\o_val_pipeline_q[0] [9]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(o_sample_q[9])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_q_1__i10.GSR = "DISABLED";
    LUT4 mux_206_Mux_2_i348_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[3]), 
         .C(index_i[2]), .D(index_i[0]), .Z(n348_adj_3421)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_2_i348_3_lut_4_lut_4_lut_4_lut.init = 16'h34c3;
    FD1S3DX o_val_pipeline_q_1__i9 (.D(\o_val_pipeline_q[0] [8]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(o_sample_q[8])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_q_1__i9.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i8 (.D(\o_val_pipeline_q[0] [7]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(o_sample_q[7])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_q_1__i8.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i7 (.D(\o_val_pipeline_q[0] [6]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(o_sample_q[6])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_q_1__i7.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i6 (.D(\o_val_pipeline_q[0] [5]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(o_sample_q[5])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_q_1__i6.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i5 (.D(\o_val_pipeline_q[0] [4]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(o_sample_q[4])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_q_1__i5.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i4 (.D(\o_val_pipeline_q[0] [3]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(o_sample_q[3])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_q_1__i4.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i3 (.D(\o_val_pipeline_q[0] [2]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(o_sample_q[2])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_q_1__i3.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i2 (.D(\o_val_pipeline_q[0] [1]), .CK(dac_clk_p_c), 
            .CD(i_sw0_c), .Q(o_sample_q[1])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam o_val_pipeline_q_1__i2.GSR = "DISABLED";
    FD1P3AX phase_q__i11 (.D(phase_q_11__N_1874[11]), .SP(dac_clk_p_c_enable_630), 
            .CK(dac_clk_p_c), .Q(phase_q[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 90[6])
    defparam phase_q__i11.GSR = "DISABLED";
    LUT4 mux_206_Mux_12_i254_4_lut (.A(n29047), .B(n22332), .C(index_i[6]), 
         .D(n29180), .Z(n254_adj_3460)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_12_i254_4_lut.init = 16'hca0a;
    LUT4 mux_206_Mux_6_i636_4_lut_4_lut (.A(index_i[1]), .B(index_i[4]), 
         .C(n635_adj_3441), .D(n16259), .Z(n636_adj_3469)) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_6_i636_4_lut_4_lut.init = 16'hf3d1;
    LUT4 i12574_3_lut_3_lut_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[0]), 
         .Z(n619)) /* synthesis lut_function=(!(A ((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12574_3_lut_3_lut_3_lut.init = 16'h5d5d;
    LUT4 mux_207_Mux_8_i542_3_lut_4_lut (.A(n29370), .B(index_q[3]), .C(index_q[4]), 
         .D(n526_adj_3247), .Z(n542_adj_3422)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_8_i542_3_lut_4_lut.init = 16'h6f60;
    LUT4 n13568_bdd_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[4]), 
         .D(index_i[2]), .Z(n26900)) /* synthesis lut_function=(A (B)+!A !(B (D)+!B !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n13568_bdd_3_lut_4_lut.init = 16'h98cc;
    PFUMX i22813 (.BLUT(n557_adj_3239), .ALUT(n572_adj_3143), .C0(index_q[4]), 
          .Z(n25314));
    LUT4 i20854_3_lut_4_lut (.A(n29370), .B(index_q[3]), .C(index_q[4]), 
         .D(n635_adj_3255), .Z(n23336)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i20854_3_lut_4_lut.init = 16'hf606;
    LUT4 n800_bdd_3_lut_26605_4_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .Z(n28101)) /* synthesis lut_function=(!(A (B)+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n800_bdd_3_lut_26605_4_lut_3_lut.init = 16'h6262;
    LUT4 mux_206_Mux_0_i490_3_lut_4_lut_4_lut_3_lut_rep_745 (.A(index_i[1]), 
         .B(index_i[2]), .C(index_i[0]), .Z(n29405)) /* synthesis lut_function=(!(A (B+(C))+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i490_3_lut_4_lut_4_lut_3_lut_rep_745.init = 16'h4242;
    LUT4 mux_206_Mux_0_i212_3_lut_rep_746 (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .Z(n29406)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i212_3_lut_rep_746.init = 16'h6464;
    LUT4 mux_206_Mux_0_i29_3_lut_rep_748 (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .Z(n29408)) /* synthesis lut_function=(A (B (C))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i29_3_lut_rep_748.init = 16'h9191;
    L6MUX21 i25737 (.D0(n27487), .D1(n27485), .SD(index_i[4]), .Z(n27488));
    PFUMX i25735 (.BLUT(n29089), .ALUT(n27486), .C0(index_i[5]), .Z(n27487));
    LUT4 mux_206_Mux_3_i859_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n859_adj_3172)) /* synthesis lut_function=(!(A (B (D)+!B !(D))+!A (B (C+(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_3_i859_3_lut_3_lut_4_lut.init = 16'h339c;
    LUT4 mux_206_Mux_0_i14_3_lut_rep_749 (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .Z(n29409)) /* synthesis lut_function=(A (B)+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i14_3_lut_rep_749.init = 16'hd9d9;
    PFUMX i25733 (.BLUT(n27484), .ALUT(n27483), .C0(index_i[5]), .Z(n27485));
    LUT4 i1_2_lut_rep_719 (.A(index_i[1]), .B(index_i[0]), .Z(n29379)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_2_lut_rep_719.init = 16'heeee;
    LUT4 mux_206_Mux_0_i15_3_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .D(index_i[3]), .Z(n15_adj_3231)) /* synthesis lut_function=(A (B)+!A ((C (D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i15_3_lut_4_lut_4_lut.init = 16'hd999;
    LUT4 mux_206_Mux_8_i93_3_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .D(index_i[3]), .Z(n93_adj_3373)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(D))+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_8_i93_3_lut_3_lut_4_lut.init = 16'h3391;
    LUT4 i20631_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n23113)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A !(B (D)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20631_3_lut_3_lut_4_lut.init = 16'ha955;
    PFUMX i25717 (.BLUT(n27466), .ALUT(n27465), .C0(index_i[4]), .Z(n27467));
    LUT4 mux_206_Mux_7_i620_3_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .D(index_i[3]), .Z(n620_adj_3416)) /* synthesis lut_function=(A (B (C+!(D)))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_7_i620_3_lut_4_lut_4_lut.init = 16'h9199;
    L6MUX21 i25713 (.D0(n27463), .D1(n27461), .SD(index_i[5]), .Z(n27464));
    LUT4 mux_207_Mux_6_i635_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n635_adj_3388)) /* synthesis lut_function=(A (B (C+(D))+!B !(D))+!A (B)) */ ;
    defparam mux_207_Mux_6_i635_3_lut_4_lut.init = 16'hcce6;
    PFUMX i25711 (.BLUT(n27462), .ALUT(n285), .C0(index_i[4]), .Z(n27463));
    LUT4 mux_206_Mux_3_i397_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n397_adj_3433)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !(B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_3_i397_3_lut_4_lut_4_lut.init = 16'ha95a;
    PFUMX i25709 (.BLUT(n875_adj_3033), .ALUT(n27460), .C0(index_i[4]), 
          .Z(n27461));
    LUT4 i20655_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n23137)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C))+!A !(B ((D)+!C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20655_3_lut_4_lut_4_lut.init = 16'h925a;
    LUT4 i12577_2_lut_rep_516_3_lut (.A(index_i[1]), .B(index_i[0]), .C(index_i[2]), 
         .Z(n29176)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12577_2_lut_rep_516_3_lut.init = 16'he0e0;
    LUT4 mux_206_Mux_3_i157_3_lut_3_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n157_adj_3248)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_3_i157_3_lut_3_lut_3_lut_4_lut.init = 16'h1ff0;
    LUT4 i14383_2_lut_rep_487_3_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n29147)) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i14383_2_lut_rep_487_3_lut_4_lut.init = 16'he000;
    LUT4 i24035_3_lut (.A(n924_adj_3445), .B(n955_adj_3267), .C(index_i[5]), 
         .Z(n25296)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24035_3_lut.init = 16'hcaca;
    LUT4 i20748_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[0]), 
         .D(index_i[3]), .Z(n23230)) /* synthesis lut_function=(!(A (B (D)+!B !(C+!(D)))+!A !(B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20748_3_lut_4_lut.init = 16'h64aa;
    LUT4 mux_206_Mux_0_i491_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .D(index_i[3]), .Z(n491_adj_3386)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !(B (C)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i491_3_lut_4_lut.init = 16'h42f0;
    PFUMX i20633 (.BLUT(n23113), .ALUT(n23114), .C0(index_i[4]), .Z(n23115));
    L6MUX21 i25669 (.D0(n27417), .D1(n27415), .SD(index_i[5]), .Z(n27418));
    LUT4 i24376_3_lut (.A(n26755), .B(n25285), .C(index_i[6]), .Z(n25299)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24376_3_lut.init = 16'hcaca;
    CCU2D unary_minus_27_add_3_7 (.A0(quarter_wave_sample_register_q[5]), 
          .B0(GND_net), .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_q[6]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n19708), .COUT(n19709), 
          .S0(o_val_pipeline_q_0__15__N_1831[5]), .S1(o_val_pipeline_q_0__15__N_1831[6]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(81[29:60])
    defparam unary_minus_27_add_3_7.INIT0 = 16'hf555;
    defparam unary_minus_27_add_3_7.INIT1 = 16'hf555;
    defparam unary_minus_27_add_3_7.INJECT1_0 = "NO";
    defparam unary_minus_27_add_3_7.INJECT1_1 = "NO";
    PFUMX i25667 (.BLUT(n572_adj_3430), .ALUT(n27416), .C0(index_i[4]), 
          .Z(n27417));
    PFUMX i25665 (.BLUT(n27414), .ALUT(n27413), .C0(index_i[4]), .Z(n27415));
    PFUMX i20723 (.BLUT(n23203), .ALUT(n23204), .C0(index_i[4]), .Z(n23205));
    LUT4 mux_207_Mux_1_i700_3_lut_4_lut (.A(n29285), .B(index_q[3]), .C(index_q[4]), 
         .D(n684_adj_2974), .Z(n700_adj_3342)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_1_i700_3_lut_4_lut.init = 16'hefe0;
    L6MUX21 i22828 (.D0(n25313), .D1(n25314), .SD(index_q[5]), .Z(n25329));
    L6MUX21 i22829 (.D0(n25315), .D1(n25316), .SD(index_q[5]), .Z(n25330));
    LUT4 mux_207_Mux_5_i781_3_lut_4_lut_4_lut_then_4_lut (.A(index_q[3]), 
         .B(index_q[0]), .C(index_q[4]), .D(index_q[2]), .Z(n29504)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_5_i781_3_lut_4_lut_4_lut_then_4_lut.init = 16'hece0;
    L6MUX21 i22830 (.D0(n25317), .D1(n25318), .SD(index_q[5]), .Z(n25331));
    L6MUX21 i22831 (.D0(n25319), .D1(n25320), .SD(index_q[5]), .Z(n25332));
    PFUMX i22814 (.BLUT(n589), .ALUT(n604), .C0(index_q[4]), .Z(n25315));
    LUT4 mux_207_Mux_0_i660_3_lut_rep_835 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n32036)) /* synthesis lut_function=(A (B)+!A (B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_0_i660_3_lut_rep_835.init = 16'hc9c9;
    L6MUX21 i22832 (.D0(n25321), .D1(n25322), .SD(index_q[5]), .Z(n25333));
    L6MUX21 i22833 (.D0(n25323), .D1(n25324), .SD(index_q[5]), .Z(n25334));
    LUT4 mux_207_Mux_5_i781_3_lut_4_lut_4_lut_else_4_lut (.A(index_q[3]), 
         .B(index_q[0]), .C(index_q[4]), .Z(n29503)) /* synthesis lut_function=(!(A (C)+!A (B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_5_i781_3_lut_4_lut_4_lut_else_4_lut.init = 16'h1f1f;
    PFUMX i22815 (.BLUT(n620_adj_3001), .ALUT(n635_adj_3449), .C0(index_q[4]), 
          .Z(n25316));
    L6MUX21 i22834 (.D0(n25325), .D1(n25326), .SD(index_q[5]), .Z(n25335));
    LUT4 i20662_3_lut (.A(n498), .B(n32024), .C(index_i[3]), .Z(n23144)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20662_3_lut.init = 16'hcaca;
    L6MUX21 i22835 (.D0(n25327), .D1(n25328), .SD(index_q[5]), .Z(n25336));
    LUT4 i24058_3_lut (.A(n286_adj_3435), .B(n317_adj_3442), .C(index_q[5]), 
         .Z(n25237)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24058_3_lut.init = 16'hcaca;
    L6MUX21 i22492 (.D0(n24979), .D1(n24980), .SD(index_q[5]), .Z(n24993));
    PFUMX i22816 (.BLUT(n653_adj_2997), .ALUT(n668_adj_3439), .C0(index_q[4]), 
          .Z(n25317));
    LUT4 i20944_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n23426)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C+(D)))+!A (B (C)+!B !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i20944_3_lut_4_lut_4_lut.init = 16'hc95a;
    LUT4 i23898_3_lut (.A(n23140), .B(n23141), .C(index_i[4]), .Z(n23142)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23898_3_lut.init = 16'hcaca;
    LUT4 i20656_3_lut (.A(n32024), .B(n29427), .C(index_i[3]), .Z(n23138)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20656_3_lut.init = 16'hcaca;
    LUT4 i23900_3_lut (.A(n23137), .B(n23138), .C(index_i[4]), .Z(n23139)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23900_3_lut.init = 16'hcaca;
    PFUMX i22817 (.BLUT(n684_adj_2980), .ALUT(n699_adj_3240), .C0(index_q[4]), 
          .Z(n25318));
    LUT4 i23903_3_lut (.A(n23134), .B(n23135), .C(index_i[4]), .Z(n23136)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i23903_3_lut.init = 16'hcaca;
    PFUMX i22753 (.BLUT(n844_adj_3454), .ALUT(n13317), .C0(index_i[4]), 
          .Z(n25254));
    LUT4 i14202_2_lut_rep_707 (.A(index_q[1]), .B(index_q[2]), .Z(n29367)) /* synthesis lut_function=(A (B)) */ ;
    defparam i14202_2_lut_rep_707.init = 16'h8888;
    LUT4 i14213_2_lut_rep_758 (.A(index_i[1]), .B(index_i[2]), .Z(n29418)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14213_2_lut_rep_758.init = 16'heeee;
    PFUMX i22822 (.BLUT(n844_adj_3410), .ALUT(n13331), .C0(index_q[4]), 
          .Z(n25323));
    LUT4 i22310_3_lut (.A(n29470), .B(n29472), .C(index_q[3]), .Z(n24811)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22310_3_lut.init = 16'hcaca;
    LUT4 i24067_3_lut (.A(n924_adj_3417), .B(n955), .C(index_q[5]), .Z(n25205)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24067_3_lut.init = 16'hcaca;
    LUT4 i13084_2_lut_rep_530_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[0]), 
         .Z(n29190)) /* synthesis lut_function=(A (C)+!A ((C)+!B)) */ ;
    defparam i13084_2_lut_rep_530_3_lut.init = 16'hf1f1;
    LUT4 i22309_3_lut (.A(n29373), .B(n29316), .C(index_q[3]), .Z(n24810)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22309_3_lut.init = 16'hcaca;
    LUT4 mux_206_Mux_0_i333_3_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n333_adj_3375)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i333_3_lut_3_lut_4_lut.init = 16'hf10e;
    LUT4 mux_206_Mux_9_i93_3_lut_3_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .Z(n93_adj_3278)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B !(C))) */ ;
    defparam mux_206_Mux_9_i93_3_lut_3_lut_3_lut.init = 16'hc1c1;
    LUT4 i22307_3_lut (.A(n29472), .B(n29181), .C(index_q[3]), .Z(n24808)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22307_3_lut.init = 16'hcaca;
    LUT4 i14161_2_lut (.A(index_q[1]), .B(index_q[3]), .Z(n541)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i14161_2_lut.init = 16'h1111;
    LUT4 i21519_3_lut_4_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n24001)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B (C+!(D))))) */ ;
    defparam i21519_3_lut_4_lut_3_lut_4_lut.init = 16'h0fe0;
    LUT4 mux_207_Mux_4_i93_3_lut_4_lut_3_lut_rep_623_4_lut (.A(index_q[1]), 
         .B(index_q[2]), .C(index_q[3]), .D(index_q[0]), .Z(n29283)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D)))) */ ;
    defparam mux_207_Mux_4_i93_3_lut_4_lut_3_lut_rep_623_4_lut.init = 16'h07f0;
    PFUMX i25018 (.BLUT(n26660), .ALUT(n29317), .C0(index_q[5]), .Z(n26661));
    LUT4 mux_206_Mux_4_i236_3_lut_4_lut_3_lut_rep_662_4_lut (.A(index_i[1]), 
         .B(index_i[2]), .C(index_i[3]), .D(index_i[0]), .Z(n29322)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B (C+!(D)))) */ ;
    defparam mux_206_Mux_4_i236_3_lut_4_lut_3_lut_rep_662_4_lut.init = 16'hf01f;
    LUT4 mux_207_Mux_0_i526_3_lut (.A(n29335), .B(n29395), .C(index_q[3]), 
         .Z(n526_adj_2940)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_0_i526_3_lut.init = 16'hcaca;
    LUT4 mux_206_Mux_8_i412_3_lut_4_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .Z(n16744)) /* synthesis lut_function=(A (B+!(C))+!A !((C)+!B)) */ ;
    defparam mux_206_Mux_8_i412_3_lut_4_lut_3_lut.init = 16'h8e8e;
    LUT4 mux_206_Mux_0_i812_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n812_adj_3467)) /* synthesis lut_function=(A (B (C+(D))+!B !(C))+!A (B (D)+!B !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i812_3_lut_4_lut_4_lut_4_lut.init = 16'hcf92;
    LUT4 i24382_3_lut (.A(n26661), .B(n25194), .C(index_q[6]), .Z(n25208)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i24382_3_lut.init = 16'hcaca;
    LUT4 i21460_3_lut_3_lut_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[3]), 
         .Z(n23942)) /* synthesis lut_function=(A (C)+!A (B+!(C))) */ ;
    defparam i21460_3_lut_3_lut_3_lut.init = 16'he5e5;
    PFUMX i22818 (.BLUT(n716_adj_2995), .ALUT(n731_adj_2998), .C0(index_q[4]), 
          .Z(n25319));
    LUT4 i12841_2_lut_rep_518_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[3]), 
         .Z(n29178)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i12841_2_lut_rep_518_3_lut.init = 16'he0e0;
    PFUMX i25016 (.BLUT(n29386), .ALUT(n26658), .C0(index_q[2]), .Z(n26659));
    LUT4 n459_bdd_3_lut_25483 (.A(n32056), .B(n29385), .C(index_i[3]), 
         .Z(n27191)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n459_bdd_3_lut_25483.init = 16'hcaca;
    LUT4 i12842_2_lut_rep_427_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[4]), .D(index_i[3]), .Z(n29087)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i12842_2_lut_rep_427_3_lut_4_lut.init = 16'hfef0;
    LUT4 n236_bdd_3_lut_26448_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[4]), .D(index_i[3]), .Z(n28360)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C+(D)))+!A (B (C (D)+!C !(D))+!B !(C))) */ ;
    defparam n236_bdd_3_lut_26448_4_lut_4_lut_4_lut.init = 16'hc10f;
    PFUMX i22819 (.BLUT(n747_adj_2988), .ALUT(n762_adj_3263), .C0(index_q[4]), 
          .Z(n25320));
    LUT4 i24413_3_lut_rep_376_4_lut (.A(n29099), .B(index_q[5]), .C(index_q[8]), 
         .D(n1021_adj_3218), .Z(n29036)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i24413_3_lut_rep_376_4_lut.init = 16'hf808;
    PFUMX i27352 (.BLUT(n29901), .ALUT(n29900), .C0(index_q[3]), .Z(n29902));
    LUT4 mux_207_Mux_0_i142_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n142_adj_3364)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C))+!A !(B (C (D)+!C !(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam mux_207_Mux_0_i142_3_lut_4_lut_4_lut.init = 16'ha569;
    LUT4 mux_206_Mux_1_i923_3_lut_4_lut_3_lut_rep_759 (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .Z(n29419)) /* synthesis lut_function=(!(A (B (C))+!A !(B+(C)))) */ ;
    defparam mux_206_Mux_1_i923_3_lut_4_lut_3_lut_rep_759.init = 16'h7e7e;
    LUT4 i11140_2_lut_3_lut (.A(index_q[1]), .B(index_q[2]), .C(index_q[3]), 
         .Z(n13436)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i11140_2_lut_3_lut.init = 16'h8080;
    LUT4 mux_206_Mux_4_i158_3_lut (.A(n142_adj_3429), .B(n157_adj_3453), 
         .C(index_i[4]), .Z(n158)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_4_i158_3_lut.init = 16'hcaca;
    L6MUX21 i27356 (.D0(n29905), .D1(n29902), .SD(index_q[5]), .Z(n29906));
    PFUMX i20726 (.BLUT(n23206), .ALUT(n23207), .C0(index_i[4]), .Z(n23208));
    PFUMX i27098 (.BLUT(n29520), .ALUT(n29521), .C0(index_i[1]), .Z(n29522));
    LUT4 i20683_3_lut_4_lut_3_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .D(index_q[0]), .Z(n23165)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D))) */ ;
    defparam i20683_3_lut_4_lut_3_lut_4_lut.init = 16'hf80f;
    PFUMX i25640 (.BLUT(n27390), .ALUT(n27389), .C0(index_q[4]), .Z(n27391));
    LUT4 n16806_bdd_3_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[3]), 
         .D(index_i[5]), .Z(n28341)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A (B (C (D))+!B (C (D)+!C !(D))))) */ ;
    defparam n16806_bdd_3_lut_3_lut_4_lut.init = 16'h0f7e;
    LUT4 i12487_2_lut_rep_760 (.A(index_i[0]), .B(index_i[1]), .Z(n29420)) /* synthesis lut_function=((B)+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12487_2_lut_rep_760.init = 16'hdddd;
    LUT4 i20761_3_lut (.A(n29429), .B(n29446), .C(index_i[3]), .Z(n23243)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20761_3_lut.init = 16'hcaca;
    LUT4 i12654_2_lut_rep_476_3_lut (.A(index_q[1]), .B(index_q[2]), .C(index_q[3]), 
         .Z(n29136)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam i12654_2_lut_rep_476_3_lut.init = 16'hf8f8;
    LUT4 i17661_3_lut_4_lut_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .D(index_q[0]), .Z(n19975)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C (D)+!C !(D)))+!A !(B (D)+!B (C (D)+!C !(D)))) */ ;
    defparam i17661_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'h83fc;
    LUT4 i1_3_lut_4_lut_adj_190 (.A(index_q[1]), .B(index_q[2]), .C(index_q[5]), 
         .D(n29369), .Z(n22170)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;
    defparam i1_3_lut_4_lut_adj_190.init = 16'hfff8;
    LUT4 i13048_2_lut_rep_505_3_lut (.A(index_q[1]), .B(index_q[2]), .C(index_q[0]), 
         .Z(n29165)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i13048_2_lut_rep_505_3_lut.init = 16'h8080;
    PFUMX i27354 (.BLUT(n29904), .ALUT(n29903), .C0(index_q[3]), .Z(n29905));
    LUT4 i13837_2_lut_rep_452_2_lut_3_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[0]), .Z(n29112)) /* synthesis lut_function=(A (B+!(C))+!A !(C)) */ ;
    defparam i13837_2_lut_rep_452_2_lut_3_lut.init = 16'h8f8f;
    L6MUX21 i25014 (.D0(n26656), .D1(n26653), .SD(index_q[5]), .Z(n26657));
    LUT4 mux_206_Mux_0_i635_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n635_adj_3462)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i635_3_lut_4_lut_4_lut.init = 16'hfd0a;
    LUT4 mux_207_Mux_9_i30_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[0]), .D(index_q[3]), .Z(n30)) /* synthesis lut_function=(A (B (C (D))+!B !(D))+!A !(B+(D))) */ ;
    defparam mux_207_Mux_9_i30_3_lut_4_lut_4_lut_4_lut.init = 16'h8033;
    LUT4 mux_206_Mux_0_i316_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n316_adj_3181)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+(D)))+!A (B (C+(D))+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i316_3_lut_4_lut_4_lut_4_lut.init = 16'h332d;
    LUT4 mux_207_Mux_8_i491_3_lut_3_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .D(index_q[0]), .Z(n491_adj_3345)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A !(C))) */ ;
    defparam mux_207_Mux_8_i491_3_lut_3_lut_4_lut.init = 16'h7870;
    PFUMX i25012 (.BLUT(n26655), .ALUT(n475_adj_3165), .C0(index_q[4]), 
          .Z(n26656));
    LUT4 i20904_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n23386)) /* synthesis lut_function=(A (B (D)+!B ((D)+!C))+!A (B (D)+!B (C+!(D)))) */ ;
    defparam i20904_3_lut_4_lut_4_lut_4_lut.init = 16'hfe13;
    PFUMX i25638 (.BLUT(n27387), .ALUT(n27386), .C0(index_i[4]), .Z(n27388));
    LUT4 i12568_2_lut_rep_408_3_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .D(index_q[0]), .Z(n29068)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;
    defparam i12568_2_lut_rep_408_3_lut_4_lut.init = 16'hf8f0;
    LUT4 i20875_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[0]), .D(index_q[3]), .Z(n23357)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(D))+!A (B+!(D)))) */ ;
    defparam i20875_3_lut_4_lut_4_lut_4_lut.init = 16'h3380;
    LUT4 n698_bdd_3_lut_25761_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n27510)) /* synthesis lut_function=(A (B (C+(D))+!B ((D)+!C))+!A !(B (C+(D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n698_bdd_3_lut_25761_4_lut.init = 16'haa96;
    LUT4 i20611_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .D(index_q[0]), .Z(n23093)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C (D)+!C !(D)))+!A !(B (D)+!B (C (D)+!C !(D))))) */ ;
    defparam i20611_3_lut_4_lut_4_lut_4_lut.init = 16'h7c03;
    LUT4 mux_206_Mux_0_i762_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n762_adj_3464)) /* synthesis lut_function=(A (B+!((D)+!C))+!A !(B (D)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i762_3_lut_4_lut_4_lut.init = 16'h98fc;
    LUT4 mux_207_Mux_3_i142_3_lut_3_lut_3_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .Z(n142_adj_3168)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B+!(C)))) */ ;
    defparam mux_207_Mux_3_i142_3_lut_3_lut_3_lut.init = 16'h3838;
    LUT4 i13045_2_lut_rep_708 (.A(index_q[1]), .B(index_q[2]), .C(index_q[0]), 
         .Z(n29368)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam i13045_2_lut_rep_708.init = 16'h7070;
    PFUMX i25009 (.BLUT(n26652), .ALUT(n23195), .C0(index_q[4]), .Z(n26653));
    LUT4 mux_207_Mux_0_i1017_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[0]), .D(index_q[3]), .Z(n1017_adj_3167)) /* synthesis lut_function=(A (B (D)+!B !((D)+!C))+!A (C+(D))) */ ;
    defparam mux_207_Mux_0_i1017_4_lut_4_lut_4_lut.init = 16'hdd70;
    LUT4 i12711_2_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[0]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n635_adj_3350)) /* synthesis lut_function=(A (C+!(D))+!A (B (C)+!B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12711_2_lut_4_lut_4_lut.init = 16'hf1fa;
    LUT4 i7699_2_lut_rep_709 (.A(index_q[3]), .B(index_q[4]), .Z(n29369)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i7699_2_lut_rep_709.init = 16'heeee;
    LUT4 i11124_3_lut_3_lut_4_lut (.A(index_q[3]), .B(index_q[4]), .C(n29395), 
         .D(index_q[0]), .Z(n605_adj_3276)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i11124_3_lut_3_lut_4_lut.init = 16'h10fe;
    LUT4 i1_3_lut_rep_439_4_lut (.A(index_q[3]), .B(index_q[4]), .C(index_q[2]), 
         .D(n29465), .Z(n29099)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(69[46:73])
    defparam i1_3_lut_rep_439_4_lut.init = 16'hfffe;
    LUT4 i20842_3_lut_then_4_lut (.A(index_q[4]), .B(index_q[1]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n29513)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)+!C !(D)))+!A !(B (C+!(D))+!B (C (D)+!C !(D))))) */ ;
    defparam i20842_3_lut_then_4_lut.init = 16'h5a65;
    LUT4 i21438_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n23920)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (D))+!A !(D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21438_3_lut_4_lut_4_lut_4_lut.init = 16'ha25d;
    LUT4 n773_bdd_3_lut_4_lut_4_lut_adj_191 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n26719)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n773_bdd_3_lut_4_lut_4_lut_adj_191.init = 16'ha5ad;
    LUT4 mux_206_Mux_0_i796_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n796_adj_3466)) /* synthesis lut_function=(A (B (C+(D))+!B (C (D)))+!A !(B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i796_3_lut_4_lut_4_lut.init = 16'hadc0;
    LUT4 mux_206_Mux_5_i475_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n475_adj_3456)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_5_i475_3_lut_4_lut_4_lut.init = 16'hd4a5;
    LUT4 i14189_2_lut_rep_710 (.A(index_q[1]), .B(index_q[2]), .Z(n29370)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i14189_2_lut_rep_710.init = 16'heeee;
    LUT4 mux_206_Mux_0_i157_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n157_adj_3363)) /* synthesis lut_function=(A (B (C+!(D))+!B !(D))+!A (B (D)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i157_3_lut_4_lut.init = 16'hd4aa;
    LUT4 i3986_2_lut_rep_762 (.A(index_i[0]), .B(index_i[2]), .Z(n29422)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i3986_2_lut_rep_762.init = 16'h6666;
    PFUMX i25626 (.BLUT(n27373), .ALUT(n27372), .C0(index_i[4]), .Z(n476_adj_3244));
    LUT4 n557_bdd_3_lut_26376_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[4]), .D(index_q[3]), .Z(n28281)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C+(D)))+!A (B (C (D)+!C !(D))+!B !(C))) */ ;
    defparam n557_bdd_3_lut_26376_4_lut_4_lut_4_lut.init = 16'hc10f;
    LUT4 mux_206_Mux_1_i62_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[4]), .D(index_i[3]), .Z(n62_adj_3455)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))+!A !(B (C)+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_1_i62_3_lut_4_lut_4_lut.init = 16'ha5a6;
    LUT4 i20610_3_lut_4_lut_3_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .D(index_q[0]), .Z(n23092)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B (C+!(D))))) */ ;
    defparam i20610_3_lut_4_lut_3_lut_4_lut.init = 16'h0fe0;
    LUT4 mux_207_Mux_4_i236_3_lut_4_lut_4_lut_3_lut_rep_621_4_lut (.A(index_q[1]), 
         .B(index_q[2]), .C(index_q[3]), .D(index_q[0]), .Z(n29281)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B (C+!(D)))) */ ;
    defparam mux_207_Mux_4_i236_3_lut_4_lut_4_lut_3_lut_rep_621_4_lut.init = 16'hf01f;
    LUT4 mux_207_Mux_9_i412_3_lut_4_lut_3_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .Z(n412_adj_3335)) /* synthesis lut_function=(!(A (B (C))+!A !(B+(C)))) */ ;
    defparam mux_207_Mux_9_i412_3_lut_4_lut_3_lut.init = 16'h7e7e;
    LUT4 mux_206_Mux_6_i572_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n572_adj_3451)) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_6_i572_3_lut_4_lut.init = 16'hccd9;
    PFUMX i17669 (.BLUT(n19981), .ALUT(n19982), .C0(index_q[4]), .Z(n19983));
    L6MUX21 i25007 (.D0(n26650), .D1(n26648), .SD(index_q[5]), .Z(n26651));
    PFUMX i25005 (.BLUT(n26649), .ALUT(n285_adj_3025), .C0(index_q[4]), 
          .Z(n26650));
    PFUMX i25003 (.BLUT(n26647), .ALUT(n26646), .C0(index_q[4]), .Z(n26648));
    L6MUX21 i25000 (.D0(n26644), .D1(n26641), .SD(index_q[5]), .Z(n26645));
    PFUMX i24998 (.BLUT(n15_adj_3339), .ALUT(n26642), .C0(index_q[4]), 
          .Z(n26644));
    LUT4 i12588_2_lut_rep_506_3_lut (.A(index_q[1]), .B(index_q[2]), .C(index_q[3]), 
         .Z(n29166)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i12588_2_lut_rep_506_3_lut.init = 16'he0e0;
    LUT4 mux_206_Mux_0_i142_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n142_adj_3362)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C))+!A !(B (C (D)+!C !(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_206_Mux_0_i142_3_lut_4_lut_4_lut.init = 16'ha569;
    LUT4 mux_207_Mux_2_i955_then_4_lut (.A(index_q[4]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n29507)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B (C+!(D))+!B !(C (D)))) */ ;
    defparam mux_207_Mux_2_i955_then_4_lut.init = 16'he95d;
    PFUMX i24995 (.BLUT(n26640), .ALUT(n26639), .C0(index_q[4]), .Z(n26641));
    PFUMX i17700 (.BLUT(n20012), .ALUT(n20013), .C0(index_i[4]), .Z(n20014));
    LUT4 mux_207_Mux_9_i93_3_lut_3_lut_3_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .Z(n93_adj_3443)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B !(C))) */ ;
    defparam mux_207_Mux_9_i93_3_lut_3_lut_3_lut.init = 16'hc1c1;
    LUT4 i13047_2_lut_rep_399_2_lut_3_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[0]), .Z(n29059)) /* synthesis lut_function=(A (C)+!A ((C)+!B)) */ ;
    defparam i13047_2_lut_rep_399_2_lut_3_lut.init = 16'hf1f1;
    LUT4 i12589_2_lut_rep_418_3_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[4]), .D(index_q[3]), .Z(n29078)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i12589_2_lut_rep_418_3_lut_4_lut.init = 16'hfef0;
    LUT4 mux_207_Mux_8_i412_3_lut_4_lut_3_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .Z(n16626)) /* synthesis lut_function=(A (B+!(C))+!A !((C)+!B)) */ ;
    defparam mux_207_Mux_8_i412_3_lut_4_lut_3_lut.init = 16'h8e8e;
    PFUMX i27094 (.BLUT(n29515), .ALUT(n29516), .C0(index_i[1]), .Z(n29517));
    LUT4 i21504_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n23986)) /* synthesis lut_function=(A (B (C (D))+!B !(C (D)))+!A !(B (D)+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21504_3_lut_4_lut_4_lut.init = 16'h9366;
    LUT4 i20947_3_lut_3_lut_3_lut (.A(index_q[1]), .B(index_q[2]), .C(index_q[3]), 
         .Z(n23429)) /* synthesis lut_function=(A (C)+!A (B+!(C))) */ ;
    defparam i20947_3_lut_3_lut_3_lut.init = 16'he5e5;
    
endmodule
//
// Verilog Description of module \nco(OW=12)_U23 
//

module \nco(OW=12)_U23  (o_phase, dac_clk_p_c, i_sw0_c, increment, GND_net) /* synthesis syn_module_defined=1 */ ;
    output [11:0]o_phase;
    input dac_clk_p_c;
    input i_sw0_c;
    input [30:0]increment;
    input GND_net;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[29:38])
    wire [31:0]n133;
    wire [31:0]n233;
    
    wire n19916, n19915, n19914, n19913, n19912, n19911, n19910, 
        n19909, n19908, n19907, n19906, n19905, n19904, n19903, 
        n19902;
    
    FD1S3DX phase_register_856__i31 (.D(n133[31]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_phase[11])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_856__i31.GSR = "DISABLED";
    FD1S3DX phase_register_856__i30 (.D(n133[30]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_phase[10])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_856__i30.GSR = "DISABLED";
    FD1S3DX phase_register_856__i29 (.D(n133[29]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_phase[9])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_856__i29.GSR = "DISABLED";
    FD1S3DX phase_register_856__i28 (.D(n133[28]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_phase[8])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_856__i28.GSR = "DISABLED";
    FD1S3DX phase_register_856__i27 (.D(n133[27]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_phase[7])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_856__i27.GSR = "DISABLED";
    FD1S3DX phase_register_856__i26 (.D(n133[26]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_phase[6])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_856__i26.GSR = "DISABLED";
    FD1S3DX phase_register_856__i25 (.D(n133[25]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_phase[5])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_856__i25.GSR = "DISABLED";
    FD1S3DX phase_register_856__i24 (.D(n133[24]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_phase[4])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_856__i24.GSR = "DISABLED";
    FD1S3DX phase_register_856__i23 (.D(n133[23]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_phase[3])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_856__i23.GSR = "DISABLED";
    FD1S3DX phase_register_856__i22 (.D(n133[22]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_phase[2])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_856__i22.GSR = "DISABLED";
    FD1S3DX phase_register_856__i21 (.D(n133[21]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_phase[1])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_856__i21.GSR = "DISABLED";
    FD1S3DX phase_register_856__i20 (.D(n133[20]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(o_phase[0])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_856__i20.GSR = "DISABLED";
    FD1S3DX phase_register_856__i19 (.D(n133[19]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[19])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_856__i19.GSR = "DISABLED";
    FD1S3DX phase_register_856__i18 (.D(n133[18]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[18])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_856__i18.GSR = "DISABLED";
    FD1S3DX phase_register_856__i17 (.D(n133[17]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[17])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_856__i17.GSR = "DISABLED";
    FD1S3DX phase_register_856__i16 (.D(n133[16]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[16])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_856__i16.GSR = "DISABLED";
    FD1S3DX phase_register_856__i15 (.D(n133[15]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[15])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_856__i15.GSR = "DISABLED";
    FD1S3DX phase_register_856__i14 (.D(n133[14]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[14])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_856__i14.GSR = "DISABLED";
    FD1S3DX phase_register_856__i13 (.D(n133[13]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[13])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_856__i13.GSR = "DISABLED";
    FD1S3DX phase_register_856__i12 (.D(n133[12]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[12])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_856__i12.GSR = "DISABLED";
    FD1S3DX phase_register_856__i11 (.D(n133[11]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[11])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_856__i11.GSR = "DISABLED";
    FD1S3DX phase_register_856__i10 (.D(n133[10]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[10])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_856__i10.GSR = "DISABLED";
    FD1S3DX phase_register_856__i9 (.D(n133[9]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[9])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_856__i9.GSR = "DISABLED";
    FD1S3DX phase_register_856__i8 (.D(n133[8]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[8])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_856__i8.GSR = "DISABLED";
    FD1S3DX phase_register_856__i7 (.D(n133[7]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[7])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_856__i7.GSR = "DISABLED";
    FD1S3DX phase_register_856__i6 (.D(n133[6]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[6])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_856__i6.GSR = "DISABLED";
    FD1S3DX phase_register_856__i5 (.D(n133[5]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[5])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_856__i5.GSR = "DISABLED";
    FD1S3DX phase_register_856__i4 (.D(n133[4]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[4])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_856__i4.GSR = "DISABLED";
    FD1S3DX phase_register_856__i3 (.D(n133[3]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[3])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_856__i3.GSR = "DISABLED";
    FD1S3DX phase_register_856__i2 (.D(n133[2]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[2])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_856__i2.GSR = "DISABLED";
    FD1S3DX phase_register_856__i1 (.D(n133[1]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[1])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_856__i1.GSR = "DISABLED";
    CCU2D phase_register_856_add_4_32 (.A0(increment[30]), .B0(o_phase[10]), 
          .C0(GND_net), .D0(GND_net), .A1(o_phase[11]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n19916), .S0(n133[30]), .S1(n133[31]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_856_add_4_32.INIT0 = 16'h5666;
    defparam phase_register_856_add_4_32.INIT1 = 16'hfaaa;
    defparam phase_register_856_add_4_32.INJECT1_0 = "NO";
    defparam phase_register_856_add_4_32.INJECT1_1 = "NO";
    CCU2D phase_register_856_add_4_30 (.A0(increment[28]), .B0(o_phase[8]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[29]), .B1(o_phase[9]), 
          .C1(GND_net), .D1(GND_net), .CIN(n19915), .COUT(n19916), .S0(n133[28]), 
          .S1(n133[29]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_856_add_4_30.INIT0 = 16'h5666;
    defparam phase_register_856_add_4_30.INIT1 = 16'h5666;
    defparam phase_register_856_add_4_30.INJECT1_0 = "NO";
    defparam phase_register_856_add_4_30.INJECT1_1 = "NO";
    CCU2D phase_register_856_add_4_28 (.A0(increment[26]), .B0(o_phase[6]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[27]), .B1(o_phase[7]), 
          .C1(GND_net), .D1(GND_net), .CIN(n19914), .COUT(n19915), .S0(n133[26]), 
          .S1(n133[27]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_856_add_4_28.INIT0 = 16'h5666;
    defparam phase_register_856_add_4_28.INIT1 = 16'h5666;
    defparam phase_register_856_add_4_28.INJECT1_0 = "NO";
    defparam phase_register_856_add_4_28.INJECT1_1 = "NO";
    CCU2D phase_register_856_add_4_26 (.A0(increment[24]), .B0(o_phase[4]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[25]), .B1(o_phase[5]), 
          .C1(GND_net), .D1(GND_net), .CIN(n19913), .COUT(n19914), .S0(n133[24]), 
          .S1(n133[25]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_856_add_4_26.INIT0 = 16'h5666;
    defparam phase_register_856_add_4_26.INIT1 = 16'h5666;
    defparam phase_register_856_add_4_26.INJECT1_0 = "NO";
    defparam phase_register_856_add_4_26.INJECT1_1 = "NO";
    CCU2D phase_register_856_add_4_24 (.A0(increment[22]), .B0(o_phase[2]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[23]), .B1(o_phase[3]), 
          .C1(GND_net), .D1(GND_net), .CIN(n19912), .COUT(n19913), .S0(n133[22]), 
          .S1(n133[23]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_856_add_4_24.INIT0 = 16'h5666;
    defparam phase_register_856_add_4_24.INIT1 = 16'h5666;
    defparam phase_register_856_add_4_24.INJECT1_0 = "NO";
    defparam phase_register_856_add_4_24.INJECT1_1 = "NO";
    CCU2D phase_register_856_add_4_22 (.A0(increment[20]), .B0(o_phase[0]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[21]), .B1(o_phase[1]), 
          .C1(GND_net), .D1(GND_net), .CIN(n19911), .COUT(n19912), .S0(n133[20]), 
          .S1(n133[21]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_856_add_4_22.INIT0 = 16'h5666;
    defparam phase_register_856_add_4_22.INIT1 = 16'h5666;
    defparam phase_register_856_add_4_22.INJECT1_0 = "NO";
    defparam phase_register_856_add_4_22.INJECT1_1 = "NO";
    CCU2D phase_register_856_add_4_20 (.A0(increment[18]), .B0(n233[18]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[19]), .B1(n233[19]), 
          .C1(GND_net), .D1(GND_net), .CIN(n19910), .COUT(n19911), .S0(n133[18]), 
          .S1(n133[19]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_856_add_4_20.INIT0 = 16'h5666;
    defparam phase_register_856_add_4_20.INIT1 = 16'h5666;
    defparam phase_register_856_add_4_20.INJECT1_0 = "NO";
    defparam phase_register_856_add_4_20.INJECT1_1 = "NO";
    CCU2D phase_register_856_add_4_18 (.A0(increment[16]), .B0(n233[16]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[17]), .B1(n233[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n19909), .COUT(n19910), .S0(n133[16]), 
          .S1(n133[17]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_856_add_4_18.INIT0 = 16'h5666;
    defparam phase_register_856_add_4_18.INIT1 = 16'h5666;
    defparam phase_register_856_add_4_18.INJECT1_0 = "NO";
    defparam phase_register_856_add_4_18.INJECT1_1 = "NO";
    CCU2D phase_register_856_add_4_16 (.A0(increment[14]), .B0(n233[14]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[15]), .B1(n233[15]), 
          .C1(GND_net), .D1(GND_net), .CIN(n19908), .COUT(n19909), .S0(n133[14]), 
          .S1(n133[15]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_856_add_4_16.INIT0 = 16'h5666;
    defparam phase_register_856_add_4_16.INIT1 = 16'h5666;
    defparam phase_register_856_add_4_16.INJECT1_0 = "NO";
    defparam phase_register_856_add_4_16.INJECT1_1 = "NO";
    CCU2D phase_register_856_add_4_14 (.A0(increment[12]), .B0(n233[12]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[13]), .B1(n233[13]), 
          .C1(GND_net), .D1(GND_net), .CIN(n19907), .COUT(n19908), .S0(n133[12]), 
          .S1(n133[13]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_856_add_4_14.INIT0 = 16'h5666;
    defparam phase_register_856_add_4_14.INIT1 = 16'h5666;
    defparam phase_register_856_add_4_14.INJECT1_0 = "NO";
    defparam phase_register_856_add_4_14.INJECT1_1 = "NO";
    CCU2D phase_register_856_add_4_12 (.A0(increment[10]), .B0(n233[10]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[11]), .B1(n233[11]), 
          .C1(GND_net), .D1(GND_net), .CIN(n19906), .COUT(n19907), .S0(n133[10]), 
          .S1(n133[11]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_856_add_4_12.INIT0 = 16'h5666;
    defparam phase_register_856_add_4_12.INIT1 = 16'h5666;
    defparam phase_register_856_add_4_12.INJECT1_0 = "NO";
    defparam phase_register_856_add_4_12.INJECT1_1 = "NO";
    CCU2D phase_register_856_add_4_10 (.A0(increment[8]), .B0(n233[8]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[9]), .B1(n233[9]), 
          .C1(GND_net), .D1(GND_net), .CIN(n19905), .COUT(n19906), .S0(n133[8]), 
          .S1(n133[9]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_856_add_4_10.INIT0 = 16'h5666;
    defparam phase_register_856_add_4_10.INIT1 = 16'h5666;
    defparam phase_register_856_add_4_10.INJECT1_0 = "NO";
    defparam phase_register_856_add_4_10.INJECT1_1 = "NO";
    CCU2D phase_register_856_add_4_8 (.A0(increment[6]), .B0(n233[6]), .C0(GND_net), 
          .D0(GND_net), .A1(increment[7]), .B1(n233[7]), .C1(GND_net), 
          .D1(GND_net), .CIN(n19904), .COUT(n19905), .S0(n133[6]), .S1(n133[7]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_856_add_4_8.INIT0 = 16'h5666;
    defparam phase_register_856_add_4_8.INIT1 = 16'h5666;
    defparam phase_register_856_add_4_8.INJECT1_0 = "NO";
    defparam phase_register_856_add_4_8.INJECT1_1 = "NO";
    CCU2D phase_register_856_add_4_6 (.A0(increment[4]), .B0(n233[4]), .C0(GND_net), 
          .D0(GND_net), .A1(increment[5]), .B1(n233[5]), .C1(GND_net), 
          .D1(GND_net), .CIN(n19903), .COUT(n19904), .S0(n133[4]), .S1(n133[5]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_856_add_4_6.INIT0 = 16'h5666;
    defparam phase_register_856_add_4_6.INIT1 = 16'h5666;
    defparam phase_register_856_add_4_6.INJECT1_0 = "NO";
    defparam phase_register_856_add_4_6.INJECT1_1 = "NO";
    CCU2D phase_register_856_add_4_4 (.A0(increment[2]), .B0(n233[2]), .C0(GND_net), 
          .D0(GND_net), .A1(increment[3]), .B1(n233[3]), .C1(GND_net), 
          .D1(GND_net), .CIN(n19902), .COUT(n19903), .S0(n133[2]), .S1(n133[3]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_856_add_4_4.INIT0 = 16'h5666;
    defparam phase_register_856_add_4_4.INIT1 = 16'h5666;
    defparam phase_register_856_add_4_4.INJECT1_0 = "NO";
    defparam phase_register_856_add_4_4.INJECT1_1 = "NO";
    LUT4 i17622_2_lut (.A(increment[0]), .B(n233[0]), .Z(n133[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i17622_2_lut.init = 16'h6666;
    CCU2D phase_register_856_add_4_2 (.A0(increment[0]), .B0(n233[0]), .C0(GND_net), 
          .D0(GND_net), .A1(increment[1]), .B1(n233[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n19902), .S1(n133[1]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_856_add_4_2.INIT0 = 16'h7000;
    defparam phase_register_856_add_4_2.INIT1 = 16'h5666;
    defparam phase_register_856_add_4_2.INJECT1_0 = "NO";
    defparam phase_register_856_add_4_2.INJECT1_1 = "NO";
    FD1S3DX phase_register_856__i0 (.D(n133[0]), .CK(dac_clk_p_c), .CD(i_sw0_c), 
            .Q(n233[0])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_856__i0.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module \txuartlite(TIMING_BITS=24,CLOCKS_PER_BAUD=10000) 
//

module \txuartlite(TIMING_BITS=24,CLOCKS_PER_BAUD=10000)  (dac_clk_p_c, o_wbu_uart_tx_c, 
            GND_net, tx_stb, tx_busy, \tx_data[0] , \tx_data[6] , 
            \tx_data[5] , \tx_data[4] , \tx_data[3] , \tx_data[2] , 
            \tx_data[1] , n32067) /* synthesis syn_module_defined=1 */ ;
    input dac_clk_p_c;
    output o_wbu_uart_tx_c;
    input GND_net;
    input tx_stb;
    output tx_busy;
    input \tx_data[0] ;
    input \tx_data[6] ;
    input \tx_data[5] ;
    input \tx_data[4] ;
    input \tx_data[3] ;
    input \tx_data[2] ;
    input \tx_data[1] ;
    input n32067;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[29:38])
    wire [7:0]lcl_data;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(84[12:20])
    
    wire dac_clk_p_c_enable_514;
    wire [7:0]lcl_data_7__N_278;
    
    wire zero_baud_counter, zero_baud_counter_N_292;
    wire [23:0]baud_counter;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(82[17:29])
    wire [23:0]baud_counter_23__N_250;
    
    wire n29211;
    wire [23:0]n133;
    
    wire n29096, zero_baud_counter_N_295;
    wire [23:0]n108;
    
    wire n29496, n29497;
    wire [3:0]state;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(83[12:17])
    
    wire n29498, n29493, n29494, n29495, n22612, n22602, n22616, 
        n29209, n19787, n29210, n29107, n19786, n19785, n19784, 
        n19783, n19782, n19781, n19780, n19779, n19778, n19777, 
        n19776, n12747;
    wire [3:0]n27;
    
    wire n22214, n22191, n22624, n22618, n22608, n22203, n9431, 
        n20035;
    
    FD1P3AY lcl_data_i0 (.D(lcl_data_7__N_278[0]), .SP(dac_clk_p_c_enable_514), 
            .CK(dac_clk_p_c), .Q(lcl_data[0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=7, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=69, LSE_RLINE=69 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(139[9] 143[40])
    defparam lcl_data_i0.GSR = "DISABLED";
    FD1S3AY zero_baud_counter_49 (.D(zero_baud_counter_N_292), .CK(dac_clk_p_c), 
            .Q(zero_baud_counter)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=7, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=69, LSE_RLINE=69 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam zero_baud_counter_49.GSR = "DISABLED";
    FD1S3AX baud_counter_i0 (.D(baud_counter_23__N_250[0]), .CK(dac_clk_p_c), 
            .Q(baud_counter[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=7, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=69, LSE_RLINE=69 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i0.GSR = "DISABLED";
    FD1P3IX o_uart_tx_48 (.D(lcl_data[0]), .SP(dac_clk_p_c_enable_514), 
            .CD(n29211), .CK(dac_clk_p_c), .Q(o_wbu_uart_tx_c)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=7, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=69, LSE_RLINE=69 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(154[9] 158[29])
    defparam o_uart_tx_48.GSR = "DISABLED";
    LUT4 baud_counter_23__I_9_i1_4_lut (.A(n29211), .B(n133[0]), .C(n29096), 
         .D(zero_baud_counter_N_295), .Z(baud_counter_23__N_250[0])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((C+(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(217[12] 224[43])
    defparam baud_counter_23__I_9_i1_4_lut.init = 16'ha0ac;
    LUT4 i12418_2_lut (.A(n108[0]), .B(zero_baud_counter), .Z(n133[0])) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(224[4:43])
    defparam i12418_2_lut.init = 16'heeee;
    PFUMX i27082 (.BLUT(n29496), .ALUT(n29497), .C0(state[3]), .Z(n29498));
    PFUMX i27080 (.BLUT(n29493), .ALUT(n29494), .C0(state[2]), .Z(n29495));
    LUT4 i1_4_lut (.A(baud_counter[14]), .B(baud_counter[15]), .C(baud_counter[18]), 
         .D(baud_counter[4]), .Z(n22612)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(207[24:43])
    defparam i1_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut (.A(baud_counter[20]), .B(baud_counter[19]), .Z(n22602)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(207[24:43])
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i1_4_lut_adj_172 (.A(baud_counter[21]), .B(baud_counter[5]), .C(baud_counter[7]), 
         .D(baud_counter[10]), .Z(n22616)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(207[24:43])
    defparam i1_4_lut_adj_172.init = 16'hfffe;
    LUT4 i1_2_lut_rep_549 (.A(state[0]), .B(state[3]), .Z(n29209)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_549.init = 16'h8888;
    CCU2D sub_36_add_2_25 (.A0(baud_counter[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n19787), .S0(n108[23]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_25.INIT0 = 16'h5555;
    defparam sub_36_add_2_25.INIT1 = 16'h0000;
    defparam sub_36_add_2_25.INJECT1_0 = "NO";
    defparam sub_36_add_2_25.INJECT1_1 = "NO";
    LUT4 i1_3_lut_rep_436_4_lut (.A(state[0]), .B(state[3]), .C(state[1]), 
         .D(state[2]), .Z(n29096)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_3_lut_rep_436_4_lut.init = 16'h8000;
    LUT4 i1_3_lut_4_lut (.A(state[0]), .B(state[3]), .C(zero_baud_counter), 
         .D(n29210), .Z(zero_baud_counter_N_295)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_3_lut_4_lut.init = 16'h0080;
    LUT4 i20552_2_lut_rep_550 (.A(state[1]), .B(state[2]), .Z(n29210)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i20552_2_lut_rep_550.init = 16'heeee;
    LUT4 i1237_3_lut_rep_447_4_lut (.A(state[1]), .B(state[2]), .C(state[0]), 
         .D(state[3]), .Z(n29107)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;
    defparam i1237_3_lut_rep_447_4_lut.init = 16'hfe00;
    LUT4 i_wr_I_0_2_lut_rep_551 (.A(tx_stb), .B(tx_busy), .Z(n29211)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(155[7:24])
    defparam i_wr_I_0_2_lut_rep_551.init = 16'h2222;
    CCU2D sub_36_add_2_23 (.A0(baud_counter[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n19786), .COUT(n19787), .S0(n108[21]), 
          .S1(n108[22]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_23.INIT0 = 16'h5555;
    defparam sub_36_add_2_23.INIT1 = 16'h5555;
    defparam sub_36_add_2_23.INJECT1_0 = "NO";
    defparam sub_36_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_36_add_2_21 (.A0(baud_counter[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n19785), .COUT(n19786), .S0(n108[19]), 
          .S1(n108[20]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_21.INIT0 = 16'h5555;
    defparam sub_36_add_2_21.INIT1 = 16'h5555;
    defparam sub_36_add_2_21.INJECT1_0 = "NO";
    defparam sub_36_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_36_add_2_19 (.A0(baud_counter[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n19784), .COUT(n19785), .S0(n108[17]), 
          .S1(n108[18]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_19.INIT0 = 16'h5555;
    defparam sub_36_add_2_19.INIT1 = 16'h5555;
    defparam sub_36_add_2_19.INJECT1_0 = "NO";
    defparam sub_36_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_36_add_2_17 (.A0(baud_counter[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n19783), .COUT(n19784), .S0(n108[15]), 
          .S1(n108[16]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_17.INIT0 = 16'h5555;
    defparam sub_36_add_2_17.INIT1 = 16'h5555;
    defparam sub_36_add_2_17.INJECT1_0 = "NO";
    defparam sub_36_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_36_add_2_15 (.A0(baud_counter[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n19782), .COUT(n19783), .S0(n108[13]), 
          .S1(n108[14]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_15.INIT0 = 16'h5555;
    defparam sub_36_add_2_15.INIT1 = 16'h5555;
    defparam sub_36_add_2_15.INJECT1_0 = "NO";
    defparam sub_36_add_2_15.INJECT1_1 = "NO";
    LUT4 lcl_data_7__I_0_i1_3_lut_4_lut (.A(tx_stb), .B(tx_busy), .C(\tx_data[0] ), 
         .D(lcl_data[1]), .Z(lcl_data_7__N_278[0])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(155[7:24])
    defparam lcl_data_7__I_0_i1_3_lut_4_lut.init = 16'hfd20;
    CCU2D sub_36_add_2_13 (.A0(baud_counter[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n19781), .COUT(n19782), .S0(n108[11]), 
          .S1(n108[12]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_13.INIT0 = 16'h5555;
    defparam sub_36_add_2_13.INIT1 = 16'h5555;
    defparam sub_36_add_2_13.INJECT1_0 = "NO";
    defparam sub_36_add_2_13.INJECT1_1 = "NO";
    LUT4 i864_2_lut_3_lut (.A(tx_stb), .B(tx_busy), .C(zero_baud_counter), 
         .Z(dac_clk_p_c_enable_514)) /* synthesis lut_function=(A ((C)+!B)+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(155[7:24])
    defparam i864_2_lut_3_lut.init = 16'hf2f2;
    CCU2D sub_36_add_2_11 (.A0(baud_counter[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n19780), .COUT(n19781), .S0(n108[9]), .S1(n108[10]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_11.INIT0 = 16'h5555;
    defparam sub_36_add_2_11.INIT1 = 16'h5555;
    defparam sub_36_add_2_11.INJECT1_0 = "NO";
    defparam sub_36_add_2_11.INJECT1_1 = "NO";
    LUT4 lcl_data_7__I_0_i7_3_lut_4_lut (.A(tx_stb), .B(tx_busy), .C(\tx_data[6] ), 
         .D(lcl_data[7]), .Z(lcl_data_7__N_278[6])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(155[7:24])
    defparam lcl_data_7__I_0_i7_3_lut_4_lut.init = 16'hfd20;
    CCU2D sub_36_add_2_9 (.A0(baud_counter[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n19779), .COUT(n19780), .S0(n108[7]), .S1(n108[8]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_9.INIT0 = 16'h5555;
    defparam sub_36_add_2_9.INIT1 = 16'h5555;
    defparam sub_36_add_2_9.INJECT1_0 = "NO";
    defparam sub_36_add_2_9.INJECT1_1 = "NO";
    LUT4 lcl_data_7__I_0_i6_3_lut_4_lut (.A(tx_stb), .B(tx_busy), .C(\tx_data[5] ), 
         .D(lcl_data[6]), .Z(lcl_data_7__N_278[5])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(155[7:24])
    defparam lcl_data_7__I_0_i6_3_lut_4_lut.init = 16'hfd20;
    LUT4 lcl_data_7__I_0_i5_3_lut_4_lut (.A(tx_stb), .B(tx_busy), .C(\tx_data[4] ), 
         .D(lcl_data[5]), .Z(lcl_data_7__N_278[4])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(155[7:24])
    defparam lcl_data_7__I_0_i5_3_lut_4_lut.init = 16'hfd20;
    CCU2D sub_36_add_2_7 (.A0(baud_counter[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n19778), .COUT(n19779), .S0(n108[5]), .S1(n108[6]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_7.INIT0 = 16'h5555;
    defparam sub_36_add_2_7.INIT1 = 16'h5555;
    defparam sub_36_add_2_7.INJECT1_0 = "NO";
    defparam sub_36_add_2_7.INJECT1_1 = "NO";
    LUT4 lcl_data_7__I_0_i4_3_lut_4_lut (.A(tx_stb), .B(tx_busy), .C(\tx_data[3] ), 
         .D(lcl_data[4]), .Z(lcl_data_7__N_278[3])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(155[7:24])
    defparam lcl_data_7__I_0_i4_3_lut_4_lut.init = 16'hfd20;
    CCU2D sub_36_add_2_5 (.A0(baud_counter[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n19777), .COUT(n19778), .S0(n108[3]), .S1(n108[4]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_5.INIT0 = 16'h5555;
    defparam sub_36_add_2_5.INIT1 = 16'h5555;
    defparam sub_36_add_2_5.INJECT1_0 = "NO";
    defparam sub_36_add_2_5.INJECT1_1 = "NO";
    LUT4 lcl_data_7__I_0_i3_3_lut_4_lut (.A(tx_stb), .B(tx_busy), .C(\tx_data[2] ), 
         .D(lcl_data[3]), .Z(lcl_data_7__N_278[2])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(155[7:24])
    defparam lcl_data_7__I_0_i3_3_lut_4_lut.init = 16'hfd20;
    CCU2D sub_36_add_2_3 (.A0(baud_counter[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n19776), .COUT(n19777), .S0(n108[1]), .S1(n108[2]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_3.INIT0 = 16'h5555;
    defparam sub_36_add_2_3.INIT1 = 16'h5555;
    defparam sub_36_add_2_3.INJECT1_0 = "NO";
    defparam sub_36_add_2_3.INJECT1_1 = "NO";
    LUT4 lcl_data_7__I_0_i2_3_lut_4_lut (.A(tx_stb), .B(tx_busy), .C(\tx_data[1] ), 
         .D(lcl_data[2]), .Z(lcl_data_7__N_278[1])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(155[7:24])
    defparam lcl_data_7__I_0_i2_3_lut_4_lut.init = 16'hfd20;
    CCU2D sub_36_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(baud_counter[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n19776), .S1(n108[0]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_1.INIT0 = 16'hF000;
    defparam sub_36_add_2_1.INIT1 = 16'h5555;
    defparam sub_36_add_2_1.INJECT1_0 = "NO";
    defparam sub_36_add_2_1.INJECT1_1 = "NO";
    LUT4 i1_2_lut_4_lut (.A(state[2]), .B(n29209), .C(state[1]), .D(zero_baud_counter), 
         .Z(n12747)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;
    defparam i1_2_lut_4_lut.init = 16'hff80;
    FD1S3IX baud_counter_i23 (.D(n108[23]), .CK(dac_clk_p_c), .CD(n12747), 
            .Q(baud_counter[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=7, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=69, LSE_RLINE=69 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i23.GSR = "DISABLED";
    FD1S3IX baud_counter_i22 (.D(n108[22]), .CK(dac_clk_p_c), .CD(n12747), 
            .Q(baud_counter[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=7, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=69, LSE_RLINE=69 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i22.GSR = "DISABLED";
    FD1S3IX baud_counter_i21 (.D(n108[21]), .CK(dac_clk_p_c), .CD(n12747), 
            .Q(baud_counter[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=7, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=69, LSE_RLINE=69 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i21.GSR = "DISABLED";
    FD1S3IX baud_counter_i20 (.D(n108[20]), .CK(dac_clk_p_c), .CD(n12747), 
            .Q(baud_counter[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=7, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=69, LSE_RLINE=69 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i20.GSR = "DISABLED";
    FD1S3IX baud_counter_i19 (.D(n108[19]), .CK(dac_clk_p_c), .CD(n12747), 
            .Q(baud_counter[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=7, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=69, LSE_RLINE=69 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i19.GSR = "DISABLED";
    FD1S3IX baud_counter_i18 (.D(n108[18]), .CK(dac_clk_p_c), .CD(n12747), 
            .Q(baud_counter[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=7, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=69, LSE_RLINE=69 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i18.GSR = "DISABLED";
    FD1S3IX baud_counter_i17 (.D(n108[17]), .CK(dac_clk_p_c), .CD(n12747), 
            .Q(baud_counter[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=7, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=69, LSE_RLINE=69 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i17.GSR = "DISABLED";
    FD1S3IX baud_counter_i16 (.D(n108[16]), .CK(dac_clk_p_c), .CD(n12747), 
            .Q(baud_counter[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=7, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=69, LSE_RLINE=69 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i16.GSR = "DISABLED";
    FD1S3IX baud_counter_i15 (.D(n108[15]), .CK(dac_clk_p_c), .CD(n12747), 
            .Q(baud_counter[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=7, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=69, LSE_RLINE=69 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i15.GSR = "DISABLED";
    FD1S3IX baud_counter_i14 (.D(n108[14]), .CK(dac_clk_p_c), .CD(n12747), 
            .Q(baud_counter[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=7, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=69, LSE_RLINE=69 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i14.GSR = "DISABLED";
    FD1S3AX baud_counter_i13 (.D(baud_counter_23__N_250[13]), .CK(dac_clk_p_c), 
            .Q(baud_counter[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=7, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=69, LSE_RLINE=69 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i13.GSR = "DISABLED";
    FD1S3IX baud_counter_i12 (.D(n108[12]), .CK(dac_clk_p_c), .CD(n12747), 
            .Q(baud_counter[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=7, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=69, LSE_RLINE=69 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i12.GSR = "DISABLED";
    FD1S3IX baud_counter_i11 (.D(n108[11]), .CK(dac_clk_p_c), .CD(n12747), 
            .Q(baud_counter[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=7, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=69, LSE_RLINE=69 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i11.GSR = "DISABLED";
    FD1S3AX baud_counter_i10 (.D(baud_counter_23__N_250[10]), .CK(dac_clk_p_c), 
            .Q(baud_counter[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=7, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=69, LSE_RLINE=69 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i10.GSR = "DISABLED";
    FD1S3AX baud_counter_i9 (.D(baud_counter_23__N_250[9]), .CK(dac_clk_p_c), 
            .Q(baud_counter[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=7, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=69, LSE_RLINE=69 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i9.GSR = "DISABLED";
    FD1S3AX baud_counter_i8 (.D(baud_counter_23__N_250[8]), .CK(dac_clk_p_c), 
            .Q(baud_counter[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=7, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=69, LSE_RLINE=69 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i8.GSR = "DISABLED";
    FD1S3IX baud_counter_i7 (.D(n108[7]), .CK(dac_clk_p_c), .CD(n12747), 
            .Q(baud_counter[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=7, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=69, LSE_RLINE=69 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i7.GSR = "DISABLED";
    FD1S3IX baud_counter_i6 (.D(n108[6]), .CK(dac_clk_p_c), .CD(n12747), 
            .Q(baud_counter[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=7, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=69, LSE_RLINE=69 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i6.GSR = "DISABLED";
    FD1S3IX baud_counter_i5 (.D(n108[5]), .CK(dac_clk_p_c), .CD(n12747), 
            .Q(baud_counter[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=7, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=69, LSE_RLINE=69 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i5.GSR = "DISABLED";
    FD1S3IX baud_counter_i4 (.D(n108[4]), .CK(dac_clk_p_c), .CD(n12747), 
            .Q(baud_counter[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=7, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=69, LSE_RLINE=69 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i4.GSR = "DISABLED";
    FD1S3AX baud_counter_i3 (.D(baud_counter_23__N_250[3]), .CK(dac_clk_p_c), 
            .Q(baud_counter[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=7, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=69, LSE_RLINE=69 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i3.GSR = "DISABLED";
    FD1S3AX baud_counter_i2 (.D(baud_counter_23__N_250[2]), .CK(dac_clk_p_c), 
            .Q(baud_counter[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=7, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=69, LSE_RLINE=69 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i2.GSR = "DISABLED";
    FD1S3AX baud_counter_i1 (.D(baud_counter_23__N_250[1]), .CK(dac_clk_p_c), 
            .Q(baud_counter[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=7, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=69, LSE_RLINE=69 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i1.GSR = "DISABLED";
    FD1P3AX state_855__i3 (.D(n29498), .SP(zero_baud_counter), .CK(dac_clk_p_c), 
            .Q(state[3]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(110[14:26])
    defparam state_855__i3.GSR = "DISABLED";
    FD1P3AX state_855__i2 (.D(n29495), .SP(zero_baud_counter), .CK(dac_clk_p_c), 
            .Q(state[2]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(110[14:26])
    defparam state_855__i2.GSR = "DISABLED";
    FD1P3AX state_855__i1 (.D(n27[1]), .SP(zero_baud_counter), .CK(dac_clk_p_c), 
            .Q(state[1]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(110[14:26])
    defparam state_855__i1.GSR = "DISABLED";
    FD1P3IX lcl_data_i7 (.D(n32067), .SP(zero_baud_counter), .CD(n29211), 
            .CK(dac_clk_p_c), .Q(lcl_data[7])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=7, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=69, LSE_RLINE=69 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(139[9] 143[40])
    defparam lcl_data_i7.GSR = "DISABLED";
    FD1P3AY lcl_data_i6 (.D(lcl_data_7__N_278[6]), .SP(dac_clk_p_c_enable_514), 
            .CK(dac_clk_p_c), .Q(lcl_data[6])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=7, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=69, LSE_RLINE=69 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(139[9] 143[40])
    defparam lcl_data_i6.GSR = "DISABLED";
    FD1P3AY lcl_data_i5 (.D(lcl_data_7__N_278[5]), .SP(dac_clk_p_c_enable_514), 
            .CK(dac_clk_p_c), .Q(lcl_data[5])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=7, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=69, LSE_RLINE=69 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(139[9] 143[40])
    defparam lcl_data_i5.GSR = "DISABLED";
    FD1P3AY lcl_data_i4 (.D(lcl_data_7__N_278[4]), .SP(dac_clk_p_c_enable_514), 
            .CK(dac_clk_p_c), .Q(lcl_data[4])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=7, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=69, LSE_RLINE=69 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(139[9] 143[40])
    defparam lcl_data_i4.GSR = "DISABLED";
    FD1P3AY lcl_data_i3 (.D(lcl_data_7__N_278[3]), .SP(dac_clk_p_c_enable_514), 
            .CK(dac_clk_p_c), .Q(lcl_data[3])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=7, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=69, LSE_RLINE=69 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(139[9] 143[40])
    defparam lcl_data_i3.GSR = "DISABLED";
    FD1P3AY lcl_data_i2 (.D(lcl_data_7__N_278[2]), .SP(dac_clk_p_c_enable_514), 
            .CK(dac_clk_p_c), .Q(lcl_data[2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=7, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=69, LSE_RLINE=69 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(139[9] 143[40])
    defparam lcl_data_i2.GSR = "DISABLED";
    FD1P3AY lcl_data_i1 (.D(lcl_data_7__N_278[1]), .SP(dac_clk_p_c_enable_514), 
            .CK(dac_clk_p_c), .Q(lcl_data[1])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=7, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=69, LSE_RLINE=69 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(139[9] 143[40])
    defparam lcl_data_i1.GSR = "DISABLED";
    LUT4 baud_counter_23__I_9_i14_4_lut (.A(n29211), .B(n133[13]), .C(n29096), 
         .D(zero_baud_counter_N_295), .Z(baud_counter_23__N_250[13])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((C+(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(217[12] 224[43])
    defparam baud_counter_23__I_9_i14_4_lut.init = 16'ha0ac;
    LUT4 i13134_2_lut (.A(n108[13]), .B(zero_baud_counter), .Z(n133[13])) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(224[4:43])
    defparam i13134_2_lut.init = 16'heeee;
    LUT4 baud_counter_23__I_9_i11_4_lut (.A(n29211), .B(n133[10]), .C(n29096), 
         .D(zero_baud_counter_N_295), .Z(baud_counter_23__N_250[10])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((C+(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(217[12] 224[43])
    defparam baud_counter_23__I_9_i11_4_lut.init = 16'ha0ac;
    LUT4 i13135_2_lut (.A(n108[10]), .B(zero_baud_counter), .Z(n133[10])) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(224[4:43])
    defparam i13135_2_lut.init = 16'heeee;
    LUT4 baud_counter_23__I_9_i10_4_lut (.A(n29211), .B(n133[9]), .C(n29096), 
         .D(zero_baud_counter_N_295), .Z(baud_counter_23__N_250[9])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((C+(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(217[12] 224[43])
    defparam baud_counter_23__I_9_i10_4_lut.init = 16'ha0ac;
    LUT4 i13136_2_lut (.A(n108[9]), .B(zero_baud_counter), .Z(n133[9])) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(224[4:43])
    defparam i13136_2_lut.init = 16'heeee;
    LUT4 baud_counter_23__I_9_i9_4_lut (.A(n29211), .B(n133[8]), .C(n29096), 
         .D(zero_baud_counter_N_295), .Z(baud_counter_23__N_250[8])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((C+(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(217[12] 224[43])
    defparam baud_counter_23__I_9_i9_4_lut.init = 16'ha0ac;
    LUT4 i13137_2_lut (.A(n108[8]), .B(zero_baud_counter), .Z(n133[8])) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(224[4:43])
    defparam i13137_2_lut.init = 16'heeee;
    LUT4 baud_counter_23__I_9_i4_4_lut (.A(n29211), .B(n133[3]), .C(n29096), 
         .D(zero_baud_counter_N_295), .Z(baud_counter_23__N_250[3])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((C+(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(217[12] 224[43])
    defparam baud_counter_23__I_9_i4_4_lut.init = 16'ha0ac;
    LUT4 i13138_2_lut (.A(n108[3]), .B(zero_baud_counter), .Z(n133[3])) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(224[4:43])
    defparam i13138_2_lut.init = 16'heeee;
    LUT4 baud_counter_23__I_9_i3_4_lut (.A(n29211), .B(n133[2]), .C(n29096), 
         .D(zero_baud_counter_N_295), .Z(baud_counter_23__N_250[2])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((C+(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(217[12] 224[43])
    defparam baud_counter_23__I_9_i3_4_lut.init = 16'ha0ac;
    LUT4 i13139_2_lut (.A(n108[2]), .B(zero_baud_counter), .Z(n133[2])) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(224[4:43])
    defparam i13139_2_lut.init = 16'heeee;
    LUT4 baud_counter_23__I_9_i2_4_lut (.A(n29211), .B(n133[1]), .C(n29096), 
         .D(zero_baud_counter_N_295), .Z(baud_counter_23__N_250[1])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((C+(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(217[12] 224[43])
    defparam baud_counter_23__I_9_i2_4_lut.init = 16'ha0ac;
    LUT4 i13140_2_lut (.A(n108[1]), .B(zero_baud_counter), .Z(n133[1])) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(224[4:43])
    defparam i13140_2_lut.init = 16'heeee;
    LUT4 state_855_mux_6_i2_4_lut (.A(state[1]), .B(n29211), .C(n29107), 
         .D(state[0]), .Z(n27[1])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(110[14:26])
    defparam state_855_mux_6_i2_4_lut.init = 16'h353a;
    LUT4 state_855_mux_6_i3_4_lut_then_4_lut (.A(n29211), .B(state[0]), 
         .C(state[1]), .D(state[3]), .Z(n29494)) /* synthesis lut_function=(!(A (B (C+(D))+!B (D))+!A !(((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(110[14:26])
    defparam state_855_mux_6_i3_4_lut_then_4_lut.init = 16'h553f;
    LUT4 zero_baud_counter_I_0_51_4_lut (.A(n29211), .B(n22214), .C(n29096), 
         .D(zero_baud_counter_N_295), .Z(zero_baud_counter_N_292)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C))+!A !((C+(D))+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(217[12] 224[43])
    defparam zero_baud_counter_I_0_51_4_lut.init = 16'h5f53;
    LUT4 i1_4_lut_adj_173 (.A(n22191), .B(n22624), .C(n22618), .D(baud_counter[0]), 
         .Z(n22214)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(207[24:43])
    defparam i1_4_lut_adj_173.init = 16'hfeff;
    LUT4 i1_4_lut_adj_174 (.A(baud_counter[6]), .B(baud_counter[9]), .C(baud_counter[8]), 
         .D(baud_counter[1]), .Z(n22191)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(207[24:43])
    defparam i1_4_lut_adj_174.init = 16'hfffe;
    LUT4 i1_4_lut_adj_175 (.A(n22608), .B(n22203), .C(n22612), .D(n22602), 
         .Z(n22624)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(207[24:43])
    defparam i1_4_lut_adj_175.init = 16'hfffe;
    LUT4 state_855_mux_6_i3_4_lut_else_4_lut (.A(n29211), .B(state[0]), 
         .C(state[1]), .D(state[3]), .Z(n29493)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A !(B (C+(D))+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(110[14:26])
    defparam state_855_mux_6_i3_4_lut_else_4_lut.init = 16'h54c0;
    LUT4 i1_4_lut_adj_176 (.A(n22616), .B(baud_counter[3]), .C(baud_counter[16]), 
         .D(baud_counter[13]), .Z(n22618)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(207[24:43])
    defparam i1_4_lut_adj_176.init = 16'hfffe;
    LUT4 state_855_mux_6_i4_4_lut_then_4_lut (.A(n29211), .B(state[2]), 
         .C(state[0]), .D(state[1]), .Z(n29497)) /* synthesis lut_function=(!(A (B+(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(110[14:26])
    defparam state_855_mux_6_i4_4_lut_then_4_lut.init = 16'h5557;
    LUT4 state_855_mux_6_i4_4_lut_else_4_lut (.A(state[2]), .B(state[0]), 
         .C(state[1]), .Z(n29496)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(110[14:26])
    defparam state_855_mux_6_i4_4_lut_else_4_lut.init = 16'h8080;
    FD1S3JX r_busy_45 (.D(n9431), .CK(dac_clk_p_c), .PD(n29211), .Q(tx_busy)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=7, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=69, LSE_RLINE=69 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(92[9] 114[5])
    defparam r_busy_45.GSR = "DISABLED";
    LUT4 i1_2_lut_adj_177 (.A(baud_counter[2]), .B(baud_counter[23]), .Z(n22608)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(207[24:43])
    defparam i1_2_lut_adj_177.init = 16'heeee;
    LUT4 i1_4_lut_adj_178 (.A(baud_counter[22]), .B(baud_counter[11]), .C(baud_counter[12]), 
         .D(baud_counter[17]), .Z(n22203)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(207[24:43])
    defparam i1_4_lut_adj_178.init = 16'hfffe;
    LUT4 i24572_2_lut_4_lut (.A(n29210), .B(state[3]), .C(state[0]), .D(zero_baud_counter), 
         .Z(n9431)) /* synthesis lut_function=(!(A (B (D))+!A (B (C (D))))) */ ;
    defparam i24572_2_lut_4_lut.init = 16'h37ff;
    LUT4 state_855_mux_6_i1_3_lut_4_lut (.A(n29210), .B(state[3]), .C(state[0]), 
         .D(n29211), .Z(n20035)) /* synthesis lut_function=(!(A (B (D)+!B (C))+!A (B (C (D))+!B (C)))) */ ;
    defparam state_855_mux_6_i1_3_lut_4_lut.init = 16'h07cf;
    FD1P3AX state_855__i0 (.D(n20035), .SP(zero_baud_counter), .CK(dac_clk_p_c), 
            .Q(state[0]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(110[14:26])
    defparam state_855__i0.GSR = "DISABLED";
    
endmodule
