// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.11.3.469
// Netlist written on Sat Feb 06 16:00:09 2021
//
// Verilog Description of module top
//

module top (i_ref_clk, i_resetb, i_wbu_uart_rx, o_wbu_uart_tx, o_dac_a, 
            o_dac_b, dac_clk_p, dac_clk_n, o_dac_cw_b, i_clk_p, i_clk_n, 
            q_clk_p, q_clk_n) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(4[8:11])
    input i_ref_clk;   // d:/documents/git_local/fm_modulator/rtl/top.v(23[12:21])
    input i_resetb;   // d:/documents/git_local/fm_modulator/rtl/top.v(23[23:31])
    input i_wbu_uart_rx;   // d:/documents/git_local/fm_modulator/rtl/top.v(25[12:25])
    output o_wbu_uart_tx;   // d:/documents/git_local/fm_modulator/rtl/top.v(26[13:26])
    output [9:0]o_dac_a;   // d:/documents/git_local/fm_modulator/rtl/top.v(28[38:45])
    output [9:0]o_dac_b;   // d:/documents/git_local/fm_modulator/rtl/top.v(28[47:54])
    output dac_clk_p;   // d:/documents/git_local/fm_modulator/rtl/top.v(29[49:58])
    output dac_clk_n;   // d:/documents/git_local/fm_modulator/rtl/top.v(29[60:69])
    output o_dac_cw_b;   // d:/documents/git_local/fm_modulator/rtl/top.v(29[71:81])
    output i_clk_p;   // d:/documents/git_local/fm_modulator/rtl/top.v(29[13:20])
    output i_clk_n;   // d:/documents/git_local/fm_modulator/rtl/top.v(29[22:29])
    output q_clk_p;   // d:/documents/git_local/fm_modulator/rtl/top.v(29[31:38])
    output q_clk_n;   // d:/documents/git_local/fm_modulator/rtl/top.v(29[40:47])
    
    wire i_ref_clk_c /* synthesis is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(23[12:21])
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(29[49:58])
    wire lo_pll_out /* synthesis is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(157[6:16])
    wire [15:0]o_sample_i /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[39:49])
    wire o_dac_b_c_15 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire o_dac_b_c_14 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire o_dac_b_c_13 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire o_dac_b_c_12 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire o_dac_b_c_11 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire o_dac_b_c_10 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire n3537 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire o_dac_b_c_8 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire o_dac_b_c_7 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire i_clk_2f_N_2250 /* synthesis is_inv_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/clock_phase_shifter.v(11[21:28])
    
    wire GND_net, VCC_net, o_dac_cw_b_c_c, i_wbu_uart_rx_c, o_wbu_uart_tx_c, 
        o_dac_a_c_9, o_dac_a_c_7, o_dac_a_c_6, o_dac_a_c_5, o_dac_a_c_4, 
        o_dac_a_c_3, o_dac_a_c_2, o_dac_a_c_1, o_dac_a_c_0, o_dac_b_c_9, 
        i_clk_p_c, q_clk_p_c, dac_clk_n_c, rx_stb;
    wire [7:0]rx_data;   // d:/documents/git_local/fm_modulator/rtl/top.v(52[12:19])
    
    wire tx_busy, wb_cyc, wb_stb, wb_we;
    wire [29:0]wb_addr;   // d:/documents/git_local/fm_modulator/rtl/top.v(69[13:20])
    wire [31:0]wb_odata;   // d:/documents/git_local/fm_modulator/rtl/top.v(70[13:21])
    
    wire wb_ack, wb_err;
    wire [31:0]wb_idata;   // d:/documents/git_local/fm_modulator/rtl/top.v(75[12:20])
    wire [29:0]bus_err_address;   // d:/documents/git_local/fm_modulator/rtl/top.v(99[12:27])
    
    wire wb_fm_ack;
    wire [31:0]wb_fm_data;   // d:/documents/git_local/fm_modulator/rtl/top.v(103[13:23])
    wire [31:0]wb_smpl_data;   // d:/documents/git_local/fm_modulator/rtl/top.v(106[12:24])
    
    wire wb_smpl_ack;
    wire [7:0]wb_lo_data;   // d:/documents/git_local/fm_modulator/rtl/top.v(135[12:22])
    
    wire wb_lo_ack, pll_clk, pll_rst, pll_stb, pll_we, pll_ack;
    wire [7:0]pll_data_i;   // d:/documents/git_local/fm_modulator/rtl/top.v(141[12:22])
    wire [7:0]pll_data_o;   // d:/documents/git_local/fm_modulator/rtl/top.v(141[24:34])
    wire [4:0]pll_addr;   // d:/documents/git_local/fm_modulator/rtl/top.v(142[12:20])
    wire [31:0]smpl_register;   // d:/documents/git_local/fm_modulator/rtl/top.v(195[13:26])
    wire [31:0]power_counter;   // d:/documents/git_local/fm_modulator/rtl/top.v(195[28:41])
    
    wire smpl_interrupt, none_sel, o_dac_a_9__N_1, wb_lo_data_7__N_96;
    wire [31:0]wb_smpl_data_31__N_64;
    wire [31:0]power_counter_31__N_232;
    wire [30:0]power_counter_31__N_201;
    wire [31:0]power_counter_31__N_129;
    
    wire wb_smpl_sel_N_311;
    wire [31:0]wb_idata_31__N_266;
    wire [31:0]wb_idata_31__N_2;
    wire [23:0]chg_counter;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(97[17:28])
    
    wire chg_counter_23__N_406, n20438;
    wire [3:0]state_adj_3087;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(83[12:17])
    wire [7:0]lcl_data;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(84[12:20])
    
    wire zero_baud_counter, o_busy_N_536, n20918;
    wire [7:0]lcl_data_7__N_511;
    
    wire n20922, n20916, n20432, i_clk_n_c, q_clk_n_c, dac_clk_p_c_enable_272, 
        n20422, n26369, n20470, n20104, n20468, n20466, n20886, 
        n26341, n20456, n2035, n2034, n2033, n2032, n26337, n2030, 
        n2029, n2028, n26342, n2025, n2024, n2023, n2022, n2021, 
        n26332, n20416, n26333, n2017, n26683, n2015, n2014, n2013, 
        n2012, n2011, n2010, n2009, n2008, n2006, n2005, n12635, 
        n2, n20412, n7, dac_clk_p_c_enable_174, n26403, n20402, 
        n9365, n20872, n17295, n26643, n17315, n17296, n17310, 
        n20774, n17314, n17309, n20770, n17301, n17308, n17307, 
        dac_clk_p_c_enable_198, n20384, n17306, n26339, n17313, n9787, 
        n20708, n20378, n20702, n26564, n26563, n26557, n26336, 
        n17324, n26540, n26535, n17305, n17323, n17299, n17312, 
        n17294, n17304, n17311, n17322, n17303, n17321, n17302, 
        n17320, n17300, n38, n34, n17598, n17319, n17298, n17318, 
        n17297, n17317, n4, n26331, n26453, dac_clk_p_c_enable_321, 
        n17316, n26428, n20912, n20910, n20864, n20904, n2_adj_3035, 
        n1, n2_adj_3036, n1_adj_3037, n2_adj_3038, n2_adj_3039, n1_adj_3040, 
        n2_adj_3041, n1_adj_3042, n2_adj_3043, n1_adj_3044, n2_adj_3045, 
        n1_adj_3046, n2_adj_3047, n1_adj_3048, n2_adj_3049, n1_adj_3050, 
        n2_adj_3051, n1_adj_3052, n2_adj_3053, n1_adj_3054, n2_adj_3055, 
        n2_adj_3056, n1_adj_3057, n2_adj_3058, n2_adj_3059, n2_adj_3060, 
        n2_adj_3061, n1_adj_3062, n2_adj_3063, n1_adj_3064, n29210, 
        n2_adj_3065, n1_adj_3066, n2_adj_3067, n1_adj_3068, n2_adj_3069, 
        n1_adj_3070, n2_adj_3071, n2_adj_3072, n2_adj_3073, n1_adj_3074, 
        n2_adj_3075, n1_adj_3076, n2_adj_3077, n1_adj_3078, n2_adj_3079, 
        n2_adj_3080, n1_adj_3081, n2_adj_3082, n1_adj_3083, n2_adj_3084, 
        n20906, n29209, n1_adj_3085, n20888;
    
    VHI i2 (.Z(VCC_net));
    GSR GSR_INST (.GSR(n26683)) /* synthesis syn_instantiated=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(34[5:28])
    \rxuartlite(CLOCKS_PER_BAUD=10000)  rxtransport (.dac_clk_p_c(dac_clk_p_c), 
            .\rx_data[0] (rx_data[0]), .rx_stb(rx_stb), .i_wbu_uart_rx_c(i_wbu_uart_rx_c), 
            .chg_counter({chg_counter}), .dac_clk_p_c_enable_174(dac_clk_p_c_enable_174), 
            .chg_counter_23__N_406(chg_counter_23__N_406), .GND_net(GND_net), 
            .\rx_data[6] (rx_data[6]), .\rx_data[5] (rx_data[5]), .\rx_data[4] (rx_data[4]), 
            .\rx_data[3] (rx_data[3]), .\rx_data[2] (rx_data[2]), .\rx_data[1] (rx_data[1])) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(54[57:105])
    hbbus genbus (.wb_odata({wb_odata}), .dac_clk_p_c(dac_clk_p_c), .wb_we(wb_we), 
          .wb_stb(wb_stb), .wb_cyc(wb_cyc), .wb_addr({wb_addr}), .GND_net(GND_net), 
          .wb_err(wb_err), .wb_ack(wb_ack), .\wb_idata[0] (wb_idata[0]), 
          .\wb_idata[2] (wb_idata[2]), .\wb_idata[3] (wb_idata[3]), .\wb_idata[4] (wb_idata[4]), 
          .\wb_idata[5] (wb_idata[5]), .\wb_idata[6] (wb_idata[6]), .\wb_idata[7] (wb_idata[7]), 
          .\wb_idata[8] (wb_idata[8]), .\wb_idata[9] (wb_idata[9]), .\wb_idata[10] (wb_idata[10]), 
          .\wb_idata[11] (wb_idata[11]), .\wb_idata[12] (wb_idata[12]), 
          .\wb_idata[13] (wb_idata[13]), .\wb_idata[14] (wb_idata[14]), 
          .\wb_idata[15] (wb_idata[15]), .\wb_idata[16] (wb_idata[16]), 
          .\wb_idata[17] (wb_idata[17]), .\wb_idata[18] (wb_idata[18]), 
          .\wb_idata[19] (wb_idata[19]), .\wb_idata[20] (wb_idata[20]), 
          .\wb_idata[21] (wb_idata[21]), .\wb_idata[22] (wb_idata[22]), 
          .\wb_idata[23] (wb_idata[23]), .\wb_idata[24] (wb_idata[24]), 
          .\wb_idata[25] (wb_idata[25]), .\wb_idata[26] (wb_idata[26]), 
          .\wb_idata[27] (wb_idata[27]), .\wb_idata[28] (wb_idata[28]), 
          .\wb_idata[29] (wb_idata[29]), .\wb_idata[30] (wb_idata[30]), 
          .\wb_idata[31] (wb_idata[31]), .n2(n2), .n12635(n12635), .n29210(n29210), 
          .VCC_net(VCC_net), .\rx_data[5] (rx_data[5]), .\rx_data[1] (rx_data[1]), 
          .rx_stb(rx_stb), .\rx_data[6] (rx_data[6]), .\rx_data[3] (rx_data[3]), 
          .\rx_data[4] (rx_data[4]), .\rx_data[0] (rx_data[0]), .\rx_data[2] (rx_data[2]), 
          .tx_busy(tx_busy), .o_busy_N_536(o_busy_N_536), .\state[0] (state_adj_3087[0]), 
          .n17598(n17598), .n26540(n26540), .\lcl_data[1] (lcl_data[1]), 
          .\lcl_data_7__N_511[0] (lcl_data_7__N_511[0]), .\lcl_data[4] (lcl_data[4]), 
          .\lcl_data_7__N_511[3] (lcl_data_7__N_511[3]), .\lcl_data[5] (lcl_data[5]), 
          .\lcl_data_7__N_511[4] (lcl_data_7__N_511[4]), .\lcl_data[6] (lcl_data[6]), 
          .\lcl_data_7__N_511[5] (lcl_data_7__N_511[5]), .\lcl_data[7] (lcl_data[7]), 
          .\lcl_data_7__N_511[6] (lcl_data_7__N_511[6]), .zero_baud_counter(zero_baud_counter), 
          .dac_clk_p_c_enable_321(dac_clk_p_c_enable_321), .\lcl_data[3] (lcl_data[3]), 
          .\lcl_data_7__N_511[2] (lcl_data_7__N_511[2]), .\lcl_data[2] (lcl_data[2]), 
          .\lcl_data_7__N_511[1] (lcl_data_7__N_511[1])) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(78[7] 94[22])
    FD1S3AX power_counter_i0 (.D(power_counter_31__N_129[0]), .CK(dac_clk_p_c), 
            .Q(power_counter[0])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(224[9] 229[54])
    defparam power_counter_i0.GSR = "DISABLED";
    FD1S3AX wb_idata_i0 (.D(wb_idata_31__N_2[0]), .CK(dac_clk_p_c), .Q(wb_idata[0]));   // d:/documents/git_local/fm_modulator/rtl/top.v(265[9] 273[53])
    defparam wb_idata_i0.GSR = "DISABLED";
    FD1S3JX wb_ack_68 (.D(n4), .CK(dac_clk_p_c), .PD(wb_smpl_ack), .Q(wb_ack)) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(262[9] 263[57])
    defparam wb_ack_68.GSR = "DISABLED";
    PUR PUR_INST (.PUR(n26683)) /* synthesis syn_instantiated=1 */ ;
    defparam PUR_INST.RST_PULSE = 1;
    FD1S3IX wb_smpl_ack_61 (.D(wb_stb), .CK(dac_clk_p_c), .CD(wb_smpl_sel_N_311), 
            .Q(wb_smpl_ack)) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(198[9] 199[44])
    defparam wb_smpl_ack_61.GSR = "DISABLED";
    \txuartlite(TIMING_BITS=24,CLOCKS_PER_BAUD=10000)  txtransport (.dac_clk_p_c(dac_clk_p_c), 
            .dac_clk_p_c_enable_321(dac_clk_p_c_enable_321), .\lcl_data_7__N_511[0] (lcl_data_7__N_511[0]), 
            .zero_baud_counter(zero_baud_counter), .o_wbu_uart_tx_c(o_wbu_uart_tx_c), 
            .n26540(n26540), .state({Open_0, Open_1, Open_2, state_adj_3087[0]}), 
            .GND_net(GND_net), .\lcl_data[7] (lcl_data[7]), .n29210(n29210), 
            .\lcl_data[6] (lcl_data[6]), .\lcl_data_7__N_511[6] (lcl_data_7__N_511[6]), 
            .\lcl_data[5] (lcl_data[5]), .\lcl_data_7__N_511[5] (lcl_data_7__N_511[5]), 
            .\lcl_data[4] (lcl_data[4]), .\lcl_data_7__N_511[4] (lcl_data_7__N_511[4]), 
            .\lcl_data[3] (lcl_data[3]), .\lcl_data_7__N_511[3] (lcl_data_7__N_511[3]), 
            .\lcl_data[2] (lcl_data[2]), .\lcl_data_7__N_511[2] (lcl_data_7__N_511[2]), 
            .\lcl_data[1] (lcl_data[1]), .\lcl_data_7__N_511[1] (lcl_data_7__N_511[1]), 
            .o_busy_N_536(o_busy_N_536), .tx_busy(tx_busy), .n17598(n17598)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(63[58:115])
    FD1P3AX smpl_register_i0_i0 (.D(wb_odata[0]), .SP(dac_clk_p_c_enable_272), 
            .CK(dac_clk_p_c), .Q(smpl_register[0]));   // d:/documents/git_local/fm_modulator/rtl/top.v(202[9] 210[6])
    defparam smpl_register_i0_i0.GSR = "DISABLED";
    FD1S3IX wb_err_66 (.D(none_sel), .CK(dac_clk_p_c), .CD(n2), .Q(wb_err));   // d:/documents/git_local/fm_modulator/rtl/top.v(251[9] 252[34])
    defparam wb_err_66.GSR = "DISABLED";
    OB o_dac_a_pad_7 (.I(o_dac_a_c_7), .O(o_dac_a[7]));   // d:/documents/git_local/fm_modulator/rtl/top.v(28[38:45])
    FD1P3AX bus_err_address_i0_i0 (.D(wb_addr[0]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[0])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(255[9] 257[31])
    defparam bus_err_address_i0_i0.GSR = "DISABLED";
    OB o_dac_a_pad_8 (.I(n26643), .O(o_dac_a[8]));   // d:/documents/git_local/fm_modulator/rtl/top.v(28[38:45])
    OB o_dac_a_pad_9 (.I(o_dac_a_c_9), .O(o_dac_a[9]));   // d:/documents/git_local/fm_modulator/rtl/top.v(28[38:45])
    OB o_wbu_uart_tx_pad (.I(o_wbu_uart_tx_c), .O(o_wbu_uart_tx));   // d:/documents/git_local/fm_modulator/rtl/top.v(26[13:26])
    CCU2D add_32_27 (.A0(power_counter[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17306), .COUT(n17307), .S0(power_counter_31__N_232[25]), 
          .S1(power_counter_31__N_232[26]));   // d:/documents/git_local/fm_modulator/rtl/top.v(227[21:41])
    defparam add_32_27.INIT0 = 16'h5aaa;
    defparam add_32_27.INIT1 = 16'h5aaa;
    defparam add_32_27.INJECT1_0 = "NO";
    defparam add_32_27.INJECT1_1 = "NO";
    CCU2D add_33_31 (.A0(power_counter[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17324), .S0(power_counter_31__N_201[29]), 
          .S1(power_counter_31__N_201[30]));   // d:/documents/git_local/fm_modulator/rtl/top.v(229[27:53])
    defparam add_33_31.INIT0 = 16'h5aaa;
    defparam add_33_31.INIT1 = 16'h5aaa;
    defparam add_33_31.INJECT1_0 = "NO";
    defparam add_33_31.INJECT1_1 = "NO";
    FD1P3AX smpl_interrupt_63 (.D(wb_odata[0]), .SP(dac_clk_p_c_enable_198), 
            .CK(dac_clk_p_c), .Q(smpl_interrupt)) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(202[9] 210[6])
    defparam smpl_interrupt_63.GSR = "DISABLED";
    CCU2D add_32_25 (.A0(power_counter[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17305), .COUT(n17306), .S0(power_counter_31__N_232[23]), 
          .S1(power_counter_31__N_232[24]));   // d:/documents/git_local/fm_modulator/rtl/top.v(227[21:41])
    defparam add_32_25.INIT0 = 16'h5aaa;
    defparam add_32_25.INIT1 = 16'h5aaa;
    defparam add_32_25.INJECT1_0 = "NO";
    defparam add_32_25.INJECT1_1 = "NO";
    CCU2D add_33_29 (.A0(power_counter[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17323), .COUT(n17324), .S0(power_counter_31__N_201[27]), 
          .S1(power_counter_31__N_201[28]));   // d:/documents/git_local/fm_modulator/rtl/top.v(229[27:53])
    defparam add_33_29.INIT0 = 16'h5aaa;
    defparam add_33_29.INIT1 = 16'h5aaa;
    defparam add_33_29.INJECT1_0 = "NO";
    defparam add_33_29.INJECT1_1 = "NO";
    CCU2D add_32_23 (.A0(power_counter[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17304), .COUT(n17305), .S0(power_counter_31__N_232[21]), 
          .S1(power_counter_31__N_232[22]));   // d:/documents/git_local/fm_modulator/rtl/top.v(227[21:41])
    defparam add_32_23.INIT0 = 16'h5aaa;
    defparam add_32_23.INIT1 = 16'h5aaa;
    defparam add_32_23.INJECT1_0 = "NO";
    defparam add_32_23.INJECT1_1 = "NO";
    CCU2D add_33_27 (.A0(power_counter[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17322), .COUT(n17323), .S0(power_counter_31__N_201[25]), 
          .S1(power_counter_31__N_201[26]));   // d:/documents/git_local/fm_modulator/rtl/top.v(229[27:53])
    defparam add_33_27.INIT0 = 16'h5aaa;
    defparam add_33_27.INIT1 = 16'h5aaa;
    defparam add_33_27.INJECT1_0 = "NO";
    defparam add_33_27.INJECT1_1 = "NO";
    CCU2D add_32_21 (.A0(power_counter[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17303), .COUT(n17304), .S0(power_counter_31__N_232[19]), 
          .S1(power_counter_31__N_232[20]));   // d:/documents/git_local/fm_modulator/rtl/top.v(227[21:41])
    defparam add_32_21.INIT0 = 16'h5aaa;
    defparam add_32_21.INIT1 = 16'h5aaa;
    defparam add_32_21.INJECT1_0 = "NO";
    defparam add_32_21.INJECT1_1 = "NO";
    CCU2D add_33_25 (.A0(power_counter[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17321), .COUT(n17322), .S0(power_counter_31__N_201[23]), 
          .S1(power_counter_31__N_201[24]));   // d:/documents/git_local/fm_modulator/rtl/top.v(229[27:53])
    defparam add_33_25.INIT0 = 16'h5aaa;
    defparam add_33_25.INIT1 = 16'h5aaa;
    defparam add_33_25.INJECT1_0 = "NO";
    defparam add_33_25.INJECT1_1 = "NO";
    LUT4 o_clk_q_I_0_1_lut (.A(q_clk_p_c), .Z(q_clk_n_c)) /* synthesis lut_function=(!(A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/clock_phase_shifter.v(18[16:24])
    defparam o_clk_q_I_0_1_lut.init = 16'h5555;
    LUT4 o_clk_i_I_0_1_lut (.A(i_clk_p_c), .Z(i_clk_n_c)) /* synthesis lut_function=(!(A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/clock_phase_shifter.v(14[16:24])
    defparam o_clk_i_I_0_1_lut.init = 16'h5555;
    LUT4 i3_4_lut (.A(wb_addr[9]), .B(wb_addr[8]), .C(wb_cyc), .D(n20104), 
         .Z(wb_lo_data_7__N_96)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i3_4_lut.init = 16'h8000;
    LUT4 i2_4_lut (.A(n34), .B(wb_addr[15]), .C(n38), .D(n26453), .Z(n20104)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i2_4_lut.init = 16'h0004;
    LUT4 i11164_2_lut (.A(smpl_register[19]), .B(wb_addr[0]), .Z(n1_adj_3057)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(213[3] 220[10])
    defparam i11164_2_lut.init = 16'h8888;
    LUT4 i1_4_lut (.A(n20916), .B(n38), .C(n26563), .D(n20384), .Z(dac_clk_p_c_enable_272)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut.init = 16'h0100;
    PFUMX mux_388_Mux_2_i3 (.BLUT(n1_adj_3085), .ALUT(n2_adj_3084), .C0(wb_addr[1]), 
          .Z(n2034));
    LUT4 i1_4_lut_adj_143 (.A(n20378), .B(wb_addr[1]), .C(wb_addr[12]), 
         .D(n26557), .Z(n20384)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_4_lut_adj_143.init = 16'h0200;
    LUT4 i1_2_lut (.A(wb_addr[0]), .B(wb_addr[15]), .Z(n20378)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i17458_2_lut (.A(wb_addr[2]), .B(wb_addr[3]), .Z(n9365)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i17458_2_lut.init = 16'heeee;
    FD1P3AX smpl_register_i0_i31 (.D(wb_odata[31]), .SP(dac_clk_p_c_enable_272), 
            .CK(dac_clk_p_c), .Q(smpl_register[31]));   // d:/documents/git_local/fm_modulator/rtl/top.v(202[9] 210[6])
    defparam smpl_register_i0_i31.GSR = "DISABLED";
    PFUMX mux_388_Mux_3_i3 (.BLUT(n1_adj_3083), .ALUT(n2_adj_3082), .C0(wb_addr[1]), 
          .Z(n2033));
    FD1P3AX smpl_register_i0_i30 (.D(wb_odata[30]), .SP(dac_clk_p_c_enable_272), 
            .CK(dac_clk_p_c), .Q(smpl_register[30]));   // d:/documents/git_local/fm_modulator/rtl/top.v(202[9] 210[6])
    defparam smpl_register_i0_i30.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i29 (.D(wb_odata[29]), .SP(dac_clk_p_c_enable_272), 
            .CK(dac_clk_p_c), .Q(smpl_register[29]));   // d:/documents/git_local/fm_modulator/rtl/top.v(202[9] 210[6])
    defparam smpl_register_i0_i29.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i28 (.D(wb_odata[28]), .SP(dac_clk_p_c_enable_272), 
            .CK(dac_clk_p_c), .Q(smpl_register[28]));   // d:/documents/git_local/fm_modulator/rtl/top.v(202[9] 210[6])
    defparam smpl_register_i0_i28.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i27 (.D(wb_odata[27]), .SP(dac_clk_p_c_enable_272), 
            .CK(dac_clk_p_c), .Q(smpl_register[27]));   // d:/documents/git_local/fm_modulator/rtl/top.v(202[9] 210[6])
    defparam smpl_register_i0_i27.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i26 (.D(wb_odata[26]), .SP(dac_clk_p_c_enable_272), 
            .CK(dac_clk_p_c), .Q(smpl_register[26]));   // d:/documents/git_local/fm_modulator/rtl/top.v(202[9] 210[6])
    defparam smpl_register_i0_i26.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i25 (.D(wb_odata[25]), .SP(dac_clk_p_c_enable_272), 
            .CK(dac_clk_p_c), .Q(smpl_register[25]));   // d:/documents/git_local/fm_modulator/rtl/top.v(202[9] 210[6])
    defparam smpl_register_i0_i25.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i24 (.D(wb_odata[24]), .SP(dac_clk_p_c_enable_272), 
            .CK(dac_clk_p_c), .Q(smpl_register[24]));   // d:/documents/git_local/fm_modulator/rtl/top.v(202[9] 210[6])
    defparam smpl_register_i0_i24.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i23 (.D(wb_odata[23]), .SP(dac_clk_p_c_enable_272), 
            .CK(dac_clk_p_c), .Q(smpl_register[23]));   // d:/documents/git_local/fm_modulator/rtl/top.v(202[9] 210[6])
    defparam smpl_register_i0_i23.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i22 (.D(wb_odata[22]), .SP(dac_clk_p_c_enable_272), 
            .CK(dac_clk_p_c), .Q(smpl_register[22]));   // d:/documents/git_local/fm_modulator/rtl/top.v(202[9] 210[6])
    defparam smpl_register_i0_i22.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i21 (.D(wb_odata[21]), .SP(dac_clk_p_c_enable_272), 
            .CK(dac_clk_p_c), .Q(smpl_register[21]));   // d:/documents/git_local/fm_modulator/rtl/top.v(202[9] 210[6])
    defparam smpl_register_i0_i21.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i20 (.D(wb_odata[20]), .SP(dac_clk_p_c_enable_272), 
            .CK(dac_clk_p_c), .Q(smpl_register[20]));   // d:/documents/git_local/fm_modulator/rtl/top.v(202[9] 210[6])
    defparam smpl_register_i0_i20.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i19 (.D(wb_odata[19]), .SP(dac_clk_p_c_enable_272), 
            .CK(dac_clk_p_c), .Q(smpl_register[19]));   // d:/documents/git_local/fm_modulator/rtl/top.v(202[9] 210[6])
    defparam smpl_register_i0_i19.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i18 (.D(wb_odata[18]), .SP(dac_clk_p_c_enable_272), 
            .CK(dac_clk_p_c), .Q(smpl_register[18]));   // d:/documents/git_local/fm_modulator/rtl/top.v(202[9] 210[6])
    defparam smpl_register_i0_i18.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i17 (.D(wb_odata[17]), .SP(dac_clk_p_c_enable_272), 
            .CK(dac_clk_p_c), .Q(smpl_register[17]));   // d:/documents/git_local/fm_modulator/rtl/top.v(202[9] 210[6])
    defparam smpl_register_i0_i17.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i16 (.D(wb_odata[16]), .SP(dac_clk_p_c_enable_272), 
            .CK(dac_clk_p_c), .Q(smpl_register[16]));   // d:/documents/git_local/fm_modulator/rtl/top.v(202[9] 210[6])
    defparam smpl_register_i0_i16.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i15 (.D(wb_odata[15]), .SP(dac_clk_p_c_enable_272), 
            .CK(dac_clk_p_c), .Q(smpl_register[15]));   // d:/documents/git_local/fm_modulator/rtl/top.v(202[9] 210[6])
    defparam smpl_register_i0_i15.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i14 (.D(wb_odata[14]), .SP(dac_clk_p_c_enable_272), 
            .CK(dac_clk_p_c), .Q(smpl_register[14]));   // d:/documents/git_local/fm_modulator/rtl/top.v(202[9] 210[6])
    defparam smpl_register_i0_i14.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i13 (.D(wb_odata[13]), .SP(dac_clk_p_c_enable_272), 
            .CK(dac_clk_p_c), .Q(smpl_register[13]));   // d:/documents/git_local/fm_modulator/rtl/top.v(202[9] 210[6])
    defparam smpl_register_i0_i13.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i12 (.D(wb_odata[12]), .SP(dac_clk_p_c_enable_272), 
            .CK(dac_clk_p_c), .Q(smpl_register[12]));   // d:/documents/git_local/fm_modulator/rtl/top.v(202[9] 210[6])
    defparam smpl_register_i0_i12.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i11 (.D(wb_odata[11]), .SP(dac_clk_p_c_enable_272), 
            .CK(dac_clk_p_c), .Q(smpl_register[11]));   // d:/documents/git_local/fm_modulator/rtl/top.v(202[9] 210[6])
    defparam smpl_register_i0_i11.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i10 (.D(wb_odata[10]), .SP(dac_clk_p_c_enable_272), 
            .CK(dac_clk_p_c), .Q(smpl_register[10]));   // d:/documents/git_local/fm_modulator/rtl/top.v(202[9] 210[6])
    defparam smpl_register_i0_i10.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i9 (.D(wb_odata[9]), .SP(dac_clk_p_c_enable_272), 
            .CK(dac_clk_p_c), .Q(smpl_register[9]));   // d:/documents/git_local/fm_modulator/rtl/top.v(202[9] 210[6])
    defparam smpl_register_i0_i9.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i8 (.D(wb_odata[8]), .SP(dac_clk_p_c_enable_272), 
            .CK(dac_clk_p_c), .Q(smpl_register[8]));   // d:/documents/git_local/fm_modulator/rtl/top.v(202[9] 210[6])
    defparam smpl_register_i0_i8.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i7 (.D(wb_odata[7]), .SP(dac_clk_p_c_enable_272), 
            .CK(dac_clk_p_c), .Q(smpl_register[7]));   // d:/documents/git_local/fm_modulator/rtl/top.v(202[9] 210[6])
    defparam smpl_register_i0_i7.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i6 (.D(wb_odata[6]), .SP(dac_clk_p_c_enable_272), 
            .CK(dac_clk_p_c), .Q(smpl_register[6]));   // d:/documents/git_local/fm_modulator/rtl/top.v(202[9] 210[6])
    defparam smpl_register_i0_i6.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i5 (.D(wb_odata[5]), .SP(dac_clk_p_c_enable_272), 
            .CK(dac_clk_p_c), .Q(smpl_register[5]));   // d:/documents/git_local/fm_modulator/rtl/top.v(202[9] 210[6])
    defparam smpl_register_i0_i5.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i4 (.D(wb_odata[4]), .SP(dac_clk_p_c_enable_272), 
            .CK(dac_clk_p_c), .Q(smpl_register[4]));   // d:/documents/git_local/fm_modulator/rtl/top.v(202[9] 210[6])
    defparam smpl_register_i0_i4.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i3 (.D(wb_odata[3]), .SP(dac_clk_p_c_enable_272), 
            .CK(dac_clk_p_c), .Q(smpl_register[3]));   // d:/documents/git_local/fm_modulator/rtl/top.v(202[9] 210[6])
    defparam smpl_register_i0_i3.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i2 (.D(wb_odata[2]), .SP(dac_clk_p_c_enable_272), 
            .CK(dac_clk_p_c), .Q(smpl_register[2]));   // d:/documents/git_local/fm_modulator/rtl/top.v(202[9] 210[6])
    defparam smpl_register_i0_i2.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i1 (.D(wb_odata[1]), .SP(dac_clk_p_c_enable_272), 
            .CK(dac_clk_p_c), .Q(smpl_register[1]));   // d:/documents/git_local/fm_modulator/rtl/top.v(202[9] 210[6])
    defparam smpl_register_i0_i1.GSR = "DISABLED";
    LUT4 i1_3_lut_4_lut (.A(wb_addr[1]), .B(n26535), .C(wb_addr[15]), 
         .D(n26563), .Z(n20402)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(241[23:49])
    defparam i1_3_lut_4_lut.init = 16'hffef;
    PFUMX mux_388_Mux_4_i3 (.BLUT(n1_adj_3081), .ALUT(n2_adj_3080), .C0(wb_addr[1]), 
          .Z(n2032));
    LUT4 i1_4_lut_adj_144 (.A(n20906), .B(n20922), .C(n20918), .D(chg_counter_23__N_406), 
         .Z(dac_clk_p_c_enable_174)) /* synthesis lut_function=((((D)+!C)+!B)+!A) */ ;
    defparam i1_4_lut_adj_144.init = 16'hff7f;
    LUT4 i18661_4_lut (.A(chg_counter[9]), .B(chg_counter[15]), .C(chg_counter[5]), 
         .D(chg_counter[6]), .Z(n20906)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i18661_4_lut.init = 16'h8000;
    LUT4 i18677_4_lut (.A(n20886), .B(n20912), .C(n20910), .D(n20888), 
         .Z(n20922)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i18677_4_lut.init = 16'h8000;
    LUT4 i18673_4_lut (.A(chg_counter[4]), .B(n20904), .C(n20872), .D(chg_counter[14]), 
         .Z(n20918)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i18673_4_lut.init = 16'h8000;
    LUT4 i18641_2_lut (.A(chg_counter[10]), .B(chg_counter[13]), .Z(n20886)) /* synthesis lut_function=(A (B)) */ ;
    defparam i18641_2_lut.init = 16'h8888;
    LUT4 i18667_4_lut (.A(chg_counter[22]), .B(chg_counter[8]), .C(chg_counter[1]), 
         .D(chg_counter[21]), .Z(n20912)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i18667_4_lut.init = 16'h8000;
    LUT4 i18665_4_lut (.A(chg_counter[16]), .B(chg_counter[11]), .C(chg_counter[23]), 
         .D(chg_counter[2]), .Z(n20910)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i18665_4_lut.init = 16'h8000;
    LUT4 i18643_2_lut (.A(chg_counter[3]), .B(chg_counter[20]), .Z(n20888)) /* synthesis lut_function=(A (B)) */ ;
    defparam i18643_2_lut.init = 16'h8888;
    LUT4 i18659_4_lut (.A(chg_counter[19]), .B(chg_counter[18]), .C(chg_counter[7]), 
         .D(chg_counter[0]), .Z(n20904)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i18659_4_lut.init = 16'h8000;
    LUT4 i18627_2_lut (.A(chg_counter[12]), .B(chg_counter[17]), .Z(n20872)) /* synthesis lut_function=(A (B)) */ ;
    defparam i18627_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_145 (.A(wb_addr[8]), .B(n26403), .C(n20774), .D(wb_addr[9]), 
         .Z(none_sel)) /* synthesis lut_function=(A (B+(C))+!A (B+(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(241[23:49])
    defparam i1_4_lut_adj_145.init = 16'hfcfd;
    PFUMX mux_388_Mux_19_i3 (.BLUT(n1_adj_3057), .ALUT(n2_adj_3056), .C0(wb_addr[1]), 
          .Z(n2017));
    LUT4 i1_4_lut_adj_146 (.A(n26563), .B(n38), .C(n34), .D(n20708), 
         .Z(o_dac_a_9__N_1)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut_adj_146.init = 16'h0100;
    LUT4 i1_4_lut_adj_147 (.A(wb_addr[8]), .B(wb_addr[12]), .C(n20702), 
         .D(wb_addr[9]), .Z(n20708)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_4_lut_adj_147.init = 16'h1000;
    LUT4 i1_2_lut_adj_148 (.A(wb_addr[15]), .B(wb_stb), .Z(n20702)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_148.init = 16'h8888;
    LUT4 mux_388_Mux_15_i2_3_lut (.A(bus_err_address[13]), .B(power_counter[15]), 
         .C(wb_addr[0]), .Z(n2_adj_3061)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(213[3] 220[10])
    defparam mux_388_Mux_15_i2_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_409_3_lut_4_lut (.A(n26563), .B(wb_addr[12]), .C(n20774), 
         .D(n38), .Z(n26369)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(241[23:49])
    defparam i1_2_lut_rep_409_3_lut_4_lut.init = 16'hfffe;
    LUT4 i11160_2_lut (.A(smpl_register[15]), .B(wb_addr[0]), .Z(n1_adj_3062)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(213[3] 220[10])
    defparam i11160_2_lut.init = 16'h8888;
    LUT4 power_counter_31__I_0_75_i1_3_lut (.A(power_counter_31__N_232[0]), 
         .B(power_counter_31__N_201[0]), .C(power_counter[31]), .Z(power_counter_31__N_129[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(229[4:54])
    defparam power_counter_31__I_0_75_i1_3_lut.init = 16'hcaca;
    LUT4 mux_388_Mux_14_i2_3_lut (.A(bus_err_address[12]), .B(power_counter[14]), 
         .C(wb_addr[0]), .Z(n2_adj_3063)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(213[3] 220[10])
    defparam mux_388_Mux_14_i2_3_lut.init = 16'hcaca;
    LUT4 i11159_2_lut (.A(smpl_register[14]), .B(wb_addr[0]), .Z(n1_adj_3064)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(213[3] 220[10])
    defparam i11159_2_lut.init = 16'h8888;
    LUT4 mux_388_Mux_13_i2_3_lut (.A(bus_err_address[11]), .B(power_counter[13]), 
         .C(wb_addr[0]), .Z(n2_adj_3065)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(213[3] 220[10])
    defparam mux_388_Mux_13_i2_3_lut.init = 16'hcaca;
    LUT4 i11158_2_lut (.A(smpl_register[13]), .B(wb_addr[0]), .Z(n1_adj_3066)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(213[3] 220[10])
    defparam i11158_2_lut.init = 16'h8888;
    LUT4 mux_388_Mux_12_i2_3_lut (.A(bus_err_address[10]), .B(power_counter[12]), 
         .C(wb_addr[0]), .Z(n2_adj_3067)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(213[3] 220[10])
    defparam mux_388_Mux_12_i2_3_lut.init = 16'hcaca;
    LUT4 i11157_2_lut (.A(smpl_register[12]), .B(wb_addr[0]), .Z(n1_adj_3068)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(213[3] 220[10])
    defparam i11157_2_lut.init = 16'h8888;
    LUT4 mux_388_Mux_11_i2_3_lut (.A(bus_err_address[9]), .B(power_counter[11]), 
         .C(wb_addr[0]), .Z(n2_adj_3069)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(213[3] 220[10])
    defparam mux_388_Mux_11_i2_3_lut.init = 16'hcaca;
    LUT4 i11156_2_lut (.A(smpl_register[11]), .B(wb_addr[0]), .Z(n1_adj_3070)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(213[3] 220[10])
    defparam i11156_2_lut.init = 16'h8888;
    LUT4 wb_idata_31__I_0_i1_3_lut (.A(wb_idata_31__N_266[0]), .B(wb_fm_data[0]), 
         .C(wb_fm_ack), .Z(wb_idata_31__N_2[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(268[8] 273[53])
    defparam wb_idata_31__I_0_i1_3_lut.init = 16'hcaca;
    LUT4 mux_57_i1_4_lut (.A(wb_lo_data[0]), .B(wb_smpl_data[0]), .C(wb_smpl_ack), 
         .D(wb_lo_ack), .Z(wb_idata_31__N_266[0])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[8] 273[53])
    defparam mux_57_i1_4_lut.init = 16'hcac0;
    LUT4 mux_388_Mux_10_i2_3_lut (.A(bus_err_address[8]), .B(power_counter[10]), 
         .C(wb_addr[0]), .Z(n2_adj_3071)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(213[3] 220[10])
    defparam mux_388_Mux_10_i2_3_lut.init = 16'hcaca;
    LUT4 mux_388_Mux_9_i2_3_lut (.A(bus_err_address[7]), .B(power_counter[9]), 
         .C(wb_addr[0]), .Z(n2_adj_3072)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(213[3] 220[10])
    defparam mux_388_Mux_9_i2_3_lut.init = 16'hcaca;
    LUT4 i22397_4_lut (.A(n26369), .B(n26564), .C(n26557), .D(n7), .Z(dac_clk_p_c_enable_198)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(202[9] 210[6])
    defparam i22397_4_lut.init = 16'h0010;
    LUT4 i1_4_lut_adj_149 (.A(wb_addr[1]), .B(wb_addr[2]), .C(wb_addr[0]), 
         .D(wb_addr[3]), .Z(n7)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(207[4:8])
    defparam i1_4_lut_adj_149.init = 16'hfffb;
    LUT4 i1_2_lut_adj_150 (.A(wb_fm_ack), .B(wb_lo_ack), .Z(n4)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(263[13:56])
    defparam i1_2_lut_adj_150.init = 16'heeee;
    LUT4 i1_2_lut_adj_151 (.A(wb_addr[15]), .B(n34), .Z(n20774)) /* synthesis lut_function=((B)+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(241[23:49])
    defparam i1_2_lut_adj_151.init = 16'hdddd;
    PFUMX mux_388_Mux_21_i3 (.BLUT(n1_adj_3054), .ALUT(n2_adj_3053), .C0(wb_addr[1]), 
          .Z(n2015));
    LUT4 i1_4_lut_adj_152 (.A(n20466), .B(n20468), .C(n20470), .D(n20456), 
         .Z(n38)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(241[23:49])
    defparam i1_4_lut_adj_152.init = 16'hfffe;
    LUT4 i1_2_lut_adj_153 (.A(wb_addr[11]), .B(wb_addr[16]), .Z(n20466)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(241[23:49])
    defparam i1_2_lut_adj_153.init = 16'heeee;
    LUT4 i1_4_lut_adj_154 (.A(wb_addr[17]), .B(wb_addr[14]), .C(wb_addr[23]), 
         .D(wb_addr[20]), .Z(n20468)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(241[23:49])
    defparam i1_4_lut_adj_154.init = 16'hfffe;
    LUT4 i1_4_lut_adj_155 (.A(wb_addr[25]), .B(wb_addr[10]), .C(wb_addr[26]), 
         .D(wb_addr[21]), .Z(n20470)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(241[23:49])
    defparam i1_4_lut_adj_155.init = 16'hfffe;
    LUT4 i1_2_lut_adj_156 (.A(wb_addr[27]), .B(wb_addr[18]), .Z(n20456)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(241[23:49])
    defparam i1_2_lut_adj_156.init = 16'heeee;
    LUT4 mux_388_Mux_8_i2_3_lut (.A(bus_err_address[6]), .B(power_counter[8]), 
         .C(wb_addr[0]), .Z(n2_adj_3073)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(213[3] 220[10])
    defparam mux_388_Mux_8_i2_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_157 (.A(wb_addr[28]), .B(wb_addr[19]), .C(wb_addr[13]), 
         .D(wb_addr[29]), .Z(n34)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(241[23:49])
    defparam i1_4_lut_adj_157.init = 16'hfffe;
    PFUMX mux_388_Mux_22_i3 (.BLUT(n1_adj_3052), .ALUT(n2_adj_3051), .C0(wb_addr[1]), 
          .Z(n2014));
    PFUMX mux_388_Mux_6_i3 (.BLUT(n1_adj_3078), .ALUT(n2_adj_3077), .C0(wb_addr[1]), 
          .Z(n2030));
    LUT4 i11153_2_lut (.A(smpl_register[8]), .B(wb_addr[0]), .Z(n1_adj_3074)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(213[3] 220[10])
    defparam i11153_2_lut.init = 16'h8888;
    PFUMX mux_388_Mux_23_i3 (.BLUT(n1_adj_3050), .ALUT(n2_adj_3049), .C0(wb_addr[1]), 
          .Z(n2013));
    PFUMX mux_388_Mux_7_i3 (.BLUT(n1_adj_3076), .ALUT(n2_adj_3075), .C0(wb_addr[1]), 
          .Z(n2029));
    PFUMX mux_388_Mux_24_i3 (.BLUT(n1_adj_3048), .ALUT(n2_adj_3047), .C0(wb_addr[1]), 
          .Z(n2012));
    PFUMX mux_388_Mux_25_i3 (.BLUT(n1_adj_3046), .ALUT(n2_adj_3045), .C0(wb_addr[1]), 
          .Z(n2011));
    LUT4 mux_388_Mux_31_i2_3_lut (.A(bus_err_address[29]), .B(power_counter[31]), 
         .C(wb_addr[0]), .Z(n2_adj_3035)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(213[3] 220[10])
    defparam mux_388_Mux_31_i2_3_lut.init = 16'hcaca;
    LUT4 i11176_2_lut (.A(smpl_register[31]), .B(wb_addr[0]), .Z(n1)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(213[3] 220[10])
    defparam i11176_2_lut.init = 16'h8888;
    LUT4 mux_388_Mux_30_i2_3_lut (.A(bus_err_address[28]), .B(power_counter[30]), 
         .C(wb_addr[0]), .Z(n2_adj_3036)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(213[3] 220[10])
    defparam mux_388_Mux_30_i2_3_lut.init = 16'hcaca;
    LUT4 i11175_2_lut (.A(smpl_register[30]), .B(wb_addr[0]), .Z(n1_adj_3037)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(213[3] 220[10])
    defparam i11175_2_lut.init = 16'h8888;
    LUT4 mux_388_Mux_29_i2_3_lut (.A(bus_err_address[27]), .B(power_counter[29]), 
         .C(wb_addr[0]), .Z(n2_adj_3038)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(213[3] 220[10])
    defparam mux_388_Mux_29_i2_3_lut.init = 16'hcaca;
    LUT4 mux_388_Mux_28_i2_3_lut (.A(bus_err_address[26]), .B(power_counter[28]), 
         .C(wb_addr[0]), .Z(n2_adj_3039)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(213[3] 220[10])
    defparam mux_388_Mux_28_i2_3_lut.init = 16'hcaca;
    PFUMX mux_388_Mux_26_i3 (.BLUT(n1_adj_3044), .ALUT(n2_adj_3043), .C0(wb_addr[1]), 
          .Z(n2010));
    LUT4 i11173_2_lut (.A(smpl_register[28]), .B(wb_addr[0]), .Z(n1_adj_3040)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(213[3] 220[10])
    defparam i11173_2_lut.init = 16'h8888;
    LUT4 mux_388_Mux_27_i2_3_lut (.A(bus_err_address[25]), .B(power_counter[27]), 
         .C(wb_addr[0]), .Z(n2_adj_3041)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(213[3] 220[10])
    defparam mux_388_Mux_27_i2_3_lut.init = 16'hcaca;
    PFUMX mux_388_Mux_27_i3 (.BLUT(n1_adj_3042), .ALUT(n2_adj_3041), .C0(wb_addr[1]), 
          .Z(n2009));
    LUT4 i11172_2_lut (.A(smpl_register[27]), .B(wb_addr[0]), .Z(n1_adj_3042)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(213[3] 220[10])
    defparam i11172_2_lut.init = 16'h8888;
    LUT4 mux_388_Mux_7_i2_3_lut (.A(bus_err_address[5]), .B(power_counter[7]), 
         .C(wb_addr[0]), .Z(n2_adj_3075)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(213[3] 220[10])
    defparam mux_388_Mux_7_i2_3_lut.init = 16'hcaca;
    LUT4 mux_388_Mux_26_i2_3_lut (.A(bus_err_address[24]), .B(power_counter[26]), 
         .C(wb_addr[0]), .Z(n2_adj_3043)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(213[3] 220[10])
    defparam mux_388_Mux_26_i2_3_lut.init = 16'hcaca;
    LUT4 i11171_2_lut (.A(smpl_register[26]), .B(wb_addr[0]), .Z(n1_adj_3044)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(213[3] 220[10])
    defparam i11171_2_lut.init = 16'h8888;
    PFUMX mux_388_Mux_28_i3 (.BLUT(n1_adj_3040), .ALUT(n2_adj_3039), .C0(wb_addr[1]), 
          .Z(n2008));
    LUT4 mux_388_Mux_25_i2_3_lut (.A(bus_err_address[23]), .B(power_counter[25]), 
         .C(wb_addr[0]), .Z(n2_adj_3045)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(213[3] 220[10])
    defparam mux_388_Mux_25_i2_3_lut.init = 16'hcaca;
    LUT4 i11170_2_lut (.A(smpl_register[25]), .B(wb_addr[0]), .Z(n1_adj_3046)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(213[3] 220[10])
    defparam i11170_2_lut.init = 16'h8888;
    LUT4 mux_388_Mux_24_i2_3_lut (.A(bus_err_address[22]), .B(power_counter[24]), 
         .C(wb_addr[0]), .Z(n2_adj_3047)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(213[3] 220[10])
    defparam mux_388_Mux_24_i2_3_lut.init = 16'hcaca;
    PFUMX mux_388_Mux_8_i3 (.BLUT(n1_adj_3074), .ALUT(n2_adj_3073), .C0(wb_addr[1]), 
          .Z(n2028));
    LUT4 i11169_2_lut (.A(smpl_register[24]), .B(wb_addr[0]), .Z(n1_adj_3048)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(213[3] 220[10])
    defparam i11169_2_lut.init = 16'h8888;
    LUT4 i11152_2_lut (.A(smpl_register[7]), .B(wb_addr[0]), .Z(n1_adj_3076)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(213[3] 220[10])
    defparam i11152_2_lut.init = 16'h8888;
    LUT4 mux_388_Mux_23_i2_3_lut (.A(bus_err_address[21]), .B(power_counter[23]), 
         .C(wb_addr[0]), .Z(n2_adj_3049)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(213[3] 220[10])
    defparam mux_388_Mux_23_i2_3_lut.init = 16'hcaca;
    LUT4 i11168_2_lut (.A(smpl_register[23]), .B(wb_addr[0]), .Z(n1_adj_3050)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(213[3] 220[10])
    defparam i11168_2_lut.init = 16'h8888;
    LUT4 mux_388_Mux_22_i2_3_lut (.A(bus_err_address[20]), .B(power_counter[22]), 
         .C(wb_addr[0]), .Z(n2_adj_3051)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(213[3] 220[10])
    defparam mux_388_Mux_22_i2_3_lut.init = 16'hcaca;
    LUT4 mux_388_Mux_6_i2_3_lut (.A(bus_err_address[4]), .B(power_counter[6]), 
         .C(wb_addr[0]), .Z(n2_adj_3077)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(213[3] 220[10])
    defparam mux_388_Mux_6_i2_3_lut.init = 16'hcaca;
    PFUMX mux_388_Mux_30_i3 (.BLUT(n1_adj_3037), .ALUT(n2_adj_3036), .C0(wb_addr[1]), 
          .Z(n2006));
    LUT4 i11167_2_lut (.A(smpl_register[22]), .B(wb_addr[0]), .Z(n1_adj_3052)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(213[3] 220[10])
    defparam i11167_2_lut.init = 16'h8888;
    LUT4 i11151_2_lut (.A(smpl_register[6]), .B(wb_addr[0]), .Z(n1_adj_3078)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(213[3] 220[10])
    defparam i11151_2_lut.init = 16'h8888;
    PFUMX mux_388_Mux_31_i3 (.BLUT(n1), .ALUT(n2_adj_3035), .C0(wb_addr[1]), 
          .Z(n2005));
    LUT4 i1_2_lut_3_lut_4_lut (.A(n38), .B(n26453), .C(n26564), .D(n20774), 
         .Z(wb_smpl_sel_N_311)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(241[23:49])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 mux_388_Mux_21_i2_3_lut (.A(bus_err_address[19]), .B(power_counter[21]), 
         .C(wb_addr[0]), .Z(n2_adj_3053)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(213[3] 220[10])
    defparam mux_388_Mux_21_i2_3_lut.init = 16'hcaca;
    LUT4 mux_388_Mux_5_i2_3_lut (.A(bus_err_address[3]), .B(power_counter[5]), 
         .C(wb_addr[0]), .Z(n2_adj_3079)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(213[3] 220[10])
    defparam mux_388_Mux_5_i2_3_lut.init = 16'hcaca;
    LUT4 i11166_2_lut (.A(smpl_register[21]), .B(wb_addr[0]), .Z(n1_adj_3054)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(213[3] 220[10])
    defparam i11166_2_lut.init = 16'h8888;
    LUT4 mux_388_Mux_20_i2_3_lut (.A(bus_err_address[18]), .B(power_counter[20]), 
         .C(wb_addr[0]), .Z(n2_adj_3055)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(213[3] 220[10])
    defparam mux_388_Mux_20_i2_3_lut.init = 16'hcaca;
    LUT4 mux_388_Mux_19_i2_3_lut (.A(bus_err_address[17]), .B(power_counter[19]), 
         .C(wb_addr[0]), .Z(n2_adj_3056)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(213[3] 220[10])
    defparam mux_388_Mux_19_i2_3_lut.init = 16'hcaca;
    LUT4 wb_idata_31__I_0_i32_4_lut (.A(wb_smpl_data[31]), .B(wb_fm_data[31]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_2[31])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(268[8] 273[53])
    defparam wb_idata_31__I_0_i32_4_lut.init = 16'hcac0;
    FD1S3AX wb_idata_i31 (.D(wb_idata_31__N_2[31]), .CK(dac_clk_p_c), .Q(wb_idata[31]));   // d:/documents/git_local/fm_modulator/rtl/top.v(265[9] 273[53])
    defparam wb_idata_i31.GSR = "DISABLED";
    LUT4 i10108_1_lut (.A(wb_idata[1]), .Z(n12635)) /* synthesis lut_function=(!(A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(265[9] 273[53])
    defparam i10108_1_lut.init = 16'h5555;
    LUT4 wb_idata_31__I_0_i31_4_lut (.A(wb_smpl_data[30]), .B(wb_fm_data[30]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_2[30])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(268[8] 273[53])
    defparam wb_idata_31__I_0_i31_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i30_4_lut (.A(wb_smpl_data[29]), .B(wb_fm_data[29]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_2[29])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(268[8] 273[53])
    defparam wb_idata_31__I_0_i30_4_lut.init = 16'hcac0;
    LUT4 mux_387_i1_4_lut (.A(smpl_interrupt), .B(n20770), .C(n7), .D(n9787), 
         .Z(wb_smpl_data_31__N_64[0])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(213[3] 220[10])
    defparam mux_387_i1_4_lut.init = 16'hca0a;
    LUT4 i1_3_lut (.A(wb_addr[3]), .B(wb_addr[2]), .C(wb_addr[0]), .Z(n20770)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_3_lut.init = 16'h1010;
    LUT4 i7406_3_lut (.A(smpl_register[0]), .B(power_counter[0]), .C(wb_addr[1]), 
         .Z(n9787)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(213[3] 220[10])
    defparam i7406_3_lut.init = 16'hcaca;
    LUT4 wb_idata_31__I_0_i29_4_lut (.A(wb_smpl_data[28]), .B(wb_fm_data[28]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_2[28])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(268[8] 273[53])
    defparam wb_idata_31__I_0_i29_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i28_4_lut (.A(wb_smpl_data[27]), .B(wb_fm_data[27]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_2[27])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(268[8] 273[53])
    defparam wb_idata_31__I_0_i28_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i27_4_lut (.A(wb_smpl_data[26]), .B(wb_fm_data[26]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_2[26])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(268[8] 273[53])
    defparam wb_idata_31__I_0_i27_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i26_4_lut (.A(wb_smpl_data[25]), .B(wb_fm_data[25]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_2[25])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(268[8] 273[53])
    defparam wb_idata_31__I_0_i26_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i25_4_lut (.A(wb_smpl_data[24]), .B(wb_fm_data[24]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_2[24])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(268[8] 273[53])
    defparam wb_idata_31__I_0_i25_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i24_4_lut (.A(wb_smpl_data[23]), .B(wb_fm_data[23]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_2[23])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(268[8] 273[53])
    defparam wb_idata_31__I_0_i24_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i23_4_lut (.A(wb_smpl_data[22]), .B(wb_fm_data[22]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_2[22])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(268[8] 273[53])
    defparam wb_idata_31__I_0_i23_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i22_4_lut (.A(wb_smpl_data[21]), .B(wb_fm_data[21]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_2[21])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(268[8] 273[53])
    defparam wb_idata_31__I_0_i22_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i21_4_lut (.A(wb_smpl_data[20]), .B(wb_fm_data[20]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_2[20])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(268[8] 273[53])
    defparam wb_idata_31__I_0_i21_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i20_4_lut (.A(wb_smpl_data[19]), .B(wb_fm_data[19]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_2[19])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(268[8] 273[53])
    defparam wb_idata_31__I_0_i20_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i19_4_lut (.A(wb_smpl_data[18]), .B(wb_fm_data[18]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_2[18])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(268[8] 273[53])
    defparam wb_idata_31__I_0_i19_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i18_4_lut (.A(wb_smpl_data[17]), .B(wb_fm_data[17]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_2[17])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(268[8] 273[53])
    defparam wb_idata_31__I_0_i18_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i17_4_lut (.A(wb_smpl_data[16]), .B(wb_fm_data[16]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_2[16])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(268[8] 273[53])
    defparam wb_idata_31__I_0_i17_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i16_4_lut (.A(wb_smpl_data[15]), .B(wb_fm_data[15]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_2[15])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(268[8] 273[53])
    defparam wb_idata_31__I_0_i16_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i15_4_lut (.A(wb_smpl_data[14]), .B(wb_fm_data[14]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_2[14])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(268[8] 273[53])
    defparam wb_idata_31__I_0_i15_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i14_4_lut (.A(wb_smpl_data[13]), .B(wb_fm_data[13]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_2[13])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(268[8] 273[53])
    defparam wb_idata_31__I_0_i14_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i13_4_lut (.A(wb_smpl_data[12]), .B(wb_fm_data[12]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_2[12])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(268[8] 273[53])
    defparam wb_idata_31__I_0_i13_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i12_4_lut (.A(wb_smpl_data[11]), .B(wb_fm_data[11]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_2[11])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(268[8] 273[53])
    defparam wb_idata_31__I_0_i12_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i11_4_lut (.A(wb_smpl_data[10]), .B(wb_fm_data[10]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_2[10])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(268[8] 273[53])
    defparam wb_idata_31__I_0_i11_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i10_4_lut (.A(wb_smpl_data[9]), .B(wb_fm_data[9]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_2[9])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(268[8] 273[53])
    defparam wb_idata_31__I_0_i10_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i9_4_lut (.A(wb_smpl_data[8]), .B(wb_fm_data[8]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_2[8])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(268[8] 273[53])
    defparam wb_idata_31__I_0_i9_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i8_3_lut (.A(wb_idata_31__N_266[7]), .B(wb_fm_data[7]), 
         .C(wb_fm_ack), .Z(wb_idata_31__N_2[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(268[8] 273[53])
    defparam wb_idata_31__I_0_i8_3_lut.init = 16'hcaca;
    LUT4 mux_57_i8_4_lut (.A(wb_lo_data[7]), .B(wb_smpl_data[7]), .C(wb_smpl_ack), 
         .D(wb_lo_ack), .Z(wb_idata_31__N_266[7])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[8] 273[53])
    defparam mux_57_i8_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i7_3_lut (.A(wb_idata_31__N_266[6]), .B(wb_fm_data[6]), 
         .C(wb_fm_ack), .Z(wb_idata_31__N_2[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(268[8] 273[53])
    defparam wb_idata_31__I_0_i7_3_lut.init = 16'hcaca;
    LUT4 mux_57_i7_4_lut (.A(wb_lo_data[6]), .B(wb_smpl_data[6]), .C(wb_smpl_ack), 
         .D(wb_lo_ack), .Z(wb_idata_31__N_266[6])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[8] 273[53])
    defparam mux_57_i7_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i6_3_lut (.A(wb_idata_31__N_266[5]), .B(wb_fm_data[5]), 
         .C(wb_fm_ack), .Z(wb_idata_31__N_2[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(268[8] 273[53])
    defparam wb_idata_31__I_0_i6_3_lut.init = 16'hcaca;
    LUT4 mux_57_i6_4_lut (.A(wb_lo_data[5]), .B(wb_smpl_data[5]), .C(wb_smpl_ack), 
         .D(wb_lo_ack), .Z(wb_idata_31__N_266[5])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[8] 273[53])
    defparam mux_57_i6_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i5_3_lut (.A(wb_idata_31__N_266[4]), .B(wb_fm_data[4]), 
         .C(wb_fm_ack), .Z(wb_idata_31__N_2[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(268[8] 273[53])
    defparam wb_idata_31__I_0_i5_3_lut.init = 16'hcaca;
    LUT4 mux_57_i5_4_lut (.A(wb_lo_data[4]), .B(wb_smpl_data[4]), .C(wb_smpl_ack), 
         .D(wb_lo_ack), .Z(wb_idata_31__N_266[4])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[8] 273[53])
    defparam mux_57_i5_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i4_3_lut (.A(wb_idata_31__N_266[3]), .B(wb_fm_data[3]), 
         .C(wb_fm_ack), .Z(wb_idata_31__N_2[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(268[8] 273[53])
    defparam wb_idata_31__I_0_i4_3_lut.init = 16'hcaca;
    LUT4 mux_57_i4_4_lut (.A(wb_lo_data[3]), .B(wb_smpl_data[3]), .C(wb_smpl_ack), 
         .D(wb_lo_ack), .Z(wb_idata_31__N_266[3])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[8] 273[53])
    defparam mux_57_i4_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i3_3_lut (.A(wb_idata_31__N_266[2]), .B(wb_fm_data[2]), 
         .C(wb_fm_ack), .Z(wb_idata_31__N_2[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(268[8] 273[53])
    defparam wb_idata_31__I_0_i3_3_lut.init = 16'hcaca;
    LUT4 mux_57_i3_4_lut (.A(wb_lo_data[2]), .B(wb_smpl_data[2]), .C(wb_smpl_ack), 
         .D(wb_lo_ack), .Z(wb_idata_31__N_266[2])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[8] 273[53])
    defparam mux_57_i3_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i2_3_lut (.A(wb_idata_31__N_266[1]), .B(wb_fm_data[1]), 
         .C(wb_fm_ack), .Z(wb_idata_31__N_2[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(268[8] 273[53])
    defparam wb_idata_31__I_0_i2_3_lut.init = 16'hcaca;
    LUT4 mux_57_i2_4_lut (.A(wb_lo_data[1]), .B(wb_smpl_data[1]), .C(wb_smpl_ack), 
         .D(wb_lo_ack), .Z(wb_idata_31__N_266[1])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[8] 273[53])
    defparam mux_57_i2_4_lut.init = 16'hcac0;
    LUT4 mux_388_Mux_4_i2_3_lut (.A(bus_err_address[2]), .B(power_counter[4]), 
         .C(wb_addr[0]), .Z(n2_adj_3080)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(213[3] 220[10])
    defparam mux_388_Mux_4_i2_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_75_i31_3_lut (.A(power_counter_31__N_232[30]), 
         .B(power_counter_31__N_201[30]), .C(power_counter[31]), .Z(power_counter_31__N_129[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(229[4:54])
    defparam power_counter_31__I_0_75_i31_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_75_i30_3_lut (.A(power_counter_31__N_232[29]), 
         .B(power_counter_31__N_201[29]), .C(power_counter[31]), .Z(power_counter_31__N_129[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(229[4:54])
    defparam power_counter_31__I_0_75_i30_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_597 (.A(wb_stb), .B(wb_we), .Z(n26557)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(203[7:30])
    defparam i1_2_lut_rep_597.init = 16'h8888;
    LUT4 i18620_2_lut_3_lut (.A(wb_stb), .B(wb_we), .C(wb_addr[0]), .Z(n20864)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(203[7:30])
    defparam i18620_2_lut_3_lut.init = 16'h8080;
    LUT4 power_counter_31__I_0_75_i29_3_lut (.A(power_counter_31__N_232[28]), 
         .B(power_counter_31__N_201[28]), .C(power_counter[31]), .Z(power_counter_31__N_129[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(229[4:54])
    defparam power_counter_31__I_0_75_i29_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_75_i28_3_lut (.A(power_counter_31__N_232[27]), 
         .B(power_counter_31__N_201[27]), .C(power_counter[31]), .Z(power_counter_31__N_129[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(229[4:54])
    defparam power_counter_31__I_0_75_i28_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_75_i27_3_lut (.A(power_counter_31__N_232[26]), 
         .B(power_counter_31__N_201[26]), .C(power_counter[31]), .Z(power_counter_31__N_129[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(229[4:54])
    defparam power_counter_31__I_0_75_i27_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_75_i26_3_lut (.A(power_counter_31__N_232[25]), 
         .B(power_counter_31__N_201[25]), .C(power_counter[31]), .Z(power_counter_31__N_129[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(229[4:54])
    defparam power_counter_31__I_0_75_i26_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_75_i25_3_lut (.A(power_counter_31__N_232[24]), 
         .B(power_counter_31__N_201[24]), .C(power_counter[31]), .Z(power_counter_31__N_129[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(229[4:54])
    defparam power_counter_31__I_0_75_i25_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_75_i24_3_lut (.A(power_counter_31__N_232[23]), 
         .B(power_counter_31__N_201[23]), .C(power_counter[31]), .Z(power_counter_31__N_129[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(229[4:54])
    defparam power_counter_31__I_0_75_i24_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_75_i23_3_lut (.A(power_counter_31__N_232[22]), 
         .B(power_counter_31__N_201[22]), .C(power_counter[31]), .Z(power_counter_31__N_129[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(229[4:54])
    defparam power_counter_31__I_0_75_i23_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_75_i22_3_lut (.A(power_counter_31__N_232[21]), 
         .B(power_counter_31__N_201[21]), .C(power_counter[31]), .Z(power_counter_31__N_129[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(229[4:54])
    defparam power_counter_31__I_0_75_i22_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_75_i21_3_lut (.A(power_counter_31__N_232[20]), 
         .B(power_counter_31__N_201[20]), .C(power_counter[31]), .Z(power_counter_31__N_129[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(229[4:54])
    defparam power_counter_31__I_0_75_i21_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_75_i20_3_lut (.A(power_counter_31__N_232[19]), 
         .B(power_counter_31__N_201[19]), .C(power_counter[31]), .Z(power_counter_31__N_129[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(229[4:54])
    defparam power_counter_31__I_0_75_i20_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_75_i19_3_lut (.A(power_counter_31__N_232[18]), 
         .B(power_counter_31__N_201[18]), .C(power_counter[31]), .Z(power_counter_31__N_129[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(229[4:54])
    defparam power_counter_31__I_0_75_i19_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_75_i18_3_lut (.A(power_counter_31__N_232[17]), 
         .B(power_counter_31__N_201[17]), .C(power_counter[31]), .Z(power_counter_31__N_129[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(229[4:54])
    defparam power_counter_31__I_0_75_i18_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_75_i17_3_lut (.A(power_counter_31__N_232[16]), 
         .B(power_counter_31__N_201[16]), .C(power_counter[31]), .Z(power_counter_31__N_129[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(229[4:54])
    defparam power_counter_31__I_0_75_i17_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_75_i16_3_lut (.A(power_counter_31__N_232[15]), 
         .B(power_counter_31__N_201[15]), .C(power_counter[31]), .Z(power_counter_31__N_129[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(229[4:54])
    defparam power_counter_31__I_0_75_i16_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_75_i15_3_lut (.A(power_counter_31__N_232[14]), 
         .B(power_counter_31__N_201[14]), .C(power_counter[31]), .Z(power_counter_31__N_129[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(229[4:54])
    defparam power_counter_31__I_0_75_i15_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_75_i14_3_lut (.A(power_counter_31__N_232[13]), 
         .B(power_counter_31__N_201[13]), .C(power_counter[31]), .Z(power_counter_31__N_129[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(229[4:54])
    defparam power_counter_31__I_0_75_i14_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_75_i13_3_lut (.A(power_counter_31__N_232[12]), 
         .B(power_counter_31__N_201[12]), .C(power_counter[31]), .Z(power_counter_31__N_129[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(229[4:54])
    defparam power_counter_31__I_0_75_i13_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_75_i12_3_lut (.A(power_counter_31__N_232[11]), 
         .B(power_counter_31__N_201[11]), .C(power_counter[31]), .Z(power_counter_31__N_129[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(229[4:54])
    defparam power_counter_31__I_0_75_i12_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_75_i11_3_lut (.A(power_counter_31__N_232[10]), 
         .B(power_counter_31__N_201[10]), .C(power_counter[31]), .Z(power_counter_31__N_129[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(229[4:54])
    defparam power_counter_31__I_0_75_i11_3_lut.init = 16'hcaca;
    LUT4 i11149_2_lut (.A(smpl_register[4]), .B(wb_addr[0]), .Z(n1_adj_3081)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(213[3] 220[10])
    defparam i11149_2_lut.init = 16'h8888;
    LUT4 power_counter_31__I_0_75_i10_3_lut (.A(power_counter_31__N_232[9]), 
         .B(power_counter_31__N_201[9]), .C(power_counter[31]), .Z(power_counter_31__N_129[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(229[4:54])
    defparam power_counter_31__I_0_75_i10_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_75_i9_3_lut (.A(power_counter_31__N_232[8]), 
         .B(power_counter_31__N_201[8]), .C(power_counter[31]), .Z(power_counter_31__N_129[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(229[4:54])
    defparam power_counter_31__I_0_75_i9_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_75_i8_3_lut (.A(power_counter_31__N_232[7]), 
         .B(power_counter_31__N_201[7]), .C(power_counter[31]), .Z(power_counter_31__N_129[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(229[4:54])
    defparam power_counter_31__I_0_75_i8_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_75_i7_3_lut (.A(power_counter_31__N_232[6]), 
         .B(power_counter_31__N_201[6]), .C(power_counter[31]), .Z(power_counter_31__N_129[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(229[4:54])
    defparam power_counter_31__I_0_75_i7_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_75_i6_3_lut (.A(power_counter_31__N_232[5]), 
         .B(power_counter_31__N_201[5]), .C(power_counter[31]), .Z(power_counter_31__N_129[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(229[4:54])
    defparam power_counter_31__I_0_75_i6_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_75_i5_3_lut (.A(power_counter_31__N_232[4]), 
         .B(power_counter_31__N_201[4]), .C(power_counter[31]), .Z(power_counter_31__N_129[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(229[4:54])
    defparam power_counter_31__I_0_75_i5_3_lut.init = 16'hcaca;
    LUT4 mux_388_Mux_3_i2_3_lut (.A(bus_err_address[1]), .B(power_counter[3]), 
         .C(wb_addr[0]), .Z(n2_adj_3082)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(213[3] 220[10])
    defparam mux_388_Mux_3_i2_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_75_i4_3_lut (.A(power_counter_31__N_232[3]), 
         .B(power_counter_31__N_201[3]), .C(power_counter[31]), .Z(power_counter_31__N_129[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(229[4:54])
    defparam power_counter_31__I_0_75_i4_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_75_i3_3_lut (.A(power_counter_31__N_232[2]), 
         .B(power_counter_31__N_201[2]), .C(power_counter[31]), .Z(power_counter_31__N_129[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(229[4:54])
    defparam power_counter_31__I_0_75_i3_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_75_i2_3_lut (.A(power_counter_31__N_232[1]), 
         .B(power_counter_31__N_201[1]), .C(power_counter[31]), .Z(power_counter_31__N_129[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(229[4:54])
    defparam power_counter_31__I_0_75_i2_3_lut.init = 16'hcaca;
    LUT4 i6_2_lut_rep_603 (.A(wb_addr[22]), .B(wb_addr[24]), .Z(n26563)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(241[23:49])
    defparam i6_2_lut_rep_603.init = 16'heeee;
    LUT4 i1_2_lut_rep_493_3_lut (.A(wb_addr[22]), .B(wb_addr[24]), .C(wb_addr[12]), 
         .Z(n26453)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(241[23:49])
    defparam i1_2_lut_rep_493_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_3_lut (.A(wb_addr[22]), .B(wb_addr[24]), .C(wb_addr[9]), 
         .Z(n20432)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(241[23:49])
    defparam i1_2_lut_3_lut.init = 16'hefef;
    LUT4 i1_2_lut_rep_443_3_lut_4_lut (.A(wb_addr[22]), .B(wb_addr[24]), 
         .C(n38), .D(wb_addr[12]), .Z(n26403)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(241[23:49])
    defparam i1_2_lut_rep_443_3_lut_4_lut.init = 16'hfffe;
    LUT4 dac_clk_p_I_0_1_lut (.A(dac_clk_p_c), .Z(dac_clk_n_c)) /* synthesis lut_function=(!(A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(47[20:30])
    defparam dac_clk_p_I_0_1_lut.init = 16'h5555;
    LUT4 i1_2_lut_rep_604 (.A(wb_addr[9]), .B(wb_addr[8]), .Z(n26564)) /* synthesis lut_function=(A+!(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(241[23:49])
    defparam i1_2_lut_rep_604.init = 16'hbbbb;
    LUT4 i18671_3_lut_4_lut (.A(wb_addr[9]), .B(wb_addr[8]), .C(n34), 
         .D(n9365), .Z(n20916)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(241[23:49])
    defparam i18671_3_lut_4_lut.init = 16'hfffb;
    LUT4 i11148_2_lut (.A(smpl_register[3]), .B(wb_addr[0]), .Z(n1_adj_3083)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(213[3] 220[10])
    defparam i11148_2_lut.init = 16'h8888;
    LUT4 mux_388_Mux_2_i2_3_lut (.A(bus_err_address[0]), .B(power_counter[2]), 
         .C(wb_addr[0]), .Z(n2_adj_3084)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(213[3] 220[10])
    defparam mux_388_Mux_2_i2_3_lut.init = 16'hcaca;
    LUT4 i11147_2_lut (.A(smpl_register[2]), .B(wb_addr[0]), .Z(n1_adj_3085)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(213[3] 220[10])
    defparam i11147_2_lut.init = 16'h8888;
    LUT4 mux_388_Mux_18_i2_3_lut (.A(bus_err_address[16]), .B(power_counter[18]), 
         .C(wb_addr[0]), .Z(n2_adj_3058)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(213[3] 220[10])
    defparam mux_388_Mux_18_i2_3_lut.init = 16'hcaca;
    PFUMX mux_388_Mux_11_i3 (.BLUT(n1_adj_3070), .ALUT(n2_adj_3069), .C0(wb_addr[1]), 
          .Z(n2025));
    PFUMX mux_388_Mux_12_i3 (.BLUT(n1_adj_3068), .ALUT(n2_adj_3067), .C0(wb_addr[1]), 
          .Z(n2024));
    PFUMX mux_388_Mux_13_i3 (.BLUT(n1_adj_3066), .ALUT(n2_adj_3065), .C0(wb_addr[1]), 
          .Z(n2023));
    PFUMX mux_388_Mux_14_i3 (.BLUT(n1_adj_3064), .ALUT(n2_adj_3063), .C0(wb_addr[1]), 
          .Z(n2022));
    PFUMX mux_388_Mux_15_i3 (.BLUT(n1_adj_3062), .ALUT(n2_adj_3061), .C0(wb_addr[1]), 
          .Z(n2021));
    LUT4 i1_2_lut_rep_575 (.A(wb_addr[12]), .B(wb_addr[8]), .Z(n26535)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(241[23:49])
    defparam i1_2_lut_rep_575.init = 16'heeee;
    VLO i1 (.Z(GND_net));
    LUT4 mux_388_Mux_17_i2_3_lut (.A(bus_err_address[15]), .B(power_counter[17]), 
         .C(wb_addr[0]), .Z(n2_adj_3059)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(213[3] 220[10])
    defparam mux_388_Mux_17_i2_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_468_3_lut (.A(wb_addr[12]), .B(wb_addr[8]), .C(wb_addr[1]), 
         .Z(n26428)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(241[23:49])
    defparam i1_2_lut_rep_468_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_3_lut_adj_158 (.A(wb_addr[12]), .B(wb_addr[8]), .C(wb_addr[0]), 
         .Z(n20412)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(241[23:49])
    defparam i1_2_lut_3_lut_adj_158.init = 16'hfefe;
    efb_inst wb_lo_data_7__I_0 (.dac_clk_p_c(dac_clk_p_c), .n26683(n26683), 
            .wb_cyc(wb_cyc), .wb_lo_data_7__N_96(wb_lo_data_7__N_96), .wb_we(wb_we), 
            .\wb_addr[7] (wb_addr[7]), .\wb_addr[6] (wb_addr[6]), .\wb_addr[5] (wb_addr[5]), 
            .\wb_addr[4] (wb_addr[4]), .\wb_addr[3] (wb_addr[3]), .\wb_addr[2] (wb_addr[2]), 
            .\wb_addr[1] (wb_addr[1]), .\wb_addr[0] (wb_addr[0]), .\wb_odata[7] (wb_odata[7]), 
            .\wb_odata[6] (wb_odata[6]), .\wb_odata[5] (wb_odata[5]), .\wb_odata[4] (wb_odata[4]), 
            .\wb_odata[3] (wb_odata[3]), .\wb_odata[2] (wb_odata[2]), .\wb_odata[1] (wb_odata[1]), 
            .\wb_odata[0] (wb_odata[0]), .pll_data_o({pll_data_o}), .pll_ack(pll_ack), 
            .wb_lo_data({wb_lo_data}), .wb_lo_ack(wb_lo_ack), .pll_clk(pll_clk), 
            .pll_rst(pll_rst), .pll_stb(pll_stb), .pll_we(pll_we), .pll_addr({pll_addr}), 
            .pll_data_i({pll_data_i}), .GND_net(GND_net), .VCC_net(VCC_net)) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(177[10] 189[3])
    LUT4 mux_388_Mux_16_i2_3_lut (.A(bus_err_address[14]), .B(power_counter[16]), 
         .C(wb_addr[0]), .Z(n2_adj_3060)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(213[3] 220[10])
    defparam mux_388_Mux_16_i2_3_lut.init = 16'hcaca;
    FD1S3AX wb_idata_i30 (.D(wb_idata_31__N_2[30]), .CK(dac_clk_p_c), .Q(wb_idata[30]));   // d:/documents/git_local/fm_modulator/rtl/top.v(265[9] 273[53])
    defparam wb_idata_i30.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_159 (.A(n26428), .B(n20432), .C(n34), .D(wb_addr[0]), 
         .Z(n20438)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(241[23:49])
    defparam i1_4_lut_adj_159.init = 16'hfffe;
    LUT4 i_resetb_I_0_1_lut_rep_723 (.A(o_dac_cw_b_c_c), .Z(n26683)) /* synthesis lut_function=(!(A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(32[16:25])
    defparam i_resetb_I_0_1_lut_rep_723.init = 16'h5555;
    LUT4 i11537_2_lut_2_lut (.A(o_dac_cw_b_c_c), .B(o_sample_i[14]), .Z(o_dac_a_c_7)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(32[16:25])
    defparam i11537_2_lut_2_lut.init = 16'h4444;
    LUT4 i11540_2_lut_2_lut (.A(o_dac_cw_b_c_c), .B(o_sample_i[11]), .Z(o_dac_a_c_4)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(32[16:25])
    defparam i11540_2_lut_2_lut.init = 16'h4444;
    LUT4 i11541_2_lut_2_lut (.A(o_dac_cw_b_c_c), .B(o_sample_i[10]), .Z(o_dac_a_c_3)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(32[16:25])
    defparam i11541_2_lut_2_lut.init = 16'h4444;
    LUT4 i11542_2_lut_2_lut (.A(o_dac_cw_b_c_c), .B(o_sample_i[9]), .Z(o_dac_a_c_2)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(32[16:25])
    defparam i11542_2_lut_2_lut.init = 16'h4444;
    LUT4 i11543_2_lut_2_lut (.A(o_dac_cw_b_c_c), .B(o_sample_i[8]), .Z(o_dac_a_c_1)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(32[16:25])
    defparam i11543_2_lut_2_lut.init = 16'h4444;
    LUT4 i11025_2_lut_2_lut (.A(o_dac_cw_b_c_c), .B(o_sample_i[7]), .Z(o_dac_a_c_0)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(32[16:25])
    defparam i11025_2_lut_2_lut.init = 16'h4444;
    LUT4 i11538_2_lut_2_lut (.A(o_dac_cw_b_c_c), .B(o_sample_i[13]), .Z(o_dac_a_c_6)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(32[16:25])
    defparam i11538_2_lut_2_lut.init = 16'h4444;
    LUT4 i1_2_lut_adj_160 (.A(n34), .B(wb_addr[9]), .Z(n20416)) /* synthesis lut_function=(A+!(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(241[23:49])
    defparam i1_2_lut_adj_160.init = 16'hbbbb;
    FD1S3AX wb_idata_i29 (.D(wb_idata_31__N_2[29]), .CK(dac_clk_p_c), .Q(wb_idata[29]));   // d:/documents/git_local/fm_modulator/rtl/top.v(265[9] 273[53])
    defparam wb_idata_i29.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_161 (.A(n26563), .B(n20416), .C(wb_addr[15]), .D(n20412), 
         .Z(n20422)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(241[23:49])
    defparam i1_4_lut_adj_161.init = 16'hffef;
    TSALL TSALL_INST (.TSALL(GND_net));
    FD1S3AX wb_smpl_data_i0 (.D(wb_smpl_data_31__N_64[0]), .CK(dac_clk_p_c), 
            .Q(wb_smpl_data[0]));   // d:/documents/git_local/fm_modulator/rtl/top.v(212[9] 220[10])
    defparam wb_smpl_data_i0.GSR = "DISABLED";
    clock_phase_shifter clock_phase_shifter_inst (.q_clk_p_c(q_clk_p_c), .i_clk_2f_N_2250(i_clk_2f_N_2250), 
            .q_clk_n_c(q_clk_n_c), .i_clk_p_c(i_clk_p_c), .lo_pll_out(lo_pll_out), 
            .i_clk_n_c(i_clk_n_c)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(158[21] 162[2])
    FD1S3AX wb_idata_i28 (.D(wb_idata_31__N_2[28]), .CK(dac_clk_p_c), .Q(wb_idata[28]));   // d:/documents/git_local/fm_modulator/rtl/top.v(265[9] 273[53])
    defparam wb_idata_i28.GSR = "DISABLED";
    CCU2D add_32_19 (.A0(power_counter[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17302), .COUT(n17303), .S0(power_counter_31__N_232[17]), 
          .S1(power_counter_31__N_232[18]));   // d:/documents/git_local/fm_modulator/rtl/top.v(227[21:41])
    defparam add_32_19.INIT0 = 16'h5aaa;
    defparam add_32_19.INIT1 = 16'h5aaa;
    defparam add_32_19.INJECT1_0 = "NO";
    defparam add_32_19.INJECT1_1 = "NO";
    CCU2D add_33_23 (.A0(power_counter[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17320), .COUT(n17321), .S0(power_counter_31__N_201[21]), 
          .S1(power_counter_31__N_201[22]));   // d:/documents/git_local/fm_modulator/rtl/top.v(229[27:53])
    defparam add_33_23.INIT0 = 16'h5aaa;
    defparam add_33_23.INIT1 = 16'h5aaa;
    defparam add_33_23.INJECT1_0 = "NO";
    defparam add_33_23.INJECT1_1 = "NO";
    CCU2D add_32_17 (.A0(power_counter[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17301), .COUT(n17302), .S0(power_counter_31__N_232[15]), 
          .S1(power_counter_31__N_232[16]));   // d:/documents/git_local/fm_modulator/rtl/top.v(227[21:41])
    defparam add_32_17.INIT0 = 16'h5aaa;
    defparam add_32_17.INIT1 = 16'h5aaa;
    defparam add_32_17.INJECT1_0 = "NO";
    defparam add_32_17.INJECT1_1 = "NO";
    FD1S3AX wb_idata_i27 (.D(wb_idata_31__N_2[27]), .CK(dac_clk_p_c), .Q(wb_idata[27]));   // d:/documents/git_local/fm_modulator/rtl/top.v(265[9] 273[53])
    defparam wb_idata_i27.GSR = "DISABLED";
    CCU2D add_33_21 (.A0(power_counter[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17319), .COUT(n17320), .S0(power_counter_31__N_201[19]), 
          .S1(power_counter_31__N_201[20]));   // d:/documents/git_local/fm_modulator/rtl/top.v(229[27:53])
    defparam add_33_21.INIT0 = 16'h5aaa;
    defparam add_33_21.INIT1 = 16'h5aaa;
    defparam add_33_21.INJECT1_0 = "NO";
    defparam add_33_21.INJECT1_1 = "NO";
    CCU2D add_32_15 (.A0(power_counter[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17300), .COUT(n17301), .S0(power_counter_31__N_232[13]), 
          .S1(power_counter_31__N_232[14]));   // d:/documents/git_local/fm_modulator/rtl/top.v(227[21:41])
    defparam add_32_15.INIT0 = 16'h5aaa;
    defparam add_32_15.INIT1 = 16'h5aaa;
    defparam add_32_15.INJECT1_0 = "NO";
    defparam add_32_15.INJECT1_1 = "NO";
    CCU2D add_33_19 (.A0(power_counter[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17318), .COUT(n17319), .S0(power_counter_31__N_201[17]), 
          .S1(power_counter_31__N_201[18]));   // d:/documents/git_local/fm_modulator/rtl/top.v(229[27:53])
    defparam add_33_19.INIT0 = 16'h5aaa;
    defparam add_33_19.INIT1 = 16'h5aaa;
    defparam add_33_19.INJECT1_0 = "NO";
    defparam add_33_19.INJECT1_1 = "NO";
    CCU2D add_32_5 (.A0(power_counter[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17295), .COUT(n17296), .S0(power_counter_31__N_232[3]), 
          .S1(power_counter_31__N_232[4]));   // d:/documents/git_local/fm_modulator/rtl/top.v(227[21:41])
    defparam add_32_5.INIT0 = 16'h5aaa;
    defparam add_32_5.INIT1 = 16'h5aaa;
    defparam add_32_5.INJECT1_0 = "NO";
    defparam add_32_5.INJECT1_1 = "NO";
    CCU2D add_33_17 (.A0(power_counter[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17317), .COUT(n17318), .S0(power_counter_31__N_201[15]), 
          .S1(power_counter_31__N_201[16]));   // d:/documents/git_local/fm_modulator/rtl/top.v(229[27:53])
    defparam add_33_17.INIT0 = 16'h5aaa;
    defparam add_33_17.INIT1 = 16'h5aaa;
    defparam add_33_17.INJECT1_0 = "NO";
    defparam add_33_17.INJECT1_1 = "NO";
    CCU2D add_33_15 (.A0(power_counter[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17316), .COUT(n17317), .S0(power_counter_31__N_201[13]), 
          .S1(power_counter_31__N_201[14]));   // d:/documents/git_local/fm_modulator/rtl/top.v(229[27:53])
    defparam add_33_15.INIT0 = 16'h5aaa;
    defparam add_33_15.INIT1 = 16'h5aaa;
    defparam add_33_15.INJECT1_0 = "NO";
    defparam add_33_15.INJECT1_1 = "NO";
    CCU2D add_33_13 (.A0(power_counter[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17315), .COUT(n17316), .S0(power_counter_31__N_201[11]), 
          .S1(power_counter_31__N_201[12]));   // d:/documents/git_local/fm_modulator/rtl/top.v(229[27:53])
    defparam add_33_13.INIT0 = 16'h5aaa;
    defparam add_33_13.INIT1 = 16'h5aaa;
    defparam add_33_13.INJECT1_0 = "NO";
    defparam add_33_13.INJECT1_1 = "NO";
    CCU2D add_33_11 (.A0(power_counter[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17314), .COUT(n17315), .S0(power_counter_31__N_201[9]), 
          .S1(power_counter_31__N_201[10]));   // d:/documents/git_local/fm_modulator/rtl/top.v(229[27:53])
    defparam add_33_11.INIT0 = 16'h5aaa;
    defparam add_33_11.INIT1 = 16'h5aaa;
    defparam add_33_11.INJECT1_0 = "NO";
    defparam add_33_11.INJECT1_1 = "NO";
    CCU2D add_32_9 (.A0(power_counter[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17297), .COUT(n17298), .S0(power_counter_31__N_232[7]), 
          .S1(power_counter_31__N_232[8]));   // d:/documents/git_local/fm_modulator/rtl/top.v(227[21:41])
    defparam add_32_9.INIT0 = 16'h5aaa;
    defparam add_32_9.INIT1 = 16'h5aaa;
    defparam add_32_9.INJECT1_0 = "NO";
    defparam add_32_9.INJECT1_1 = "NO";
    CCU2D add_33_9 (.A0(power_counter[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17313), .COUT(n17314), .S0(power_counter_31__N_201[7]), 
          .S1(power_counter_31__N_201[8]));   // d:/documents/git_local/fm_modulator/rtl/top.v(229[27:53])
    defparam add_33_9.INIT0 = 16'h5aaa;
    defparam add_33_9.INIT1 = 16'h5aaa;
    defparam add_33_9.INJECT1_0 = "NO";
    defparam add_33_9.INJECT1_1 = "NO";
    OB o_dac_a_pad_6 (.I(o_dac_a_c_6), .O(o_dac_a[6]));   // d:/documents/git_local/fm_modulator/rtl/top.v(28[38:45])
    FD1S3AX wb_idata_i26 (.D(wb_idata_31__N_2[26]), .CK(dac_clk_p_c), .Q(wb_idata[26]));   // d:/documents/git_local/fm_modulator/rtl/top.v(265[9] 273[53])
    defparam wb_idata_i26.GSR = "DISABLED";
    FD1S3AX wb_idata_i25 (.D(wb_idata_31__N_2[25]), .CK(dac_clk_p_c), .Q(wb_idata[25]));   // d:/documents/git_local/fm_modulator/rtl/top.v(265[9] 273[53])
    defparam wb_idata_i25.GSR = "DISABLED";
    FD1S3AX wb_idata_i24 (.D(wb_idata_31__N_2[24]), .CK(dac_clk_p_c), .Q(wb_idata[24]));   // d:/documents/git_local/fm_modulator/rtl/top.v(265[9] 273[53])
    defparam wb_idata_i24.GSR = "DISABLED";
    FD1S3AX wb_idata_i23 (.D(wb_idata_31__N_2[23]), .CK(dac_clk_p_c), .Q(wb_idata[23]));   // d:/documents/git_local/fm_modulator/rtl/top.v(265[9] 273[53])
    defparam wb_idata_i23.GSR = "DISABLED";
    FD1S3AX wb_idata_i22 (.D(wb_idata_31__N_2[22]), .CK(dac_clk_p_c), .Q(wb_idata[22]));   // d:/documents/git_local/fm_modulator/rtl/top.v(265[9] 273[53])
    defparam wb_idata_i22.GSR = "DISABLED";
    FD1S3AX wb_idata_i21 (.D(wb_idata_31__N_2[21]), .CK(dac_clk_p_c), .Q(wb_idata[21]));   // d:/documents/git_local/fm_modulator/rtl/top.v(265[9] 273[53])
    defparam wb_idata_i21.GSR = "DISABLED";
    FD1S3AX wb_idata_i20 (.D(wb_idata_31__N_2[20]), .CK(dac_clk_p_c), .Q(wb_idata[20]));   // d:/documents/git_local/fm_modulator/rtl/top.v(265[9] 273[53])
    defparam wb_idata_i20.GSR = "DISABLED";
    FD1S3AX wb_idata_i19 (.D(wb_idata_31__N_2[19]), .CK(dac_clk_p_c), .Q(wb_idata[19]));   // d:/documents/git_local/fm_modulator/rtl/top.v(265[9] 273[53])
    defparam wb_idata_i19.GSR = "DISABLED";
    FD1S3AX wb_idata_i18 (.D(wb_idata_31__N_2[18]), .CK(dac_clk_p_c), .Q(wb_idata[18]));   // d:/documents/git_local/fm_modulator/rtl/top.v(265[9] 273[53])
    defparam wb_idata_i18.GSR = "DISABLED";
    FD1S3AX wb_idata_i17 (.D(wb_idata_31__N_2[17]), .CK(dac_clk_p_c), .Q(wb_idata[17]));   // d:/documents/git_local/fm_modulator/rtl/top.v(265[9] 273[53])
    defparam wb_idata_i17.GSR = "DISABLED";
    FD1S3AX wb_idata_i16 (.D(wb_idata_31__N_2[16]), .CK(dac_clk_p_c), .Q(wb_idata[16]));   // d:/documents/git_local/fm_modulator/rtl/top.v(265[9] 273[53])
    defparam wb_idata_i16.GSR = "DISABLED";
    FD1S3AX wb_idata_i15 (.D(wb_idata_31__N_2[15]), .CK(dac_clk_p_c), .Q(wb_idata[15]));   // d:/documents/git_local/fm_modulator/rtl/top.v(265[9] 273[53])
    defparam wb_idata_i15.GSR = "DISABLED";
    FD1S3AX wb_idata_i14 (.D(wb_idata_31__N_2[14]), .CK(dac_clk_p_c), .Q(wb_idata[14]));   // d:/documents/git_local/fm_modulator/rtl/top.v(265[9] 273[53])
    defparam wb_idata_i14.GSR = "DISABLED";
    FD1S3AX wb_idata_i13 (.D(wb_idata_31__N_2[13]), .CK(dac_clk_p_c), .Q(wb_idata[13]));   // d:/documents/git_local/fm_modulator/rtl/top.v(265[9] 273[53])
    defparam wb_idata_i13.GSR = "DISABLED";
    FD1S3AX wb_idata_i12 (.D(wb_idata_31__N_2[12]), .CK(dac_clk_p_c), .Q(wb_idata[12]));   // d:/documents/git_local/fm_modulator/rtl/top.v(265[9] 273[53])
    defparam wb_idata_i12.GSR = "DISABLED";
    FD1S3AX wb_idata_i11 (.D(wb_idata_31__N_2[11]), .CK(dac_clk_p_c), .Q(wb_idata[11]));   // d:/documents/git_local/fm_modulator/rtl/top.v(265[9] 273[53])
    defparam wb_idata_i11.GSR = "DISABLED";
    FD1S3AX wb_idata_i10 (.D(wb_idata_31__N_2[10]), .CK(dac_clk_p_c), .Q(wb_idata[10]));   // d:/documents/git_local/fm_modulator/rtl/top.v(265[9] 273[53])
    defparam wb_idata_i10.GSR = "DISABLED";
    FD1S3AX wb_idata_i9 (.D(wb_idata_31__N_2[9]), .CK(dac_clk_p_c), .Q(wb_idata[9]));   // d:/documents/git_local/fm_modulator/rtl/top.v(265[9] 273[53])
    defparam wb_idata_i9.GSR = "DISABLED";
    FD1S3AX wb_idata_i8 (.D(wb_idata_31__N_2[8]), .CK(dac_clk_p_c), .Q(wb_idata[8]));   // d:/documents/git_local/fm_modulator/rtl/top.v(265[9] 273[53])
    defparam wb_idata_i8.GSR = "DISABLED";
    FD1S3AX wb_idata_i7 (.D(wb_idata_31__N_2[7]), .CK(dac_clk_p_c), .Q(wb_idata[7]));   // d:/documents/git_local/fm_modulator/rtl/top.v(265[9] 273[53])
    defparam wb_idata_i7.GSR = "DISABLED";
    FD1S3AX wb_idata_i6 (.D(wb_idata_31__N_2[6]), .CK(dac_clk_p_c), .Q(wb_idata[6]));   // d:/documents/git_local/fm_modulator/rtl/top.v(265[9] 273[53])
    defparam wb_idata_i6.GSR = "DISABLED";
    FD1S3AX wb_idata_i5 (.D(wb_idata_31__N_2[5]), .CK(dac_clk_p_c), .Q(wb_idata[5]));   // d:/documents/git_local/fm_modulator/rtl/top.v(265[9] 273[53])
    defparam wb_idata_i5.GSR = "DISABLED";
    FD1S3AX wb_idata_i4 (.D(wb_idata_31__N_2[4]), .CK(dac_clk_p_c), .Q(wb_idata[4]));   // d:/documents/git_local/fm_modulator/rtl/top.v(265[9] 273[53])
    defparam wb_idata_i4.GSR = "DISABLED";
    FD1S3AX wb_idata_i3 (.D(wb_idata_31__N_2[3]), .CK(dac_clk_p_c), .Q(wb_idata[3]));   // d:/documents/git_local/fm_modulator/rtl/top.v(265[9] 273[53])
    defparam wb_idata_i3.GSR = "DISABLED";
    FD1S3AX wb_idata_i2 (.D(wb_idata_31__N_2[2]), .CK(dac_clk_p_c), .Q(wb_idata[2]));   // d:/documents/git_local/fm_modulator/rtl/top.v(265[9] 273[53])
    defparam wb_idata_i2.GSR = "DISABLED";
    FD1S3AX wb_idata_i1 (.D(wb_idata_31__N_2[1]), .CK(dac_clk_p_c), .Q(wb_idata[1]));   // d:/documents/git_local/fm_modulator/rtl/top.v(265[9] 273[53])
    defparam wb_idata_i1.GSR = "DISABLED";
    CCU2D add_33_7 (.A0(power_counter[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17312), .COUT(n17313), .S0(power_counter_31__N_201[5]), 
          .S1(power_counter_31__N_201[6]));   // d:/documents/git_local/fm_modulator/rtl/top.v(229[27:53])
    defparam add_33_7.INIT0 = 16'h5aaa;
    defparam add_33_7.INIT1 = 16'h5aaa;
    defparam add_33_7.INJECT1_0 = "NO";
    defparam add_33_7.INJECT1_1 = "NO";
    CCU2D add_32_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(power_counter[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n17294), .S1(power_counter_31__N_232[0]));   // d:/documents/git_local/fm_modulator/rtl/top.v(227[21:41])
    defparam add_32_1.INIT0 = 16'hF000;
    defparam add_32_1.INIT1 = 16'h5555;
    defparam add_32_1.INJECT1_0 = "NO";
    defparam add_32_1.INJECT1_1 = "NO";
    CCU2D add_33_5 (.A0(power_counter[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17311), .COUT(n17312), .S0(power_counter_31__N_201[3]), 
          .S1(power_counter_31__N_201[4]));   // d:/documents/git_local/fm_modulator/rtl/top.v(229[27:53])
    defparam add_33_5.INIT0 = 16'h5aaa;
    defparam add_33_5.INIT1 = 16'h5aaa;
    defparam add_33_5.INJECT1_0 = "NO";
    defparam add_33_5.INJECT1_1 = "NO";
    CCU2D add_33_3 (.A0(power_counter[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17310), .COUT(n17311), .S0(power_counter_31__N_201[1]), 
          .S1(power_counter_31__N_201[2]));   // d:/documents/git_local/fm_modulator/rtl/top.v(229[27:53])
    defparam add_33_3.INIT0 = 16'h5aaa;
    defparam add_33_3.INIT1 = 16'h5aaa;
    defparam add_33_3.INJECT1_0 = "NO";
    defparam add_33_3.INJECT1_1 = "NO";
    CCU2D add_32_3 (.A0(power_counter[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17294), .COUT(n17295), .S0(power_counter_31__N_232[1]), 
          .S1(power_counter_31__N_232[2]));   // d:/documents/git_local/fm_modulator/rtl/top.v(227[21:41])
    defparam add_32_3.INIT0 = 16'h5aaa;
    defparam add_32_3.INIT1 = 16'h5aaa;
    defparam add_32_3.INJECT1_0 = "NO";
    defparam add_32_3.INJECT1_1 = "NO";
    CCU2D add_33_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(power_counter[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n17310), .S1(power_counter_31__N_201[0]));   // d:/documents/git_local/fm_modulator/rtl/top.v(229[27:53])
    defparam add_33_1.INIT0 = 16'hF000;
    defparam add_33_1.INIT1 = 16'h5555;
    defparam add_33_1.INJECT1_0 = "NO";
    defparam add_33_1.INJECT1_1 = "NO";
    CCU2D add_32_13 (.A0(power_counter[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17299), .COUT(n17300), .S0(power_counter_31__N_232[11]), 
          .S1(power_counter_31__N_232[12]));   // d:/documents/git_local/fm_modulator/rtl/top.v(227[21:41])
    defparam add_32_13.INIT0 = 16'h5aaa;
    defparam add_32_13.INIT1 = 16'h5aaa;
    defparam add_32_13.INJECT1_0 = "NO";
    defparam add_32_13.INJECT1_1 = "NO";
    CCU2D add_32_33 (.A0(power_counter[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n17309), .S0(power_counter_31__N_232[31]));   // d:/documents/git_local/fm_modulator/rtl/top.v(227[21:41])
    defparam add_32_33.INIT0 = 16'h5aaa;
    defparam add_32_33.INIT1 = 16'h0000;
    defparam add_32_33.INJECT1_0 = "NO";
    defparam add_32_33.INJECT1_1 = "NO";
    CCU2D add_32_7 (.A0(power_counter[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17296), .COUT(n17297), .S0(power_counter_31__N_232[5]), 
          .S1(power_counter_31__N_232[6]));   // d:/documents/git_local/fm_modulator/rtl/top.v(227[21:41])
    defparam add_32_7.INIT0 = 16'h5aaa;
    defparam add_32_7.INIT1 = 16'h5aaa;
    defparam add_32_7.INJECT1_0 = "NO";
    defparam add_32_7.INJECT1_1 = "NO";
    CCU2D add_32_31 (.A0(power_counter[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17308), .COUT(n17309), .S0(power_counter_31__N_232[29]), 
          .S1(power_counter_31__N_232[30]));   // d:/documents/git_local/fm_modulator/rtl/top.v(227[21:41])
    defparam add_32_31.INIT0 = 16'h5aaa;
    defparam add_32_31.INIT1 = 16'h5aaa;
    defparam add_32_31.INJECT1_0 = "NO";
    defparam add_32_31.INJECT1_1 = "NO";
    CCU2D add_32_11 (.A0(power_counter[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17298), .COUT(n17299), .S0(power_counter_31__N_232[9]), 
          .S1(power_counter_31__N_232[10]));   // d:/documents/git_local/fm_modulator/rtl/top.v(227[21:41])
    defparam add_32_11.INIT0 = 16'h5aaa;
    defparam add_32_11.INIT1 = 16'h5aaa;
    defparam add_32_11.INJECT1_0 = "NO";
    defparam add_32_11.INJECT1_1 = "NO";
    CCU2D add_32_29 (.A0(power_counter[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17307), .COUT(n17308), .S0(power_counter_31__N_232[27]), 
          .S1(power_counter_31__N_232[28]));   // d:/documents/git_local/fm_modulator/rtl/top.v(227[21:41])
    defparam add_32_29.INIT0 = 16'h5aaa;
    defparam add_32_29.INIT1 = 16'h5aaa;
    defparam add_32_29.INJECT1_0 = "NO";
    defparam add_32_29.INJECT1_1 = "NO";
    FD1P3AX power_counter_i31 (.D(n29210), .SP(power_counter_31__N_232[31]), 
            .CK(dac_clk_p_c), .Q(power_counter[31])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(224[9] 229[54])
    defparam power_counter_i31.GSR = "DISABLED";
    sys_clk sys_clk_inst (.i_ref_clk_c(i_ref_clk_c), .dac_clk_p_c(dac_clk_p_c), 
            .GND_net(GND_net)) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(38[10:54])
    FD1S3AX power_counter_i30 (.D(power_counter_31__N_129[30]), .CK(dac_clk_p_c), 
            .Q(power_counter[30])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(224[9] 229[54])
    defparam power_counter_i30.GSR = "DISABLED";
    FD1S3AX power_counter_i29 (.D(power_counter_31__N_129[29]), .CK(dac_clk_p_c), 
            .Q(power_counter[29])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(224[9] 229[54])
    defparam power_counter_i29.GSR = "DISABLED";
    LUT4 m1_lut (.Z(n29210)) /* synthesis lut_function=1, syn_instantiated=1 */ ;
    defparam m1_lut.init = 16'hffff;
    FD1S3AX power_counter_i28 (.D(power_counter_31__N_129[28]), .CK(dac_clk_p_c), 
            .Q(power_counter[28])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(224[9] 229[54])
    defparam power_counter_i28.GSR = "DISABLED";
    FD1S3AX power_counter_i27 (.D(power_counter_31__N_129[27]), .CK(dac_clk_p_c), 
            .Q(power_counter[27])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(224[9] 229[54])
    defparam power_counter_i27.GSR = "DISABLED";
    FD1S3AX power_counter_i26 (.D(power_counter_31__N_129[26]), .CK(dac_clk_p_c), 
            .Q(power_counter[26])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(224[9] 229[54])
    defparam power_counter_i26.GSR = "DISABLED";
    FD1S3AX power_counter_i25 (.D(power_counter_31__N_129[25]), .CK(dac_clk_p_c), 
            .Q(power_counter[25])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(224[9] 229[54])
    defparam power_counter_i25.GSR = "DISABLED";
    FD1S3AX power_counter_i24 (.D(power_counter_31__N_129[24]), .CK(dac_clk_p_c), 
            .Q(power_counter[24])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(224[9] 229[54])
    defparam power_counter_i24.GSR = "DISABLED";
    FD1S3AX power_counter_i23 (.D(power_counter_31__N_129[23]), .CK(dac_clk_p_c), 
            .Q(power_counter[23])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(224[9] 229[54])
    defparam power_counter_i23.GSR = "DISABLED";
    FD1S3AX power_counter_i22 (.D(power_counter_31__N_129[22]), .CK(dac_clk_p_c), 
            .Q(power_counter[22])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(224[9] 229[54])
    defparam power_counter_i22.GSR = "DISABLED";
    FD1S3AX power_counter_i21 (.D(power_counter_31__N_129[21]), .CK(dac_clk_p_c), 
            .Q(power_counter[21])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(224[9] 229[54])
    defparam power_counter_i21.GSR = "DISABLED";
    FD1S3AX power_counter_i20 (.D(power_counter_31__N_129[20]), .CK(dac_clk_p_c), 
            .Q(power_counter[20])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(224[9] 229[54])
    defparam power_counter_i20.GSR = "DISABLED";
    FD1S3AX power_counter_i19 (.D(power_counter_31__N_129[19]), .CK(dac_clk_p_c), 
            .Q(power_counter[19])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(224[9] 229[54])
    defparam power_counter_i19.GSR = "DISABLED";
    FD1S3AX power_counter_i18 (.D(power_counter_31__N_129[18]), .CK(dac_clk_p_c), 
            .Q(power_counter[18])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(224[9] 229[54])
    defparam power_counter_i18.GSR = "DISABLED";
    FD1S3AX power_counter_i17 (.D(power_counter_31__N_129[17]), .CK(dac_clk_p_c), 
            .Q(power_counter[17])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(224[9] 229[54])
    defparam power_counter_i17.GSR = "DISABLED";
    FD1S3AX power_counter_i16 (.D(power_counter_31__N_129[16]), .CK(dac_clk_p_c), 
            .Q(power_counter[16])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(224[9] 229[54])
    defparam power_counter_i16.GSR = "DISABLED";
    FD1S3AX power_counter_i15 (.D(power_counter_31__N_129[15]), .CK(dac_clk_p_c), 
            .Q(power_counter[15])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(224[9] 229[54])
    defparam power_counter_i15.GSR = "DISABLED";
    FD1S3AX power_counter_i14 (.D(power_counter_31__N_129[14]), .CK(dac_clk_p_c), 
            .Q(power_counter[14])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(224[9] 229[54])
    defparam power_counter_i14.GSR = "DISABLED";
    FD1S3AX power_counter_i13 (.D(power_counter_31__N_129[13]), .CK(dac_clk_p_c), 
            .Q(power_counter[13])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(224[9] 229[54])
    defparam power_counter_i13.GSR = "DISABLED";
    FD1S3AX power_counter_i12 (.D(power_counter_31__N_129[12]), .CK(dac_clk_p_c), 
            .Q(power_counter[12])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(224[9] 229[54])
    defparam power_counter_i12.GSR = "DISABLED";
    FD1S3AX power_counter_i11 (.D(power_counter_31__N_129[11]), .CK(dac_clk_p_c), 
            .Q(power_counter[11])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(224[9] 229[54])
    defparam power_counter_i11.GSR = "DISABLED";
    FD1S3AX power_counter_i10 (.D(power_counter_31__N_129[10]), .CK(dac_clk_p_c), 
            .Q(power_counter[10])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(224[9] 229[54])
    defparam power_counter_i10.GSR = "DISABLED";
    FD1S3AX power_counter_i9 (.D(power_counter_31__N_129[9]), .CK(dac_clk_p_c), 
            .Q(power_counter[9])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(224[9] 229[54])
    defparam power_counter_i9.GSR = "DISABLED";
    FD1S3AX power_counter_i8 (.D(power_counter_31__N_129[8]), .CK(dac_clk_p_c), 
            .Q(power_counter[8])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(224[9] 229[54])
    defparam power_counter_i8.GSR = "DISABLED";
    FD1S3AX power_counter_i7 (.D(power_counter_31__N_129[7]), .CK(dac_clk_p_c), 
            .Q(power_counter[7])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(224[9] 229[54])
    defparam power_counter_i7.GSR = "DISABLED";
    FD1S3AX power_counter_i6 (.D(power_counter_31__N_129[6]), .CK(dac_clk_p_c), 
            .Q(power_counter[6])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(224[9] 229[54])
    defparam power_counter_i6.GSR = "DISABLED";
    FD1S3AX power_counter_i5 (.D(power_counter_31__N_129[5]), .CK(dac_clk_p_c), 
            .Q(power_counter[5])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(224[9] 229[54])
    defparam power_counter_i5.GSR = "DISABLED";
    FD1S3AX power_counter_i4 (.D(power_counter_31__N_129[4]), .CK(dac_clk_p_c), 
            .Q(power_counter[4])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(224[9] 229[54])
    defparam power_counter_i4.GSR = "DISABLED";
    FD1S3AX power_counter_i3 (.D(power_counter_31__N_129[3]), .CK(dac_clk_p_c), 
            .Q(power_counter[3])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(224[9] 229[54])
    defparam power_counter_i3.GSR = "DISABLED";
    FD1S3AX power_counter_i2 (.D(power_counter_31__N_129[2]), .CK(dac_clk_p_c), 
            .Q(power_counter[2])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(224[9] 229[54])
    defparam power_counter_i2.GSR = "DISABLED";
    FD1S3AX power_counter_i1 (.D(power_counter_31__N_129[1]), .CK(dac_clk_p_c), 
            .Q(power_counter[1])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(224[9] 229[54])
    defparam power_counter_i1.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i31 (.D(n2005), .CK(dac_clk_p_c), .CD(n9365), 
            .Q(wb_smpl_data[31]));   // d:/documents/git_local/fm_modulator/rtl/top.v(212[9] 220[10])
    defparam wb_smpl_data_i31.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i29 (.D(wb_addr[29]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[29])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(255[9] 257[31])
    defparam bus_err_address_i0_i29.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i28 (.D(wb_addr[28]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[28])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(255[9] 257[31])
    defparam bus_err_address_i0_i28.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i27 (.D(wb_addr[27]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[27])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(255[9] 257[31])
    defparam bus_err_address_i0_i27.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i26 (.D(wb_addr[26]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[26])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(255[9] 257[31])
    defparam bus_err_address_i0_i26.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i25 (.D(wb_addr[25]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[25])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(255[9] 257[31])
    defparam bus_err_address_i0_i25.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i24 (.D(wb_addr[24]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[24])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(255[9] 257[31])
    defparam bus_err_address_i0_i24.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i23 (.D(wb_addr[23]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[23])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(255[9] 257[31])
    defparam bus_err_address_i0_i23.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i22 (.D(wb_addr[22]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[22])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(255[9] 257[31])
    defparam bus_err_address_i0_i22.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i21 (.D(wb_addr[21]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[21])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(255[9] 257[31])
    defparam bus_err_address_i0_i21.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i20 (.D(wb_addr[20]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[20])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(255[9] 257[31])
    defparam bus_err_address_i0_i20.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i19 (.D(wb_addr[19]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[19])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(255[9] 257[31])
    defparam bus_err_address_i0_i19.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i18 (.D(wb_addr[18]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[18])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(255[9] 257[31])
    defparam bus_err_address_i0_i18.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i17 (.D(wb_addr[17]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[17])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(255[9] 257[31])
    defparam bus_err_address_i0_i17.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i16 (.D(wb_addr[16]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[16])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(255[9] 257[31])
    defparam bus_err_address_i0_i16.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i15 (.D(wb_addr[15]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[15])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(255[9] 257[31])
    defparam bus_err_address_i0_i15.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i14 (.D(wb_addr[14]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[14])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(255[9] 257[31])
    defparam bus_err_address_i0_i14.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i13 (.D(wb_addr[13]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[13])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(255[9] 257[31])
    defparam bus_err_address_i0_i13.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i12 (.D(wb_addr[12]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[12])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(255[9] 257[31])
    defparam bus_err_address_i0_i12.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i11 (.D(wb_addr[11]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[11])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(255[9] 257[31])
    defparam bus_err_address_i0_i11.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i10 (.D(wb_addr[10]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[10])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(255[9] 257[31])
    defparam bus_err_address_i0_i10.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i9 (.D(wb_addr[9]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[9])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(255[9] 257[31])
    defparam bus_err_address_i0_i9.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i8 (.D(wb_addr[8]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[8])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(255[9] 257[31])
    defparam bus_err_address_i0_i8.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i7 (.D(wb_addr[7]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[7])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(255[9] 257[31])
    defparam bus_err_address_i0_i7.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i6 (.D(wb_addr[6]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[6])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(255[9] 257[31])
    defparam bus_err_address_i0_i6.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i5 (.D(wb_addr[5]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[5])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(255[9] 257[31])
    defparam bus_err_address_i0_i5.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i4 (.D(wb_addr[4]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[4])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(255[9] 257[31])
    defparam bus_err_address_i0_i4.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i3 (.D(wb_addr[3]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[3])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(255[9] 257[31])
    defparam bus_err_address_i0_i3.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i2 (.D(wb_addr[2]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[2])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(255[9] 257[31])
    defparam bus_err_address_i0_i2.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i1 (.D(wb_addr[1]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[1])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(255[9] 257[31])
    defparam bus_err_address_i0_i1.GSR = "DISABLED";
    LUT4 m0_lut (.Z(n29209)) /* synthesis lut_function=0, syn_instantiated=1 */ ;
    defparam m0_lut.init = 16'h0000;
    FD1S3IX wb_smpl_data_i30 (.D(n2006), .CK(dac_clk_p_c), .CD(n9365), 
            .Q(wb_smpl_data[30]));   // d:/documents/git_local/fm_modulator/rtl/top.v(212[9] 220[10])
    defparam wb_smpl_data_i30.GSR = "DISABLED";
    OB o_dac_a_pad_5 (.I(o_dac_a_c_5), .O(o_dac_a[5]));   // d:/documents/git_local/fm_modulator/rtl/top.v(28[38:45])
    OB o_dac_a_pad_4 (.I(o_dac_a_c_4), .O(o_dac_a[4]));   // d:/documents/git_local/fm_modulator/rtl/top.v(28[38:45])
    OB o_dac_a_pad_3 (.I(o_dac_a_c_3), .O(o_dac_a[3]));   // d:/documents/git_local/fm_modulator/rtl/top.v(28[38:45])
    OB o_dac_a_pad_2 (.I(o_dac_a_c_2), .O(o_dac_a[2]));   // d:/documents/git_local/fm_modulator/rtl/top.v(28[38:45])
    OB o_dac_a_pad_1 (.I(o_dac_a_c_1), .O(o_dac_a[1]));   // d:/documents/git_local/fm_modulator/rtl/top.v(28[38:45])
    OB o_dac_a_pad_0 (.I(o_dac_a_c_0), .O(o_dac_a[0]));   // d:/documents/git_local/fm_modulator/rtl/top.v(28[38:45])
    OB o_dac_b_pad_9 (.I(o_dac_b_c_9), .O(o_dac_b[9]));   // d:/documents/git_local/fm_modulator/rtl/top.v(28[47:54])
    OB o_dac_b_pad_8 (.I(o_dac_b_c_15), .O(o_dac_b[8]));   // d:/documents/git_local/fm_modulator/rtl/top.v(28[47:54])
    OB o_dac_b_pad_7 (.I(o_dac_b_c_14), .O(o_dac_b[7]));   // d:/documents/git_local/fm_modulator/rtl/top.v(28[47:54])
    OB o_dac_b_pad_6 (.I(o_dac_b_c_13), .O(o_dac_b[6]));   // d:/documents/git_local/fm_modulator/rtl/top.v(28[47:54])
    OB o_dac_b_pad_5 (.I(o_dac_b_c_12), .O(o_dac_b[5]));   // d:/documents/git_local/fm_modulator/rtl/top.v(28[47:54])
    OB o_dac_b_pad_4 (.I(o_dac_b_c_11), .O(o_dac_b[4]));   // d:/documents/git_local/fm_modulator/rtl/top.v(28[47:54])
    OB o_dac_b_pad_3 (.I(o_dac_b_c_10), .O(o_dac_b[3]));   // d:/documents/git_local/fm_modulator/rtl/top.v(28[47:54])
    OB o_dac_b_pad_2 (.I(n3537), .O(o_dac_b[2]));   // d:/documents/git_local/fm_modulator/rtl/top.v(28[47:54])
    OB o_dac_b_pad_1 (.I(o_dac_b_c_8), .O(o_dac_b[1]));   // d:/documents/git_local/fm_modulator/rtl/top.v(28[47:54])
    OB o_dac_b_pad_0 (.I(o_dac_b_c_7), .O(o_dac_b[0]));   // d:/documents/git_local/fm_modulator/rtl/top.v(28[47:54])
    OB dac_clk_p_pad (.I(dac_clk_p_c), .O(dac_clk_p));   // d:/documents/git_local/fm_modulator/rtl/top.v(29[49:58])
    OB dac_clk_n_pad (.I(dac_clk_n_c), .O(dac_clk_n));   // d:/documents/git_local/fm_modulator/rtl/top.v(29[60:69])
    OB o_dac_cw_b_pad (.I(o_dac_cw_b_c_c), .O(o_dac_cw_b));   // d:/documents/git_local/fm_modulator/rtl/top.v(29[71:81])
    OB i_clk_p_pad (.I(i_clk_p_c), .O(i_clk_p));   // d:/documents/git_local/fm_modulator/rtl/top.v(29[13:20])
    OB i_clk_n_pad (.I(i_clk_n_c), .O(i_clk_n));   // d:/documents/git_local/fm_modulator/rtl/top.v(29[22:29])
    OB q_clk_p_pad (.I(q_clk_p_c), .O(q_clk_p));   // d:/documents/git_local/fm_modulator/rtl/top.v(29[31:38])
    OB q_clk_n_pad (.I(q_clk_n_c), .O(q_clk_n));   // d:/documents/git_local/fm_modulator/rtl/top.v(29[40:47])
    IB i_ref_clk_pad (.I(i_ref_clk), .O(i_ref_clk_c));   // d:/documents/git_local/fm_modulator/rtl/top.v(23[12:21])
    IB o_dac_cw_b_c_pad (.I(i_resetb), .O(o_dac_cw_b_c_c));   // d:/documents/git_local/fm_modulator/rtl/top.v(23[23:31])
    IB i_wbu_uart_rx_pad (.I(i_wbu_uart_rx), .O(i_wbu_uart_rx_c));   // d:/documents/git_local/fm_modulator/rtl/top.v(25[12:25])
    FD1S3IX wb_smpl_data_i11 (.D(n2025), .CK(dac_clk_p_c), .CD(n9365), 
            .Q(wb_smpl_data[11]));   // d:/documents/git_local/fm_modulator/rtl/top.v(212[9] 220[10])
    defparam wb_smpl_data_i11.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i29 (.D(n26339), .CK(dac_clk_p_c), .CD(n9365), 
            .Q(wb_smpl_data[29]));   // d:/documents/git_local/fm_modulator/rtl/top.v(212[9] 220[10])
    defparam wb_smpl_data_i29.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i10 (.D(n26342), .CK(dac_clk_p_c), .CD(n9365), 
            .Q(wb_smpl_data[10]));   // d:/documents/git_local/fm_modulator/rtl/top.v(212[9] 220[10])
    defparam wb_smpl_data_i10.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i28 (.D(n2008), .CK(dac_clk_p_c), .CD(n9365), 
            .Q(wb_smpl_data[28]));   // d:/documents/git_local/fm_modulator/rtl/top.v(212[9] 220[10])
    defparam wb_smpl_data_i28.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i9 (.D(n26341), .CK(dac_clk_p_c), .CD(n9365), 
            .Q(wb_smpl_data[9]));   // d:/documents/git_local/fm_modulator/rtl/top.v(212[9] 220[10])
    defparam wb_smpl_data_i9.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i27 (.D(n2009), .CK(dac_clk_p_c), .CD(n9365), 
            .Q(wb_smpl_data[27]));   // d:/documents/git_local/fm_modulator/rtl/top.v(212[9] 220[10])
    defparam wb_smpl_data_i27.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i8 (.D(n2028), .CK(dac_clk_p_c), .CD(n9365), 
            .Q(wb_smpl_data[8]));   // d:/documents/git_local/fm_modulator/rtl/top.v(212[9] 220[10])
    defparam wb_smpl_data_i8.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i26 (.D(n2010), .CK(dac_clk_p_c), .CD(n9365), 
            .Q(wb_smpl_data[26]));   // d:/documents/git_local/fm_modulator/rtl/top.v(212[9] 220[10])
    defparam wb_smpl_data_i26.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i7 (.D(n2029), .CK(dac_clk_p_c), .CD(n9365), 
            .Q(wb_smpl_data[7]));   // d:/documents/git_local/fm_modulator/rtl/top.v(212[9] 220[10])
    defparam wb_smpl_data_i7.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i25 (.D(n2011), .CK(dac_clk_p_c), .CD(n9365), 
            .Q(wb_smpl_data[25]));   // d:/documents/git_local/fm_modulator/rtl/top.v(212[9] 220[10])
    defparam wb_smpl_data_i25.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i6 (.D(n2030), .CK(dac_clk_p_c), .CD(n9365), 
            .Q(wb_smpl_data[6]));   // d:/documents/git_local/fm_modulator/rtl/top.v(212[9] 220[10])
    defparam wb_smpl_data_i6.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i24 (.D(n2012), .CK(dac_clk_p_c), .CD(n9365), 
            .Q(wb_smpl_data[24]));   // d:/documents/git_local/fm_modulator/rtl/top.v(212[9] 220[10])
    defparam wb_smpl_data_i24.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i5 (.D(n26336), .CK(dac_clk_p_c), .CD(n9365), 
            .Q(wb_smpl_data[5]));   // d:/documents/git_local/fm_modulator/rtl/top.v(212[9] 220[10])
    defparam wb_smpl_data_i5.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i23 (.D(n2013), .CK(dac_clk_p_c), .CD(n9365), 
            .Q(wb_smpl_data[23]));   // d:/documents/git_local/fm_modulator/rtl/top.v(212[9] 220[10])
    defparam wb_smpl_data_i23.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i4 (.D(n2032), .CK(dac_clk_p_c), .CD(n9365), 
            .Q(wb_smpl_data[4]));   // d:/documents/git_local/fm_modulator/rtl/top.v(212[9] 220[10])
    defparam wb_smpl_data_i4.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i22 (.D(n2014), .CK(dac_clk_p_c), .CD(n9365), 
            .Q(wb_smpl_data[22]));   // d:/documents/git_local/fm_modulator/rtl/top.v(212[9] 220[10])
    defparam wb_smpl_data_i22.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i3 (.D(n2033), .CK(dac_clk_p_c), .CD(n9365), 
            .Q(wb_smpl_data[3]));   // d:/documents/git_local/fm_modulator/rtl/top.v(212[9] 220[10])
    defparam wb_smpl_data_i3.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i21 (.D(n2015), .CK(dac_clk_p_c), .CD(n9365), 
            .Q(wb_smpl_data[21]));   // d:/documents/git_local/fm_modulator/rtl/top.v(212[9] 220[10])
    defparam wb_smpl_data_i21.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i2 (.D(n2034), .CK(dac_clk_p_c), .CD(n9365), 
            .Q(wb_smpl_data[2]));   // d:/documents/git_local/fm_modulator/rtl/top.v(212[9] 220[10])
    defparam wb_smpl_data_i2.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i20 (.D(n26337), .CK(dac_clk_p_c), .CD(n9365), 
            .Q(wb_smpl_data[20]));   // d:/documents/git_local/fm_modulator/rtl/top.v(212[9] 220[10])
    defparam wb_smpl_data_i20.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i1 (.D(n2035), .CK(dac_clk_p_c), .CD(n9365), 
            .Q(wb_smpl_data[1]));   // d:/documents/git_local/fm_modulator/rtl/top.v(212[9] 220[10])
    defparam wb_smpl_data_i1.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i19 (.D(n2017), .CK(dac_clk_p_c), .CD(n9365), 
            .Q(wb_smpl_data[19]));   // d:/documents/git_local/fm_modulator/rtl/top.v(212[9] 220[10])
    defparam wb_smpl_data_i19.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i18 (.D(n26333), .CK(dac_clk_p_c), .CD(n9365), 
            .Q(wb_smpl_data[18]));   // d:/documents/git_local/fm_modulator/rtl/top.v(212[9] 220[10])
    defparam wb_smpl_data_i18.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i17 (.D(n26332), .CK(dac_clk_p_c), .CD(n9365), 
            .Q(wb_smpl_data[17]));   // d:/documents/git_local/fm_modulator/rtl/top.v(212[9] 220[10])
    defparam wb_smpl_data_i17.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i16 (.D(n26331), .CK(dac_clk_p_c), .CD(n9365), 
            .Q(wb_smpl_data[16]));   // d:/documents/git_local/fm_modulator/rtl/top.v(212[9] 220[10])
    defparam wb_smpl_data_i16.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i15 (.D(n2021), .CK(dac_clk_p_c), .CD(n9365), 
            .Q(wb_smpl_data[15]));   // d:/documents/git_local/fm_modulator/rtl/top.v(212[9] 220[10])
    defparam wb_smpl_data_i15.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i14 (.D(n2022), .CK(dac_clk_p_c), .CD(n9365), 
            .Q(wb_smpl_data[14]));   // d:/documents/git_local/fm_modulator/rtl/top.v(212[9] 220[10])
    defparam wb_smpl_data_i14.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i13 (.D(n2023), .CK(dac_clk_p_c), .CD(n9365), 
            .Q(wb_smpl_data[13]));   // d:/documents/git_local/fm_modulator/rtl/top.v(212[9] 220[10])
    defparam wb_smpl_data_i13.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i12 (.D(n2024), .CK(dac_clk_p_c), .CD(n9365), 
            .Q(wb_smpl_data[12]));   // d:/documents/git_local/fm_modulator/rtl/top.v(212[9] 220[10])
    defparam wb_smpl_data_i12.GSR = "DISABLED";
    fm_generator_wb_slave o_dac_a_9__I_0 (.dac_clk_p_c(dac_clk_p_c), .wb_odata({wb_odata}), 
            .n26683(n26683), .wb_fm_data({wb_fm_data}), .\wb_addr[1] (wb_addr[1]), 
            .wb_fm_ack(wb_fm_ack), .o_dac_a_9__N_1(o_dac_a_9__N_1), .GND_net(GND_net), 
            .\wb_addr[0] (wb_addr[0]), .\power_counter[1] (power_counter[1]), 
            .\smpl_register[1] (smpl_register[1]), .n2035(n2035), .n26563(n26563), 
            .n38(n38), .n34(n34), .\wb_addr[8] (wb_addr[8]), .\wb_addr[12] (wb_addr[12]), 
            .n26557(n26557), .\wb_addr[15] (wb_addr[15]), .\wb_addr[9] (wb_addr[9]), 
            .o_dac_cw_b_c_c(o_dac_cw_b_c_c), .n2(n2_adj_3060), .\smpl_register[16] (smpl_register[16]), 
            .n26331(n26331), .n2_adj_1(n2_adj_3071), .\smpl_register[10] (smpl_register[10]), 
            .n26342(n26342), .n2_adj_2(n2_adj_3072), .\smpl_register[9] (smpl_register[9]), 
            .n26341(n26341), .n2_adj_3(n2_adj_3038), .\smpl_register[29] (smpl_register[29]), 
            .n26339(n26339), .n2_adj_4(n2_adj_3055), .\smpl_register[20] (smpl_register[20]), 
            .n26337(n26337), .n2_adj_5(n2_adj_3079), .\smpl_register[5] (smpl_register[5]), 
            .n26336(n26336), .n2_adj_6(n2_adj_3058), .\smpl_register[18] (smpl_register[18]), 
            .n26333(n26333), .n2_adj_7(n2_adj_3059), .\smpl_register[17] (smpl_register[17]), 
            .n26332(n26332), .o_dac_a_c_5(o_dac_a_c_5), .o_dac_b_c_15(o_dac_b_c_15), 
            .o_dac_b_c_9(o_dac_b_c_9), .n26643(n26643), .o_dac_a_c_9(o_dac_a_c_9), 
            .n20438(n20438), .n20864(n20864), .n20416(n20416), .n20402(n20402), 
            .n20422(n20422), .o_dac_b_c_7(o_dac_b_c_7), .\o_sample_i[7] (o_sample_i[7]), 
            .\o_sample_i[14] (o_sample_i[14]), .\o_sample_i[13] (o_sample_i[13]), 
            .\o_sample_i[11] (o_sample_i[11]), .\o_sample_i[10] (o_sample_i[10]), 
            .\o_sample_i[9] (o_sample_i[9]), .\o_sample_i[8] (o_sample_i[8]), 
            .n29209(n29209), .o_dac_b_c_14(o_dac_b_c_14), .o_dac_b_c_13(o_dac_b_c_13), 
            .o_dac_b_c_12(o_dac_b_c_12), .o_dac_b_c_11(o_dac_b_c_11), .o_dac_b_c_10(o_dac_b_c_10), 
            .n3537(n3537), .o_dac_b_c_8(o_dac_b_c_8)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(120[2] 132[2])
    dynamic_pll lo_gen (.i_clk_2f_N_2250(i_clk_2f_N_2250), .lo_pll_out(lo_pll_out), 
            .i_ref_clk_c(i_ref_clk_c), .pll_clk(pll_clk), .pll_rst(pll_rst), 
            .pll_stb(pll_stb), .pll_we(pll_we), .pll_data_i({pll_data_i}), 
            .pll_addr({pll_addr}), .pll_data_o({pll_data_o}), .pll_ack(pll_ack), 
            .GND_net(GND_net)) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(164[13] 175[5])
    
endmodule
//
// Verilog Description of module \rxuartlite(CLOCKS_PER_BAUD=10000) 
//

module \rxuartlite(CLOCKS_PER_BAUD=10000)  (dac_clk_p_c, \rx_data[0] , rx_stb, 
            i_wbu_uart_rx_c, chg_counter, dac_clk_p_c_enable_174, chg_counter_23__N_406, 
            GND_net, \rx_data[6] , \rx_data[5] , \rx_data[4] , \rx_data[3] , 
            \rx_data[2] , \rx_data[1] ) /* synthesis syn_module_defined=1 */ ;
    input dac_clk_p_c;
    output \rx_data[0] ;
    output rx_stb;
    input i_wbu_uart_rx_c;
    output [23:0]chg_counter;
    input dac_clk_p_c_enable_174;
    output chg_counter_23__N_406;
    input GND_net;
    output \rx_data[6] ;
    output \rx_data[5] ;
    output \rx_data[4] ;
    output \rx_data[3] ;
    output \rx_data[2] ;
    output \rx_data[1] ;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(29[49:58])
    
    wire qq_uart, q_uart, ck_uart, o_data_7__N_418;
    wire [7:0]data_reg;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(142[12:20])
    wire [3:0]state;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(75[13:18])
    
    wire dac_clk_p_c_enable_347;
    wire [3:0]state_3__N_322;
    
    wire half_baud_time, half_baud_time_N_457;
    wire [23:0]baud_counter;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(78[17:29])
    
    wire dac_clk_p_c_enable_412, baud_counter_23__N_445;
    wire [23:0]baud_counter_23__N_421;
    wire [23:0]n8;
    
    wire zero_baud_counter, dac_clk_p_c_enable_144, n14838, n17388, 
        n17389, n17331, n17332, n17387, n17330, n17329, n17386, 
        n17385, n17384, n17383, n17382, n17381, n17328, n17380, 
        n17379, n17327, n17326, n164;
    wire [3:0]n174;
    
    wire state_3__N_415, n171, n26444, zero_baud_counter_N_454;
    wire [23:0]n254;
    
    wire n11580, n17422, n17421, n17420, n17419, n20107, n26420, 
        n20676, n20684, n20682, n20674, n20660, n20670, n20672, 
        n20662, n17418, n17417, n17416, n26788, n26787, n26554, 
        n17415, n25473, n25472, data_reg_7__N_416, n17414, n17413, 
        n17412, n17411, half_baud_time_N_458, dac_clk_p_c_enable_343, 
        n17337, n17336, n17335, n17334, n17333, n17390;
    
    FD1S3AY qq_uart_70 (.D(q_uart), .CK(dac_clk_p_c), .Q(qq_uart)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(90[9] 91[66])
    defparam qq_uart_70.GSR = "DISABLED";
    FD1S3AY ck_uart_71 (.D(qq_uart), .CK(dac_clk_p_c), .Q(ck_uart)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(90[9] 91[66])
    defparam ck_uart_71.GSR = "DISABLED";
    FD1P3AX o_data__i1 (.D(data_reg[0]), .SP(o_data_7__N_418), .CK(dac_clk_p_c), 
            .Q(\rx_data[0] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(155[9] 161[18])
    defparam o_data__i1.GSR = "DISABLED";
    FD1P3AY state_i0 (.D(state_3__N_322[0]), .SP(dac_clk_p_c_enable_347), 
            .CK(dac_clk_p_c), .Q(state[0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(116[9] 134[5])
    defparam state_i0.GSR = "DISABLED";
    FD1S3AX half_baud_time_73 (.D(half_baud_time_N_457), .CK(dac_clk_p_c), 
            .Q(half_baud_time)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(111[9] 112[70])
    defparam half_baud_time_73.GSR = "DISABLED";
    FD1S3AX o_wr_76 (.D(o_data_7__N_418), .CK(dac_clk_p_c), .Q(rx_stb)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(155[9] 161[18])
    defparam o_wr_76.GSR = "DISABLED";
    FD1S3AY q_uart_69 (.D(i_wbu_uart_rx_c), .CK(dac_clk_p_c), .Q(q_uart)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(90[9] 91[66])
    defparam q_uart_69.GSR = "DISABLED";
    FD1P3JX baud_counter_i1 (.D(baud_counter_23__N_421[1]), .SP(dac_clk_p_c_enable_412), 
            .PD(baud_counter_23__N_445), .CK(dac_clk_p_c), .Q(baud_counter[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i1.GSR = "DISABLED";
    FD1P3IX chg_counter__i0 (.D(n8[0]), .SP(dac_clk_p_c_enable_174), .CD(chg_counter_23__N_406), 
            .CK(dac_clk_p_c), .Q(chg_counter[0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i0.GSR = "DISABLED";
    FD1P3JX baud_counter_i2 (.D(baud_counter_23__N_421[2]), .SP(dac_clk_p_c_enable_412), 
            .PD(baud_counter_23__N_445), .CK(dac_clk_p_c), .Q(baud_counter[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i2.GSR = "DISABLED";
    FD1P3JX baud_counter_i3 (.D(baud_counter_23__N_421[3]), .SP(dac_clk_p_c_enable_412), 
            .PD(baud_counter_23__N_445), .CK(dac_clk_p_c), .Q(baud_counter[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i3.GSR = "DISABLED";
    FD1P3AY zero_baud_counter_79 (.D(n14838), .SP(dac_clk_p_c_enable_144), 
            .CK(dac_clk_p_c), .Q(zero_baud_counter)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(187[9] 195[29])
    defparam zero_baud_counter_79.GSR = "DISABLED";
    CCU2D sub_389_add_2_22 (.A0(chg_counter[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17388), .COUT(n17389));
    defparam sub_389_add_2_22.INIT0 = 16'h5555;
    defparam sub_389_add_2_22.INIT1 = 16'h5555;
    defparam sub_389_add_2_22.INJECT1_0 = "NO";
    defparam sub_389_add_2_22.INJECT1_1 = "NO";
    CCU2D add_8_13 (.A0(chg_counter[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17331), .COUT(n17332), .S0(n8[11]), .S1(n8[12]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:36])
    defparam add_8_13.INIT0 = 16'h5aaa;
    defparam add_8_13.INIT1 = 16'h5aaa;
    defparam add_8_13.INJECT1_0 = "NO";
    defparam add_8_13.INJECT1_1 = "NO";
    CCU2D sub_389_add_2_20 (.A0(chg_counter[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17387), .COUT(n17388));
    defparam sub_389_add_2_20.INIT0 = 16'h5555;
    defparam sub_389_add_2_20.INIT1 = 16'h5555;
    defparam sub_389_add_2_20.INJECT1_0 = "NO";
    defparam sub_389_add_2_20.INJECT1_1 = "NO";
    CCU2D add_8_11 (.A0(chg_counter[9]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(chg_counter[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n17330), .COUT(n17331), .S0(n8[9]), .S1(n8[10]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:36])
    defparam add_8_11.INIT0 = 16'h5aaa;
    defparam add_8_11.INIT1 = 16'h5aaa;
    defparam add_8_11.INJECT1_0 = "NO";
    defparam add_8_11.INJECT1_1 = "NO";
    CCU2D add_8_9 (.A0(chg_counter[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(chg_counter[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n17329), .COUT(n17330), .S0(n8[7]), .S1(n8[8]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:36])
    defparam add_8_9.INIT0 = 16'h5aaa;
    defparam add_8_9.INIT1 = 16'h5aaa;
    defparam add_8_9.INJECT1_0 = "NO";
    defparam add_8_9.INJECT1_1 = "NO";
    CCU2D sub_389_add_2_18 (.A0(chg_counter[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17386), .COUT(n17387));
    defparam sub_389_add_2_18.INIT0 = 16'h5555;
    defparam sub_389_add_2_18.INIT1 = 16'h5555;
    defparam sub_389_add_2_18.INJECT1_0 = "NO";
    defparam sub_389_add_2_18.INJECT1_1 = "NO";
    CCU2D sub_389_add_2_16 (.A0(chg_counter[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17385), .COUT(n17386));
    defparam sub_389_add_2_16.INIT0 = 16'h5555;
    defparam sub_389_add_2_16.INIT1 = 16'h5555;
    defparam sub_389_add_2_16.INJECT1_0 = "NO";
    defparam sub_389_add_2_16.INJECT1_1 = "NO";
    CCU2D sub_389_add_2_14 (.A0(chg_counter[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17384), .COUT(n17385));
    defparam sub_389_add_2_14.INIT0 = 16'h5aaa;
    defparam sub_389_add_2_14.INIT1 = 16'h5555;
    defparam sub_389_add_2_14.INJECT1_0 = "NO";
    defparam sub_389_add_2_14.INJECT1_1 = "NO";
    CCU2D sub_389_add_2_12 (.A0(chg_counter[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17383), .COUT(n17384));
    defparam sub_389_add_2_12.INIT0 = 16'h5555;
    defparam sub_389_add_2_12.INIT1 = 16'h5555;
    defparam sub_389_add_2_12.INJECT1_0 = "NO";
    defparam sub_389_add_2_12.INJECT1_1 = "NO";
    CCU2D sub_389_add_2_10 (.A0(chg_counter[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17382), .COUT(n17383));
    defparam sub_389_add_2_10.INIT0 = 16'h5aaa;
    defparam sub_389_add_2_10.INIT1 = 16'h5aaa;
    defparam sub_389_add_2_10.INJECT1_0 = "NO";
    defparam sub_389_add_2_10.INJECT1_1 = "NO";
    CCU2D sub_389_add_2_8 (.A0(chg_counter[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17381), .COUT(n17382));
    defparam sub_389_add_2_8.INIT0 = 16'h5555;
    defparam sub_389_add_2_8.INIT1 = 16'h5aaa;
    defparam sub_389_add_2_8.INJECT1_0 = "NO";
    defparam sub_389_add_2_8.INJECT1_1 = "NO";
    CCU2D add_8_7 (.A0(chg_counter[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(chg_counter[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n17328), .COUT(n17329), .S0(n8[5]), .S1(n8[6]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:36])
    defparam add_8_7.INIT0 = 16'h5aaa;
    defparam add_8_7.INIT1 = 16'h5aaa;
    defparam add_8_7.INJECT1_0 = "NO";
    defparam add_8_7.INJECT1_1 = "NO";
    CCU2D sub_389_add_2_6 (.A0(chg_counter[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17380), .COUT(n17381));
    defparam sub_389_add_2_6.INIT0 = 16'h5555;
    defparam sub_389_add_2_6.INIT1 = 16'h5555;
    defparam sub_389_add_2_6.INJECT1_0 = "NO";
    defparam sub_389_add_2_6.INJECT1_1 = "NO";
    CCU2D sub_389_add_2_4 (.A0(chg_counter[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17379), .COUT(n17380));
    defparam sub_389_add_2_4.INIT0 = 16'h5aaa;
    defparam sub_389_add_2_4.INIT1 = 16'h5555;
    defparam sub_389_add_2_4.INJECT1_0 = "NO";
    defparam sub_389_add_2_4.INJECT1_1 = "NO";
    CCU2D sub_389_add_2_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(chg_counter[1]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n17379));
    defparam sub_389_add_2_2.INIT0 = 16'h0000;
    defparam sub_389_add_2_2.INIT1 = 16'h5aaa;
    defparam sub_389_add_2_2.INJECT1_0 = "NO";
    defparam sub_389_add_2_2.INJECT1_1 = "NO";
    CCU2D add_8_5 (.A0(chg_counter[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(chg_counter[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n17327), .COUT(n17328), .S0(n8[3]), .S1(n8[4]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:36])
    defparam add_8_5.INIT0 = 16'h5aaa;
    defparam add_8_5.INIT1 = 16'h5aaa;
    defparam add_8_5.INJECT1_0 = "NO";
    defparam add_8_5.INJECT1_1 = "NO";
    CCU2D add_8_3 (.A0(chg_counter[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(chg_counter[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n17326), .COUT(n17327), .S0(n8[1]), .S1(n8[2]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:36])
    defparam add_8_3.INIT0 = 16'h5aaa;
    defparam add_8_3.INIT1 = 16'h5aaa;
    defparam add_8_3.INJECT1_0 = "NO";
    defparam add_8_3.INJECT1_1 = "NO";
    CCU2D add_8_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(chg_counter[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n17326), .S1(n8[0]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:36])
    defparam add_8_1.INIT0 = 16'hF000;
    defparam add_8_1.INIT1 = 16'h5555;
    defparam add_8_1.INJECT1_0 = "NO";
    defparam add_8_1.INJECT1_1 = "NO";
    FD1P3IX chg_counter__i23 (.D(n8[23]), .SP(dac_clk_p_c_enable_174), .CD(chg_counter_23__N_406), 
            .CK(dac_clk_p_c), .Q(chg_counter[23])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i23.GSR = "DISABLED";
    LUT4 state_3__I_0_80_i3_4_lut (.A(n164), .B(n174[2]), .C(state_3__N_415), 
         .D(n171), .Z(state_3__N_322[2])) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A !(B+(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(125[11] 134[5])
    defparam state_3__I_0_80_i3_4_lut.init = 16'h5f5c;
    FD1P3JX baud_counter_i8 (.D(baud_counter_23__N_421[8]), .SP(dac_clk_p_c_enable_412), 
            .PD(baud_counter_23__N_445), .CK(dac_clk_p_c), .Q(baud_counter[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i8.GSR = "DISABLED";
    FD1P3IX chg_counter__i22 (.D(n8[22]), .SP(dac_clk_p_c_enable_174), .CD(chg_counter_23__N_406), 
            .CK(dac_clk_p_c), .Q(chg_counter[22])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i22.GSR = "DISABLED";
    FD1P3IX chg_counter__i21 (.D(n8[21]), .SP(dac_clk_p_c_enable_174), .CD(chg_counter_23__N_406), 
            .CK(dac_clk_p_c), .Q(chg_counter[21])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i21.GSR = "DISABLED";
    FD1P3IX chg_counter__i20 (.D(n8[20]), .SP(dac_clk_p_c_enable_174), .CD(chg_counter_23__N_406), 
            .CK(dac_clk_p_c), .Q(chg_counter[20])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i20.GSR = "DISABLED";
    FD1P3IX chg_counter__i19 (.D(n8[19]), .SP(dac_clk_p_c_enable_174), .CD(chg_counter_23__N_406), 
            .CK(dac_clk_p_c), .Q(chg_counter[19])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i19.GSR = "DISABLED";
    FD1P3IX chg_counter__i18 (.D(n8[18]), .SP(dac_clk_p_c_enable_174), .CD(chg_counter_23__N_406), 
            .CK(dac_clk_p_c), .Q(chg_counter[18])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i18.GSR = "DISABLED";
    FD1P3IX chg_counter__i17 (.D(n8[17]), .SP(dac_clk_p_c_enable_174), .CD(chg_counter_23__N_406), 
            .CK(dac_clk_p_c), .Q(chg_counter[17])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i17.GSR = "DISABLED";
    FD1P3IX chg_counter__i16 (.D(n8[16]), .SP(dac_clk_p_c_enable_174), .CD(chg_counter_23__N_406), 
            .CK(dac_clk_p_c), .Q(chg_counter[16])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i16.GSR = "DISABLED";
    FD1P3IX chg_counter__i15 (.D(n8[15]), .SP(dac_clk_p_c_enable_174), .CD(chg_counter_23__N_406), 
            .CK(dac_clk_p_c), .Q(chg_counter[15])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i15.GSR = "DISABLED";
    FD1P3IX chg_counter__i14 (.D(n8[14]), .SP(dac_clk_p_c_enable_174), .CD(chg_counter_23__N_406), 
            .CK(dac_clk_p_c), .Q(chg_counter[14])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i14.GSR = "DISABLED";
    LUT4 state_3__I_0_80_i2_4_lut (.A(n164), .B(n174[1]), .C(state_3__N_415), 
         .D(n171), .Z(state_3__N_322[1])) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A !(B+(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(125[11] 134[5])
    defparam state_3__I_0_80_i2_4_lut.init = 16'h5f5c;
    FD1P3IX chg_counter__i13 (.D(n8[13]), .SP(dac_clk_p_c_enable_174), .CD(chg_counter_23__N_406), 
            .CK(dac_clk_p_c), .Q(chg_counter[13])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i13.GSR = "DISABLED";
    FD1P3IX chg_counter__i12 (.D(n8[12]), .SP(dac_clk_p_c_enable_174), .CD(chg_counter_23__N_406), 
            .CK(dac_clk_p_c), .Q(chg_counter[12])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i12.GSR = "DISABLED";
    FD1P3IX chg_counter__i11 (.D(n8[11]), .SP(dac_clk_p_c_enable_174), .CD(chg_counter_23__N_406), 
            .CK(dac_clk_p_c), .Q(chg_counter[11])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i11.GSR = "DISABLED";
    FD1P3IX chg_counter__i10 (.D(n8[10]), .SP(dac_clk_p_c_enable_174), .CD(chg_counter_23__N_406), 
            .CK(dac_clk_p_c), .Q(chg_counter[10])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i10.GSR = "DISABLED";
    FD1P3IX chg_counter__i9 (.D(n8[9]), .SP(dac_clk_p_c_enable_174), .CD(chg_counter_23__N_406), 
            .CK(dac_clk_p_c), .Q(chg_counter[9])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i9.GSR = "DISABLED";
    FD1P3IX chg_counter__i8 (.D(n8[8]), .SP(dac_clk_p_c_enable_174), .CD(chg_counter_23__N_406), 
            .CK(dac_clk_p_c), .Q(chg_counter[8])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i8.GSR = "DISABLED";
    FD1P3IX chg_counter__i7 (.D(n8[7]), .SP(dac_clk_p_c_enable_174), .CD(chg_counter_23__N_406), 
            .CK(dac_clk_p_c), .Q(chg_counter[7])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i7.GSR = "DISABLED";
    FD1P3IX chg_counter__i6 (.D(n8[6]), .SP(dac_clk_p_c_enable_174), .CD(chg_counter_23__N_406), 
            .CK(dac_clk_p_c), .Q(chg_counter[6])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i6.GSR = "DISABLED";
    FD1P3IX chg_counter__i5 (.D(n8[5]), .SP(dac_clk_p_c_enable_174), .CD(chg_counter_23__N_406), 
            .CK(dac_clk_p_c), .Q(chg_counter[5])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i5.GSR = "DISABLED";
    FD1P3IX chg_counter__i4 (.D(n8[4]), .SP(dac_clk_p_c_enable_174), .CD(chg_counter_23__N_406), 
            .CK(dac_clk_p_c), .Q(chg_counter[4])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i4.GSR = "DISABLED";
    FD1P3IX chg_counter__i3 (.D(n8[3]), .SP(dac_clk_p_c_enable_174), .CD(chg_counter_23__N_406), 
            .CK(dac_clk_p_c), .Q(chg_counter[3])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i3.GSR = "DISABLED";
    FD1P3IX chg_counter__i2 (.D(n8[2]), .SP(dac_clk_p_c_enable_174), .CD(chg_counter_23__N_406), 
            .CK(dac_clk_p_c), .Q(chg_counter[2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i2.GSR = "DISABLED";
    FD1P3IX chg_counter__i1 (.D(n8[1]), .SP(dac_clk_p_c_enable_174), .CD(chg_counter_23__N_406), 
            .CK(dac_clk_p_c), .Q(chg_counter[1])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[37])
    defparam chg_counter__i1.GSR = "DISABLED";
    FD1P3JX baud_counter_i9 (.D(baud_counter_23__N_421[9]), .SP(dac_clk_p_c_enable_412), 
            .PD(baud_counter_23__N_445), .CK(dac_clk_p_c), .Q(baud_counter[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i9.GSR = "DISABLED";
    FD1P3JX baud_counter_i10 (.D(baud_counter_23__N_421[10]), .SP(dac_clk_p_c_enable_412), 
            .PD(baud_counter_23__N_445), .CK(dac_clk_p_c), .Q(baud_counter[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i10.GSR = "DISABLED";
    FD1P3JX baud_counter_i13 (.D(baud_counter_23__N_421[13]), .SP(dac_clk_p_c_enable_412), 
            .PD(baud_counter_23__N_445), .CK(dac_clk_p_c), .Q(baud_counter[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i13.GSR = "DISABLED";
    LUT4 i11577_3_lut_4_lut (.A(state[0]), .B(n26444), .C(zero_baud_counter_N_454), 
         .D(n254[1]), .Z(baud_counter_23__N_421[1])) /* synthesis lut_function=(A (B (C+(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(144[27:48])
    defparam i11577_3_lut_4_lut.init = 16'hddd0;
    LUT4 i1_2_lut_3_lut_4_lut (.A(state[0]), .B(n26444), .C(zero_baud_counter_N_454), 
         .D(baud_counter_23__N_445), .Z(n11580)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(144[27:48])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfff2;
    LUT4 i11576_3_lut_4_lut (.A(state[0]), .B(n26444), .C(zero_baud_counter_N_454), 
         .D(n254[2]), .Z(baud_counter_23__N_421[2])) /* synthesis lut_function=(A (B (C+(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(144[27:48])
    defparam i11576_3_lut_4_lut.init = 16'hddd0;
    LUT4 i11575_3_lut_4_lut (.A(state[0]), .B(n26444), .C(zero_baud_counter_N_454), 
         .D(n254[3]), .Z(baud_counter_23__N_421[3])) /* synthesis lut_function=(A (B (C+(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(144[27:48])
    defparam i11575_3_lut_4_lut.init = 16'hddd0;
    LUT4 i22475_3_lut_4_lut (.A(state[0]), .B(n26444), .C(baud_counter_23__N_445), 
         .D(zero_baud_counter_N_454), .Z(n14838)) /* synthesis lut_function=(!(A (B (C+(D))+!B (C))+!A (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(144[27:48])
    defparam i22475_3_lut_4_lut.init = 16'h020f;
    LUT4 i11573_3_lut_4_lut (.A(state[0]), .B(n26444), .C(zero_baud_counter_N_454), 
         .D(n254[8]), .Z(baud_counter_23__N_421[8])) /* synthesis lut_function=(A (B (C+(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(144[27:48])
    defparam i11573_3_lut_4_lut.init = 16'hddd0;
    LUT4 i11572_3_lut_4_lut (.A(state[0]), .B(n26444), .C(zero_baud_counter_N_454), 
         .D(n254[9]), .Z(baud_counter_23__N_421[9])) /* synthesis lut_function=(A (B (C+(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(144[27:48])
    defparam i11572_3_lut_4_lut.init = 16'hddd0;
    LUT4 i11571_3_lut_4_lut (.A(state[0]), .B(n26444), .C(zero_baud_counter_N_454), 
         .D(n254[10]), .Z(baud_counter_23__N_421[10])) /* synthesis lut_function=(A (B (C+(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(144[27:48])
    defparam i11571_3_lut_4_lut.init = 16'hddd0;
    LUT4 i11570_3_lut_4_lut (.A(state[0]), .B(n26444), .C(zero_baud_counter_N_454), 
         .D(n254[13]), .Z(baud_counter_23__N_421[13])) /* synthesis lut_function=(A (B (C+(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(144[27:48])
    defparam i11570_3_lut_4_lut.init = 16'hddd0;
    LUT4 i11018_3_lut_4_lut (.A(state[0]), .B(n26444), .C(zero_baud_counter_N_454), 
         .D(n254[0]), .Z(baud_counter_23__N_421[0])) /* synthesis lut_function=(A (B (C+(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(144[27:48])
    defparam i11018_3_lut_4_lut.init = 16'hddd0;
    LUT4 i1_3_lut (.A(ck_uart), .B(state_3__N_415), .C(half_baud_time), 
         .Z(baud_counter_23__N_445)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(171[6:57])
    defparam i1_3_lut.init = 16'h4040;
    CCU2D sub_49_add_2_25 (.A0(baud_counter[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n17422), .S0(n254[23]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_25.INIT0 = 16'h5555;
    defparam sub_49_add_2_25.INIT1 = 16'h0000;
    defparam sub_49_add_2_25.INJECT1_0 = "NO";
    defparam sub_49_add_2_25.INJECT1_1 = "NO";
    LUT4 zero_baud_counter_I_0_2_lut (.A(zero_baud_counter), .B(state[3]), 
         .Z(zero_baud_counter_N_454)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(175[11:52])
    defparam zero_baud_counter_I_0_2_lut.init = 16'h2222;
    LUT4 qq_uart_I_0_2_lut (.A(qq_uart), .B(ck_uart), .Z(chg_counter_23__N_406)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(100[6:24])
    defparam qq_uart_I_0_2_lut.init = 16'h6666;
    CCU2D sub_49_add_2_23 (.A0(baud_counter[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17421), .COUT(n17422), .S0(n254[21]), 
          .S1(n254[22]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_23.INIT0 = 16'h5555;
    defparam sub_49_add_2_23.INIT1 = 16'h5555;
    defparam sub_49_add_2_23.INJECT1_0 = "NO";
    defparam sub_49_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_49_add_2_21 (.A0(baud_counter[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17420), .COUT(n17421), .S0(n254[19]), 
          .S1(n254[20]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_21.INIT0 = 16'h5555;
    defparam sub_49_add_2_21.INIT1 = 16'h5555;
    defparam sub_49_add_2_21.INJECT1_0 = "NO";
    defparam sub_49_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_49_add_2_19 (.A0(baud_counter[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17419), .COUT(n17420), .S0(n254[17]), 
          .S1(n254[18]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_19.INIT0 = 16'h5555;
    defparam sub_49_add_2_19.INIT1 = 16'h5555;
    defparam sub_49_add_2_19.INJECT1_0 = "NO";
    defparam sub_49_add_2_19.INJECT1_1 = "NO";
    LUT4 i1_4_lut (.A(n20107), .B(n26420), .C(baud_counter_23__N_445), 
         .D(zero_baud_counter_N_454), .Z(dac_clk_p_c_enable_144)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;
    defparam i1_4_lut.init = 16'hfff7;
    LUT4 i1_4_lut_adj_131 (.A(n20676), .B(n20684), .C(n20682), .D(n20674), 
         .Z(n20107)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(194[11:28])
    defparam i1_4_lut_adj_131.init = 16'hfffe;
    LUT4 i1_4_lut_adj_132 (.A(baud_counter[14]), .B(baud_counter[21]), .C(baud_counter[20]), 
         .D(baud_counter[3]), .Z(n20676)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(194[11:28])
    defparam i1_4_lut_adj_132.init = 16'hfffe;
    LUT4 i1_4_lut_adj_133 (.A(n20660), .B(baud_counter[0]), .C(n20670), 
         .D(baud_counter[8]), .Z(n20684)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(194[11:28])
    defparam i1_4_lut_adj_133.init = 16'hfffb;
    LUT4 i1_4_lut_adj_134 (.A(baud_counter[7]), .B(n20672), .C(n20662), 
         .D(baud_counter[22]), .Z(n20682)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(194[11:28])
    defparam i1_4_lut_adj_134.init = 16'hfffe;
    LUT4 i1_4_lut_adj_135 (.A(baud_counter[6]), .B(baud_counter[12]), .C(baud_counter[13]), 
         .D(baud_counter[5]), .Z(n20674)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(194[11:28])
    defparam i1_4_lut_adj_135.init = 16'hfffe;
    LUT4 i1_2_lut (.A(baud_counter[19]), .B(baud_counter[1]), .Z(n20660)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(194[11:28])
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i1_4_lut_adj_136 (.A(baud_counter[15]), .B(baud_counter[9]), .C(baud_counter[17]), 
         .D(baud_counter[23]), .Z(n20670)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(194[11:28])
    defparam i1_4_lut_adj_136.init = 16'hfffe;
    LUT4 i1_4_lut_adj_137 (.A(baud_counter[4]), .B(baud_counter[16]), .C(baud_counter[18]), 
         .D(baud_counter[2]), .Z(n20672)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(194[11:28])
    defparam i1_4_lut_adj_137.init = 16'hfffe;
    LUT4 i1_2_lut_adj_138 (.A(baud_counter[11]), .B(baud_counter[10]), .Z(n20662)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(194[11:28])
    defparam i1_2_lut_adj_138.init = 16'heeee;
    CCU2D sub_49_add_2_17 (.A0(baud_counter[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17418), .COUT(n17419), .S0(n254[15]), 
          .S1(n254[16]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_17.INIT0 = 16'h5555;
    defparam sub_49_add_2_17.INIT1 = 16'h5555;
    defparam sub_49_add_2_17.INJECT1_0 = "NO";
    defparam sub_49_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_49_add_2_15 (.A0(baud_counter[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17417), .COUT(n17418), .S0(n254[13]), 
          .S1(n254[14]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_15.INIT0 = 16'h5555;
    defparam sub_49_add_2_15.INIT1 = 16'h5555;
    defparam sub_49_add_2_15.INJECT1_0 = "NO";
    defparam sub_49_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_49_add_2_13 (.A0(baud_counter[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17416), .COUT(n17417), .S0(n254[11]), 
          .S1(n254[12]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_13.INIT0 = 16'h5555;
    defparam sub_49_add_2_13.INIT1 = 16'h5555;
    defparam sub_49_add_2_13.INJECT1_0 = "NO";
    defparam sub_49_add_2_13.INJECT1_1 = "NO";
    LUT4 state_3__I_0_80_i4_4_lut_then_4_lut (.A(n164), .B(state[0]), .C(state[2]), 
         .D(state[1]), .Z(n26788)) /* synthesis lut_function=(!(A (B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(125[11] 134[5])
    defparam state_3__I_0_80_i4_4_lut_then_4_lut.init = 16'h7fff;
    LUT4 state_3__I_0_80_i4_4_lut_else_4_lut (.A(state[0]), .B(n171), .C(state[2]), 
         .D(state[1]), .Z(n26787)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(125[11] 134[5])
    defparam state_3__I_0_80_i4_4_lut_else_4_lut.init = 16'heccc;
    LUT4 i1_3_lut_4_lut (.A(state[0]), .B(n26554), .C(ck_uart), .D(state[3]), 
         .Z(n171)) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(144[27:48])
    defparam i1_3_lut_4_lut.init = 16'he000;
    CCU2D sub_49_add_2_11 (.A0(baud_counter[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17415), .COUT(n17416), .S0(n254[9]), .S1(n254[10]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_11.INIT0 = 16'h5555;
    defparam sub_49_add_2_11.INIT1 = 16'h5555;
    defparam sub_49_add_2_11.INJECT1_0 = "NO";
    defparam sub_49_add_2_11.INJECT1_1 = "NO";
    LUT4 state_3__N_415_bdd_4_lut (.A(state[0]), .B(state[3]), .C(n26554), 
         .D(ck_uart), .Z(n25473)) /* synthesis lut_function=(A (B)+!A (((D)+!C)+!B)) */ ;
    defparam state_3__N_415_bdd_4_lut.init = 16'hdd9d;
    LUT4 state_3__N_415_bdd_2_lut (.A(half_baud_time), .B(ck_uart), .Z(n25472)) /* synthesis lut_function=((B)+!A) */ ;
    defparam state_3__N_415_bdd_2_lut.init = 16'hdddd;
    LUT4 zero_baud_counter_I_0_82_2_lut_3_lut_4_lut (.A(state[3]), .B(n26554), 
         .C(zero_baud_counter), .D(state[0]), .Z(data_reg_7__N_416)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(144[27:48])
    defparam zero_baud_counter_I_0_82_2_lut_3_lut_4_lut.init = 16'hf0d0;
    CCU2D sub_49_add_2_9 (.A0(baud_counter[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17414), .COUT(n17415), .S0(n254[7]), .S1(n254[8]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_9.INIT0 = 16'h5555;
    defparam sub_49_add_2_9.INIT1 = 16'h5555;
    defparam sub_49_add_2_9.INJECT1_0 = "NO";
    defparam sub_49_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_49_add_2_7 (.A0(baud_counter[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17413), .COUT(n17414), .S0(n254[5]), .S1(n254[6]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_7.INIT0 = 16'h5555;
    defparam sub_49_add_2_7.INIT1 = 16'h5555;
    defparam sub_49_add_2_7.INJECT1_0 = "NO";
    defparam sub_49_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_49_add_2_5 (.A0(baud_counter[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17412), .COUT(n17413), .S0(n254[3]), .S1(n254[4]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_5.INIT0 = 16'h5555;
    defparam sub_49_add_2_5.INIT1 = 16'h5555;
    defparam sub_49_add_2_5.INJECT1_0 = "NO";
    defparam sub_49_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_49_add_2_3 (.A0(baud_counter[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17411), .COUT(n17412), .S0(n254[1]), .S1(n254[2]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_3.INIT0 = 16'h5555;
    defparam sub_49_add_2_3.INIT1 = 16'h5555;
    defparam sub_49_add_2_3.INJECT1_0 = "NO";
    defparam sub_49_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_49_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(baud_counter[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n17411), .S1(n254[0]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_1.INIT0 = 16'hF000;
    defparam sub_49_add_2_1.INIT1 = 16'h5555;
    defparam sub_49_add_2_1.INJECT1_0 = "NO";
    defparam sub_49_add_2_1.INJECT1_1 = "NO";
    LUT4 i1_3_lut_4_lut_adj_139 (.A(state[0]), .B(n26444), .C(ck_uart), 
         .D(zero_baud_counter), .Z(o_data_7__N_418)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(144[27:48])
    defparam i1_3_lut_4_lut_adj_139.init = 16'h1000;
    LUT4 i1_3_lut_adj_140 (.A(state_3__N_415), .B(n171), .C(zero_baud_counter), 
         .Z(dac_clk_p_c_enable_347)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_3_lut_adj_140.init = 16'hfefe;
    LUT4 i21_2_lut (.A(ck_uart), .B(half_baud_time), .Z(n164)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(121[7:35])
    defparam i21_2_lut.init = 16'h4444;
    LUT4 i1_4_lut_adj_141 (.A(state[0]), .B(state[2]), .C(state[3]), .D(state[1]), 
         .Z(state_3__N_415)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_141.init = 16'h8000;
    LUT4 ck_uart_N_448_I_0_2_lut (.A(ck_uart), .B(half_baud_time_N_458), 
         .Z(half_baud_time_N_457)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(112[21:69])
    defparam ck_uart_N_448_I_0_2_lut.init = 16'h4444;
    FD1P3IX baud_counter_i23 (.D(n254[23]), .SP(dac_clk_p_c_enable_343), 
            .CD(n11580), .CK(dac_clk_p_c), .Q(baud_counter[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i23.GSR = "DISABLED";
    LUT4 i1_3_lut_4_lut_adj_142 (.A(baud_counter_23__N_445), .B(n26420), 
         .C(state[3]), .D(zero_baud_counter), .Z(dac_clk_p_c_enable_412)) /* synthesis lut_function=(A+!(B (C (D)))) */ ;
    defparam i1_3_lut_4_lut_adj_142.init = 16'hbfff;
    LUT4 i9663_1_lut (.A(zero_baud_counter), .Z(dac_clk_p_c_enable_343)) /* synthesis lut_function=(!(A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(187[9] 195[29])
    defparam i9663_1_lut.init = 16'h5555;
    FD1P3IX baud_counter_i22 (.D(n254[22]), .SP(dac_clk_p_c_enable_343), 
            .CD(n11580), .CK(dac_clk_p_c), .Q(baud_counter[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i22.GSR = "DISABLED";
    FD1P3IX baud_counter_i21 (.D(n254[21]), .SP(dac_clk_p_c_enable_343), 
            .CD(n11580), .CK(dac_clk_p_c), .Q(baud_counter[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i21.GSR = "DISABLED";
    FD1P3IX baud_counter_i20 (.D(n254[20]), .SP(dac_clk_p_c_enable_343), 
            .CD(n11580), .CK(dac_clk_p_c), .Q(baud_counter[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i20.GSR = "DISABLED";
    FD1P3IX baud_counter_i19 (.D(n254[19]), .SP(dac_clk_p_c_enable_343), 
            .CD(n11580), .CK(dac_clk_p_c), .Q(baud_counter[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i19.GSR = "DISABLED";
    FD1P3IX baud_counter_i18 (.D(n254[18]), .SP(dac_clk_p_c_enable_343), 
            .CD(n11580), .CK(dac_clk_p_c), .Q(baud_counter[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i18.GSR = "DISABLED";
    FD1P3IX baud_counter_i17 (.D(n254[17]), .SP(dac_clk_p_c_enable_343), 
            .CD(n11580), .CK(dac_clk_p_c), .Q(baud_counter[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i17.GSR = "DISABLED";
    FD1P3IX baud_counter_i16 (.D(n254[16]), .SP(dac_clk_p_c_enable_343), 
            .CD(n11580), .CK(dac_clk_p_c), .Q(baud_counter[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i16.GSR = "DISABLED";
    FD1P3IX baud_counter_i15 (.D(n254[15]), .SP(dac_clk_p_c_enable_343), 
            .CD(n11580), .CK(dac_clk_p_c), .Q(baud_counter[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i15.GSR = "DISABLED";
    FD1P3IX baud_counter_i14 (.D(n254[14]), .SP(dac_clk_p_c_enable_343), 
            .CD(n11580), .CK(dac_clk_p_c), .Q(baud_counter[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i14.GSR = "DISABLED";
    FD1P3IX baud_counter_i12 (.D(n254[12]), .SP(dac_clk_p_c_enable_343), 
            .CD(n11580), .CK(dac_clk_p_c), .Q(baud_counter[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i12.GSR = "DISABLED";
    FD1P3IX baud_counter_i11 (.D(n254[11]), .SP(dac_clk_p_c_enable_343), 
            .CD(n11580), .CK(dac_clk_p_c), .Q(baud_counter[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i11.GSR = "DISABLED";
    FD1P3IX baud_counter_i7 (.D(n254[7]), .SP(dac_clk_p_c_enable_343), .CD(n11580), 
            .CK(dac_clk_p_c), .Q(baud_counter[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i7.GSR = "DISABLED";
    FD1P3IX baud_counter_i6 (.D(n254[6]), .SP(dac_clk_p_c_enable_343), .CD(n11580), 
            .CK(dac_clk_p_c), .Q(baud_counter[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i6.GSR = "DISABLED";
    FD1P3IX baud_counter_i5 (.D(n254[5]), .SP(dac_clk_p_c_enable_343), .CD(n11580), 
            .CK(dac_clk_p_c), .Q(baud_counter[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i5.GSR = "DISABLED";
    FD1P3IX baud_counter_i4 (.D(n254[4]), .SP(dac_clk_p_c_enable_343), .CD(n11580), 
            .CK(dac_clk_p_c), .Q(baud_counter[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i4.GSR = "DISABLED";
    FD1P3AY state_i3 (.D(state_3__N_322[3]), .SP(dac_clk_p_c_enable_347), 
            .CK(dac_clk_p_c), .Q(state[3])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(116[9] 134[5])
    defparam state_i3.GSR = "DISABLED";
    CCU2D add_8_25 (.A0(chg_counter[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n17337), .S0(n8[23]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:36])
    defparam add_8_25.INIT0 = 16'h5aaa;
    defparam add_8_25.INIT1 = 16'h0000;
    defparam add_8_25.INJECT1_0 = "NO";
    defparam add_8_25.INJECT1_1 = "NO";
    FD1P3AY state_i2 (.D(state_3__N_322[2]), .SP(dac_clk_p_c_enable_347), 
            .CK(dac_clk_p_c), .Q(state[2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(116[9] 134[5])
    defparam state_i2.GSR = "DISABLED";
    FD1P3AY state_i1 (.D(state_3__N_322[1]), .SP(dac_clk_p_c_enable_347), 
            .CK(dac_clk_p_c), .Q(state[1])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(116[9] 134[5])
    defparam state_i1.GSR = "DISABLED";
    FD1P3AX o_data__i7 (.D(data_reg[6]), .SP(o_data_7__N_418), .CK(dac_clk_p_c), 
            .Q(\rx_data[6] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(155[9] 161[18])
    defparam o_data__i7.GSR = "DISABLED";
    FD1P3AX o_data__i6 (.D(data_reg[5]), .SP(o_data_7__N_418), .CK(dac_clk_p_c), 
            .Q(\rx_data[5] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(155[9] 161[18])
    defparam o_data__i6.GSR = "DISABLED";
    FD1P3AX o_data__i5 (.D(data_reg[4]), .SP(o_data_7__N_418), .CK(dac_clk_p_c), 
            .Q(\rx_data[4] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(155[9] 161[18])
    defparam o_data__i5.GSR = "DISABLED";
    FD1P3AX o_data__i4 (.D(data_reg[3]), .SP(o_data_7__N_418), .CK(dac_clk_p_c), 
            .Q(\rx_data[3] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(155[9] 161[18])
    defparam o_data__i4.GSR = "DISABLED";
    FD1P3AX o_data__i3 (.D(data_reg[2]), .SP(o_data_7__N_418), .CK(dac_clk_p_c), 
            .Q(\rx_data[2] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(155[9] 161[18])
    defparam o_data__i3.GSR = "DISABLED";
    FD1P3AX o_data__i2 (.D(data_reg[1]), .SP(o_data_7__N_418), .CK(dac_clk_p_c), 
            .Q(\rx_data[1] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(155[9] 161[18])
    defparam o_data__i2.GSR = "DISABLED";
    CCU2D add_8_23 (.A0(chg_counter[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17336), .COUT(n17337), .S0(n8[21]), .S1(n8[22]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:36])
    defparam add_8_23.INIT0 = 16'h5aaa;
    defparam add_8_23.INIT1 = 16'h5aaa;
    defparam add_8_23.INJECT1_0 = "NO";
    defparam add_8_23.INJECT1_1 = "NO";
    LUT4 i6508_2_lut_rep_594 (.A(state[1]), .B(state[2]), .Z(n26554)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(129[7:26])
    defparam i6508_2_lut_rep_594.init = 16'heeee;
    LUT4 i1_2_lut_rep_484_3_lut (.A(state[1]), .B(state[2]), .C(state[3]), 
         .Z(n26444)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(129[7:26])
    defparam i1_2_lut_rep_484_3_lut.init = 16'hefef;
    LUT4 i1_2_lut_rep_460_3_lut_4_lut (.A(state[1]), .B(state[2]), .C(state[0]), 
         .D(state[3]), .Z(n26420)) /* synthesis lut_function=(A+(B+!(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(129[7:26])
    defparam i1_2_lut_rep_460_3_lut_4_lut.init = 16'hefff;
    CCU2D add_8_21 (.A0(chg_counter[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17335), .COUT(n17336), .S0(n8[19]), .S1(n8[20]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:36])
    defparam add_8_21.INIT0 = 16'h5aaa;
    defparam add_8_21.INIT1 = 16'h5aaa;
    defparam add_8_21.INJECT1_0 = "NO";
    defparam add_8_21.INJECT1_1 = "NO";
    LUT4 i764_2_lut_3_lut (.A(state[0]), .B(state[3]), .C(state[1]), .Z(n174[1])) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(133[13:25])
    defparam i764_2_lut_3_lut.init = 16'hd2d2;
    LUT4 i771_2_lut_3_lut_4_lut (.A(state[0]), .B(state[3]), .C(state[2]), 
         .D(state[1]), .Z(n174[2])) /* synthesis lut_function=(A (B (C)+!B !(C (D)+!C !(D)))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(133[13:25])
    defparam i771_2_lut_3_lut_4_lut.init = 16'hd2f0;
    PFUMX i23792 (.BLUT(n25473), .ALUT(n25472), .C0(state_3__N_415), .Z(state_3__N_322[0]));
    PFUMX i24495 (.BLUT(n26787), .ALUT(n26788), .C0(state[3]), .Z(state_3__N_322[3]));
    CCU2D add_8_19 (.A0(chg_counter[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17334), .COUT(n17335), .S0(n8[17]), .S1(n8[18]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:36])
    defparam add_8_19.INIT0 = 16'h5aaa;
    defparam add_8_19.INIT1 = 16'h5aaa;
    defparam add_8_19.INJECT1_0 = "NO";
    defparam add_8_19.INJECT1_1 = "NO";
    FD1P3JX baud_counter_i0 (.D(baud_counter_23__N_421[0]), .SP(dac_clk_p_c_enable_412), 
            .PD(baud_counter_23__N_445), .CK(dac_clk_p_c), .Q(baud_counter[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i0.GSR = "DISABLED";
    CCU2D add_8_17 (.A0(chg_counter[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17333), .COUT(n17334), .S0(n8[15]), .S1(n8[16]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:36])
    defparam add_8_17.INIT0 = 16'h5aaa;
    defparam add_8_17.INIT1 = 16'h5aaa;
    defparam add_8_17.INJECT1_0 = "NO";
    defparam add_8_17.INJECT1_1 = "NO";
    CCU2D sub_389_add_2_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n17390), .S0(half_baud_time_N_458));
    defparam sub_389_add_2_cout.INIT0 = 16'h0000;
    defparam sub_389_add_2_cout.INIT1 = 16'h0000;
    defparam sub_389_add_2_cout.INJECT1_0 = "NO";
    defparam sub_389_add_2_cout.INJECT1_1 = "NO";
    CCU2D add_8_15 (.A0(chg_counter[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17332), .COUT(n17333), .S0(n8[13]), .S1(n8[14]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:36])
    defparam add_8_15.INIT0 = 16'h5aaa;
    defparam add_8_15.INIT1 = 16'h5aaa;
    defparam add_8_15.INJECT1_0 = "NO";
    defparam add_8_15.INJECT1_1 = "NO";
    CCU2D sub_389_add_2_24 (.A0(chg_counter[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17389), .COUT(n17390));
    defparam sub_389_add_2_24.INIT0 = 16'h5555;
    defparam sub_389_add_2_24.INIT1 = 16'h5555;
    defparam sub_389_add_2_24.INJECT1_0 = "NO";
    defparam sub_389_add_2_24.INJECT1_1 = "NO";
    FD1P3AX data_reg_i0_i7 (.D(qq_uart), .SP(data_reg_7__N_416), .CK(dac_clk_p_c), 
            .Q(data_reg[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(143[9] 145[42])
    defparam data_reg_i0_i7.GSR = "DISABLED";
    FD1P3AX data_reg_i0_i6 (.D(data_reg[7]), .SP(data_reg_7__N_416), .CK(dac_clk_p_c), 
            .Q(data_reg[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(143[9] 145[42])
    defparam data_reg_i0_i6.GSR = "DISABLED";
    FD1P3AX data_reg_i0_i5 (.D(data_reg[6]), .SP(data_reg_7__N_416), .CK(dac_clk_p_c), 
            .Q(data_reg[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(143[9] 145[42])
    defparam data_reg_i0_i5.GSR = "DISABLED";
    FD1P3AX data_reg_i0_i4 (.D(data_reg[5]), .SP(data_reg_7__N_416), .CK(dac_clk_p_c), 
            .Q(data_reg[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(143[9] 145[42])
    defparam data_reg_i0_i4.GSR = "DISABLED";
    FD1P3AX data_reg_i0_i3 (.D(data_reg[4]), .SP(data_reg_7__N_416), .CK(dac_clk_p_c), 
            .Q(data_reg[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(143[9] 145[42])
    defparam data_reg_i0_i3.GSR = "DISABLED";
    FD1P3AX data_reg_i0_i2 (.D(data_reg[3]), .SP(data_reg_7__N_416), .CK(dac_clk_p_c), 
            .Q(data_reg[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(143[9] 145[42])
    defparam data_reg_i0_i2.GSR = "DISABLED";
    FD1P3AX data_reg_i0_i1 (.D(data_reg[2]), .SP(data_reg_7__N_416), .CK(dac_clk_p_c), 
            .Q(data_reg[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(143[9] 145[42])
    defparam data_reg_i0_i1.GSR = "DISABLED";
    FD1P3AX data_reg_i0_i0 (.D(data_reg[1]), .SP(data_reg_7__N_416), .CK(dac_clk_p_c), 
            .Q(data_reg[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(143[9] 145[42])
    defparam data_reg_i0_i0.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module hbbus
//

module hbbus (wb_odata, dac_clk_p_c, wb_we, wb_stb, wb_cyc, wb_addr, 
            GND_net, wb_err, wb_ack, \wb_idata[0] , \wb_idata[2] , 
            \wb_idata[3] , \wb_idata[4] , \wb_idata[5] , \wb_idata[6] , 
            \wb_idata[7] , \wb_idata[8] , \wb_idata[9] , \wb_idata[10] , 
            \wb_idata[11] , \wb_idata[12] , \wb_idata[13] , \wb_idata[14] , 
            \wb_idata[15] , \wb_idata[16] , \wb_idata[17] , \wb_idata[18] , 
            \wb_idata[19] , \wb_idata[20] , \wb_idata[21] , \wb_idata[22] , 
            \wb_idata[23] , \wb_idata[24] , \wb_idata[25] , \wb_idata[26] , 
            \wb_idata[27] , \wb_idata[28] , \wb_idata[29] , \wb_idata[30] , 
            \wb_idata[31] , n2, n12635, n29210, VCC_net, \rx_data[5] , 
            \rx_data[1] , rx_stb, \rx_data[6] , \rx_data[3] , \rx_data[4] , 
            \rx_data[0] , \rx_data[2] , tx_busy, o_busy_N_536, \state[0] , 
            n17598, n26540, \lcl_data[1] , \lcl_data_7__N_511[0] , \lcl_data[4] , 
            \lcl_data_7__N_511[3] , \lcl_data[5] , \lcl_data_7__N_511[4] , 
            \lcl_data[6] , \lcl_data_7__N_511[5] , \lcl_data[7] , \lcl_data_7__N_511[6] , 
            zero_baud_counter, dac_clk_p_c_enable_321, \lcl_data[3] , 
            \lcl_data_7__N_511[2] , \lcl_data[2] , \lcl_data_7__N_511[1] ) /* synthesis syn_module_defined=1 */ ;
    output [31:0]wb_odata;
    input dac_clk_p_c;
    output wb_we;
    output wb_stb;
    output wb_cyc;
    output [29:0]wb_addr;
    input GND_net;
    input wb_err;
    input wb_ack;
    input \wb_idata[0] ;
    input \wb_idata[2] ;
    input \wb_idata[3] ;
    input \wb_idata[4] ;
    input \wb_idata[5] ;
    input \wb_idata[6] ;
    input \wb_idata[7] ;
    input \wb_idata[8] ;
    input \wb_idata[9] ;
    input \wb_idata[10] ;
    input \wb_idata[11] ;
    input \wb_idata[12] ;
    input \wb_idata[13] ;
    input \wb_idata[14] ;
    input \wb_idata[15] ;
    input \wb_idata[16] ;
    input \wb_idata[17] ;
    input \wb_idata[18] ;
    input \wb_idata[19] ;
    input \wb_idata[20] ;
    input \wb_idata[21] ;
    input \wb_idata[22] ;
    input \wb_idata[23] ;
    input \wb_idata[24] ;
    input \wb_idata[25] ;
    input \wb_idata[26] ;
    input \wb_idata[27] ;
    input \wb_idata[28] ;
    input \wb_idata[29] ;
    input \wb_idata[30] ;
    input \wb_idata[31] ;
    output n2;
    input n12635;
    input n29210;
    input VCC_net;
    input \rx_data[5] ;
    input \rx_data[1] ;
    input rx_stb;
    input \rx_data[6] ;
    input \rx_data[3] ;
    input \rx_data[4] ;
    input \rx_data[0] ;
    input \rx_data[2] ;
    input tx_busy;
    input o_busy_N_536;
    input \state[0] ;
    output n17598;
    output n26540;
    input \lcl_data[1] ;
    output \lcl_data_7__N_511[0] ;
    input \lcl_data[4] ;
    output \lcl_data_7__N_511[3] ;
    input \lcl_data[5] ;
    output \lcl_data_7__N_511[4] ;
    input \lcl_data[6] ;
    output \lcl_data_7__N_511[5] ;
    input \lcl_data[7] ;
    output \lcl_data_7__N_511[6] ;
    input zero_baud_counter;
    output dac_clk_p_c_enable_321;
    input \lcl_data[3] ;
    output \lcl_data_7__N_511[2] ;
    input \lcl_data[2] ;
    output \lcl_data_7__N_511[1] ;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(29[49:58])
    wire [33:0]iw_word;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(71[14:21])
    
    wire inc, dac_clk_p_c_enable_136, ow_stb;
    wire [33:0]ow_word;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(73[14:21])
    
    wire n29269, i_cmd_wr, n21860, newaddr_N_990, n17206, n29268, 
        n26716, n26715, dac_clk_p_c_enable_446, dac_clk_p_c_enable_307;
    wire [4:0]hb_bits;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(79[13:20])
    
    wire dac_clk_p_c_enable_193;
    wire [33:0]idl_word;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(77[14:22])
    
    wire hb_busy, w_reset, n26536, idl_stb, nl_busy, hx_stb, dac_clk_p_c_enable_380, 
        o_pck_stb_N_765, cmd_loaded, dac_clk_p_c_enable_196, cmd_loaded_N_768;
    wire [4:0]dec_bits;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(69[13:21])
    
    wire dac_clk_p_c_enable_349;
    wire [33:0]n14;
    wire [7:0]w_gx_char;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbgenhex.v(80[12:21])
    
    wire n11652;
    wire [33:0]int_word;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(75[14:22])
    
    wire n26742, int_stb;
    
    hbexec wbexec (.wb_odata({wb_odata}), .dac_clk_p_c(dac_clk_p_c), .\iw_word[0] (iw_word[0]), 
           .inc(inc), .dac_clk_p_c_enable_136(dac_clk_p_c_enable_136), .ow_stb(ow_stb), 
           .ow_word({ow_word}), .n29269(n29269), .wb_we(wb_we), .i_cmd_wr(i_cmd_wr), 
           .wb_stb(wb_stb), .n21860(n21860), .wb_cyc(wb_cyc), .newaddr_N_990(newaddr_N_990), 
           .\iw_word[1] (iw_word[1]), .\iw_word[30] (iw_word[30]), .\iw_word[31] (iw_word[31]), 
           .\iw_word[28] (iw_word[28]), .\iw_word[29] (iw_word[29]), .\iw_word[26] (iw_word[26]), 
           .\iw_word[27] (iw_word[27]), .\iw_word[24] (iw_word[24]), .\iw_word[25] (iw_word[25]), 
           .\iw_word[22] (iw_word[22]), .\iw_word[23] (iw_word[23]), .\iw_word[20] (iw_word[20]), 
           .\iw_word[21] (iw_word[21]), .\iw_word[18] (iw_word[18]), .\iw_word[19] (iw_word[19]), 
           .\iw_word[16] (iw_word[16]), .\iw_word[17] (iw_word[17]), .\iw_word[14] (iw_word[14]), 
           .\iw_word[15] (iw_word[15]), .\iw_word[12] (iw_word[12]), .\iw_word[13] (iw_word[13]), 
           .\iw_word[10] (iw_word[10]), .\iw_word[11] (iw_word[11]), .\iw_word[8] (iw_word[8]), 
           .\iw_word[9] (iw_word[9]), .\iw_word[6] (iw_word[6]), .\iw_word[7] (iw_word[7]), 
           .\iw_word[4] (iw_word[4]), .\iw_word[5] (iw_word[5]), .n17206(n17206), 
           .wb_addr({wb_addr}), .\iw_word[3] (iw_word[3]), .GND_net(GND_net), 
           .\iw_word[2] (iw_word[2]), .wb_err(wb_err), .n29268(n29268), 
           .wb_ack(wb_ack), .\wb_idata[0] (\wb_idata[0] ), .\wb_idata[2] (\wb_idata[2] ), 
           .\wb_idata[3] (\wb_idata[3] ), .\wb_idata[4] (\wb_idata[4] ), 
           .\wb_idata[5] (\wb_idata[5] ), .\wb_idata[6] (\wb_idata[6] ), 
           .\wb_idata[7] (\wb_idata[7] ), .\wb_idata[8] (\wb_idata[8] ), 
           .\wb_idata[9] (\wb_idata[9] ), .\wb_idata[10] (\wb_idata[10] ), 
           .\wb_idata[11] (\wb_idata[11] ), .\wb_idata[12] (\wb_idata[12] ), 
           .\wb_idata[13] (\wb_idata[13] ), .\wb_idata[14] (\wb_idata[14] ), 
           .\wb_idata[15] (\wb_idata[15] ), .\wb_idata[16] (\wb_idata[16] ), 
           .\wb_idata[17] (\wb_idata[17] ), .\wb_idata[18] (\wb_idata[18] ), 
           .\wb_idata[19] (\wb_idata[19] ), .\wb_idata[20] (\wb_idata[20] ), 
           .\wb_idata[21] (\wb_idata[21] ), .\wb_idata[22] (\wb_idata[22] ), 
           .\wb_idata[23] (\wb_idata[23] ), .\wb_idata[24] (\wb_idata[24] ), 
           .\wb_idata[25] (\wb_idata[25] ), .\wb_idata[26] (\wb_idata[26] ), 
           .\wb_idata[27] (\wb_idata[27] ), .\wb_idata[28] (\wb_idata[28] ), 
           .\wb_idata[29] (\wb_idata[29] ), .\wb_idata[30] (\wb_idata[30] ), 
           .\wb_idata[31] (\wb_idata[31] ), .n2(n2), .n26716(n26716), 
           .\iw_word[32] (iw_word[32]), .n26715(n26715), .n12635(n12635), 
           .dac_clk_p_c_enable_446(dac_clk_p_c_enable_446)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(105[15] 109[15])
    hbdeword unpackx (.dac_clk_p_c(dac_clk_p_c), .dac_clk_p_c_enable_307(dac_clk_p_c_enable_307), 
            .hb_bits({hb_bits}), .dac_clk_p_c_enable_193(dac_clk_p_c_enable_193), 
            .n29269(n29269), .idl_word({idl_word}), .n29210(n29210), .hb_busy(hb_busy), 
            .w_reset(w_reset), .n26536(n26536), .idl_stb(idl_stb), .n29268(n29268), 
            .nl_busy(nl_busy), .hx_stb(hx_stb)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(127[11] 129[29])
    hbpack packxi (.dac_clk_p_c(dac_clk_p_c), .dac_clk_p_c_enable_380(dac_clk_p_c_enable_380), 
           .n29269(n29269), .iw_word({Open_3, Open_4, Open_5, Open_6, 
           Open_7, Open_8, Open_9, Open_10, Open_11, Open_12, Open_13, 
           Open_14, Open_15, Open_16, Open_17, Open_18, Open_19, 
           Open_20, Open_21, Open_22, Open_23, Open_24, Open_25, 
           Open_26, Open_27, Open_28, Open_29, Open_30, Open_31, 
           Open_32, Open_33, iw_word[2], Open_34, iw_word[0]}), .w_reset(w_reset), 
           .o_pck_stb_N_765(o_pck_stb_N_765), .cmd_loaded(cmd_loaded), .dac_clk_p_c_enable_196(dac_clk_p_c_enable_196), 
           .cmd_loaded_N_768(cmd_loaded_N_768), .\dec_bits[4] (dec_bits[4]), 
           .wb_cyc(wb_cyc), .inc(inc), .n17206(n17206), .\iw_word[32] (iw_word[32]), 
           .\iw_word[31] (iw_word[31]), .\iw_word[30] (iw_word[30]), .\iw_word[29] (iw_word[29]), 
           .\iw_word[28] (iw_word[28]), .\iw_word[27] (iw_word[27]), .\iw_word[26] (iw_word[26]), 
           .\iw_word[25] (iw_word[25]), .\iw_word[24] (iw_word[24]), .\iw_word[23] (iw_word[23]), 
           .\iw_word[22] (iw_word[22]), .\iw_word[21] (iw_word[21]), .\iw_word[20] (iw_word[20]), 
           .\iw_word[19] (iw_word[19]), .\iw_word[18] (iw_word[18]), .\iw_word[17] (iw_word[17]), 
           .\iw_word[16] (iw_word[16]), .\iw_word[15] (iw_word[15]), .\iw_word[14] (iw_word[14]), 
           .\iw_word[13] (iw_word[13]), .\iw_word[12] (iw_word[12]), .\iw_word[11] (iw_word[11]), 
           .\iw_word[10] (iw_word[10]), .\iw_word[9] (iw_word[9]), .\iw_word[8] (iw_word[8]), 
           .\iw_word[7] (iw_word[7]), .\iw_word[6] (iw_word[6]), .\iw_word[5] (iw_word[5]), 
           .\iw_word[4] (iw_word[4]), .\iw_word[3] (iw_word[3]), .\iw_word[1] (iw_word[1]), 
           .\dec_bits[0] (dec_bits[0]), .\dec_bits[1] (dec_bits[1]), .dac_clk_p_c_enable_349(dac_clk_p_c_enable_349), 
           .n26716(n26716), .wb_stb(wb_stb), .dac_clk_p_c_enable_446(dac_clk_p_c_enable_446), 
           .n45(n14[3]), .n46(n14[2]), .n26715(n26715), .i_cmd_wr(i_cmd_wr), 
           .n21860(n21860), .dac_clk_p_c_enable_136(dac_clk_p_c_enable_136), 
           .n29268(n29268), .newaddr_N_990(newaddr_N_990)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(99[9] 100[38])
    hbgenhex genhex (.hb_bits({hb_bits}), .\w_gx_char[0] (w_gx_char[0]), 
            .\w_gx_char[1] (w_gx_char[1]), .\w_gx_char[2] (w_gx_char[2]), 
            .\w_gx_char[3] (w_gx_char[3]), .\w_gx_char[4] (w_gx_char[4]), 
            .\w_gx_char[5] (w_gx_char[5]), .\w_gx_char[6] (w_gx_char[6]), 
            .dac_clk_p_c(dac_clk_p_c), .dac_clk_p_c_enable_307(dac_clk_p_c_enable_307), 
            .GND_net(GND_net), .VCC_net(VCC_net), .hx_stb(hx_stb), .w_reset(w_reset), 
            .hb_busy(hb_busy), .nl_busy(nl_busy), .n29268(n29268), .n26536(n26536), 
            .dac_clk_p_c_enable_193(dac_clk_p_c_enable_193), .n11652(n11652)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(132[11] 133[29])
    hbdechex dechxi (.dac_clk_p_c(dac_clk_p_c), .dec_bits({dec_bits[4], 
            Open_35, Open_36, Open_37, dec_bits[0]}), .w_reset(w_reset), 
            .\rx_data[5] (\rx_data[5] ), .\rx_data[1] (\rx_data[1] ), .rx_stb(rx_stb), 
            .\rx_data[6] (\rx_data[6] ), .\rx_data[3] (\rx_data[3] ), .\rx_data[4] (\rx_data[4] ), 
            .\rx_data[0] (\rx_data[0] ), .\rx_data[2] (\rx_data[2] ), .\dec_bits[1] (dec_bits[1]), 
            .n29269(n29269), .n29268(n29268), .n45(n14[3]), .n46(n14[2]), 
            .dac_clk_p_c_enable_380(dac_clk_p_c_enable_380), .dac_clk_p_c_enable_349(dac_clk_p_c_enable_349), 
            .cmd_loaded(cmd_loaded), .o_pck_stb_N_765(o_pck_stb_N_765), 
            .dac_clk_p_c_enable_196(dac_clk_p_c_enable_196), .cmd_loaded_N_768(cmd_loaded_N_768)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(93[11] 95[30])
    hbnewline addnl (.tx_busy(tx_busy), .o_busy_N_536(o_busy_N_536), .\state[0] (\state[0] ), 
            .n17598(n17598), .dac_clk_p_c(dac_clk_p_c), .n29269(n29269), 
            .w_reset(w_reset), .hx_stb(hx_stb), .nl_busy(nl_busy), .\w_gx_char[2] (w_gx_char[2]), 
            .\w_gx_char[0] (w_gx_char[0]), .n26540(n26540), .\lcl_data[1] (\lcl_data[1] ), 
            .\lcl_data_7__N_511[0] (\lcl_data_7__N_511[0] ), .\lcl_data[4] (\lcl_data[4] ), 
            .\lcl_data_7__N_511[3] (\lcl_data_7__N_511[3] ), .\lcl_data[5] (\lcl_data[5] ), 
            .\lcl_data_7__N_511[4] (\lcl_data_7__N_511[4] ), .\lcl_data[6] (\lcl_data[6] ), 
            .\lcl_data_7__N_511[5] (\lcl_data_7__N_511[5] ), .\lcl_data[7] (\lcl_data[7] ), 
            .\lcl_data_7__N_511[6] (\lcl_data_7__N_511[6] ), .zero_baud_counter(zero_baud_counter), 
            .dac_clk_p_c_enable_321(dac_clk_p_c_enable_321), .\lcl_data[3] (\lcl_data[3] ), 
            .\lcl_data_7__N_511[2] (\lcl_data_7__N_511[2] ), .\lcl_data[2] (\lcl_data[2] ), 
            .\lcl_data_7__N_511[1] (\lcl_data_7__N_511[1] ), .\w_gx_char[4] (w_gx_char[4]), 
            .n29268(n29268), .\w_gx_char[3] (w_gx_char[3]), .\w_gx_char[5] (w_gx_char[5]), 
            .\w_gx_char[1] (w_gx_char[1]), .\w_gx_char[6] (w_gx_char[6]), 
            .n11652(n11652)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(138[12] 139[40])
    hbints addints (.int_word({int_word}), .dac_clk_p_c(dac_clk_p_c), .ow_word({ow_word}), 
           .n29268(n29268), .n26742(n26742), .int_stb(int_stb), .ow_stb(ow_stb), 
           .n29269(n29269)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(114[9] 116[32])
    hbidle addidles (.idl_word({idl_word}), .dac_clk_p_c(dac_clk_p_c), .int_word({int_word}), 
           .hb_busy(hb_busy), .int_stb(int_stb), .idl_stb(idl_stb), .n29268(n29268), 
           .w_reset(w_reset), .n26742(n26742)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(121[9] 123[31])
    
endmodule
//
// Verilog Description of module hbexec
//

module hbexec (wb_odata, dac_clk_p_c, \iw_word[0] , inc, dac_clk_p_c_enable_136, 
            ow_stb, ow_word, n29269, wb_we, i_cmd_wr, wb_stb, n21860, 
            wb_cyc, newaddr_N_990, \iw_word[1] , \iw_word[30] , \iw_word[31] , 
            \iw_word[28] , \iw_word[29] , \iw_word[26] , \iw_word[27] , 
            \iw_word[24] , \iw_word[25] , \iw_word[22] , \iw_word[23] , 
            \iw_word[20] , \iw_word[21] , \iw_word[18] , \iw_word[19] , 
            \iw_word[16] , \iw_word[17] , \iw_word[14] , \iw_word[15] , 
            \iw_word[12] , \iw_word[13] , \iw_word[10] , \iw_word[11] , 
            \iw_word[8] , \iw_word[9] , \iw_word[6] , \iw_word[7] , 
            \iw_word[4] , \iw_word[5] , n17206, wb_addr, \iw_word[3] , 
            GND_net, \iw_word[2] , wb_err, n29268, wb_ack, \wb_idata[0] , 
            \wb_idata[2] , \wb_idata[3] , \wb_idata[4] , \wb_idata[5] , 
            \wb_idata[6] , \wb_idata[7] , \wb_idata[8] , \wb_idata[9] , 
            \wb_idata[10] , \wb_idata[11] , \wb_idata[12] , \wb_idata[13] , 
            \wb_idata[14] , \wb_idata[15] , \wb_idata[16] , \wb_idata[17] , 
            \wb_idata[18] , \wb_idata[19] , \wb_idata[20] , \wb_idata[21] , 
            \wb_idata[22] , \wb_idata[23] , \wb_idata[24] , \wb_idata[25] , 
            \wb_idata[26] , \wb_idata[27] , \wb_idata[28] , \wb_idata[29] , 
            \wb_idata[30] , \wb_idata[31] , n2, n26716, \iw_word[32] , 
            n26715, n12635, dac_clk_p_c_enable_446) /* synthesis syn_module_defined=1 */ ;
    output [31:0]wb_odata;
    input dac_clk_p_c;
    input \iw_word[0] ;
    output inc;
    input dac_clk_p_c_enable_136;
    output ow_stb;
    output [33:0]ow_word;
    input n29269;
    output wb_we;
    input i_cmd_wr;
    output wb_stb;
    input n21860;
    output wb_cyc;
    input newaddr_N_990;
    input \iw_word[1] ;
    input \iw_word[30] ;
    input \iw_word[31] ;
    input \iw_word[28] ;
    input \iw_word[29] ;
    input \iw_word[26] ;
    input \iw_word[27] ;
    input \iw_word[24] ;
    input \iw_word[25] ;
    input \iw_word[22] ;
    input \iw_word[23] ;
    input \iw_word[20] ;
    input \iw_word[21] ;
    input \iw_word[18] ;
    input \iw_word[19] ;
    input \iw_word[16] ;
    input \iw_word[17] ;
    input \iw_word[14] ;
    input \iw_word[15] ;
    input \iw_word[12] ;
    input \iw_word[13] ;
    input \iw_word[10] ;
    input \iw_word[11] ;
    input \iw_word[8] ;
    input \iw_word[9] ;
    input \iw_word[6] ;
    input \iw_word[7] ;
    input \iw_word[4] ;
    input \iw_word[5] ;
    input n17206;
    output [29:0]wb_addr;
    input \iw_word[3] ;
    input GND_net;
    input \iw_word[2] ;
    input wb_err;
    input n29268;
    input wb_ack;
    input \wb_idata[0] ;
    input \wb_idata[2] ;
    input \wb_idata[3] ;
    input \wb_idata[4] ;
    input \wb_idata[5] ;
    input \wb_idata[6] ;
    input \wb_idata[7] ;
    input \wb_idata[8] ;
    input \wb_idata[9] ;
    input \wb_idata[10] ;
    input \wb_idata[11] ;
    input \wb_idata[12] ;
    input \wb_idata[13] ;
    input \wb_idata[14] ;
    input \wb_idata[15] ;
    input \wb_idata[16] ;
    input \wb_idata[17] ;
    input \wb_idata[18] ;
    input \wb_idata[19] ;
    input \wb_idata[20] ;
    input \wb_idata[21] ;
    input \wb_idata[22] ;
    input \wb_idata[23] ;
    input \wb_idata[24] ;
    input \wb_idata[25] ;
    input \wb_idata[26] ;
    input \wb_idata[27] ;
    input \wb_idata[28] ;
    input \wb_idata[29] ;
    input \wb_idata[30] ;
    input \wb_idata[31] ;
    output n2;
    input n26716;
    input \iw_word[32] ;
    input n26715;
    input n12635;
    input dac_clk_p_c_enable_446;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(29[49:58])
    
    wire i_cmd_word_0__N_995, n8903, o_rsp_stb_N_987;
    wire [33:0]n338;
    wire [33:0]o_rsp_word_33__N_951;
    
    wire o_cmd_busy_N_931, n19567, newaddr, n17464, n17151, n17149;
    wire [29:0]n125;
    
    wire n17463, n17155, n17153, n17462, n17159, n17157, n17461, 
        n17163, n17161, n17460, n17167, n17165, n17459, n17171, 
        n17169, n17458, n17175, n17173, n17457, n17179, n17177, 
        n17456, n17183, n17181, n17455, n17187, n17185, n17454, 
        n17191, n17189, n17453, n17195, n17193, n17452, n17199, 
        n17197, n17451, n17203, n17201, n17450, n17205;
    wire [32:0]n2123;
    
    wire n3, n20131, o_cmd_busy_N_941, o_cmd_busy_N_933, dac_clk_p_c_enable_414;
    
    FD1S3AX o_wb_data_i0 (.D(\iw_word[0] ), .CK(dac_clk_p_c), .Q(wb_odata[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i0.GSR = "DISABLED";
    FD1P3AX inc_71 (.D(i_cmd_word_0__N_995), .SP(dac_clk_p_c_enable_136), 
            .CK(dac_clk_p_c), .Q(inc)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(192[9] 236[5])
    defparam inc_71.GSR = "DISABLED";
    FD1S3JX o_rsp_stb_74 (.D(o_rsp_stb_N_987), .CK(dac_clk_p_c), .PD(n8903), 
            .Q(ow_stb)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_stb_74.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i0 (.D(n338[0]), .CK(dac_clk_p_c), .CD(n8903), 
            .Q(ow_word[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i0.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i2 (.D(n338[2]), .CK(dac_clk_p_c), .CD(n8903), 
            .Q(ow_word[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i2.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i3 (.D(n338[3]), .CK(dac_clk_p_c), .CD(n8903), 
            .Q(ow_word[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i3.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i4 (.D(n338[4]), .CK(dac_clk_p_c), .CD(n8903), 
            .Q(ow_word[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i4.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i5 (.D(n338[5]), .CK(dac_clk_p_c), .CD(n8903), 
            .Q(ow_word[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i5.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i6 (.D(n338[6]), .CK(dac_clk_p_c), .CD(n8903), 
            .Q(ow_word[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i6.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i7 (.D(n338[7]), .CK(dac_clk_p_c), .CD(n8903), 
            .Q(ow_word[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i7.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i8 (.D(n338[8]), .CK(dac_clk_p_c), .CD(n8903), 
            .Q(ow_word[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i8.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i9 (.D(n338[9]), .CK(dac_clk_p_c), .CD(n8903), 
            .Q(ow_word[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i9.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i10 (.D(n338[10]), .CK(dac_clk_p_c), .CD(n8903), 
            .Q(ow_word[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i10.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i11 (.D(n338[11]), .CK(dac_clk_p_c), .CD(n8903), 
            .Q(ow_word[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i11.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i12 (.D(n338[12]), .CK(dac_clk_p_c), .CD(n8903), 
            .Q(ow_word[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i12.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i13 (.D(n338[13]), .CK(dac_clk_p_c), .CD(n8903), 
            .Q(ow_word[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i13.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i14 (.D(n338[14]), .CK(dac_clk_p_c), .CD(n8903), 
            .Q(ow_word[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i14.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i15 (.D(n338[15]), .CK(dac_clk_p_c), .CD(n8903), 
            .Q(ow_word[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i15.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i16 (.D(n338[16]), .CK(dac_clk_p_c), .CD(n8903), 
            .Q(ow_word[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i16.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i17 (.D(n338[17]), .CK(dac_clk_p_c), .CD(n8903), 
            .Q(ow_word[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i17.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i18 (.D(n338[18]), .CK(dac_clk_p_c), .CD(n8903), 
            .Q(ow_word[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i18.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i19 (.D(n338[19]), .CK(dac_clk_p_c), .CD(n8903), 
            .Q(ow_word[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i19.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i20 (.D(n338[20]), .CK(dac_clk_p_c), .CD(n8903), 
            .Q(ow_word[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i20.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i21 (.D(n338[21]), .CK(dac_clk_p_c), .CD(n8903), 
            .Q(ow_word[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i21.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i22 (.D(n338[22]), .CK(dac_clk_p_c), .CD(n8903), 
            .Q(ow_word[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i22.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i23 (.D(n338[23]), .CK(dac_clk_p_c), .CD(n8903), 
            .Q(ow_word[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i23.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i24 (.D(n338[24]), .CK(dac_clk_p_c), .CD(n8903), 
            .Q(ow_word[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i24.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i25 (.D(n338[25]), .CK(dac_clk_p_c), .CD(n8903), 
            .Q(ow_word[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i25.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i26 (.D(n338[26]), .CK(dac_clk_p_c), .CD(n8903), 
            .Q(ow_word[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i26.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i27 (.D(n338[27]), .CK(dac_clk_p_c), .CD(n8903), 
            .Q(ow_word[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i27.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i28 (.D(n338[28]), .CK(dac_clk_p_c), .CD(n8903), 
            .Q(ow_word[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i28.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i29 (.D(o_rsp_word_33__N_951[29]), .CK(dac_clk_p_c), 
            .CD(n29269), .Q(ow_word[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i29.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i30 (.D(n338[30]), .CK(dac_clk_p_c), .CD(n8903), 
            .Q(ow_word[30])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i30.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i31 (.D(n338[31]), .CK(dac_clk_p_c), .CD(n8903), 
            .Q(ow_word[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i31.GSR = "DISABLED";
    FD1S3JX o_rsp_word_i32 (.D(n338[32]), .CK(dac_clk_p_c), .PD(n8903), 
            .Q(ow_word[32])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i32.GSR = "DISABLED";
    FD1S3JX o_rsp_word_i33 (.D(o_cmd_busy_N_931), .CK(dac_clk_p_c), .PD(n8903), 
            .Q(ow_word[33])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i33.GSR = "DISABLED";
    FD1P3AX o_wb_we_69 (.D(i_cmd_wr), .SP(o_cmd_busy_N_931), .CK(dac_clk_p_c), 
            .Q(wb_we)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(184[9] 186[26])
    defparam o_wb_we_69.GSR = "DISABLED";
    FD1P3IX o_wb_stb_68 (.D(n21860), .SP(o_cmd_busy_N_931), .CD(n19567), 
            .CK(dac_clk_p_c), .Q(wb_stb)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(121[9] 168[5])
    defparam o_wb_stb_68.GSR = "DISABLED";
    FD1S3IX newaddr_72 (.D(newaddr_N_990), .CK(dac_clk_p_c), .CD(wb_cyc), 
            .Q(newaddr)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(192[9] 236[5])
    defparam newaddr_72.GSR = "DISABLED";
    CCU2D o_wb_addr_546_add_4_31 (.A0(n17151), .B0(\iw_word[1] ), .C0(dac_clk_p_c_enable_136), 
          .D0(\iw_word[30] ), .A1(n17149), .B1(\iw_word[1] ), .C1(dac_clk_p_c_enable_136), 
          .D1(\iw_word[31] ), .CIN(n17464), .S0(n125[28]), .S1(n125[29]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_546_add_4_31.INIT0 = 16'h5aaa;
    defparam o_wb_addr_546_add_4_31.INIT1 = 16'h5aaa;
    defparam o_wb_addr_546_add_4_31.INJECT1_0 = "NO";
    defparam o_wb_addr_546_add_4_31.INJECT1_1 = "NO";
    CCU2D o_wb_addr_546_add_4_29 (.A0(n17155), .B0(\iw_word[1] ), .C0(dac_clk_p_c_enable_136), 
          .D0(\iw_word[28] ), .A1(n17153), .B1(\iw_word[1] ), .C1(dac_clk_p_c_enable_136), 
          .D1(\iw_word[29] ), .CIN(n17463), .COUT(n17464), .S0(n125[26]), 
          .S1(n125[27]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_546_add_4_29.INIT0 = 16'h5aaa;
    defparam o_wb_addr_546_add_4_29.INIT1 = 16'h5aaa;
    defparam o_wb_addr_546_add_4_29.INJECT1_0 = "NO";
    defparam o_wb_addr_546_add_4_29.INJECT1_1 = "NO";
    CCU2D o_wb_addr_546_add_4_27 (.A0(n17159), .B0(\iw_word[1] ), .C0(dac_clk_p_c_enable_136), 
          .D0(\iw_word[26] ), .A1(n17157), .B1(\iw_word[1] ), .C1(dac_clk_p_c_enable_136), 
          .D1(\iw_word[27] ), .CIN(n17462), .COUT(n17463), .S0(n125[24]), 
          .S1(n125[25]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_546_add_4_27.INIT0 = 16'h5aaa;
    defparam o_wb_addr_546_add_4_27.INIT1 = 16'h5aaa;
    defparam o_wb_addr_546_add_4_27.INJECT1_0 = "NO";
    defparam o_wb_addr_546_add_4_27.INJECT1_1 = "NO";
    CCU2D o_wb_addr_546_add_4_25 (.A0(n17163), .B0(\iw_word[1] ), .C0(dac_clk_p_c_enable_136), 
          .D0(\iw_word[24] ), .A1(n17161), .B1(\iw_word[1] ), .C1(dac_clk_p_c_enable_136), 
          .D1(\iw_word[25] ), .CIN(n17461), .COUT(n17462), .S0(n125[22]), 
          .S1(n125[23]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_546_add_4_25.INIT0 = 16'h5aaa;
    defparam o_wb_addr_546_add_4_25.INIT1 = 16'h5aaa;
    defparam o_wb_addr_546_add_4_25.INJECT1_0 = "NO";
    defparam o_wb_addr_546_add_4_25.INJECT1_1 = "NO";
    CCU2D o_wb_addr_546_add_4_23 (.A0(n17167), .B0(\iw_word[1] ), .C0(dac_clk_p_c_enable_136), 
          .D0(\iw_word[22] ), .A1(n17165), .B1(\iw_word[1] ), .C1(dac_clk_p_c_enable_136), 
          .D1(\iw_word[23] ), .CIN(n17460), .COUT(n17461), .S0(n125[20]), 
          .S1(n125[21]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_546_add_4_23.INIT0 = 16'h5aaa;
    defparam o_wb_addr_546_add_4_23.INIT1 = 16'h5aaa;
    defparam o_wb_addr_546_add_4_23.INJECT1_0 = "NO";
    defparam o_wb_addr_546_add_4_23.INJECT1_1 = "NO";
    CCU2D o_wb_addr_546_add_4_21 (.A0(n17171), .B0(\iw_word[1] ), .C0(dac_clk_p_c_enable_136), 
          .D0(\iw_word[20] ), .A1(n17169), .B1(\iw_word[1] ), .C1(dac_clk_p_c_enable_136), 
          .D1(\iw_word[21] ), .CIN(n17459), .COUT(n17460), .S0(n125[18]), 
          .S1(n125[19]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_546_add_4_21.INIT0 = 16'h5aaa;
    defparam o_wb_addr_546_add_4_21.INIT1 = 16'h5aaa;
    defparam o_wb_addr_546_add_4_21.INJECT1_0 = "NO";
    defparam o_wb_addr_546_add_4_21.INJECT1_1 = "NO";
    CCU2D o_wb_addr_546_add_4_19 (.A0(n17175), .B0(\iw_word[1] ), .C0(dac_clk_p_c_enable_136), 
          .D0(\iw_word[18] ), .A1(n17173), .B1(\iw_word[1] ), .C1(dac_clk_p_c_enable_136), 
          .D1(\iw_word[19] ), .CIN(n17458), .COUT(n17459), .S0(n125[16]), 
          .S1(n125[17]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_546_add_4_19.INIT0 = 16'h5aaa;
    defparam o_wb_addr_546_add_4_19.INIT1 = 16'h5aaa;
    defparam o_wb_addr_546_add_4_19.INJECT1_0 = "NO";
    defparam o_wb_addr_546_add_4_19.INJECT1_1 = "NO";
    CCU2D o_wb_addr_546_add_4_17 (.A0(n17179), .B0(\iw_word[1] ), .C0(dac_clk_p_c_enable_136), 
          .D0(\iw_word[16] ), .A1(n17177), .B1(\iw_word[1] ), .C1(dac_clk_p_c_enable_136), 
          .D1(\iw_word[17] ), .CIN(n17457), .COUT(n17458), .S0(n125[14]), 
          .S1(n125[15]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_546_add_4_17.INIT0 = 16'h5aaa;
    defparam o_wb_addr_546_add_4_17.INIT1 = 16'h5aaa;
    defparam o_wb_addr_546_add_4_17.INJECT1_0 = "NO";
    defparam o_wb_addr_546_add_4_17.INJECT1_1 = "NO";
    CCU2D o_wb_addr_546_add_4_15 (.A0(n17183), .B0(\iw_word[1] ), .C0(dac_clk_p_c_enable_136), 
          .D0(\iw_word[14] ), .A1(n17181), .B1(\iw_word[1] ), .C1(dac_clk_p_c_enable_136), 
          .D1(\iw_word[15] ), .CIN(n17456), .COUT(n17457), .S0(n125[12]), 
          .S1(n125[13]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_546_add_4_15.INIT0 = 16'h5aaa;
    defparam o_wb_addr_546_add_4_15.INIT1 = 16'h5aaa;
    defparam o_wb_addr_546_add_4_15.INJECT1_0 = "NO";
    defparam o_wb_addr_546_add_4_15.INJECT1_1 = "NO";
    CCU2D o_wb_addr_546_add_4_13 (.A0(n17187), .B0(\iw_word[1] ), .C0(dac_clk_p_c_enable_136), 
          .D0(\iw_word[12] ), .A1(n17185), .B1(\iw_word[1] ), .C1(dac_clk_p_c_enable_136), 
          .D1(\iw_word[13] ), .CIN(n17455), .COUT(n17456), .S0(n125[10]), 
          .S1(n125[11]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_546_add_4_13.INIT0 = 16'h5aaa;
    defparam o_wb_addr_546_add_4_13.INIT1 = 16'h5aaa;
    defparam o_wb_addr_546_add_4_13.INJECT1_0 = "NO";
    defparam o_wb_addr_546_add_4_13.INJECT1_1 = "NO";
    CCU2D o_wb_addr_546_add_4_11 (.A0(n17191), .B0(\iw_word[1] ), .C0(dac_clk_p_c_enable_136), 
          .D0(\iw_word[10] ), .A1(n17189), .B1(\iw_word[1] ), .C1(dac_clk_p_c_enable_136), 
          .D1(\iw_word[11] ), .CIN(n17454), .COUT(n17455), .S0(n125[8]), 
          .S1(n125[9]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_546_add_4_11.INIT0 = 16'h5aaa;
    defparam o_wb_addr_546_add_4_11.INIT1 = 16'h5aaa;
    defparam o_wb_addr_546_add_4_11.INJECT1_0 = "NO";
    defparam o_wb_addr_546_add_4_11.INJECT1_1 = "NO";
    CCU2D o_wb_addr_546_add_4_9 (.A0(n17195), .B0(\iw_word[1] ), .C0(dac_clk_p_c_enable_136), 
          .D0(\iw_word[8] ), .A1(n17193), .B1(\iw_word[1] ), .C1(dac_clk_p_c_enable_136), 
          .D1(\iw_word[9] ), .CIN(n17453), .COUT(n17454), .S0(n125[6]), 
          .S1(n125[7]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_546_add_4_9.INIT0 = 16'h5aaa;
    defparam o_wb_addr_546_add_4_9.INIT1 = 16'h5aaa;
    defparam o_wb_addr_546_add_4_9.INJECT1_0 = "NO";
    defparam o_wb_addr_546_add_4_9.INJECT1_1 = "NO";
    CCU2D o_wb_addr_546_add_4_7 (.A0(n17199), .B0(\iw_word[1] ), .C0(dac_clk_p_c_enable_136), 
          .D0(\iw_word[6] ), .A1(n17197), .B1(\iw_word[1] ), .C1(dac_clk_p_c_enable_136), 
          .D1(\iw_word[7] ), .CIN(n17452), .COUT(n17453), .S0(n125[4]), 
          .S1(n125[5]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_546_add_4_7.INIT0 = 16'h5aaa;
    defparam o_wb_addr_546_add_4_7.INIT1 = 16'h5aaa;
    defparam o_wb_addr_546_add_4_7.INJECT1_0 = "NO";
    defparam o_wb_addr_546_add_4_7.INJECT1_1 = "NO";
    CCU2D o_wb_addr_546_add_4_5 (.A0(n17203), .B0(\iw_word[1] ), .C0(dac_clk_p_c_enable_136), 
          .D0(\iw_word[4] ), .A1(n17201), .B1(\iw_word[1] ), .C1(dac_clk_p_c_enable_136), 
          .D1(\iw_word[5] ), .CIN(n17451), .COUT(n17452), .S0(n125[2]), 
          .S1(n125[3]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_546_add_4_5.INIT0 = 16'h5aaa;
    defparam o_wb_addr_546_add_4_5.INIT1 = 16'h5aaa;
    defparam o_wb_addr_546_add_4_5.INJECT1_0 = "NO";
    defparam o_wb_addr_546_add_4_5.INJECT1_1 = "NO";
    CCU2D o_wb_addr_546_add_4_3 (.A0(n17206), .B0(dac_clk_p_c_enable_136), 
          .C0(\iw_word[1] ), .D0(wb_addr[0]), .A1(n17205), .B1(\iw_word[1] ), 
          .C1(dac_clk_p_c_enable_136), .D1(\iw_word[3] ), .CIN(n17450), 
          .COUT(n17451), .S0(n125[0]), .S1(n125[1]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_546_add_4_3.INIT0 = 16'h59aa;
    defparam o_wb_addr_546_add_4_3.INIT1 = 16'h5aaa;
    defparam o_wb_addr_546_add_4_3.INJECT1_0 = "NO";
    defparam o_wb_addr_546_add_4_3.INJECT1_1 = "NO";
    CCU2D o_wb_addr_546_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\iw_word[1] ), .B1(dac_clk_p_c_enable_136), 
          .C1(GND_net), .D1(GND_net), .COUT(n17450));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_546_add_4_1.INIT0 = 16'hF000;
    defparam o_wb_addr_546_add_4_1.INIT1 = 16'hffff;
    defparam o_wb_addr_546_add_4_1.INJECT1_0 = "NO";
    defparam o_wb_addr_546_add_4_1.INJECT1_1 = "NO";
    FD1S3AX o_wb_data_i31 (.D(\iw_word[31] ), .CK(dac_clk_p_c), .Q(wb_odata[31])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i31.GSR = "DISABLED";
    FD1S3AX o_wb_data_i30 (.D(\iw_word[30] ), .CK(dac_clk_p_c), .Q(wb_odata[30])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i30.GSR = "DISABLED";
    FD1S3AX o_wb_data_i29 (.D(\iw_word[29] ), .CK(dac_clk_p_c), .Q(wb_odata[29])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i29.GSR = "DISABLED";
    FD1S3AX o_wb_data_i28 (.D(\iw_word[28] ), .CK(dac_clk_p_c), .Q(wb_odata[28])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i28.GSR = "DISABLED";
    FD1S3AX o_wb_data_i27 (.D(\iw_word[27] ), .CK(dac_clk_p_c), .Q(wb_odata[27])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i27.GSR = "DISABLED";
    FD1S3AX o_wb_data_i26 (.D(\iw_word[26] ), .CK(dac_clk_p_c), .Q(wb_odata[26])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i26.GSR = "DISABLED";
    FD1S3AX o_wb_data_i25 (.D(\iw_word[25] ), .CK(dac_clk_p_c), .Q(wb_odata[25])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i25.GSR = "DISABLED";
    FD1S3AX o_wb_data_i24 (.D(\iw_word[24] ), .CK(dac_clk_p_c), .Q(wb_odata[24])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i24.GSR = "DISABLED";
    FD1S3AX o_wb_data_i23 (.D(\iw_word[23] ), .CK(dac_clk_p_c), .Q(wb_odata[23])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i23.GSR = "DISABLED";
    FD1S3AX o_wb_data_i22 (.D(\iw_word[22] ), .CK(dac_clk_p_c), .Q(wb_odata[22])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i22.GSR = "DISABLED";
    FD1S3AX o_wb_data_i21 (.D(\iw_word[21] ), .CK(dac_clk_p_c), .Q(wb_odata[21])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i21.GSR = "DISABLED";
    FD1S3AX o_wb_data_i20 (.D(\iw_word[20] ), .CK(dac_clk_p_c), .Q(wb_odata[20])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i20.GSR = "DISABLED";
    FD1S3AX o_wb_data_i19 (.D(\iw_word[19] ), .CK(dac_clk_p_c), .Q(wb_odata[19])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i19.GSR = "DISABLED";
    FD1S3AX o_wb_data_i18 (.D(\iw_word[18] ), .CK(dac_clk_p_c), .Q(wb_odata[18])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i18.GSR = "DISABLED";
    FD1S3AX o_wb_data_i17 (.D(\iw_word[17] ), .CK(dac_clk_p_c), .Q(wb_odata[17])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i17.GSR = "DISABLED";
    FD1S3AX o_wb_data_i16 (.D(\iw_word[16] ), .CK(dac_clk_p_c), .Q(wb_odata[16])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i16.GSR = "DISABLED";
    FD1S3AX o_wb_data_i15 (.D(\iw_word[15] ), .CK(dac_clk_p_c), .Q(wb_odata[15])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i15.GSR = "DISABLED";
    FD1S3AX o_wb_data_i14 (.D(\iw_word[14] ), .CK(dac_clk_p_c), .Q(wb_odata[14])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i14.GSR = "DISABLED";
    FD1S3AX o_wb_data_i13 (.D(\iw_word[13] ), .CK(dac_clk_p_c), .Q(wb_odata[13])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i13.GSR = "DISABLED";
    FD1S3AX o_wb_data_i12 (.D(\iw_word[12] ), .CK(dac_clk_p_c), .Q(wb_odata[12])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i12.GSR = "DISABLED";
    FD1S3AX o_wb_data_i11 (.D(\iw_word[11] ), .CK(dac_clk_p_c), .Q(wb_odata[11])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i11.GSR = "DISABLED";
    FD1S3AX o_wb_data_i10 (.D(\iw_word[10] ), .CK(dac_clk_p_c), .Q(wb_odata[10])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i10.GSR = "DISABLED";
    FD1S3AX o_wb_data_i9 (.D(\iw_word[9] ), .CK(dac_clk_p_c), .Q(wb_odata[9])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i9.GSR = "DISABLED";
    FD1S3AX o_wb_data_i8 (.D(\iw_word[8] ), .CK(dac_clk_p_c), .Q(wb_odata[8])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i8.GSR = "DISABLED";
    FD1S3AX o_wb_data_i7 (.D(\iw_word[7] ), .CK(dac_clk_p_c), .Q(wb_odata[7])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i7.GSR = "DISABLED";
    FD1S3AX o_wb_data_i6 (.D(\iw_word[6] ), .CK(dac_clk_p_c), .Q(wb_odata[6])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i6.GSR = "DISABLED";
    FD1S3AX o_wb_data_i5 (.D(\iw_word[5] ), .CK(dac_clk_p_c), .Q(wb_odata[5])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i5.GSR = "DISABLED";
    FD1S3AX o_wb_data_i4 (.D(\iw_word[4] ), .CK(dac_clk_p_c), .Q(wb_odata[4])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i4.GSR = "DISABLED";
    FD1S3AX o_wb_data_i3 (.D(\iw_word[3] ), .CK(dac_clk_p_c), .Q(wb_odata[3])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i3.GSR = "DISABLED";
    FD1S3AX o_wb_data_i2 (.D(\iw_word[2] ), .CK(dac_clk_p_c), .Q(wb_odata[2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i2.GSR = "DISABLED";
    FD1S3AX o_wb_data_i1 (.D(\iw_word[1] ), .CK(dac_clk_p_c), .Q(wb_odata[1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i1.GSR = "DISABLED";
    LUT4 i_cmd_word_0__I_0_1_lut (.A(\iw_word[0] ), .Z(i_cmd_word_0__N_995)) /* synthesis lut_function=(!(A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(214[11:25])
    defparam i_cmd_word_0__I_0_1_lut.init = 16'h5555;
    LUT4 i6522_2_lut (.A(wb_err), .B(n29268), .Z(n8903)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(283[11] 309[5])
    defparam i6522_2_lut.init = 16'heeee;
    LUT4 newaddr_I_0_3_lut (.A(newaddr), .B(wb_ack), .C(wb_cyc), .Z(o_rsp_stb_N_987)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam newaddr_I_0_3_lut.init = 16'hcaca;
    LUT4 mux_59_i1_4_lut (.A(inc), .B(\wb_idata[0] ), .C(wb_cyc), .D(wb_we), 
         .Z(n338[0])) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A (B (C (D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i1_4_lut.init = 16'h05c5;
    LUT4 mux_59_i3_4_lut (.A(wb_addr[0]), .B(\wb_idata[2] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[2])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i3_4_lut.init = 16'h0aca;
    LUT4 mux_59_i4_4_lut (.A(wb_addr[1]), .B(\wb_idata[3] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[3])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i4_4_lut.init = 16'h0aca;
    LUT4 mux_59_i5_4_lut (.A(wb_addr[2]), .B(\wb_idata[4] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[4])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i5_4_lut.init = 16'h0aca;
    LUT4 mux_59_i6_4_lut (.A(wb_addr[3]), .B(\wb_idata[5] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[5])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i6_4_lut.init = 16'h0aca;
    LUT4 mux_59_i7_4_lut (.A(wb_addr[4]), .B(\wb_idata[6] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[6])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i7_4_lut.init = 16'h0aca;
    LUT4 mux_59_i8_4_lut (.A(wb_addr[5]), .B(\wb_idata[7] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[7])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i8_4_lut.init = 16'h0aca;
    LUT4 mux_59_i9_4_lut (.A(wb_addr[6]), .B(\wb_idata[8] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[8])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i9_4_lut.init = 16'h0aca;
    LUT4 mux_59_i10_4_lut (.A(wb_addr[7]), .B(\wb_idata[9] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[9])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i10_4_lut.init = 16'h0aca;
    LUT4 mux_59_i11_4_lut (.A(wb_addr[8]), .B(\wb_idata[10] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[10])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i11_4_lut.init = 16'h0aca;
    LUT4 mux_59_i12_4_lut (.A(wb_addr[9]), .B(\wb_idata[11] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[11])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i12_4_lut.init = 16'h0aca;
    LUT4 mux_59_i13_4_lut (.A(wb_addr[10]), .B(\wb_idata[12] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[12])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i13_4_lut.init = 16'h0aca;
    LUT4 mux_59_i14_4_lut (.A(wb_addr[11]), .B(\wb_idata[13] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[13])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i14_4_lut.init = 16'h0aca;
    LUT4 mux_59_i15_4_lut (.A(wb_addr[12]), .B(\wb_idata[14] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[14])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i15_4_lut.init = 16'h0aca;
    LUT4 mux_59_i16_4_lut (.A(wb_addr[13]), .B(\wb_idata[15] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[15])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i16_4_lut.init = 16'h0aca;
    LUT4 mux_59_i17_4_lut (.A(wb_addr[14]), .B(\wb_idata[16] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[16])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i17_4_lut.init = 16'h0aca;
    LUT4 mux_59_i18_4_lut (.A(wb_addr[15]), .B(\wb_idata[17] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[17])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i18_4_lut.init = 16'h0aca;
    LUT4 mux_59_i19_4_lut (.A(wb_addr[16]), .B(\wb_idata[18] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[18])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i19_4_lut.init = 16'h0aca;
    LUT4 mux_59_i20_4_lut (.A(wb_addr[17]), .B(\wb_idata[19] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[19])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i20_4_lut.init = 16'h0aca;
    LUT4 mux_59_i21_4_lut (.A(wb_addr[18]), .B(\wb_idata[20] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[20])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i21_4_lut.init = 16'h0aca;
    LUT4 mux_59_i22_4_lut (.A(wb_addr[19]), .B(\wb_idata[21] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[21])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i22_4_lut.init = 16'h0aca;
    LUT4 mux_59_i23_4_lut (.A(wb_addr[20]), .B(\wb_idata[22] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[22])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i23_4_lut.init = 16'h0aca;
    LUT4 mux_59_i24_4_lut (.A(wb_addr[21]), .B(\wb_idata[23] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[23])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i24_4_lut.init = 16'h0aca;
    LUT4 mux_59_i25_4_lut (.A(wb_addr[22]), .B(\wb_idata[24] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[24])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i25_4_lut.init = 16'h0aca;
    LUT4 mux_59_i26_4_lut (.A(wb_addr[23]), .B(\wb_idata[25] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[25])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i26_4_lut.init = 16'h0aca;
    LUT4 mux_59_i27_4_lut (.A(wb_addr[24]), .B(\wb_idata[26] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[26])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i27_4_lut.init = 16'h0aca;
    LUT4 mux_59_i28_4_lut (.A(wb_addr[25]), .B(\wb_idata[27] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[27])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i28_4_lut.init = 16'h0aca;
    LUT4 mux_59_i29_4_lut (.A(wb_addr[26]), .B(\wb_idata[28] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[28])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i29_4_lut.init = 16'h0aca;
    LUT4 i11311_4_lut (.A(wb_addr[27]), .B(wb_err), .C(n2123[29]), .D(wb_cyc), 
         .Z(o_rsp_word_33__N_951[29])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(287[11] 309[5])
    defparam i11311_4_lut.init = 16'hfcee;
    LUT4 i11373_2_lut (.A(\wb_idata[29] ), .B(wb_we), .Z(n2123[29])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(299[4:47])
    defparam i11373_2_lut.init = 16'h2222;
    LUT4 mux_59_i31_4_lut (.A(wb_addr[28]), .B(\wb_idata[30] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[30])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i31_4_lut.init = 16'h0aca;
    LUT4 mux_59_i32_4_lut (.A(wb_addr[29]), .B(\wb_idata[31] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[31])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i32_4_lut.init = 16'h0aca;
    LUT4 i11317_2_lut (.A(wb_we), .B(wb_cyc), .Z(n338[32])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam i11317_2_lut.init = 16'h8888;
    LUT4 o_cmd_busy_I_0_1_lut (.A(wb_cyc), .Z(o_cmd_busy_N_931)) /* synthesis lut_function=(!(A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(194[21:34])
    defparam o_cmd_busy_I_0_1_lut.init = 16'h5555;
    LUT4 i2_1_lut (.A(wb_stb), .Z(n2)) /* synthesis lut_function=(!(A)) */ ;
    defparam i2_1_lut.init = 16'h5555;
    LUT4 i15453_2_lut (.A(wb_addr[28]), .B(n3), .Z(n17151)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15453_2_lut.init = 16'h8888;
    LUT4 i15454_2_lut (.A(wb_addr[29]), .B(n3), .Z(n17149)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15454_2_lut.init = 16'h8888;
    LUT4 i1_4_lut (.A(\iw_word[1] ), .B(n26716), .C(wb_cyc), .D(\iw_word[32] ), 
         .Z(n3)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;
    defparam i1_4_lut.init = 16'hfffb;
    LUT4 i15447_2_lut (.A(wb_addr[26]), .B(n3), .Z(n17155)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15447_2_lut.init = 16'h8888;
    LUT4 i15452_2_lut (.A(wb_addr[27]), .B(n3), .Z(n17153)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15452_2_lut.init = 16'h8888;
    LUT4 i15445_2_lut (.A(wb_addr[24]), .B(n3), .Z(n17159)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15445_2_lut.init = 16'h8888;
    LUT4 i15446_2_lut (.A(wb_addr[25]), .B(n3), .Z(n17157)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15446_2_lut.init = 16'h8888;
    LUT4 i15436_2_lut (.A(wb_addr[22]), .B(n3), .Z(n17163)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15436_2_lut.init = 16'h8888;
    LUT4 i15440_2_lut (.A(wb_addr[23]), .B(n3), .Z(n17161)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15440_2_lut.init = 16'h8888;
    LUT4 i15451_2_lut (.A(wb_addr[20]), .B(n3), .Z(n17167)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15451_2_lut.init = 16'h8888;
    LUT4 i15415_2_lut (.A(wb_addr[21]), .B(n3), .Z(n17165)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15415_2_lut.init = 16'h8888;
    LUT4 i15404_2_lut (.A(wb_addr[18]), .B(n3), .Z(n17171)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15404_2_lut.init = 16'h8888;
    LUT4 i15414_2_lut (.A(wb_addr[19]), .B(n3), .Z(n17169)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15414_2_lut.init = 16'h8888;
    LUT4 i15422_2_lut (.A(wb_addr[16]), .B(n3), .Z(n17175)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15422_2_lut.init = 16'h8888;
    LUT4 i15449_2_lut (.A(wb_addr[17]), .B(n3), .Z(n17173)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15449_2_lut.init = 16'h8888;
    LUT4 i15412_2_lut (.A(wb_addr[14]), .B(n3), .Z(n17179)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15412_2_lut.init = 16'h8888;
    LUT4 i15421_2_lut (.A(wb_addr[15]), .B(n3), .Z(n17177)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15421_2_lut.init = 16'h8888;
    LUT4 i15405_2_lut (.A(wb_addr[12]), .B(n3), .Z(n17183)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15405_2_lut.init = 16'h8888;
    LUT4 i15406_2_lut (.A(wb_addr[13]), .B(n3), .Z(n17181)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15406_2_lut.init = 16'h8888;
    LUT4 i15402_2_lut (.A(wb_addr[10]), .B(n3), .Z(n17187)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15402_2_lut.init = 16'h8888;
    LUT4 i15403_2_lut (.A(wb_addr[11]), .B(n3), .Z(n17185)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15403_2_lut.init = 16'h8888;
    LUT4 i15439_2_lut (.A(wb_addr[8]), .B(n3), .Z(n17191)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15439_2_lut.init = 16'h8888;
    LUT4 i15450_2_lut (.A(wb_addr[9]), .B(n3), .Z(n17189)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15450_2_lut.init = 16'h8888;
    LUT4 i15420_2_lut (.A(wb_addr[6]), .B(n3), .Z(n17195)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15420_2_lut.init = 16'h8888;
    LUT4 i15426_2_lut (.A(wb_addr[7]), .B(n3), .Z(n17193)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15426_2_lut.init = 16'h8888;
    LUT4 i15413_2_lut (.A(wb_addr[4]), .B(n3), .Z(n17199)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15413_2_lut.init = 16'h8888;
    LUT4 i15416_2_lut (.A(wb_addr[5]), .B(n3), .Z(n17197)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15416_2_lut.init = 16'h8888;
    LUT4 i15410_2_lut (.A(wb_addr[2]), .B(n3), .Z(n17203)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15410_2_lut.init = 16'h8888;
    LUT4 i15411_2_lut (.A(wb_addr[3]), .B(n3), .Z(n17201)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15411_2_lut.init = 16'h8888;
    LUT4 i15409_2_lut (.A(wb_addr[1]), .B(n3), .Z(n17205)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15409_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_129 (.A(wb_err), .B(n29268), .C(wb_we), .D(wb_cyc), 
         .Z(n20131)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut_adj_129.init = 16'h0100;
    LUT4 i1_4_lut_adj_130 (.A(n26715), .B(o_cmd_busy_N_941), .C(wb_ack), 
         .D(o_cmd_busy_N_933), .Z(dac_clk_p_c_enable_414)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+!((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(122[6:41])
    defparam i1_4_lut_adj_130.init = 16'heefc;
    LUT4 i22392_2_lut (.A(wb_cyc), .B(wb_stb), .Z(o_cmd_busy_N_933)) /* synthesis lut_function=(!(A+(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(149[11] 168[5])
    defparam i22392_2_lut.init = 16'h1111;
    LUT4 i1_2_lut_3_lut_4_lut (.A(wb_err), .B(wb_cyc), .C(wb_stb), .D(n29268), 
         .Z(n19567)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(122[17:41])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfff8;
    LUT4 i1_2_lut_rep_556_3_lut (.A(wb_err), .B(wb_cyc), .C(n29268), .Z(o_cmd_busy_N_941)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(122[17:41])
    defparam i1_2_lut_rep_556_3_lut.init = 16'hf8f8;
    FD1S3IX o_rsp_word_i1 (.D(n20131), .CK(dac_clk_p_c), .CD(n12635), 
            .Q(ow_word[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i1.GSR = "DISABLED";
    FD1P3IX o_wb_cyc_67 (.D(o_cmd_busy_N_933), .SP(dac_clk_p_c_enable_414), 
            .CD(o_cmd_busy_N_941), .CK(dac_clk_p_c), .Q(wb_cyc)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(121[9] 168[5])
    defparam o_wb_cyc_67.GSR = "DISABLED";
    FD1P3AX o_wb_addr_546__i29 (.D(n125[29]), .SP(dac_clk_p_c_enable_446), 
            .CK(dac_clk_p_c), .Q(wb_addr[29])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_546__i29.GSR = "DISABLED";
    FD1P3AX o_wb_addr_546__i28 (.D(n125[28]), .SP(dac_clk_p_c_enable_446), 
            .CK(dac_clk_p_c), .Q(wb_addr[28])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_546__i28.GSR = "DISABLED";
    FD1P3AX o_wb_addr_546__i27 (.D(n125[27]), .SP(dac_clk_p_c_enable_446), 
            .CK(dac_clk_p_c), .Q(wb_addr[27])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_546__i27.GSR = "DISABLED";
    FD1P3AX o_wb_addr_546__i26 (.D(n125[26]), .SP(dac_clk_p_c_enable_446), 
            .CK(dac_clk_p_c), .Q(wb_addr[26])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_546__i26.GSR = "DISABLED";
    FD1P3AX o_wb_addr_546__i25 (.D(n125[25]), .SP(dac_clk_p_c_enable_446), 
            .CK(dac_clk_p_c), .Q(wb_addr[25])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_546__i25.GSR = "DISABLED";
    FD1P3AX o_wb_addr_546__i24 (.D(n125[24]), .SP(dac_clk_p_c_enable_446), 
            .CK(dac_clk_p_c), .Q(wb_addr[24])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_546__i24.GSR = "DISABLED";
    FD1P3AX o_wb_addr_546__i23 (.D(n125[23]), .SP(dac_clk_p_c_enable_446), 
            .CK(dac_clk_p_c), .Q(wb_addr[23])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_546__i23.GSR = "DISABLED";
    FD1P3AX o_wb_addr_546__i22 (.D(n125[22]), .SP(dac_clk_p_c_enable_446), 
            .CK(dac_clk_p_c), .Q(wb_addr[22])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_546__i22.GSR = "DISABLED";
    FD1P3AX o_wb_addr_546__i21 (.D(n125[21]), .SP(dac_clk_p_c_enable_446), 
            .CK(dac_clk_p_c), .Q(wb_addr[21])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_546__i21.GSR = "DISABLED";
    FD1P3AX o_wb_addr_546__i20 (.D(n125[20]), .SP(dac_clk_p_c_enable_446), 
            .CK(dac_clk_p_c), .Q(wb_addr[20])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_546__i20.GSR = "DISABLED";
    FD1P3AX o_wb_addr_546__i19 (.D(n125[19]), .SP(dac_clk_p_c_enable_446), 
            .CK(dac_clk_p_c), .Q(wb_addr[19])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_546__i19.GSR = "DISABLED";
    FD1P3AX o_wb_addr_546__i18 (.D(n125[18]), .SP(dac_clk_p_c_enable_446), 
            .CK(dac_clk_p_c), .Q(wb_addr[18])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_546__i18.GSR = "DISABLED";
    FD1P3AX o_wb_addr_546__i17 (.D(n125[17]), .SP(dac_clk_p_c_enable_446), 
            .CK(dac_clk_p_c), .Q(wb_addr[17])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_546__i17.GSR = "DISABLED";
    FD1P3AX o_wb_addr_546__i16 (.D(n125[16]), .SP(dac_clk_p_c_enable_446), 
            .CK(dac_clk_p_c), .Q(wb_addr[16])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_546__i16.GSR = "DISABLED";
    FD1P3AX o_wb_addr_546__i15 (.D(n125[15]), .SP(dac_clk_p_c_enable_446), 
            .CK(dac_clk_p_c), .Q(wb_addr[15])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_546__i15.GSR = "DISABLED";
    FD1P3AX o_wb_addr_546__i14 (.D(n125[14]), .SP(dac_clk_p_c_enable_446), 
            .CK(dac_clk_p_c), .Q(wb_addr[14])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_546__i14.GSR = "DISABLED";
    FD1P3AX o_wb_addr_546__i13 (.D(n125[13]), .SP(dac_clk_p_c_enable_446), 
            .CK(dac_clk_p_c), .Q(wb_addr[13])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_546__i13.GSR = "DISABLED";
    FD1P3AX o_wb_addr_546__i12 (.D(n125[12]), .SP(dac_clk_p_c_enable_446), 
            .CK(dac_clk_p_c), .Q(wb_addr[12])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_546__i12.GSR = "DISABLED";
    FD1P3AX o_wb_addr_546__i11 (.D(n125[11]), .SP(dac_clk_p_c_enable_446), 
            .CK(dac_clk_p_c), .Q(wb_addr[11])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_546__i11.GSR = "DISABLED";
    FD1P3AX o_wb_addr_546__i10 (.D(n125[10]), .SP(dac_clk_p_c_enable_446), 
            .CK(dac_clk_p_c), .Q(wb_addr[10])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_546__i10.GSR = "DISABLED";
    FD1P3AX o_wb_addr_546__i9 (.D(n125[9]), .SP(dac_clk_p_c_enable_446), 
            .CK(dac_clk_p_c), .Q(wb_addr[9])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_546__i9.GSR = "DISABLED";
    FD1P3AX o_wb_addr_546__i8 (.D(n125[8]), .SP(dac_clk_p_c_enable_446), 
            .CK(dac_clk_p_c), .Q(wb_addr[8])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_546__i8.GSR = "DISABLED";
    FD1P3AX o_wb_addr_546__i7 (.D(n125[7]), .SP(dac_clk_p_c_enable_446), 
            .CK(dac_clk_p_c), .Q(wb_addr[7])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_546__i7.GSR = "DISABLED";
    FD1P3AX o_wb_addr_546__i6 (.D(n125[6]), .SP(dac_clk_p_c_enable_446), 
            .CK(dac_clk_p_c), .Q(wb_addr[6])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_546__i6.GSR = "DISABLED";
    FD1P3AX o_wb_addr_546__i5 (.D(n125[5]), .SP(dac_clk_p_c_enable_446), 
            .CK(dac_clk_p_c), .Q(wb_addr[5])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_546__i5.GSR = "DISABLED";
    FD1P3AX o_wb_addr_546__i4 (.D(n125[4]), .SP(dac_clk_p_c_enable_446), 
            .CK(dac_clk_p_c), .Q(wb_addr[4])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_546__i4.GSR = "DISABLED";
    FD1P3AX o_wb_addr_546__i3 (.D(n125[3]), .SP(dac_clk_p_c_enable_446), 
            .CK(dac_clk_p_c), .Q(wb_addr[3])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_546__i3.GSR = "DISABLED";
    FD1P3AX o_wb_addr_546__i2 (.D(n125[2]), .SP(dac_clk_p_c_enable_446), 
            .CK(dac_clk_p_c), .Q(wb_addr[2])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_546__i2.GSR = "DISABLED";
    FD1P3AX o_wb_addr_546__i1 (.D(n125[1]), .SP(dac_clk_p_c_enable_446), 
            .CK(dac_clk_p_c), .Q(wb_addr[1])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_546__i1.GSR = "DISABLED";
    FD1P3AX o_wb_addr_546__i0 (.D(n125[0]), .SP(dac_clk_p_c_enable_446), 
            .CK(dac_clk_p_c), .Q(wb_addr[0])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_546__i0.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module hbdeword
//

module hbdeword (dac_clk_p_c, dac_clk_p_c_enable_307, hb_bits, dac_clk_p_c_enable_193, 
            n29269, idl_word, n29210, hb_busy, w_reset, n26536, 
            idl_stb, n29268, nl_busy, hx_stb) /* synthesis syn_module_defined=1 */ ;
    input dac_clk_p_c;
    input dac_clk_p_c_enable_307;
    output [4:0]hb_bits;
    input dac_clk_p_c_enable_193;
    input n29269;
    input [33:0]idl_word;
    input n29210;
    output hb_busy;
    input w_reset;
    output n26536;
    input idl_stb;
    input n29268;
    input nl_busy;
    input hx_stb;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(29[49:58])
    wire [3:0]r_len;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(58[12:17])
    
    wire n26423;
    wire [3:0]n13;
    
    wire dac_clk_p_c_enable_236;
    wire [4:0]o_dw_bits_4__N_1188;
    wire [31:0]r_word;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(59[13:19])
    wire [31:0]r_word_31__N_1197;
    wire [3:0]r_len_3__N_1229;
    
    wire n12707, o_dw_busy_N_1269, n11468;
    wire [4:0]o_dw_bits_4__N_1279;
    
    wire n11464, n19914, n25745, n26207, n26532;
    
    FD1P3IX r_len__i0 (.D(n13[0]), .SP(dac_clk_p_c_enable_307), .CD(n26423), 
            .CK(dac_clk_p_c), .Q(r_len[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(64[9] 81[6])
    defparam r_len__i0.GSR = "DISABLED";
    FD1P3AX o_dw_bits_i0 (.D(o_dw_bits_4__N_1188[0]), .SP(dac_clk_p_c_enable_236), 
            .CK(dac_clk_p_c), .Q(hb_bits[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(95[9] 103[41])
    defparam o_dw_bits_i0.GSR = "DISABLED";
    FD1P3AX o_dw_bits_i3 (.D(o_dw_bits_4__N_1188[3]), .SP(dac_clk_p_c_enable_236), 
            .CK(dac_clk_p_c), .Q(hb_bits[3])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(95[9] 103[41])
    defparam o_dw_bits_i3.GSR = "DISABLED";
    FD1P3AX o_dw_bits_i2 (.D(o_dw_bits_4__N_1188[2]), .SP(dac_clk_p_c_enable_236), 
            .CK(dac_clk_p_c), .Q(hb_bits[2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(95[9] 103[41])
    defparam o_dw_bits_i2.GSR = "DISABLED";
    FD1P3AX o_dw_bits_i1 (.D(o_dw_bits_4__N_1188[1]), .SP(dac_clk_p_c_enable_236), 
            .CK(dac_clk_p_c), .Q(hb_bits[1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(95[9] 103[41])
    defparam o_dw_bits_i1.GSR = "DISABLED";
    FD1P3AX r_word_i31 (.D(r_word_31__N_1197[31]), .SP(dac_clk_p_c_enable_236), 
            .CK(dac_clk_p_c), .Q(r_word[31])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i31.GSR = "DISABLED";
    FD1P3IX r_len__i3 (.D(r_len_3__N_1229[3]), .SP(dac_clk_p_c_enable_193), 
            .CD(n29269), .CK(dac_clk_p_c), .Q(r_len[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(64[9] 81[6])
    defparam r_len__i3.GSR = "DISABLED";
    FD1P3IX r_word_i1 (.D(idl_word[1]), .SP(dac_clk_p_c_enable_236), .CD(n12707), 
            .CK(dac_clk_p_c), .Q(r_word[1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i1.GSR = "DISABLED";
    FD1P3IX r_word_i2 (.D(idl_word[2]), .SP(dac_clk_p_c_enable_236), .CD(n12707), 
            .CK(dac_clk_p_c), .Q(r_word[2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i2.GSR = "DISABLED";
    FD1P3IX r_word_i3 (.D(idl_word[3]), .SP(dac_clk_p_c_enable_236), .CD(n12707), 
            .CK(dac_clk_p_c), .Q(r_word[3])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i3.GSR = "DISABLED";
    FD1P3IX o_dw_bits_i4 (.D(n29210), .SP(dac_clk_p_c_enable_236), .CD(n12707), 
            .CK(dac_clk_p_c), .Q(hb_bits[4])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(95[9] 103[41])
    defparam o_dw_bits_i4.GSR = "DISABLED";
    FD1P3IX o_dw_stb_36 (.D(o_dw_busy_N_1269), .SP(dac_clk_p_c_enable_193), 
            .CD(w_reset), .CK(dac_clk_p_c), .Q(hb_busy)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(64[9] 81[6])
    defparam o_dw_stb_36.GSR = "DISABLED";
    FD1P3IX r_word_i0 (.D(idl_word[0]), .SP(dac_clk_p_c_enable_236), .CD(n12707), 
            .CK(dac_clk_p_c), .Q(r_word[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i0.GSR = "DISABLED";
    FD1P3AX r_word_i30 (.D(r_word_31__N_1197[30]), .SP(dac_clk_p_c_enable_236), 
            .CK(dac_clk_p_c), .Q(r_word[30])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i30.GSR = "DISABLED";
    FD1P3AX r_word_i29 (.D(r_word_31__N_1197[29]), .SP(dac_clk_p_c_enable_236), 
            .CK(dac_clk_p_c), .Q(r_word[29])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i29.GSR = "DISABLED";
    FD1P3AX r_word_i28 (.D(r_word_31__N_1197[28]), .SP(dac_clk_p_c_enable_236), 
            .CK(dac_clk_p_c), .Q(r_word[28])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i28.GSR = "DISABLED";
    FD1P3AX r_word_i27 (.D(r_word_31__N_1197[27]), .SP(dac_clk_p_c_enable_236), 
            .CK(dac_clk_p_c), .Q(r_word[27])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i27.GSR = "DISABLED";
    FD1P3AX r_word_i26 (.D(r_word_31__N_1197[26]), .SP(dac_clk_p_c_enable_236), 
            .CK(dac_clk_p_c), .Q(r_word[26])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i26.GSR = "DISABLED";
    FD1P3AX r_word_i25 (.D(r_word_31__N_1197[25]), .SP(dac_clk_p_c_enable_236), 
            .CK(dac_clk_p_c), .Q(r_word[25])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i25.GSR = "DISABLED";
    FD1P3AX r_word_i24 (.D(r_word_31__N_1197[24]), .SP(dac_clk_p_c_enable_236), 
            .CK(dac_clk_p_c), .Q(r_word[24])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i24.GSR = "DISABLED";
    FD1P3AX r_word_i23 (.D(r_word_31__N_1197[23]), .SP(dac_clk_p_c_enable_236), 
            .CK(dac_clk_p_c), .Q(r_word[23])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i23.GSR = "DISABLED";
    FD1P3AX r_word_i22 (.D(r_word_31__N_1197[22]), .SP(dac_clk_p_c_enable_236), 
            .CK(dac_clk_p_c), .Q(r_word[22])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i22.GSR = "DISABLED";
    FD1P3AX r_word_i21 (.D(r_word_31__N_1197[21]), .SP(dac_clk_p_c_enable_236), 
            .CK(dac_clk_p_c), .Q(r_word[21])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i21.GSR = "DISABLED";
    FD1P3AX r_word_i20 (.D(r_word_31__N_1197[20]), .SP(dac_clk_p_c_enable_236), 
            .CK(dac_clk_p_c), .Q(r_word[20])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i20.GSR = "DISABLED";
    FD1P3AX r_word_i19 (.D(r_word_31__N_1197[19]), .SP(dac_clk_p_c_enable_236), 
            .CK(dac_clk_p_c), .Q(r_word[19])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i19.GSR = "DISABLED";
    FD1P3AX r_word_i18 (.D(r_word_31__N_1197[18]), .SP(dac_clk_p_c_enable_236), 
            .CK(dac_clk_p_c), .Q(r_word[18])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i18.GSR = "DISABLED";
    FD1P3AX r_word_i17 (.D(r_word_31__N_1197[17]), .SP(dac_clk_p_c_enable_236), 
            .CK(dac_clk_p_c), .Q(r_word[17])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i17.GSR = "DISABLED";
    FD1P3AX r_word_i16 (.D(r_word_31__N_1197[16]), .SP(dac_clk_p_c_enable_236), 
            .CK(dac_clk_p_c), .Q(r_word[16])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i16.GSR = "DISABLED";
    FD1P3AX r_word_i15 (.D(r_word_31__N_1197[15]), .SP(dac_clk_p_c_enable_236), 
            .CK(dac_clk_p_c), .Q(r_word[15])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i15.GSR = "DISABLED";
    FD1P3AX r_word_i14 (.D(r_word_31__N_1197[14]), .SP(dac_clk_p_c_enable_236), 
            .CK(dac_clk_p_c), .Q(r_word[14])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i14.GSR = "DISABLED";
    FD1P3AX r_word_i13 (.D(r_word_31__N_1197[13]), .SP(dac_clk_p_c_enable_236), 
            .CK(dac_clk_p_c), .Q(r_word[13])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i13.GSR = "DISABLED";
    FD1P3AX r_word_i12 (.D(r_word_31__N_1197[12]), .SP(dac_clk_p_c_enable_236), 
            .CK(dac_clk_p_c), .Q(r_word[12])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i12.GSR = "DISABLED";
    FD1P3AX r_word_i11 (.D(r_word_31__N_1197[11]), .SP(dac_clk_p_c_enable_236), 
            .CK(dac_clk_p_c), .Q(r_word[11])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i11.GSR = "DISABLED";
    FD1P3AX r_word_i10 (.D(r_word_31__N_1197[10]), .SP(dac_clk_p_c_enable_236), 
            .CK(dac_clk_p_c), .Q(r_word[10])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i10.GSR = "DISABLED";
    FD1P3AX r_word_i9 (.D(r_word_31__N_1197[9]), .SP(dac_clk_p_c_enable_236), 
            .CK(dac_clk_p_c), .Q(r_word[9])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i9.GSR = "DISABLED";
    FD1P3AX r_word_i8 (.D(r_word_31__N_1197[8]), .SP(dac_clk_p_c_enable_236), 
            .CK(dac_clk_p_c), .Q(r_word[8])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i8.GSR = "DISABLED";
    FD1P3AX r_word_i7 (.D(r_word_31__N_1197[7]), .SP(dac_clk_p_c_enable_236), 
            .CK(dac_clk_p_c), .Q(r_word[7])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i7.GSR = "DISABLED";
    FD1P3AX r_word_i6 (.D(r_word_31__N_1197[6]), .SP(dac_clk_p_c_enable_236), 
            .CK(dac_clk_p_c), .Q(r_word[6])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i6.GSR = "DISABLED";
    FD1P3AX r_word_i5 (.D(r_word_31__N_1197[5]), .SP(dac_clk_p_c_enable_236), 
            .CK(dac_clk_p_c), .Q(r_word[5])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i5.GSR = "DISABLED";
    FD1P3AX r_word_i4 (.D(r_word_31__N_1197[4]), .SP(dac_clk_p_c_enable_236), 
            .CK(dac_clk_p_c), .Q(r_word[4])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i4.GSR = "DISABLED";
    LUT4 i1_3_lut_4_lut_3_lut_4_lut (.A(r_len[0]), .B(r_len[1]), .C(r_len[2]), 
         .D(r_len[3]), .Z(n11468)) /* synthesis lut_function=(A (B)+!A !(B+!(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(80[14:26])
    defparam i1_3_lut_4_lut_3_lut_4_lut.init = 16'h9998;
    LUT4 i11042_2_lut (.A(idl_word[32]), .B(idl_word[33]), .Z(o_dw_bits_4__N_1279[3])) /* synthesis lut_function=(A (B)) */ ;
    defparam i11042_2_lut.init = 16'h8888;
    FD1P3IX r_len__i2 (.D(n11464), .SP(dac_clk_p_c_enable_307), .CD(n26423), 
            .CK(dac_clk_p_c), .Q(r_len[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(64[9] 81[6])
    defparam r_len__i2.GSR = "DISABLED";
    FD1P3IX r_len__i1 (.D(n11468), .SP(dac_clk_p_c_enable_307), .CD(n26423), 
            .CK(dac_clk_p_c), .Q(r_len[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(64[9] 81[6])
    defparam r_len__i1.GSR = "DISABLED";
    LUT4 o_dw_bits_4__I_0_i3_4_lut (.A(r_word[30]), .B(idl_word[31]), .C(n26536), 
         .D(o_dw_bits_4__N_1279[3]), .Z(o_dw_bits_4__N_1188[2])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(102[12] 103[41])
    defparam o_dw_bits_4__I_0_i3_4_lut.init = 16'hca0a;
    LUT4 mux_15_i4_4_lut (.A(r_len[3]), .B(o_dw_bits_4__N_1279[3]), .C(n26536), 
         .D(n19914), .Z(r_len_3__N_1229[3])) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(76[12] 81[6])
    defparam mux_15_i4_4_lut.init = 16'h3a35;
    LUT4 r_word_29__bdd_3_lut_24012 (.A(idl_word[30]), .B(idl_word[33]), 
         .C(idl_word[32]), .Z(n25745)) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam r_word_29__bdd_3_lut_24012.init = 16'h8c8c;
    LUT4 r_word_28__bdd_3_lut_24355 (.A(idl_word[29]), .B(idl_word[32]), 
         .C(idl_word[33]), .Z(n26207)) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam r_word_28__bdd_3_lut_24355.init = 16'h8c8c;
    LUT4 r_word_31__I_0_i21_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[20]), 
         .D(r_word[16]), .Z(r_word_31__N_1197[20])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i21_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i20_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[19]), 
         .D(r_word[15]), .Z(r_word_31__N_1197[19])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i20_3_lut_4_lut.init = 16'hfd20;
    LUT4 i1_3_lut_3_lut_4_lut (.A(r_len[0]), .B(r_len[1]), .C(r_len[3]), 
         .D(r_len[2]), .Z(n11464)) /* synthesis lut_function=(A (D)+!A (B (D)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(80[14:26])
    defparam i1_3_lut_3_lut_4_lut.init = 16'hee10;
    LUT4 i1_4_lut_4_lut (.A(r_len[0]), .B(r_len[1]), .C(r_len[3]), .D(r_len[2]), 
         .Z(n19914)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(80[14:26])
    defparam i1_4_lut_4_lut.init = 16'hffef;
    LUT4 r_word_31__I_0_i19_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[18]), 
         .D(r_word[14]), .Z(r_word_31__N_1197[18])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i19_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i18_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[17]), 
         .D(r_word[13]), .Z(r_word_31__N_1197[17])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i18_3_lut_4_lut.init = 16'hfd20;
    LUT4 i3_4_lut_rep_572 (.A(r_len[0]), .B(r_len[1]), .C(r_len[2]), .D(r_len[3]), 
         .Z(n26532)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(78[16:31])
    defparam i3_4_lut_rep_572.init = 16'hfffe;
    LUT4 i1_2_lut_4_lut (.A(r_len[0]), .B(r_len[1]), .C(r_len[2]), .D(r_len[3]), 
         .Z(n13[0])) /* synthesis lut_function=(!(A+!(B+(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(78[16:31])
    defparam i1_2_lut_4_lut.init = 16'h5554;
    LUT4 r_word_31__I_0_i17_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[16]), 
         .D(r_word[12]), .Z(r_word_31__N_1197[16])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i17_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i16_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[15]), 
         .D(r_word[11]), .Z(r_word_31__N_1197[15])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i16_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i15_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[14]), 
         .D(r_word[10]), .Z(r_word_31__N_1197[14])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i15_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i14_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[13]), 
         .D(r_word[9]), .Z(r_word_31__N_1197[13])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i14_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i13_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[12]), 
         .D(r_word[8]), .Z(r_word_31__N_1197[12])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i13_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i12_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[11]), 
         .D(r_word[7]), .Z(r_word_31__N_1197[11])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i12_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i11_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[10]), 
         .D(r_word[6]), .Z(r_word_31__N_1197[10])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i11_3_lut_4_lut.init = 16'hfd20;
    LUT4 i_stb_I_0_2_lut_rep_576 (.A(idl_stb), .B(hb_busy), .Z(n26536)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam i_stb_I_0_2_lut_rep_576.init = 16'h2222;
    LUT4 r_word_31__I_0_i10_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[9]), 
         .D(r_word[5]), .Z(r_word_31__N_1197[9])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i10_3_lut_4_lut.init = 16'hfd20;
    LUT4 i11049_2_lut_3_lut (.A(idl_stb), .B(hb_busy), .C(n26532), .Z(o_dw_busy_N_1269)) /* synthesis lut_function=(A ((C)+!B)+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam i11049_2_lut_3_lut.init = 16'hf2f2;
    LUT4 r_word_31__I_0_i9_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[8]), 
         .D(r_word[4]), .Z(r_word_31__N_1197[8])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i9_3_lut_4_lut.init = 16'hfd20;
    LUT4 o_dw_bits_4__I_0_i4_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(o_dw_bits_4__N_1279[3]), 
         .D(r_word[31]), .Z(o_dw_bits_4__N_1188[3])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam o_dw_bits_4__I_0_i4_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_28__bdd_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(n26207), 
         .D(r_word[28]), .Z(o_dw_bits_4__N_1188[0])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_28__bdd_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i8_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[7]), 
         .D(r_word[3]), .Z(r_word_31__N_1197[7])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i8_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i7_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[6]), 
         .D(r_word[2]), .Z(r_word_31__N_1197[6])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i7_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i6_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[5]), 
         .D(r_word[1]), .Z(r_word_31__N_1197[5])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i6_3_lut_4_lut.init = 16'hfd20;
    LUT4 i7025_2_lut_rep_463_3_lut (.A(idl_stb), .B(hb_busy), .C(n29268), 
         .Z(n26423)) /* synthesis lut_function=(A ((C)+!B)+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam i7025_2_lut_rep_463_3_lut.init = 16'hf2f2;
    LUT4 i22405_2_lut_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(nl_busy), 
         .D(hx_stb), .Z(n12707)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam i22405_2_lut_3_lut_4_lut.init = 16'h0ddd;
    LUT4 i1_2_lut_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(nl_busy), 
         .D(hx_stb), .Z(dac_clk_p_c_enable_236)) /* synthesis lut_function=(!(A (B (C (D)))+!A (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h2fff;
    LUT4 r_word_31__I_0_i32_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[31]), 
         .D(r_word[27]), .Z(r_word_31__N_1197[31])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i32_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i5_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[4]), 
         .D(r_word[0]), .Z(r_word_31__N_1197[4])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i5_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i31_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[30]), 
         .D(r_word[26]), .Z(r_word_31__N_1197[30])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i31_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i30_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[29]), 
         .D(r_word[25]), .Z(r_word_31__N_1197[29])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i30_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_29__bdd_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(n25745), 
         .D(r_word[29]), .Z(o_dw_bits_4__N_1188[1])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_29__bdd_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i29_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[28]), 
         .D(r_word[24]), .Z(r_word_31__N_1197[28])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i29_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i28_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[27]), 
         .D(r_word[23]), .Z(r_word_31__N_1197[27])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i28_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i27_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[26]), 
         .D(r_word[22]), .Z(r_word_31__N_1197[26])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i27_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i26_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[25]), 
         .D(r_word[21]), .Z(r_word_31__N_1197[25])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i26_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i25_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[24]), 
         .D(r_word[20]), .Z(r_word_31__N_1197[24])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i25_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i24_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[23]), 
         .D(r_word[19]), .Z(r_word_31__N_1197[23])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i24_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i23_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[22]), 
         .D(r_word[18]), .Z(r_word_31__N_1197[22])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i23_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i22_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[21]), 
         .D(r_word[17]), .Z(r_word_31__N_1197[21])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i22_3_lut_4_lut.init = 16'hfd20;
    
endmodule
//
// Verilog Description of module hbpack
//

module hbpack (dac_clk_p_c, dac_clk_p_c_enable_380, n29269, iw_word, 
            w_reset, o_pck_stb_N_765, cmd_loaded, dac_clk_p_c_enable_196, 
            cmd_loaded_N_768, \dec_bits[4] , wb_cyc, inc, n17206, 
            \iw_word[32] , \iw_word[31] , \iw_word[30] , \iw_word[29] , 
            \iw_word[28] , \iw_word[27] , \iw_word[26] , \iw_word[25] , 
            \iw_word[24] , \iw_word[23] , \iw_word[22] , \iw_word[21] , 
            \iw_word[20] , \iw_word[19] , \iw_word[18] , \iw_word[17] , 
            \iw_word[16] , \iw_word[15] , \iw_word[14] , \iw_word[13] , 
            \iw_word[12] , \iw_word[11] , \iw_word[10] , \iw_word[9] , 
            \iw_word[8] , \iw_word[7] , \iw_word[6] , \iw_word[5] , 
            \iw_word[4] , \iw_word[3] , \iw_word[1] , \dec_bits[0] , 
            \dec_bits[1] , dac_clk_p_c_enable_349, n26716, wb_stb, dac_clk_p_c_enable_446, 
            n45, n46, n26715, i_cmd_wr, n21860, dac_clk_p_c_enable_136, 
            n29268, newaddr_N_990) /* synthesis syn_module_defined=1 */ ;
    input dac_clk_p_c;
    input dac_clk_p_c_enable_380;
    input n29269;
    output [33:0]iw_word;
    input w_reset;
    input o_pck_stb_N_765;
    output cmd_loaded;
    input dac_clk_p_c_enable_196;
    input cmd_loaded_N_768;
    input \dec_bits[4] ;
    input wb_cyc;
    input inc;
    output n17206;
    output \iw_word[32] ;
    output \iw_word[31] ;
    output \iw_word[30] ;
    output \iw_word[29] ;
    output \iw_word[28] ;
    output \iw_word[27] ;
    output \iw_word[26] ;
    output \iw_word[25] ;
    output \iw_word[24] ;
    output \iw_word[23] ;
    output \iw_word[22] ;
    output \iw_word[21] ;
    output \iw_word[20] ;
    output \iw_word[19] ;
    output \iw_word[18] ;
    output \iw_word[17] ;
    output \iw_word[16] ;
    output \iw_word[15] ;
    output \iw_word[14] ;
    output \iw_word[13] ;
    output \iw_word[12] ;
    output \iw_word[11] ;
    output \iw_word[10] ;
    output \iw_word[9] ;
    output \iw_word[8] ;
    output \iw_word[7] ;
    output \iw_word[6] ;
    output \iw_word[5] ;
    output \iw_word[4] ;
    output \iw_word[3] ;
    output \iw_word[1] ;
    input \dec_bits[0] ;
    input \dec_bits[1] ;
    input dac_clk_p_c_enable_349;
    output n26716;
    input wb_stb;
    output dac_clk_p_c_enable_446;
    input n45;
    input n46;
    output n26715;
    output i_cmd_wr;
    output n21860;
    output dac_clk_p_c_enable_136;
    input n29268;
    output newaddr_N_990;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(29[49:58])
    wire [33:0]r_word;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(71[13:19])
    wire [33:0]n14;
    
    wire iw_stb, n26525;
    wire [33:0]iw_word_c;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(71[14:21])
    
    FD1P3IX r_word__i0 (.D(n14[0]), .SP(dac_clk_p_c_enable_380), .CD(n29269), 
            .CK(dac_clk_p_c), .Q(r_word[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i0.GSR = "DISABLED";
    FD1P3IX o_pck_word__i0 (.D(r_word[0]), .SP(dac_clk_p_c_enable_380), 
            .CD(n29269), .CK(dac_clk_p_c), .Q(iw_word[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i0.GSR = "DISABLED";
    FD1S3IX o_pck_stb_24 (.D(o_pck_stb_N_765), .CK(dac_clk_p_c), .CD(w_reset), 
            .Q(iw_stb)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(83[9] 84[65])
    defparam o_pck_stb_24.GSR = "DISABLED";
    FD1P3IX cmd_loaded_23 (.D(cmd_loaded_N_768), .SP(dac_clk_p_c_enable_196), 
            .CD(n29269), .CK(dac_clk_p_c), .Q(cmd_loaded)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(74[9] 80[23])
    defparam cmd_loaded_23.GSR = "DISABLED";
    LUT4 i11325_2_lut (.A(r_word[27]), .B(\dec_bits[4] ), .Z(n14[31])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11325_2_lut.init = 16'h2222;
    LUT4 i11326_2_lut (.A(r_word[26]), .B(\dec_bits[4] ), .Z(n14[30])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11326_2_lut.init = 16'h2222;
    LUT4 i11327_2_lut (.A(r_word[25]), .B(\dec_bits[4] ), .Z(n14[29])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11327_2_lut.init = 16'h2222;
    LUT4 i11328_2_lut (.A(r_word[24]), .B(\dec_bits[4] ), .Z(n14[28])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11328_2_lut.init = 16'h2222;
    LUT4 i15408_3_lut_4_lut (.A(n26525), .B(wb_cyc), .C(iw_word[2]), .D(inc), 
         .Z(n17206)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(83[9] 84[65])
    defparam i15408_3_lut_4_lut.init = 16'hfd20;
    FD1P3IX o_pck_word__i33 (.D(r_word[33]), .SP(dac_clk_p_c_enable_380), 
            .CD(w_reset), .CK(dac_clk_p_c), .Q(iw_word_c[33])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i33.GSR = "DISABLED";
    FD1P3IX o_pck_word__i32 (.D(r_word[32]), .SP(dac_clk_p_c_enable_380), 
            .CD(w_reset), .CK(dac_clk_p_c), .Q(\iw_word[32] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i32.GSR = "DISABLED";
    FD1P3IX o_pck_word__i31 (.D(r_word[31]), .SP(dac_clk_p_c_enable_380), 
            .CD(w_reset), .CK(dac_clk_p_c), .Q(\iw_word[31] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i31.GSR = "DISABLED";
    FD1P3IX o_pck_word__i30 (.D(r_word[30]), .SP(dac_clk_p_c_enable_380), 
            .CD(w_reset), .CK(dac_clk_p_c), .Q(\iw_word[30] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i30.GSR = "DISABLED";
    FD1P3IX o_pck_word__i29 (.D(r_word[29]), .SP(dac_clk_p_c_enable_380), 
            .CD(w_reset), .CK(dac_clk_p_c), .Q(\iw_word[29] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i29.GSR = "DISABLED";
    FD1P3IX o_pck_word__i28 (.D(r_word[28]), .SP(dac_clk_p_c_enable_380), 
            .CD(w_reset), .CK(dac_clk_p_c), .Q(\iw_word[28] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i28.GSR = "DISABLED";
    FD1P3IX o_pck_word__i27 (.D(r_word[27]), .SP(dac_clk_p_c_enable_380), 
            .CD(w_reset), .CK(dac_clk_p_c), .Q(\iw_word[27] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i27.GSR = "DISABLED";
    FD1P3IX o_pck_word__i26 (.D(r_word[26]), .SP(dac_clk_p_c_enable_380), 
            .CD(w_reset), .CK(dac_clk_p_c), .Q(\iw_word[26] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i26.GSR = "DISABLED";
    FD1P3IX o_pck_word__i25 (.D(r_word[25]), .SP(dac_clk_p_c_enable_380), 
            .CD(w_reset), .CK(dac_clk_p_c), .Q(\iw_word[25] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i25.GSR = "DISABLED";
    FD1P3IX o_pck_word__i24 (.D(r_word[24]), .SP(dac_clk_p_c_enable_380), 
            .CD(n29269), .CK(dac_clk_p_c), .Q(\iw_word[24] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i24.GSR = "DISABLED";
    FD1P3IX o_pck_word__i23 (.D(r_word[23]), .SP(dac_clk_p_c_enable_380), 
            .CD(w_reset), .CK(dac_clk_p_c), .Q(\iw_word[23] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i23.GSR = "DISABLED";
    FD1P3IX o_pck_word__i22 (.D(r_word[22]), .SP(dac_clk_p_c_enable_380), 
            .CD(w_reset), .CK(dac_clk_p_c), .Q(\iw_word[22] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i22.GSR = "DISABLED";
    FD1P3IX o_pck_word__i21 (.D(r_word[21]), .SP(dac_clk_p_c_enable_380), 
            .CD(n29269), .CK(dac_clk_p_c), .Q(\iw_word[21] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i21.GSR = "DISABLED";
    FD1P3IX o_pck_word__i20 (.D(r_word[20]), .SP(dac_clk_p_c_enable_380), 
            .CD(n29269), .CK(dac_clk_p_c), .Q(\iw_word[20] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i20.GSR = "DISABLED";
    FD1P3IX o_pck_word__i19 (.D(r_word[19]), .SP(dac_clk_p_c_enable_380), 
            .CD(n29269), .CK(dac_clk_p_c), .Q(\iw_word[19] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i19.GSR = "DISABLED";
    FD1P3IX o_pck_word__i18 (.D(r_word[18]), .SP(dac_clk_p_c_enable_380), 
            .CD(n29269), .CK(dac_clk_p_c), .Q(\iw_word[18] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i18.GSR = "DISABLED";
    FD1P3IX o_pck_word__i17 (.D(r_word[17]), .SP(dac_clk_p_c_enable_380), 
            .CD(n29269), .CK(dac_clk_p_c), .Q(\iw_word[17] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i17.GSR = "DISABLED";
    FD1P3IX o_pck_word__i16 (.D(r_word[16]), .SP(dac_clk_p_c_enable_380), 
            .CD(n29269), .CK(dac_clk_p_c), .Q(\iw_word[16] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i16.GSR = "DISABLED";
    FD1P3IX o_pck_word__i15 (.D(r_word[15]), .SP(dac_clk_p_c_enable_380), 
            .CD(n29269), .CK(dac_clk_p_c), .Q(\iw_word[15] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i15.GSR = "DISABLED";
    FD1P3IX o_pck_word__i14 (.D(r_word[14]), .SP(dac_clk_p_c_enable_380), 
            .CD(n29269), .CK(dac_clk_p_c), .Q(\iw_word[14] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i14.GSR = "DISABLED";
    FD1P3IX o_pck_word__i13 (.D(r_word[13]), .SP(dac_clk_p_c_enable_380), 
            .CD(n29269), .CK(dac_clk_p_c), .Q(\iw_word[13] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i13.GSR = "DISABLED";
    FD1P3IX o_pck_word__i12 (.D(r_word[12]), .SP(dac_clk_p_c_enable_380), 
            .CD(n29269), .CK(dac_clk_p_c), .Q(\iw_word[12] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i12.GSR = "DISABLED";
    FD1P3IX o_pck_word__i11 (.D(r_word[11]), .SP(dac_clk_p_c_enable_380), 
            .CD(n29269), .CK(dac_clk_p_c), .Q(\iw_word[11] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i11.GSR = "DISABLED";
    FD1P3IX o_pck_word__i10 (.D(r_word[10]), .SP(dac_clk_p_c_enable_380), 
            .CD(n29269), .CK(dac_clk_p_c), .Q(\iw_word[10] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i10.GSR = "DISABLED";
    FD1P3IX o_pck_word__i9 (.D(r_word[9]), .SP(dac_clk_p_c_enable_380), 
            .CD(n29269), .CK(dac_clk_p_c), .Q(\iw_word[9] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i9.GSR = "DISABLED";
    FD1P3IX o_pck_word__i8 (.D(r_word[8]), .SP(dac_clk_p_c_enable_380), 
            .CD(n29269), .CK(dac_clk_p_c), .Q(\iw_word[8] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i8.GSR = "DISABLED";
    FD1P3IX o_pck_word__i7 (.D(r_word[7]), .SP(dac_clk_p_c_enable_380), 
            .CD(n29269), .CK(dac_clk_p_c), .Q(\iw_word[7] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i7.GSR = "DISABLED";
    FD1P3IX o_pck_word__i6 (.D(r_word[6]), .SP(dac_clk_p_c_enable_380), 
            .CD(n29269), .CK(dac_clk_p_c), .Q(\iw_word[6] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i6.GSR = "DISABLED";
    FD1P3IX o_pck_word__i5 (.D(r_word[5]), .SP(dac_clk_p_c_enable_380), 
            .CD(n29269), .CK(dac_clk_p_c), .Q(\iw_word[5] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i5.GSR = "DISABLED";
    FD1P3IX o_pck_word__i4 (.D(r_word[4]), .SP(dac_clk_p_c_enable_380), 
            .CD(n29269), .CK(dac_clk_p_c), .Q(\iw_word[4] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i4.GSR = "DISABLED";
    FD1P3IX o_pck_word__i3 (.D(r_word[3]), .SP(dac_clk_p_c_enable_380), 
            .CD(n29269), .CK(dac_clk_p_c), .Q(\iw_word[3] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i3.GSR = "DISABLED";
    FD1P3IX o_pck_word__i2 (.D(r_word[2]), .SP(dac_clk_p_c_enable_380), 
            .CD(n29269), .CK(dac_clk_p_c), .Q(iw_word[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i2.GSR = "DISABLED";
    FD1P3IX o_pck_word__i1 (.D(r_word[1]), .SP(dac_clk_p_c_enable_380), 
            .CD(n29269), .CK(dac_clk_p_c), .Q(\iw_word[1] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i1.GSR = "DISABLED";
    LUT4 i11329_2_lut (.A(r_word[23]), .B(\dec_bits[4] ), .Z(n14[27])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11329_2_lut.init = 16'h2222;
    LUT4 i11330_2_lut (.A(r_word[22]), .B(\dec_bits[4] ), .Z(n14[26])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11330_2_lut.init = 16'h2222;
    LUT4 i11331_2_lut (.A(r_word[21]), .B(\dec_bits[4] ), .Z(n14[25])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11331_2_lut.init = 16'h2222;
    LUT4 i11037_2_lut (.A(\dec_bits[0] ), .B(\dec_bits[4] ), .Z(n14[0])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11037_2_lut.init = 16'h2222;
    LUT4 i11332_2_lut (.A(r_word[20]), .B(\dec_bits[4] ), .Z(n14[24])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11332_2_lut.init = 16'h2222;
    LUT4 i11333_2_lut (.A(r_word[19]), .B(\dec_bits[4] ), .Z(n14[23])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11333_2_lut.init = 16'h2222;
    LUT4 i11334_2_lut (.A(r_word[18]), .B(\dec_bits[4] ), .Z(n14[22])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11334_2_lut.init = 16'h2222;
    LUT4 i11335_2_lut (.A(r_word[17]), .B(\dec_bits[4] ), .Z(n14[21])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11335_2_lut.init = 16'h2222;
    LUT4 i11336_2_lut (.A(r_word[16]), .B(\dec_bits[4] ), .Z(n14[20])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11336_2_lut.init = 16'h2222;
    LUT4 i11337_2_lut (.A(r_word[15]), .B(\dec_bits[4] ), .Z(n14[19])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11337_2_lut.init = 16'h2222;
    LUT4 i11338_2_lut (.A(r_word[14]), .B(\dec_bits[4] ), .Z(n14[18])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11338_2_lut.init = 16'h2222;
    LUT4 i11339_2_lut (.A(r_word[13]), .B(\dec_bits[4] ), .Z(n14[17])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11339_2_lut.init = 16'h2222;
    LUT4 i11340_2_lut (.A(r_word[12]), .B(\dec_bits[4] ), .Z(n14[16])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11340_2_lut.init = 16'h2222;
    LUT4 i11341_2_lut (.A(r_word[11]), .B(\dec_bits[4] ), .Z(n14[15])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11341_2_lut.init = 16'h2222;
    LUT4 i11342_2_lut (.A(r_word[10]), .B(\dec_bits[4] ), .Z(n14[14])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11342_2_lut.init = 16'h2222;
    LUT4 i11343_2_lut (.A(r_word[9]), .B(\dec_bits[4] ), .Z(n14[13])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11343_2_lut.init = 16'h2222;
    LUT4 i11345_2_lut (.A(r_word[8]), .B(\dec_bits[4] ), .Z(n14[12])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11345_2_lut.init = 16'h2222;
    LUT4 i11346_2_lut (.A(r_word[7]), .B(\dec_bits[4] ), .Z(n14[11])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11346_2_lut.init = 16'h2222;
    LUT4 i11347_2_lut (.A(r_word[6]), .B(\dec_bits[4] ), .Z(n14[10])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11347_2_lut.init = 16'h2222;
    LUT4 i11348_2_lut (.A(r_word[5]), .B(\dec_bits[4] ), .Z(n14[9])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11348_2_lut.init = 16'h2222;
    LUT4 i11349_2_lut (.A(r_word[4]), .B(\dec_bits[4] ), .Z(n14[8])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11349_2_lut.init = 16'h2222;
    LUT4 i11350_2_lut (.A(r_word[3]), .B(\dec_bits[4] ), .Z(n14[7])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11350_2_lut.init = 16'h2222;
    LUT4 i11351_2_lut (.A(r_word[2]), .B(\dec_bits[4] ), .Z(n14[6])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11351_2_lut.init = 16'h2222;
    LUT4 i11352_2_lut (.A(r_word[1]), .B(\dec_bits[4] ), .Z(n14[5])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11352_2_lut.init = 16'h2222;
    LUT4 i11353_2_lut (.A(r_word[0]), .B(\dec_bits[4] ), .Z(n14[4])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11353_2_lut.init = 16'h2222;
    LUT4 i11354_2_lut (.A(\dec_bits[1] ), .B(\dec_bits[4] ), .Z(n14[1])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11354_2_lut.init = 16'h2222;
    FD1P3IX r_word__i33 (.D(\dec_bits[1] ), .SP(dac_clk_p_c_enable_349), 
            .CD(n29269), .CK(dac_clk_p_c), .Q(r_word[33])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i33.GSR = "DISABLED";
    FD1P3IX r_word__i32 (.D(\dec_bits[0] ), .SP(dac_clk_p_c_enable_349), 
            .CD(n29269), .CK(dac_clk_p_c), .Q(r_word[32])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i32.GSR = "DISABLED";
    FD1P3IX r_word__i31 (.D(n14[31]), .SP(dac_clk_p_c_enable_380), .CD(n29269), 
            .CK(dac_clk_p_c), .Q(r_word[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i31.GSR = "DISABLED";
    FD1P3IX r_word__i30 (.D(n14[30]), .SP(dac_clk_p_c_enable_380), .CD(n29269), 
            .CK(dac_clk_p_c), .Q(r_word[30])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i30.GSR = "DISABLED";
    FD1P3IX r_word__i29 (.D(n14[29]), .SP(dac_clk_p_c_enable_380), .CD(n29269), 
            .CK(dac_clk_p_c), .Q(r_word[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i29.GSR = "DISABLED";
    FD1P3IX r_word__i28 (.D(n14[28]), .SP(dac_clk_p_c_enable_380), .CD(n29269), 
            .CK(dac_clk_p_c), .Q(r_word[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i28.GSR = "DISABLED";
    FD1P3IX r_word__i27 (.D(n14[27]), .SP(dac_clk_p_c_enable_380), .CD(n29269), 
            .CK(dac_clk_p_c), .Q(r_word[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i27.GSR = "DISABLED";
    FD1P3IX r_word__i26 (.D(n14[26]), .SP(dac_clk_p_c_enable_380), .CD(n29269), 
            .CK(dac_clk_p_c), .Q(r_word[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i26.GSR = "DISABLED";
    FD1P3IX r_word__i25 (.D(n14[25]), .SP(dac_clk_p_c_enable_380), .CD(n29269), 
            .CK(dac_clk_p_c), .Q(r_word[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i25.GSR = "DISABLED";
    FD1P3IX r_word__i24 (.D(n14[24]), .SP(dac_clk_p_c_enable_380), .CD(n29269), 
            .CK(dac_clk_p_c), .Q(r_word[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i24.GSR = "DISABLED";
    FD1P3IX r_word__i23 (.D(n14[23]), .SP(dac_clk_p_c_enable_380), .CD(n29269), 
            .CK(dac_clk_p_c), .Q(r_word[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i23.GSR = "DISABLED";
    LUT4 i11031_2_lut_3_lut_4_lut (.A(\iw_word[32] ), .B(n26716), .C(wb_stb), 
         .D(wb_cyc), .Z(dac_clk_p_c_enable_446)) /* synthesis lut_function=(A (C)+!A (B (C+!(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(83[9] 84[65])
    defparam i11031_2_lut_3_lut_4_lut.init = 16'hf0f4;
    FD1P3IX r_word__i22 (.D(n14[22]), .SP(dac_clk_p_c_enable_380), .CD(n29269), 
            .CK(dac_clk_p_c), .Q(r_word[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i22.GSR = "DISABLED";
    FD1P3IX r_word__i21 (.D(n14[21]), .SP(dac_clk_p_c_enable_380), .CD(n29269), 
            .CK(dac_clk_p_c), .Q(r_word[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i21.GSR = "DISABLED";
    FD1P3IX r_word__i20 (.D(n14[20]), .SP(dac_clk_p_c_enable_380), .CD(n29269), 
            .CK(dac_clk_p_c), .Q(r_word[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i20.GSR = "DISABLED";
    FD1P3IX r_word__i19 (.D(n14[19]), .SP(dac_clk_p_c_enable_380), .CD(n29269), 
            .CK(dac_clk_p_c), .Q(r_word[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i19.GSR = "DISABLED";
    FD1P3IX r_word__i18 (.D(n14[18]), .SP(dac_clk_p_c_enable_380), .CD(n29269), 
            .CK(dac_clk_p_c), .Q(r_word[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i18.GSR = "DISABLED";
    FD1P3IX r_word__i17 (.D(n14[17]), .SP(dac_clk_p_c_enable_380), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i17.GSR = "DISABLED";
    FD1P3IX r_word__i16 (.D(n14[16]), .SP(dac_clk_p_c_enable_380), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i16.GSR = "DISABLED";
    FD1P3IX r_word__i15 (.D(n14[15]), .SP(dac_clk_p_c_enable_380), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i15.GSR = "DISABLED";
    FD1P3IX r_word__i14 (.D(n14[14]), .SP(dac_clk_p_c_enable_380), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i14.GSR = "DISABLED";
    FD1P3IX r_word__i13 (.D(n14[13]), .SP(dac_clk_p_c_enable_380), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i13.GSR = "DISABLED";
    FD1P3IX r_word__i12 (.D(n14[12]), .SP(dac_clk_p_c_enable_380), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i12.GSR = "DISABLED";
    FD1P3IX r_word__i11 (.D(n14[11]), .SP(dac_clk_p_c_enable_380), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i11.GSR = "DISABLED";
    FD1P3IX r_word__i10 (.D(n14[10]), .SP(dac_clk_p_c_enable_380), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i10.GSR = "DISABLED";
    FD1P3IX r_word__i9 (.D(n14[9]), .SP(dac_clk_p_c_enable_380), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i9.GSR = "DISABLED";
    FD1P3IX r_word__i8 (.D(n14[8]), .SP(dac_clk_p_c_enable_380), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i8.GSR = "DISABLED";
    FD1P3IX r_word__i7 (.D(n14[7]), .SP(dac_clk_p_c_enable_380), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i7.GSR = "DISABLED";
    FD1P3IX r_word__i6 (.D(n14[6]), .SP(dac_clk_p_c_enable_380), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i6.GSR = "DISABLED";
    FD1P3IX r_word__i5 (.D(n14[5]), .SP(dac_clk_p_c_enable_380), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i5.GSR = "DISABLED";
    FD1P3IX r_word__i4 (.D(n14[4]), .SP(dac_clk_p_c_enable_380), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i4.GSR = "DISABLED";
    FD1P3IX r_word__i3 (.D(n45), .SP(dac_clk_p_c_enable_380), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i3.GSR = "DISABLED";
    FD1P3IX r_word__i2 (.D(n46), .SP(dac_clk_p_c_enable_380), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i2.GSR = "DISABLED";
    FD1P3IX r_word__i1 (.D(n14[1]), .SP(dac_clk_p_c_enable_380), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i1.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_755 (.A(iw_stb), .B(iw_word_c[33]), .Z(n26715)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(83[9] 84[65])
    defparam i1_2_lut_rep_755.init = 16'h2222;
    LUT4 i1_2_lut_3_lut (.A(iw_stb), .B(iw_word_c[33]), .C(\iw_word[32] ), 
         .Z(i_cmd_wr)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(83[9] 84[65])
    defparam i1_2_lut_3_lut.init = 16'h2020;
    LUT4 i19540_3_lut_3_lut (.A(iw_stb), .B(iw_word_c[33]), .C(wb_stb), 
         .Z(n21860)) /* synthesis lut_function=(A ((C)+!B)+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(83[9] 84[65])
    defparam i19540_3_lut_3_lut.init = 16'hf2f2;
    LUT4 i1_2_lut_rep_756 (.A(iw_word_c[33]), .B(iw_stb), .Z(n26716)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(83[9] 84[65])
    defparam i1_2_lut_rep_756.init = 16'h8888;
    LUT4 i1_2_lut_rep_565_3_lut (.A(iw_word_c[33]), .B(iw_stb), .C(\iw_word[32] ), 
         .Z(n26525)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(83[9] 84[65])
    defparam i1_2_lut_rep_565_3_lut.init = 16'h0808;
    LUT4 i1_2_lut_rep_461_3_lut_4_lut (.A(iw_word_c[33]), .B(iw_stb), .C(wb_cyc), 
         .D(\iw_word[32] ), .Z(dac_clk_p_c_enable_136)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(83[9] 84[65])
    defparam i1_2_lut_rep_461_3_lut_4_lut.init = 16'h0008;
    LUT4 i1_2_lut_3_lut_4_lut (.A(iw_word_c[33]), .B(iw_stb), .C(n29268), 
         .D(\iw_word[32] ), .Z(newaddr_N_990)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(83[9] 84[65])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0008;
    
endmodule
//
// Verilog Description of module hbgenhex
//

module hbgenhex (hb_bits, \w_gx_char[0] , \w_gx_char[1] , \w_gx_char[2] , 
            \w_gx_char[3] , \w_gx_char[4] , \w_gx_char[5] , \w_gx_char[6] , 
            dac_clk_p_c, dac_clk_p_c_enable_307, GND_net, VCC_net, hx_stb, 
            w_reset, hb_busy, nl_busy, n29268, n26536, dac_clk_p_c_enable_193, 
            n11652) /* synthesis syn_module_defined=1 */ ;
    input [4:0]hb_bits;
    output \w_gx_char[0] ;
    output \w_gx_char[1] ;
    output \w_gx_char[2] ;
    output \w_gx_char[3] ;
    output \w_gx_char[4] ;
    output \w_gx_char[5] ;
    output \w_gx_char[6] ;
    input dac_clk_p_c;
    output dac_clk_p_c_enable_307;
    input GND_net;
    input VCC_net;
    output hx_stb;
    input w_reset;
    input hb_busy;
    input nl_busy;
    input n29268;
    input n26536;
    output dac_clk_p_c_enable_193;
    output n11652;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(29[49:58])
    
    wire dac_clk_p_c_enable_145, n20240;
    
    SP8KC mux_100 (.DI0(GND_net), .DI1(GND_net), .DI2(GND_net), .DI3(GND_net), 
          .DI4(GND_net), .DI5(GND_net), .DI6(GND_net), .DI7(GND_net), 
          .DI8(GND_net), .AD0(GND_net), .AD1(GND_net), .AD2(GND_net), 
          .AD3(hb_bits[0]), .AD4(hb_bits[1]), .AD5(hb_bits[2]), .AD6(hb_bits[3]), 
          .AD7(hb_bits[4]), .AD8(GND_net), .AD9(GND_net), .AD10(GND_net), 
          .AD11(GND_net), .AD12(GND_net), .CE(dac_clk_p_c_enable_307), 
          .OCE(VCC_net), .CLK(dac_clk_p_c), .WE(GND_net), .CS0(GND_net), 
          .CS1(GND_net), .CS2(GND_net), .RST(GND_net), .DO0(\w_gx_char[0] ), 
          .DO1(\w_gx_char[1] ), .DO2(\w_gx_char[2] ), .DO3(\w_gx_char[3] ), 
          .DO4(\w_gx_char[4] ), .DO5(\w_gx_char[5] ), .DO6(\w_gx_char[6] ));
    defparam mux_100.DATA_WIDTH = 9;
    defparam mux_100.REGMODE = "NOREG";
    defparam mux_100.CSDECODE = "0b000";
    defparam mux_100.WRITEMODE = "NORMAL";
    defparam mux_100.GSR = "DISABLED";
    defparam mux_100.RESETMODE = "ASYNC";
    defparam mux_100.ASYNC_RESET_RELEASE = "SYNC";
    defparam mux_100.INIT_DATA = "STATIC";
    defparam mux_100.INITVAL_00 = "0x01A0D01A0D0B44908A5401A0D01A0D0A641096520CC650C8630C4610723806E3606A340663206230";
    defparam mux_100.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_100.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_100.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_100.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_100.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_100.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_100.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_100.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_100.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_100.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_100.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_100.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_100.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_100.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_100.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_100.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_100.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_100.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_100.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_100.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_100.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_100.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_100.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_100.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_100.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_100.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_100.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_100.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_100.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_100.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_100.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    FD1P3IX o_gx_stb_13 (.D(hb_busy), .SP(dac_clk_p_c_enable_145), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(hx_stb)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=132, LSE_RLINE=133 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbgenhex.v(74[9] 78[21])
    defparam o_gx_stb_13.GSR = "DISABLED";
    LUT4 i22388_2_lut_rep_464 (.A(hx_stb), .B(nl_busy), .Z(dac_clk_p_c_enable_307)) /* synthesis lut_function=(!(A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(76[16:26])
    defparam i22388_2_lut_rep_464.init = 16'h7777;
    LUT4 i632_2_lut_3_lut (.A(hx_stb), .B(nl_busy), .C(n29268), .Z(dac_clk_p_c_enable_145)) /* synthesis lut_function=(((C)+!B)+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(76[16:26])
    defparam i632_2_lut_3_lut.init = 16'hf7f7;
    LUT4 i1_2_lut_3_lut_4_lut (.A(hx_stb), .B(nl_busy), .C(n29268), .D(n26536), 
         .Z(dac_clk_p_c_enable_193)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(76[16:26])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfff7;
    LUT4 i1_4_lut (.A(\w_gx_char[3] ), .B(\w_gx_char[0] ), .C(\w_gx_char[2] ), 
         .D(n20240), .Z(n11652)) /* synthesis lut_function=((((D)+!C)+!B)+!A) */ ;
    defparam i1_4_lut.init = 16'hff7f;
    LUT4 i1_4_lut_adj_128 (.A(\w_gx_char[1] ), .B(\w_gx_char[6] ), .C(\w_gx_char[4] ), 
         .D(\w_gx_char[5] ), .Z(n20240)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_128.init = 16'hfffe;
    
endmodule
//
// Verilog Description of module hbdechex
//

module hbdechex (dac_clk_p_c, dec_bits, w_reset, \rx_data[5] , \rx_data[1] , 
            rx_stb, \rx_data[6] , \rx_data[3] , \rx_data[4] , \rx_data[0] , 
            \rx_data[2] , \dec_bits[1] , n29269, n29268, n45, n46, 
            dac_clk_p_c_enable_380, dac_clk_p_c_enable_349, cmd_loaded, 
            o_pck_stb_N_765, dac_clk_p_c_enable_196, cmd_loaded_N_768) /* synthesis syn_module_defined=1 */ ;
    input dac_clk_p_c;
    output [4:0]dec_bits;
    output w_reset;
    input \rx_data[5] ;
    input \rx_data[1] ;
    input rx_stb;
    input \rx_data[6] ;
    input \rx_data[3] ;
    input \rx_data[4] ;
    input \rx_data[0] ;
    input \rx_data[2] ;
    output \dec_bits[1] ;
    output n29269;
    output n29268;
    output n45;
    output n46;
    output dac_clk_p_c_enable_380;
    output dac_clk_p_c_enable_349;
    input cmd_loaded;
    output o_pck_stb_N_765;
    output dac_clk_p_c_enable_196;
    output cmd_loaded_N_768;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(29[49:58])
    
    wire dec_stb, o_dh_stb_N_623;
    wire [4:0]o_dh_bits_4__N_596;
    
    wire o_reset_N_625, n24305, n24304, n24306, n26852, n26853, 
        n26854, n26838, n26839, n26840, n19617, n14504, n20538, 
        n52, n19683, n26829, n26830, n26831, n13, n20568, n24302, 
        n24300, n24303, n25658;
    wire [4:0]dec_bits_c;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(69[13:21])
    
    wire n64, n4, n25600, n25602, n25644, n25645, n20446, n25643, 
        n28305, n28307, n28306, n20194, n26530, n28308, n20190, 
        n36, n43, n19950, n26343, n47, n26729;
    
    FD1S3AX o_dh_stb_35 (.D(o_dh_stb_N_623), .CK(dac_clk_p_c), .Q(dec_stb)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=30, LSE_LLINE=93, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(57[9] 58[47])
    defparam o_dh_stb_35.GSR = "DISABLED";
    FD1S3AX o_dh_bits_i0 (.D(o_dh_bits_4__N_596[0]), .CK(dac_clk_p_c), .Q(dec_bits[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=30, LSE_LLINE=93, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(60[9] 100[5])
    defparam o_dh_bits_i0.GSR = "DISABLED";
    FD1S3AY o_reset_34 (.D(o_reset_N_625), .CK(dac_clk_p_c), .Q(w_reset)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=30, LSE_LLINE=93, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(53[9] 54[46])
    defparam o_reset_34.GSR = "DISABLED";
    PFUMX i22729 (.BLUT(n24305), .ALUT(n24304), .C0(\rx_data[5] ), .Z(n24306));
    PFUMX i24537 (.BLUT(n26852), .ALUT(n26853), .C0(\rx_data[1] ), .Z(n26854));
    PFUMX i24528 (.BLUT(n26838), .ALUT(n26839), .C0(\rx_data[1] ), .Z(n26840));
    LUT4 i_stb_I_0_58_4_lut (.A(rx_stb), .B(n19617), .C(n14504), .D(n20538), 
         .Z(o_dh_stb_N_623)) /* synthesis lut_function=(!((B (C (D)))+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(58[15:46])
    defparam i_stb_I_0_58_4_lut.init = 16'h2aaa;
    LUT4 i1_2_lut (.A(\rx_data[6] ), .B(\rx_data[3] ), .Z(n20538)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i17436_2_lut (.A(\rx_data[5] ), .B(\rx_data[4] ), .Z(n19617)) /* synthesis lut_function=(A (B)) */ ;
    defparam i17436_2_lut.init = 16'h8888;
    LUT4 i1_4_lut (.A(n26854), .B(n52), .C(n19683), .D(n24306), .Z(o_dh_bits_4__N_596[0])) /* synthesis lut_function=((B+((D)+!C))+!A) */ ;
    defparam i1_4_lut.init = 16'hffdf;
    PFUMX i24522 (.BLUT(n26829), .ALUT(n26830), .C0(\rx_data[0] ), .Z(n26831));
    LUT4 i_stb_I_0_2_lut (.A(rx_stb), .B(n13), .Z(o_reset_N_625)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(54[14:45])
    defparam i_stb_I_0_2_lut.init = 16'h2222;
    LUT4 i1_4_lut_adj_117 (.A(\rx_data[4] ), .B(\rx_data[2] ), .C(\rx_data[6] ), 
         .D(n20568), .Z(n13)) /* synthesis lut_function=((((D)+!C)+!B)+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(72[3:8])
    defparam i1_4_lut_adj_117.init = 16'hff7f;
    LUT4 i1_4_lut_adj_118 (.A(\rx_data[5] ), .B(\rx_data[3] ), .C(\rx_data[0] ), 
         .D(\rx_data[1] ), .Z(n20568)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(72[3:8])
    defparam i1_4_lut_adj_118.init = 16'hfffe;
    PFUMX i22726 (.BLUT(n24302), .ALUT(n24300), .C0(\rx_data[2] ), .Z(n24303));
    FD1S3AX o_dh_bits_i4 (.D(o_dh_bits_4__N_596[4]), .CK(dac_clk_p_c), .Q(dec_bits[4])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=30, LSE_LLINE=93, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(60[9] 100[5])
    defparam o_dh_bits_i4.GSR = "DISABLED";
    LUT4 n26840_bdd_4_lut (.A(n26840), .B(\rx_data[3] ), .C(n25658), .D(\rx_data[6] ), 
         .Z(o_dh_bits_4__N_596[4])) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !((D)+!C))) */ ;
    defparam n26840_bdd_4_lut.init = 16'heef0;
    FD1S3AX o_dh_bits_i3 (.D(o_dh_bits_4__N_596[3]), .CK(dac_clk_p_c), .Q(dec_bits_c[3])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=30, LSE_LLINE=93, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(60[9] 100[5])
    defparam o_dh_bits_i3.GSR = "DISABLED";
    FD1S3AX o_dh_bits_i2 (.D(o_dh_bits_4__N_596[2]), .CK(dac_clk_p_c), .Q(dec_bits_c[2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=30, LSE_LLINE=93, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(60[9] 100[5])
    defparam o_dh_bits_i2.GSR = "DISABLED";
    FD1S3AX o_dh_bits_i1 (.D(o_dh_bits_4__N_596[1]), .CK(dac_clk_p_c), .Q(\dec_bits[1] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=30, LSE_LLINE=93, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(60[9] 100[5])
    defparam o_dh_bits_i1.GSR = "DISABLED";
    LUT4 i1_2_lut_4_lut_4_lut (.A(\rx_data[5] ), .B(\rx_data[2] ), .C(\rx_data[1] ), 
         .D(\rx_data[0] ), .Z(n64)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C+(D)))+!A (B+(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(65[3] 99[10])
    defparam i1_2_lut_4_lut_4_lut.init = 16'h2ba8;
    LUT4 i22491_2_lut (.A(\rx_data[3] ), .B(\rx_data[6] ), .Z(n4)) /* synthesis lut_function=(!(A+(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(72[3:8])
    defparam i22491_2_lut.init = 16'h1111;
    LUT4 rx_data_3__bdd_4_lut_23900 (.A(\rx_data[1] ), .B(\rx_data[6] ), 
         .C(\rx_data[0] ), .D(\rx_data[4] ), .Z(n25600)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(D))+!A (((D)+!C)+!B))) */ ;
    defparam rx_data_3__bdd_4_lut_23900.init = 16'h2248;
    LUT4 rx_data_3__bdd_4_lut_25456 (.A(\rx_data[1] ), .B(\rx_data[0] ), 
         .C(\rx_data[4] ), .D(\rx_data[2] ), .Z(n25602)) /* synthesis lut_function=(!(A+(B (C+(D))+!B !(C (D))))) */ ;
    defparam rx_data_3__bdd_4_lut_25456.init = 16'h1004;
    LUT4 n888_bdd_2_lut_23930 (.A(n25644), .B(\rx_data[5] ), .Z(n25645)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam n888_bdd_2_lut_23930.init = 16'hbbbb;
    LUT4 rx_data_4__bdd_4_lut_23929 (.A(\rx_data[4] ), .B(\rx_data[2] ), 
         .C(\rx_data[1] ), .D(\rx_data[3] ), .Z(n25644)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;
    defparam rx_data_4__bdd_4_lut_23929.init = 16'hfe00;
    LUT4 n20446_bdd_4_lut_24017 (.A(n20446), .B(\rx_data[0] ), .C(\rx_data[1] ), 
         .D(\rx_data[2] ), .Z(n25643)) /* synthesis lut_function=(!((B (C (D))+!B !(C+(D)))+!A)) */ ;
    defparam n20446_bdd_4_lut_24017.init = 16'h2aa8;
    LUT4 rx_data_0__bdd_4_lut_25624 (.A(\rx_data[0] ), .B(\rx_data[6] ), 
         .C(\rx_data[2] ), .D(\rx_data[1] ), .Z(n28305)) /* synthesis lut_function=(!(A ((D)+!B)+!A !(B (C+!(D))+!B !((D)+!C)))) */ ;
    defparam rx_data_0__bdd_4_lut_25624.init = 16'h40dc;
    LUT4 rx_data_4__bdd_4_lut (.A(\rx_data[0] ), .B(\rx_data[2] ), .C(\rx_data[1] ), 
         .D(\rx_data[5] ), .Z(n28307)) /* synthesis lut_function=(A (B (C+!(D))+!B !((D)+!C))+!A !(B (D)+!B (C (D)))) */ ;
    defparam rx_data_4__bdd_4_lut.init = 16'h81fd;
    LUT4 n28305_bdd_3_lut (.A(n28305), .B(\rx_data[6] ), .C(\rx_data[5] ), 
         .Z(n28306)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n28305_bdd_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_119 (.A(n20194), .B(n25645), .C(n26530), .D(\rx_data[6] ), 
         .Z(o_dh_bits_4__N_596[3])) /* synthesis lut_function=(A+(B (C+!(D))+!B (C (D)))) */ ;
    defparam i1_4_lut_adj_119.init = 16'hfaee;
    LUT4 i1_4_lut_adj_120 (.A(\rx_data[4] ), .B(n25643), .C(n64), .D(\rx_data[6] ), 
         .Z(n20194)) /* synthesis lut_function=(A (B)+!A (B+!(C (D)))) */ ;
    defparam i1_4_lut_adj_120.init = 16'hcddd;
    LUT4 i1_4_lut_adj_121 (.A(n20446), .B(n28308), .C(n20190), .D(n36), 
         .Z(o_dh_bits_4__N_596[2])) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_121.init = 16'hfefc;
    LUT4 i1_4_lut_adj_122 (.A(n43), .B(n19950), .C(\rx_data[6] ), .D(n19617), 
         .Z(n20190)) /* synthesis lut_function=(A+(B+!(C+(D)))) */ ;
    defparam i1_4_lut_adj_122.init = 16'heeef;
    LUT4 i20838_3_lut (.A(\rx_data[2] ), .B(\rx_data[0] ), .C(\rx_data[1] ), 
         .Z(n36)) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;
    defparam i20838_3_lut.init = 16'h6a6a;
    LUT4 i1_4_lut_adj_123 (.A(\rx_data[5] ), .B(n4), .C(\rx_data[4] ), 
         .D(\rx_data[2] ), .Z(n19950)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_123.init = 16'h8000;
    LUT4 i1_4_lut_adj_124 (.A(n26831), .B(n52), .C(n26343), .D(n19683), 
         .Z(o_dh_bits_4__N_596[1])) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;
    defparam i1_4_lut_adj_124.init = 16'hfeff;
    FD1S3AY o_reset_34_rep_823 (.D(o_reset_N_625), .CK(dac_clk_p_c), .Q(n29269)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=30, LSE_LLINE=93, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(53[9] 54[46])
    defparam o_reset_34_rep_823.GSR = "DISABLED";
    LUT4 n25600_bdd_4_lut (.A(n25600), .B(\rx_data[3] ), .C(n25602), .D(\rx_data[5] ), 
         .Z(n26343)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A ((D)+!C))) */ ;
    defparam n25600_bdd_4_lut.init = 16'h22f0;
    FD1S3AY o_reset_34_rep_822 (.D(o_reset_N_625), .CK(dac_clk_p_c), .Q(n29268)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=30, LSE_LLINE=93, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(53[9] 54[46])
    defparam o_reset_34_rep_822.GSR = "DISABLED";
    LUT4 rx_data_5__bdd_4_lut_25621 (.A(\rx_data[5] ), .B(\rx_data[0] ), 
         .C(\rx_data[1] ), .D(\rx_data[2] ), .Z(n47)) /* synthesis lut_function=(!(A+!(B (C)+!B !(C (D)+!C !(D))))) */ ;
    defparam rx_data_5__bdd_4_lut_25621.init = 16'h4150;
    LUT4 rx_data_3__bdd_3_lut (.A(\rx_data[0] ), .B(\rx_data[4] ), .C(\rx_data[1] ), 
         .Z(n24305)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam rx_data_3__bdd_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_adj_125 (.A(dec_bits[4]), .B(dec_bits_c[3]), .Z(n45)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(60[9] 100[5])
    defparam i1_2_lut_adj_125.init = 16'h4444;
    LUT4 i1_2_lut_adj_126 (.A(dec_bits[4]), .B(dec_bits_c[2]), .Z(n46)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(60[9] 100[5])
    defparam i1_2_lut_adj_126.init = 16'h4444;
    LUT4 n24303_bdd_3_lut (.A(n24303), .B(n24300), .C(\rx_data[1] ), .Z(n24304)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n24303_bdd_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_769 (.A(\rx_data[2] ), .B(\rx_data[1] ), .Z(n26729)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(65[3] 99[10])
    defparam i1_2_lut_rep_769.init = 16'heeee;
    LUT4 n47_bdd_1_lut_2_lut_3_lut_4_lut (.A(\rx_data[2] ), .B(\rx_data[1] ), 
         .C(n19617), .D(\rx_data[3] ), .Z(n25658)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(65[3] 99[10])
    defparam n47_bdd_1_lut_2_lut_3_lut_4_lut.init = 16'hef0f;
    LUT4 i1_2_lut_rep_606 (.A(n29268), .B(dec_stb), .Z(dac_clk_p_c_enable_380)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(53[9] 54[46])
    defparam i1_2_lut_rep_606.init = 16'heeee;
    LUT4 i8111_2_lut_3_lut (.A(n29268), .B(dec_stb), .C(dec_bits[4]), 
         .Z(dac_clk_p_c_enable_349)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(53[9] 54[46])
    defparam i8111_2_lut_3_lut.init = 16'he0e0;
    LUT4 i83_4_lut_then_4_lut (.A(\rx_data[2] ), .B(\rx_data[4] ), .C(\rx_data[5] ), 
         .D(\rx_data[1] ), .Z(n26830)) /* synthesis lut_function=(!(A (B+!((D)+!C))+!A (C+!(D)))) */ ;
    defparam i83_4_lut_then_4_lut.init = 16'h2702;
    PFUMX i25622 (.BLUT(n28307), .ALUT(n28306), .C0(\rx_data[4] ), .Z(n28308));
    LUT4 i83_4_lut_else_4_lut (.A(\rx_data[2] ), .B(\rx_data[4] ), .C(\rx_data[5] ), 
         .D(\rx_data[1] ), .Z(n26829)) /* synthesis lut_function=(!(A (B+(C))+!A (B+(C (D))))) */ ;
    defparam i83_4_lut_else_4_lut.init = 16'h0313;
    LUT4 n47_bdd_4_lut_then_4_lut (.A(\rx_data[4] ), .B(\rx_data[5] ), .C(\rx_data[2] ), 
         .D(\rx_data[0] ), .Z(n26839)) /* synthesis lut_function=(A+((C (D))+!B)) */ ;
    defparam n47_bdd_4_lut_then_4_lut.init = 16'hfbbb;
    LUT4 n47_bdd_4_lut_else_4_lut (.A(\rx_data[4] ), .B(\rx_data[5] ), .C(\rx_data[2] ), 
         .D(\rx_data[0] ), .Z(n26838)) /* synthesis lut_function=(A+!(B (C+(D)))) */ ;
    defparam n47_bdd_4_lut_else_4_lut.init = 16'hbbbf;
    LUT4 i17498_2_lut_3_lut_4_lut (.A(\rx_data[3] ), .B(n26729), .C(\rx_data[6] ), 
         .D(n19617), .Z(n19683)) /* synthesis lut_function=(A (B (C)+!B (C+(D)))+!A (C+(D))) */ ;
    defparam i17498_2_lut_3_lut_4_lut.init = 16'hf7f0;
    LUT4 i1_2_lut_3_lut (.A(dec_stb), .B(dec_bits[4]), .C(cmd_loaded), 
         .Z(o_pck_stb_N_765)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(60[9] 100[5])
    defparam i1_2_lut_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_127 (.A(dec_stb), .B(dec_bits[4]), .C(n29268), 
         .Z(dac_clk_p_c_enable_196)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(60[9] 100[5])
    defparam i1_2_lut_3_lut_adj_127.init = 16'hf8f8;
    LUT4 i2_3_lut_4_lut (.A(dec_stb), .B(dec_bits[4]), .C(dec_bits_c[2]), 
         .D(dec_bits_c[3]), .Z(cmd_loaded_N_768)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(60[9] 100[5])
    defparam i2_3_lut_4_lut.init = 16'h0008;
    LUT4 i1_3_lut_rep_570 (.A(n47), .B(\rx_data[3] ), .C(\rx_data[4] ), 
         .Z(n26530)) /* synthesis lut_function=(A (B)+!A (B+(C))) */ ;
    defparam i1_3_lut_rep_570.init = 16'hdcdc;
    LUT4 i1_3_lut_4_lut (.A(\rx_data[2] ), .B(\rx_data[1] ), .C(\rx_data[6] ), 
         .D(\rx_data[3] ), .Z(n43)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(65[3] 99[10])
    defparam i1_3_lut_4_lut.init = 16'hfe00;
    LUT4 i11944_2_lut_3_lut (.A(\rx_data[1] ), .B(\rx_data[2] ), .C(\rx_data[0] ), 
         .Z(n14504)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i11944_2_lut_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_4_lut (.A(n47), .B(\rx_data[3] ), .C(\rx_data[4] ), 
         .D(\rx_data[6] ), .Z(n52)) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C (D)))) */ ;
    defparam i1_2_lut_4_lut.init = 16'hdc00;
    LUT4 i1_3_lut_then_4_lut (.A(\rx_data[4] ), .B(\rx_data[2] ), .C(\rx_data[0] ), 
         .D(\rx_data[5] ), .Z(n26853)) /* synthesis lut_function=(A+!(B (C+!(D))+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(65[3] 99[10])
    defparam i1_3_lut_then_4_lut.init = 16'hbfaa;
    LUT4 i1_3_lut_else_4_lut (.A(\rx_data[4] ), .B(\rx_data[2] ), .C(\rx_data[0] ), 
         .D(\rx_data[5] ), .Z(n26852)) /* synthesis lut_function=(A+(B (D)+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(65[3] 99[10])
    defparam i1_3_lut_else_4_lut.init = 16'hfeba;
    LUT4 rx_data_3__bdd_3_lut_22728 (.A(\rx_data[0] ), .B(\rx_data[6] ), 
         .C(\rx_data[4] ), .Z(n24302)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam rx_data_3__bdd_3_lut_22728.init = 16'h2020;
    LUT4 rx_data_4__bdd_3_lut_4_lut (.A(\rx_data[5] ), .B(\rx_data[6] ), 
         .C(\rx_data[3] ), .D(\rx_data[4] ), .Z(n20446)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam rx_data_4__bdd_3_lut_4_lut.init = 16'h0008;
    LUT4 rx_data_3__bdd_4_lut_22725 (.A(\rx_data[3] ), .B(\rx_data[0] ), 
         .C(\rx_data[6] ), .D(\rx_data[4] ), .Z(n24300)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B ((D)+!C)))) */ ;
    defparam rx_data_3__bdd_4_lut_22725.init = 16'h0410;
    
endmodule
//
// Verilog Description of module hbnewline
//

module hbnewline (tx_busy, o_busy_N_536, \state[0] , n17598, dac_clk_p_c, 
            n29269, w_reset, hx_stb, nl_busy, \w_gx_char[2] , \w_gx_char[0] , 
            n26540, \lcl_data[1] , \lcl_data_7__N_511[0] , \lcl_data[4] , 
            \lcl_data_7__N_511[3] , \lcl_data[5] , \lcl_data_7__N_511[4] , 
            \lcl_data[6] , \lcl_data_7__N_511[5] , \lcl_data[7] , \lcl_data_7__N_511[6] , 
            zero_baud_counter, dac_clk_p_c_enable_321, \lcl_data[3] , 
            \lcl_data_7__N_511[2] , \lcl_data[2] , \lcl_data_7__N_511[1] , 
            \w_gx_char[4] , n29268, \w_gx_char[3] , \w_gx_char[5] , 
            \w_gx_char[1] , \w_gx_char[6] , n11652) /* synthesis syn_module_defined=1 */ ;
    input tx_busy;
    input o_busy_N_536;
    input \state[0] ;
    output n17598;
    input dac_clk_p_c;
    input n29269;
    input w_reset;
    input hx_stb;
    output nl_busy;
    input \w_gx_char[2] ;
    input \w_gx_char[0] ;
    output n26540;
    input \lcl_data[1] ;
    output \lcl_data_7__N_511[0] ;
    input \lcl_data[4] ;
    output \lcl_data_7__N_511[3] ;
    input \lcl_data[5] ;
    output \lcl_data_7__N_511[4] ;
    input \lcl_data[6] ;
    output \lcl_data_7__N_511[5] ;
    input \lcl_data[7] ;
    output \lcl_data_7__N_511[6] ;
    input zero_baud_counter;
    output dac_clk_p_c_enable_321;
    input \lcl_data[3] ;
    output \lcl_data_7__N_511[2] ;
    input \lcl_data[2] ;
    output \lcl_data_7__N_511[1] ;
    input \w_gx_char[4] ;
    input n29268;
    input \w_gx_char[3] ;
    input \w_gx_char[5] ;
    input \w_gx_char[1] ;
    input \w_gx_char[6] ;
    input n11652;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(29[49:58])
    
    wire tx_stb, last_cr, last_cr_N_1323, o_nl_stb_N_1315;
    wire [7:0]tx_data;   // d:/documents/git_local/fm_modulator/rtl/top.v(60[12:19])
    
    wire dac_clk_p_c_enable_199;
    wire [6:0]o_nl_byte_6__N_1302;
    wire [6:0]o_nl_byte_6__N_1295;
    
    wire cr_state, cr_state_N_1331, loaded, n26404, n26846, n26847, 
        n25431, n25430;
    wire [6:0]n32;
    
    wire n26520;
    
    LUT4 state_544_mux_6_i1_3_lut_4_lut (.A(tx_stb), .B(tx_busy), .C(o_busy_N_536), 
         .D(\state[0] ), .Z(n17598)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam state_544_mux_6_i1_3_lut_4_lut.init = 16'hd0df;
    FD1S3JX last_cr_45 (.D(last_cr_N_1323), .CK(dac_clk_p_c), .PD(n29269), 
            .Q(last_cr)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=12, LSE_RCOL=40, LSE_LLINE=138, LSE_RLINE=139 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam last_cr_45.GSR = "DISABLED";
    FD1S3IX o_nl_stb_46 (.D(o_nl_stb_N_1315), .CK(dac_clk_p_c), .CD(n29269), 
            .Q(tx_stb)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=12, LSE_RCOL=40, LSE_LLINE=138, LSE_RLINE=139 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam o_nl_stb_46.GSR = "DISABLED";
    FD1P3JX o_nl_byte_i2 (.D(o_nl_byte_6__N_1302[1]), .SP(dac_clk_p_c_enable_199), 
            .PD(w_reset), .CK(dac_clk_p_c), .Q(tx_data[1])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=12, LSE_RCOL=40, LSE_LLINE=138, LSE_RLINE=139 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam o_nl_byte_i2.GSR = "DISABLED";
    FD1P3JX o_nl_byte_i3 (.D(o_nl_byte_6__N_1302[2]), .SP(dac_clk_p_c_enable_199), 
            .PD(w_reset), .CK(dac_clk_p_c), .Q(tx_data[2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=12, LSE_RCOL=40, LSE_LLINE=138, LSE_RLINE=139 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam o_nl_byte_i3.GSR = "DISABLED";
    FD1P3AY o_nl_byte_i4 (.D(o_nl_byte_6__N_1295[3]), .SP(dac_clk_p_c_enable_199), 
            .CK(dac_clk_p_c), .Q(tx_data[3])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=12, LSE_RCOL=40, LSE_LLINE=138, LSE_RLINE=139 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam o_nl_byte_i4.GSR = "DISABLED";
    FD1P3JX o_nl_byte_i5 (.D(o_nl_byte_6__N_1302[4]), .SP(dac_clk_p_c_enable_199), 
            .PD(w_reset), .CK(dac_clk_p_c), .Q(tx_data[4])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=12, LSE_RCOL=40, LSE_LLINE=138, LSE_RLINE=139 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam o_nl_byte_i5.GSR = "DISABLED";
    FD1P3JX o_nl_byte_i6 (.D(o_nl_byte_6__N_1302[5]), .SP(dac_clk_p_c_enable_199), 
            .PD(w_reset), .CK(dac_clk_p_c), .Q(tx_data[5])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=12, LSE_RCOL=40, LSE_LLINE=138, LSE_RLINE=139 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam o_nl_byte_i6.GSR = "DISABLED";
    FD1P3JX o_nl_byte_i7 (.D(o_nl_byte_6__N_1302[6]), .SP(dac_clk_p_c_enable_199), 
            .PD(w_reset), .CK(dac_clk_p_c), .Q(tx_data[6])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=12, LSE_RCOL=40, LSE_LLINE=138, LSE_RLINE=139 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam o_nl_byte_i7.GSR = "DISABLED";
    FD1P3IX cr_state_44 (.D(cr_state_N_1331), .SP(dac_clk_p_c_enable_199), 
            .CD(n29269), .CK(dac_clk_p_c), .Q(cr_state)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=12, LSE_RCOL=40, LSE_LLINE=138, LSE_RLINE=139 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam cr_state_44.GSR = "DISABLED";
    FD1P3IX loaded_47 (.D(n26404), .SP(dac_clk_p_c_enable_199), .CD(n29269), 
            .CK(dac_clk_p_c), .Q(loaded)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=12, LSE_RCOL=40, LSE_LLINE=138, LSE_RLINE=139 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam loaded_47.GSR = "DISABLED";
    FD1P3JX o_nl_byte_i1 (.D(o_nl_byte_6__N_1302[0]), .SP(dac_clk_p_c_enable_199), 
            .PD(n29269), .CK(dac_clk_p_c), .Q(tx_data[0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=12, LSE_RCOL=40, LSE_LLINE=138, LSE_RLINE=139 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam o_nl_byte_i1.GSR = "DISABLED";
    PFUMX i24533 (.BLUT(n26846), .ALUT(n26847), .C0(last_cr), .Z(last_cr_N_1323));
    LUT4 tx_stb_bdd_3_lut (.A(hx_stb), .B(last_cr), .C(cr_state), .Z(n25431)) /* synthesis lut_function=(A (B+!(C))+!A ((C)+!B)) */ ;
    defparam tx_stb_bdd_3_lut.init = 16'hdbdb;
    LUT4 tx_stb_bdd_2_lut (.A(tx_stb), .B(hx_stb), .Z(n25430)) /* synthesis lut_function=(A+(B)) */ ;
    defparam tx_stb_bdd_2_lut.init = 16'heeee;
    LUT4 i1_2_lut (.A(last_cr), .B(cr_state), .Z(n32[4])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam i1_2_lut.init = 16'h2222;
    LUT4 i_stb_I_0_2_lut_rep_560 (.A(hx_stb), .B(nl_busy), .Z(n26520)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(90[16:37])
    defparam i_stb_I_0_2_lut_rep_560.init = 16'h2222;
    LUT4 i1_3_lut_4_lut (.A(last_cr), .B(n26520), .C(cr_state), .D(\w_gx_char[2] ), 
         .Z(o_nl_byte_6__N_1302[2])) /* synthesis lut_function=(A (B (D)+!B !(C))+!A ((D)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(97[12] 120[6])
    defparam i1_3_lut_4_lut.init = 16'hdf13;
    LUT4 i1_3_lut_4_lut_adj_114 (.A(last_cr), .B(n26520), .C(cr_state), 
         .D(\w_gx_char[0] ), .Z(o_nl_byte_6__N_1302[0])) /* synthesis lut_function=(A (B (D)+!B !(C))+!A ((D)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(97[12] 120[6])
    defparam i1_3_lut_4_lut_adj_114.init = 16'hdf13;
    LUT4 i1_2_lut_rep_580 (.A(tx_stb), .B(tx_busy), .Z(n26540)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam i1_2_lut_rep_580.init = 16'h2222;
    LUT4 lcl_data_7__I_0_i1_3_lut_4_lut (.A(tx_stb), .B(tx_busy), .C(tx_data[0]), 
         .D(\lcl_data[1] ), .Z(\lcl_data_7__N_511[0] )) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam lcl_data_7__I_0_i1_3_lut_4_lut.init = 16'hfd20;
    LUT4 lcl_data_7__I_0_i4_3_lut_4_lut (.A(tx_stb), .B(tx_busy), .C(tx_data[3]), 
         .D(\lcl_data[4] ), .Z(\lcl_data_7__N_511[3] )) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam lcl_data_7__I_0_i4_3_lut_4_lut.init = 16'hfd20;
    LUT4 lcl_data_7__I_0_i5_3_lut_4_lut (.A(tx_stb), .B(tx_busy), .C(tx_data[4]), 
         .D(\lcl_data[5] ), .Z(\lcl_data_7__N_511[4] )) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam lcl_data_7__I_0_i5_3_lut_4_lut.init = 16'hfd20;
    LUT4 lcl_data_7__I_0_i6_3_lut_4_lut (.A(tx_stb), .B(tx_busy), .C(tx_data[5]), 
         .D(\lcl_data[6] ), .Z(\lcl_data_7__N_511[5] )) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam lcl_data_7__I_0_i6_3_lut_4_lut.init = 16'hfd20;
    LUT4 lcl_data_7__I_0_i7_3_lut_4_lut (.A(tx_stb), .B(tx_busy), .C(tx_data[6]), 
         .D(\lcl_data[7] ), .Z(\lcl_data_7__N_511[6] )) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam lcl_data_7__I_0_i7_3_lut_4_lut.init = 16'hfd20;
    LUT4 i559_2_lut_3_lut (.A(tx_stb), .B(tx_busy), .C(zero_baud_counter), 
         .Z(dac_clk_p_c_enable_321)) /* synthesis lut_function=(A ((C)+!B)+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam i559_2_lut_3_lut.init = 16'hf2f2;
    LUT4 lcl_data_7__I_0_i3_3_lut_4_lut (.A(tx_stb), .B(tx_busy), .C(tx_data[2]), 
         .D(\lcl_data[3] ), .Z(\lcl_data_7__N_511[2] )) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam lcl_data_7__I_0_i3_3_lut_4_lut.init = 16'hfd20;
    LUT4 lcl_data_7__I_0_i2_3_lut_4_lut (.A(tx_stb), .B(tx_busy), .C(tx_data[1]), 
         .D(\lcl_data[2] ), .Z(\lcl_data_7__N_511[1] )) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam lcl_data_7__I_0_i2_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_24_i5_3_lut_4_lut (.A(hx_stb), .B(nl_busy), .C(\w_gx_char[4] ), 
         .D(n32[4]), .Z(o_nl_byte_6__N_1302[4])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(90[16:37])
    defparam mux_24_i5_3_lut_4_lut.init = 16'hfd20;
    LUT4 i1_3_lut_4_lut_adj_115 (.A(hx_stb), .B(nl_busy), .C(n29268), 
         .D(\w_gx_char[3] ), .Z(o_nl_byte_6__N_1295[3])) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(90[16:37])
    defparam i1_3_lut_4_lut_adj_115.init = 16'hfffd;
    LUT4 i1_3_lut_4_lut_adj_116 (.A(hx_stb), .B(nl_busy), .C(n29268), 
         .D(tx_busy), .Z(dac_clk_p_c_enable_199)) /* synthesis lut_function=(A ((C+!(D))+!B)+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(90[16:37])
    defparam i1_3_lut_4_lut_adj_116.init = 16'hf2ff;
    LUT4 i11050_3_lut_rep_444_4_lut (.A(hx_stb), .B(nl_busy), .C(cr_state), 
         .D(last_cr), .Z(n26404)) /* synthesis lut_function=(A ((C (D))+!B)+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(90[16:37])
    defparam i11050_3_lut_rep_444_4_lut.init = 16'hf222;
    LUT4 i10804_3_lut_4_lut (.A(hx_stb), .B(nl_busy), .C(\w_gx_char[5] ), 
         .D(n32[4]), .Z(o_nl_byte_6__N_1302[5])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(90[16:37])
    defparam i10804_3_lut_4_lut.init = 16'hfd20;
    LUT4 i10807_3_lut_4_lut (.A(hx_stb), .B(nl_busy), .C(\w_gx_char[1] ), 
         .D(last_cr), .Z(o_nl_byte_6__N_1302[1])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(90[16:37])
    defparam i10807_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_24_i7_3_lut_4_lut (.A(hx_stb), .B(nl_busy), .C(\w_gx_char[6] ), 
         .D(n32[4]), .Z(o_nl_byte_6__N_1302[6])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(90[16:37])
    defparam mux_24_i7_3_lut_4_lut.init = 16'hfd20;
    LUT4 cr_state_I_41_3_lut_4_lut (.A(hx_stb), .B(nl_busy), .C(n11652), 
         .D(last_cr), .Z(cr_state_N_1331)) /* synthesis lut_function=(!(A (B (D)+!B (C))+!A (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(90[16:37])
    defparam cr_state_I_41_3_lut_4_lut.init = 16'h02df;
    LUT4 i20837_4_lut (.A(cr_state), .B(tx_stb), .C(tx_busy), .D(loaded), 
         .Z(nl_busy)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(123[21] 124[30])
    defparam i20837_4_lut.init = 16'hca0a;
    LUT4 last_cr_I_39_4_lut_then_3_lut (.A(n11652), .B(hx_stb), .C(nl_busy), 
         .Z(n26847)) /* synthesis lut_function=(((C)+!B)+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(97[12] 120[6])
    defparam last_cr_I_39_4_lut_then_3_lut.init = 16'hf7f7;
    LUT4 last_cr_I_39_4_lut_else_3_lut (.A(n11652), .B(tx_busy), .C(hx_stb), 
         .D(nl_busy), .Z(n26846)) /* synthesis lut_function=(!(A (B+(C))+!A (B ((D)+!C)+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(97[12] 120[6])
    defparam last_cr_I_39_4_lut_else_3_lut.init = 16'h0353;
    PFUMX i23748 (.BLUT(n25431), .ALUT(n25430), .C0(tx_busy), .Z(o_nl_stb_N_1315));
    
endmodule
//
// Verilog Description of module hbints
//

module hbints (int_word, dac_clk_p_c, ow_word, n29268, n26742, int_stb, 
            ow_stb, n29269) /* synthesis syn_module_defined=1 */ ;
    output [33:0]int_word;
    input dac_clk_p_c;
    input [33:0]ow_word;
    input n29268;
    input n26742;
    output int_stb;
    input ow_stb;
    input n29269;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(29[49:58])
    
    wire dac_clk_p_c_enable_416, n12645, n26574, dac_clk_p_c_enable_410, 
        loaded, dac_clk_p_c_enable_409;
    
    FD1P3IX o_int_word_i10 (.D(ow_word[10]), .SP(dac_clk_p_c_enable_416), 
            .CD(n12645), .CK(dac_clk_p_c), .Q(int_word[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i10.GSR = "DISABLED";
    FD1P3JX o_int_word_i33 (.D(ow_word[33]), .SP(dac_clk_p_c_enable_416), 
            .PD(n12645), .CK(dac_clk_p_c), .Q(int_word[33])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i33.GSR = "DISABLED";
    LUT4 i1_2_lut_3_lut_4_lut (.A(n29268), .B(n26574), .C(n26742), .D(int_stb), 
         .Z(dac_clk_p_c_enable_410)) /* synthesis lut_function=(A+(B+!(C+!(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'hefee;
    LUT4 i1_3_lut_4_lut (.A(n29268), .B(n26574), .C(loaded), .D(n26742), 
         .Z(dac_clk_p_c_enable_409)) /* synthesis lut_function=(A+(B+!(C (D)))) */ ;
    defparam i1_3_lut_4_lut.init = 16'hefff;
    FD1P3JX o_int_word_i32 (.D(ow_word[32]), .SP(dac_clk_p_c_enable_416), 
            .PD(n12645), .CK(dac_clk_p_c), .Q(int_word[32])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i32.GSR = "DISABLED";
    LUT4 i_stb_I_0_3_lut_rep_614 (.A(ow_stb), .B(int_stb), .C(loaded), 
         .Z(n26574)) /* synthesis lut_function=(!((B (C))+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(93[12:34])
    defparam i_stb_I_0_3_lut_rep_614.init = 16'h2a2a;
    LUT4 i1_2_lut_3_lut_4_lut_adj_113 (.A(ow_stb), .B(int_stb), .C(loaded), 
         .D(n26742), .Z(dac_clk_p_c_enable_416)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(93[12:34])
    defparam i1_2_lut_3_lut_4_lut_adj_113.init = 16'h3bff;
    LUT4 i22384_2_lut_3_lut_4_lut (.A(ow_stb), .B(int_stb), .C(loaded), 
         .D(n26742), .Z(n12645)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A (B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(93[12:34])
    defparam i22384_2_lut_3_lut_4_lut.init = 16'h11d5;
    FD1P3IX o_int_word_i9 (.D(ow_word[9]), .SP(dac_clk_p_c_enable_416), 
            .CD(n12645), .CK(dac_clk_p_c), .Q(int_word[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i9.GSR = "DISABLED";
    FD1P3IX o_int_word_i31 (.D(ow_word[31]), .SP(dac_clk_p_c_enable_416), 
            .CD(n12645), .CK(dac_clk_p_c), .Q(int_word[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i31.GSR = "DISABLED";
    FD1P3JX o_int_word_i30 (.D(ow_word[30]), .SP(dac_clk_p_c_enable_416), 
            .PD(n12645), .CK(dac_clk_p_c), .Q(int_word[30])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i30.GSR = "DISABLED";
    FD1P3IX o_int_word_i29 (.D(ow_word[29]), .SP(dac_clk_p_c_enable_416), 
            .CD(n12645), .CK(dac_clk_p_c), .Q(int_word[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i29.GSR = "DISABLED";
    FD1P3IX o_int_word_i8 (.D(ow_word[8]), .SP(dac_clk_p_c_enable_416), 
            .CD(n12645), .CK(dac_clk_p_c), .Q(int_word[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i8.GSR = "DISABLED";
    FD1P3IX o_int_word_i28 (.D(ow_word[28]), .SP(dac_clk_p_c_enable_416), 
            .CD(n12645), .CK(dac_clk_p_c), .Q(int_word[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i28.GSR = "DISABLED";
    FD1P3IX o_int_word_i7 (.D(ow_word[7]), .SP(dac_clk_p_c_enable_416), 
            .CD(n12645), .CK(dac_clk_p_c), .Q(int_word[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i7.GSR = "DISABLED";
    FD1P3IX o_int_word_i27 (.D(ow_word[27]), .SP(dac_clk_p_c_enable_416), 
            .CD(n12645), .CK(dac_clk_p_c), .Q(int_word[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i27.GSR = "DISABLED";
    FD1P3IX o_int_word_i6 (.D(ow_word[6]), .SP(dac_clk_p_c_enable_416), 
            .CD(n12645), .CK(dac_clk_p_c), .Q(int_word[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i6.GSR = "DISABLED";
    FD1P3IX o_int_word_i5 (.D(ow_word[5]), .SP(dac_clk_p_c_enable_416), 
            .CD(n12645), .CK(dac_clk_p_c), .Q(int_word[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i5.GSR = "DISABLED";
    FD1P3IX o_int_word_i26 (.D(ow_word[26]), .SP(dac_clk_p_c_enable_416), 
            .CD(n12645), .CK(dac_clk_p_c), .Q(int_word[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i26.GSR = "DISABLED";
    FD1P3IX o_int_word_i25 (.D(ow_word[25]), .SP(dac_clk_p_c_enable_416), 
            .CD(n12645), .CK(dac_clk_p_c), .Q(int_word[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i25.GSR = "DISABLED";
    FD1P3IX o_int_word_i4 (.D(ow_word[4]), .SP(dac_clk_p_c_enable_416), 
            .CD(n12645), .CK(dac_clk_p_c), .Q(int_word[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i4.GSR = "DISABLED";
    FD1P3IX o_int_word_i24 (.D(ow_word[24]), .SP(dac_clk_p_c_enable_416), 
            .CD(n12645), .CK(dac_clk_p_c), .Q(int_word[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i24.GSR = "DISABLED";
    FD1P3IX o_int_word_i3 (.D(ow_word[3]), .SP(dac_clk_p_c_enable_416), 
            .CD(n12645), .CK(dac_clk_p_c), .Q(int_word[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i3.GSR = "DISABLED";
    FD1P3IX o_int_word_i23 (.D(ow_word[23]), .SP(dac_clk_p_c_enable_416), 
            .CD(n12645), .CK(dac_clk_p_c), .Q(int_word[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i23.GSR = "DISABLED";
    FD1P3IX o_int_word_i2 (.D(ow_word[2]), .SP(dac_clk_p_c_enable_416), 
            .CD(n12645), .CK(dac_clk_p_c), .Q(int_word[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i2.GSR = "DISABLED";
    FD1P3IX o_int_word_i1 (.D(ow_word[1]), .SP(dac_clk_p_c_enable_416), 
            .CD(n12645), .CK(dac_clk_p_c), .Q(int_word[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i1.GSR = "DISABLED";
    FD1P3IX o_int_word_i22 (.D(ow_word[22]), .SP(dac_clk_p_c_enable_416), 
            .CD(n12645), .CK(dac_clk_p_c), .Q(int_word[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i22.GSR = "DISABLED";
    FD1P3IX o_int_word_i21 (.D(ow_word[21]), .SP(dac_clk_p_c_enable_416), 
            .CD(n12645), .CK(dac_clk_p_c), .Q(int_word[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i21.GSR = "DISABLED";
    FD1P3IX o_int_word_i0 (.D(ow_word[0]), .SP(dac_clk_p_c_enable_416), 
            .CD(n12645), .CK(dac_clk_p_c), .Q(int_word[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i0.GSR = "DISABLED";
    FD1P3IX o_int_word_i20 (.D(ow_word[20]), .SP(dac_clk_p_c_enable_416), 
            .CD(n12645), .CK(dac_clk_p_c), .Q(int_word[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i20.GSR = "DISABLED";
    FD1P3IX o_int_word_i19 (.D(ow_word[19]), .SP(dac_clk_p_c_enable_416), 
            .CD(n12645), .CK(dac_clk_p_c), .Q(int_word[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i19.GSR = "DISABLED";
    FD1P3IX o_int_word_i18 (.D(ow_word[18]), .SP(dac_clk_p_c_enable_416), 
            .CD(n12645), .CK(dac_clk_p_c), .Q(int_word[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i18.GSR = "DISABLED";
    FD1P3IX o_int_word_i17 (.D(ow_word[17]), .SP(dac_clk_p_c_enable_416), 
            .CD(n12645), .CK(dac_clk_p_c), .Q(int_word[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i17.GSR = "DISABLED";
    FD1P3IX o_int_word_i16 (.D(ow_word[16]), .SP(dac_clk_p_c_enable_416), 
            .CD(n12645), .CK(dac_clk_p_c), .Q(int_word[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i16.GSR = "DISABLED";
    FD1P3IX o_int_word_i15 (.D(ow_word[15]), .SP(dac_clk_p_c_enable_416), 
            .CD(n12645), .CK(dac_clk_p_c), .Q(int_word[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i15.GSR = "DISABLED";
    FD1P3IX o_int_stb_58 (.D(n26574), .SP(dac_clk_p_c_enable_409), .CD(n29269), 
            .CK(dac_clk_p_c), .Q(int_stb)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(90[9] 98[22])
    defparam o_int_stb_58.GSR = "DISABLED";
    FD1P3IX loaded_57 (.D(n26574), .SP(dac_clk_p_c_enable_410), .CD(n29269), 
            .CK(dac_clk_p_c), .Q(loaded)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(81[9] 87[19])
    defparam loaded_57.GSR = "DISABLED";
    FD1P3IX o_int_word_i14 (.D(ow_word[14]), .SP(dac_clk_p_c_enable_416), 
            .CD(n12645), .CK(dac_clk_p_c), .Q(int_word[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i14.GSR = "DISABLED";
    FD1P3IX o_int_word_i13 (.D(ow_word[13]), .SP(dac_clk_p_c_enable_416), 
            .CD(n12645), .CK(dac_clk_p_c), .Q(int_word[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i13.GSR = "DISABLED";
    FD1P3IX o_int_word_i12 (.D(ow_word[12]), .SP(dac_clk_p_c_enable_416), 
            .CD(n12645), .CK(dac_clk_p_c), .Q(int_word[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i12.GSR = "DISABLED";
    FD1P3IX o_int_word_i11 (.D(ow_word[11]), .SP(dac_clk_p_c_enable_416), 
            .CD(n12645), .CK(dac_clk_p_c), .Q(int_word[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i11.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module hbidle
//

module hbidle (idl_word, dac_clk_p_c, int_word, hb_busy, int_stb, 
            idl_stb, n29268, w_reset, n26742) /* synthesis syn_module_defined=1 */ ;
    output [33:0]idl_word;
    input dac_clk_p_c;
    input [33:0]int_word;
    input hb_busy;
    input int_stb;
    output idl_stb;
    input n29268;
    input w_reset;
    output n26742;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(29[49:58])
    
    wire dac_clk_p_c_enable_403, n12674, dac_clk_p_c_enable_194, n26422;
    
    FD1P3IX o_idl_word_i10 (.D(int_word[10]), .SP(dac_clk_p_c_enable_403), 
            .CD(n12674), .CK(dac_clk_p_c), .Q(idl_word[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i10.GSR = "DISABLED";
    FD1P3IX o_idl_word_i9 (.D(int_word[9]), .SP(dac_clk_p_c_enable_403), 
            .CD(n12674), .CK(dac_clk_p_c), .Q(idl_word[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i9.GSR = "DISABLED";
    LUT4 i22417_2_lut (.A(hb_busy), .B(int_stb), .Z(n12674)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i22417_2_lut.init = 16'h1111;
    FD1P3IX o_idl_word_i8 (.D(int_word[8]), .SP(dac_clk_p_c_enable_403), 
            .CD(n12674), .CK(dac_clk_p_c), .Q(idl_word[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i8.GSR = "DISABLED";
    LUT4 i1_3_lut_4_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(n29268), .D(int_stb), 
         .Z(dac_clk_p_c_enable_194)) /* synthesis lut_function=(A ((C)+!B)+!A ((C+(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(97[22:43])
    defparam i1_3_lut_4_lut_4_lut.init = 16'hf7f3;
    FD1P3IX o_idl_word_i7 (.D(int_word[7]), .SP(dac_clk_p_c_enable_403), 
            .CD(n12674), .CK(dac_clk_p_c), .Q(idl_word[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i7.GSR = "DISABLED";
    FD1P3IX o_idl_word_i6 (.D(int_word[6]), .SP(dac_clk_p_c_enable_403), 
            .CD(n12674), .CK(dac_clk_p_c), .Q(idl_word[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i6.GSR = "DISABLED";
    FD1P3IX o_idl_word_i5 (.D(int_word[5]), .SP(dac_clk_p_c_enable_403), 
            .CD(n12674), .CK(dac_clk_p_c), .Q(idl_word[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i5.GSR = "DISABLED";
    LUT4 i1_2_lut_3_lut_3_lut (.A(idl_stb), .B(hb_busy), .C(int_stb), 
         .Z(dac_clk_p_c_enable_403)) /* synthesis lut_function=(!(A (B)+!A !((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(97[22:43])
    defparam i1_2_lut_3_lut_3_lut.init = 16'h7373;
    FD1P3IX o_idl_stb_28 (.D(n26422), .SP(dac_clk_p_c_enable_194), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(idl_stb)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(80[9] 88[22])
    defparam o_idl_stb_28.GSR = "DISABLED";
    FD1P3JX o_idl_word_i33 (.D(int_word[33]), .SP(dac_clk_p_c_enable_403), 
            .PD(n12674), .CK(dac_clk_p_c), .Q(idl_word[33])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i33.GSR = "DISABLED";
    FD1P3JX o_idl_word_i32 (.D(int_word[32]), .SP(dac_clk_p_c_enable_403), 
            .PD(n12674), .CK(dac_clk_p_c), .Q(idl_word[32])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i32.GSR = "DISABLED";
    FD1P3IX o_idl_word_i31 (.D(int_word[31]), .SP(dac_clk_p_c_enable_403), 
            .CD(n12674), .CK(dac_clk_p_c), .Q(idl_word[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i31.GSR = "DISABLED";
    FD1P3JX o_idl_word_i30 (.D(int_word[30]), .SP(dac_clk_p_c_enable_403), 
            .PD(n12674), .CK(dac_clk_p_c), .Q(idl_word[30])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i30.GSR = "DISABLED";
    FD1P3JX o_idl_word_i29 (.D(int_word[29]), .SP(dac_clk_p_c_enable_403), 
            .PD(n12674), .CK(dac_clk_p_c), .Q(idl_word[29])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i29.GSR = "DISABLED";
    FD1P3IX o_idl_word_i28 (.D(int_word[28]), .SP(dac_clk_p_c_enable_403), 
            .CD(n12674), .CK(dac_clk_p_c), .Q(idl_word[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i28.GSR = "DISABLED";
    FD1P3IX o_idl_word_i27 (.D(int_word[27]), .SP(dac_clk_p_c_enable_403), 
            .CD(n12674), .CK(dac_clk_p_c), .Q(idl_word[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i27.GSR = "DISABLED";
    FD1P3IX o_idl_word_i26 (.D(int_word[26]), .SP(dac_clk_p_c_enable_403), 
            .CD(n12674), .CK(dac_clk_p_c), .Q(idl_word[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i26.GSR = "DISABLED";
    FD1P3IX o_idl_word_i4 (.D(int_word[4]), .SP(dac_clk_p_c_enable_403), 
            .CD(n12674), .CK(dac_clk_p_c), .Q(idl_word[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i4.GSR = "DISABLED";
    FD1P3IX o_idl_word_i3 (.D(int_word[3]), .SP(dac_clk_p_c_enable_403), 
            .CD(n12674), .CK(dac_clk_p_c), .Q(idl_word[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i3.GSR = "DISABLED";
    FD1P3IX o_idl_word_i2 (.D(int_word[2]), .SP(dac_clk_p_c_enable_403), 
            .CD(n12674), .CK(dac_clk_p_c), .Q(idl_word[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i2.GSR = "DISABLED";
    FD1P3IX o_idl_word_i1 (.D(int_word[1]), .SP(dac_clk_p_c_enable_403), 
            .CD(n12674), .CK(dac_clk_p_c), .Q(idl_word[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i1.GSR = "DISABLED";
    FD1P3IX o_idl_word_i0 (.D(int_word[0]), .SP(dac_clk_p_c_enable_403), 
            .CD(n12674), .CK(dac_clk_p_c), .Q(idl_word[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i0.GSR = "DISABLED";
    LUT4 o_idl_stb_I_0_30_2_lut_rep_782 (.A(idl_stb), .B(hb_busy), .Z(n26742)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(97[22:43])
    defparam o_idl_stb_I_0_30_2_lut_rep_782.init = 16'h8888;
    LUT4 o_int_stb_I_0_66_2_lut_rep_462_3_lut (.A(idl_stb), .B(hb_busy), 
         .C(int_stb), .Z(n26422)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(97[22:43])
    defparam o_int_stb_I_0_66_2_lut_rep_462_3_lut.init = 16'h7070;
    FD1P3IX o_idl_word_i13 (.D(int_word[13]), .SP(dac_clk_p_c_enable_403), 
            .CD(n12674), .CK(dac_clk_p_c), .Q(idl_word[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i13.GSR = "DISABLED";
    FD1P3IX o_idl_word_i25 (.D(int_word[25]), .SP(dac_clk_p_c_enable_403), 
            .CD(n12674), .CK(dac_clk_p_c), .Q(idl_word[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i25.GSR = "DISABLED";
    FD1P3IX o_idl_word_i24 (.D(int_word[24]), .SP(dac_clk_p_c_enable_403), 
            .CD(n12674), .CK(dac_clk_p_c), .Q(idl_word[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i24.GSR = "DISABLED";
    FD1P3IX o_idl_word_i23 (.D(int_word[23]), .SP(dac_clk_p_c_enable_403), 
            .CD(n12674), .CK(dac_clk_p_c), .Q(idl_word[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i23.GSR = "DISABLED";
    FD1P3IX o_idl_word_i22 (.D(int_word[22]), .SP(dac_clk_p_c_enable_403), 
            .CD(n12674), .CK(dac_clk_p_c), .Q(idl_word[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i22.GSR = "DISABLED";
    FD1P3IX o_idl_word_i21 (.D(int_word[21]), .SP(dac_clk_p_c_enable_403), 
            .CD(n12674), .CK(dac_clk_p_c), .Q(idl_word[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i21.GSR = "DISABLED";
    FD1P3IX o_idl_word_i20 (.D(int_word[20]), .SP(dac_clk_p_c_enable_403), 
            .CD(n12674), .CK(dac_clk_p_c), .Q(idl_word[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i20.GSR = "DISABLED";
    FD1P3IX o_idl_word_i19 (.D(int_word[19]), .SP(dac_clk_p_c_enable_403), 
            .CD(n12674), .CK(dac_clk_p_c), .Q(idl_word[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i19.GSR = "DISABLED";
    FD1P3IX o_idl_word_i18 (.D(int_word[18]), .SP(dac_clk_p_c_enable_403), 
            .CD(n12674), .CK(dac_clk_p_c), .Q(idl_word[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i18.GSR = "DISABLED";
    FD1P3IX o_idl_word_i17 (.D(int_word[17]), .SP(dac_clk_p_c_enable_403), 
            .CD(n12674), .CK(dac_clk_p_c), .Q(idl_word[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i17.GSR = "DISABLED";
    FD1P3IX o_idl_word_i16 (.D(int_word[16]), .SP(dac_clk_p_c_enable_403), 
            .CD(n12674), .CK(dac_clk_p_c), .Q(idl_word[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i16.GSR = "DISABLED";
    FD1P3IX o_idl_word_i15 (.D(int_word[15]), .SP(dac_clk_p_c_enable_403), 
            .CD(n12674), .CK(dac_clk_p_c), .Q(idl_word[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i15.GSR = "DISABLED";
    FD1P3IX o_idl_word_i14 (.D(int_word[14]), .SP(dac_clk_p_c_enable_403), 
            .CD(n12674), .CK(dac_clk_p_c), .Q(idl_word[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i14.GSR = "DISABLED";
    FD1P3IX o_idl_word_i12 (.D(int_word[12]), .SP(dac_clk_p_c_enable_403), 
            .CD(n12674), .CK(dac_clk_p_c), .Q(idl_word[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i12.GSR = "DISABLED";
    FD1P3IX o_idl_word_i11 (.D(int_word[11]), .SP(dac_clk_p_c_enable_403), 
            .CD(n12674), .CK(dac_clk_p_c), .Q(idl_word[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i11.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module \txuartlite(TIMING_BITS=24,CLOCKS_PER_BAUD=10000) 
//

module \txuartlite(TIMING_BITS=24,CLOCKS_PER_BAUD=10000)  (dac_clk_p_c, dac_clk_p_c_enable_321, 
            \lcl_data_7__N_511[0] , zero_baud_counter, o_wbu_uart_tx_c, 
            n26540, state, GND_net, \lcl_data[7] , n29210, \lcl_data[6] , 
            \lcl_data_7__N_511[6] , \lcl_data[5] , \lcl_data_7__N_511[5] , 
            \lcl_data[4] , \lcl_data_7__N_511[4] , \lcl_data[3] , \lcl_data_7__N_511[3] , 
            \lcl_data[2] , \lcl_data_7__N_511[2] , \lcl_data[1] , \lcl_data_7__N_511[1] , 
            o_busy_N_536, tx_busy, n17598) /* synthesis syn_module_defined=1 */ ;
    input dac_clk_p_c;
    input dac_clk_p_c_enable_321;
    input \lcl_data_7__N_511[0] ;
    output zero_baud_counter;
    output o_wbu_uart_tx_c;
    input n26540;
    output [3:0]state;
    input GND_net;
    output \lcl_data[7] ;
    input n29210;
    output \lcl_data[6] ;
    input \lcl_data_7__N_511[6] ;
    output \lcl_data[5] ;
    input \lcl_data_7__N_511[5] ;
    output \lcl_data[4] ;
    input \lcl_data_7__N_511[4] ;
    output \lcl_data[3] ;
    input \lcl_data_7__N_511[3] ;
    output \lcl_data[2] ;
    input \lcl_data_7__N_511[2] ;
    output \lcl_data[1] ;
    input \lcl_data_7__N_511[1] ;
    output o_busy_N_536;
    output tx_busy;
    input n17598;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(29[49:58])
    wire [7:0]lcl_data;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(84[12:20])
    
    wire zero_baud_counter_N_525;
    wire [23:0]baud_counter;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(82[17:29])
    wire [23:0]baud_counter_23__N_483;
    wire [3:0]state_c;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(83[12:17])
    
    wire n26779, n26778, n26534, n11421, n26782, n26781;
    wire [23:0]n108;
    
    wire n17410, n17409, n17408, n17407, n17406, n17405, n17404, 
        n17403, n17402;
    wire [23:0]n133;
    
    wire n26427, zero_baud_counter_N_528, n17401, n17400, n17399, 
        n8876;
    wire [3:0]n27;
    
    wire n20118, n20526, n20534, n20532, n20524, n20510, n20520, 
        n20522, n20512, n26783, n26780;
    
    FD1P3AY lcl_data_i0 (.D(\lcl_data_7__N_511[0] ), .SP(dac_clk_p_c_enable_321), 
            .CK(dac_clk_p_c), .Q(lcl_data[0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(139[9] 143[40])
    defparam lcl_data_i0.GSR = "DISABLED";
    FD1S3AY zero_baud_counter_49 (.D(zero_baud_counter_N_525), .CK(dac_clk_p_c), 
            .Q(zero_baud_counter)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam zero_baud_counter_49.GSR = "DISABLED";
    FD1S3AX baud_counter_i0 (.D(baud_counter_23__N_483[0]), .CK(dac_clk_p_c), 
            .Q(baud_counter[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i0.GSR = "DISABLED";
    FD1P3IX o_uart_tx_48 (.D(lcl_data[0]), .SP(dac_clk_p_c_enable_321), 
            .CD(n26540), .CK(dac_clk_p_c), .Q(o_wbu_uart_tx_c)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(154[9] 158[29])
    defparam o_uart_tx_48.GSR = "DISABLED";
    LUT4 state_544_mux_6_i3_4_lut_then_4_lut (.A(n26540), .B(state[0]), 
         .C(state_c[1]), .D(state_c[3]), .Z(n26779)) /* synthesis lut_function=(!(A (B (C+(D))+!B (D))+!A !(((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(110[14:26])
    defparam state_544_mux_6_i3_4_lut_then_4_lut.init = 16'h553f;
    LUT4 state_544_mux_6_i3_4_lut_else_4_lut (.A(n26540), .B(state[0]), 
         .C(state_c[1]), .D(state_c[3]), .Z(n26778)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A !(B (C+(D))+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(110[14:26])
    defparam state_544_mux_6_i3_4_lut_else_4_lut.init = 16'h54c0;
    LUT4 i1_2_lut_4_lut (.A(state_c[2]), .B(n26534), .C(state_c[1]), .D(zero_baud_counter), 
         .Z(n11421)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(110[14:26])
    defparam i1_2_lut_4_lut.init = 16'hff80;
    LUT4 state_544_mux_6_i4_4_lut_then_4_lut (.A(n26540), .B(state_c[2]), 
         .C(state[0]), .D(state_c[1]), .Z(n26782)) /* synthesis lut_function=(!(A (B+(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(110[14:26])
    defparam state_544_mux_6_i4_4_lut_then_4_lut.init = 16'h5557;
    LUT4 state_544_mux_6_i4_4_lut_else_4_lut (.A(state_c[2]), .B(state[0]), 
         .C(state_c[1]), .Z(n26781)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(110[14:26])
    defparam state_544_mux_6_i4_4_lut_else_4_lut.init = 16'h8080;
    FD1S3IX baud_counter_i23 (.D(n108[23]), .CK(dac_clk_p_c), .CD(n11421), 
            .Q(baud_counter[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i23.GSR = "DISABLED";
    CCU2D sub_36_add_2_25 (.A0(baud_counter[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n17410), .S0(n108[23]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_25.INIT0 = 16'h5555;
    defparam sub_36_add_2_25.INIT1 = 16'h0000;
    defparam sub_36_add_2_25.INJECT1_0 = "NO";
    defparam sub_36_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_36_add_2_23 (.A0(baud_counter[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17409), .COUT(n17410), .S0(n108[21]), 
          .S1(n108[22]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_23.INIT0 = 16'h5555;
    defparam sub_36_add_2_23.INIT1 = 16'h5555;
    defparam sub_36_add_2_23.INJECT1_0 = "NO";
    defparam sub_36_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_36_add_2_21 (.A0(baud_counter[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17408), .COUT(n17409), .S0(n108[19]), 
          .S1(n108[20]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_21.INIT0 = 16'h5555;
    defparam sub_36_add_2_21.INIT1 = 16'h5555;
    defparam sub_36_add_2_21.INJECT1_0 = "NO";
    defparam sub_36_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_36_add_2_19 (.A0(baud_counter[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17407), .COUT(n17408), .S0(n108[17]), 
          .S1(n108[18]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_19.INIT0 = 16'h5555;
    defparam sub_36_add_2_19.INIT1 = 16'h5555;
    defparam sub_36_add_2_19.INJECT1_0 = "NO";
    defparam sub_36_add_2_19.INJECT1_1 = "NO";
    FD1S3IX baud_counter_i22 (.D(n108[22]), .CK(dac_clk_p_c), .CD(n11421), 
            .Q(baud_counter[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i22.GSR = "DISABLED";
    FD1S3IX baud_counter_i21 (.D(n108[21]), .CK(dac_clk_p_c), .CD(n11421), 
            .Q(baud_counter[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i21.GSR = "DISABLED";
    FD1S3IX baud_counter_i20 (.D(n108[20]), .CK(dac_clk_p_c), .CD(n11421), 
            .Q(baud_counter[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i20.GSR = "DISABLED";
    FD1S3IX baud_counter_i19 (.D(n108[19]), .CK(dac_clk_p_c), .CD(n11421), 
            .Q(baud_counter[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i19.GSR = "DISABLED";
    FD1S3IX baud_counter_i18 (.D(n108[18]), .CK(dac_clk_p_c), .CD(n11421), 
            .Q(baud_counter[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i18.GSR = "DISABLED";
    FD1S3IX baud_counter_i17 (.D(n108[17]), .CK(dac_clk_p_c), .CD(n11421), 
            .Q(baud_counter[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i17.GSR = "DISABLED";
    FD1S3IX baud_counter_i16 (.D(n108[16]), .CK(dac_clk_p_c), .CD(n11421), 
            .Q(baud_counter[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i16.GSR = "DISABLED";
    FD1S3IX baud_counter_i15 (.D(n108[15]), .CK(dac_clk_p_c), .CD(n11421), 
            .Q(baud_counter[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i15.GSR = "DISABLED";
    FD1S3IX baud_counter_i14 (.D(n108[14]), .CK(dac_clk_p_c), .CD(n11421), 
            .Q(baud_counter[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i14.GSR = "DISABLED";
    FD1S3AX baud_counter_i13 (.D(baud_counter_23__N_483[13]), .CK(dac_clk_p_c), 
            .Q(baud_counter[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i13.GSR = "DISABLED";
    FD1S3IX baud_counter_i12 (.D(n108[12]), .CK(dac_clk_p_c), .CD(n11421), 
            .Q(baud_counter[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i12.GSR = "DISABLED";
    FD1S3IX baud_counter_i11 (.D(n108[11]), .CK(dac_clk_p_c), .CD(n11421), 
            .Q(baud_counter[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i11.GSR = "DISABLED";
    FD1S3AX baud_counter_i10 (.D(baud_counter_23__N_483[10]), .CK(dac_clk_p_c), 
            .Q(baud_counter[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i10.GSR = "DISABLED";
    FD1S3AX baud_counter_i9 (.D(baud_counter_23__N_483[9]), .CK(dac_clk_p_c), 
            .Q(baud_counter[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i9.GSR = "DISABLED";
    FD1S3AX baud_counter_i8 (.D(baud_counter_23__N_483[8]), .CK(dac_clk_p_c), 
            .Q(baud_counter[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i8.GSR = "DISABLED";
    FD1S3IX baud_counter_i7 (.D(n108[7]), .CK(dac_clk_p_c), .CD(n11421), 
            .Q(baud_counter[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i7.GSR = "DISABLED";
    FD1S3IX baud_counter_i6 (.D(n108[6]), .CK(dac_clk_p_c), .CD(n11421), 
            .Q(baud_counter[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i6.GSR = "DISABLED";
    FD1S3IX baud_counter_i5 (.D(n108[5]), .CK(dac_clk_p_c), .CD(n11421), 
            .Q(baud_counter[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i5.GSR = "DISABLED";
    FD1S3IX baud_counter_i4 (.D(n108[4]), .CK(dac_clk_p_c), .CD(n11421), 
            .Q(baud_counter[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i4.GSR = "DISABLED";
    FD1S3AX baud_counter_i3 (.D(baud_counter_23__N_483[3]), .CK(dac_clk_p_c), 
            .Q(baud_counter[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i3.GSR = "DISABLED";
    FD1S3AX baud_counter_i2 (.D(baud_counter_23__N_483[2]), .CK(dac_clk_p_c), 
            .Q(baud_counter[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i2.GSR = "DISABLED";
    FD1S3AX baud_counter_i1 (.D(baud_counter_23__N_483[1]), .CK(dac_clk_p_c), 
            .Q(baud_counter[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i1.GSR = "DISABLED";
    FD1P3IX lcl_data_i7 (.D(n29210), .SP(zero_baud_counter), .CD(n26540), 
            .CK(dac_clk_p_c), .Q(\lcl_data[7] )) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(139[9] 143[40])
    defparam lcl_data_i7.GSR = "DISABLED";
    CCU2D sub_36_add_2_17 (.A0(baud_counter[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17406), .COUT(n17407), .S0(n108[15]), 
          .S1(n108[16]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_17.INIT0 = 16'h5555;
    defparam sub_36_add_2_17.INIT1 = 16'h5555;
    defparam sub_36_add_2_17.INJECT1_0 = "NO";
    defparam sub_36_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_36_add_2_15 (.A0(baud_counter[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17405), .COUT(n17406), .S0(n108[13]), 
          .S1(n108[14]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_15.INIT0 = 16'h5555;
    defparam sub_36_add_2_15.INIT1 = 16'h5555;
    defparam sub_36_add_2_15.INJECT1_0 = "NO";
    defparam sub_36_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_36_add_2_13 (.A0(baud_counter[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17404), .COUT(n17405), .S0(n108[11]), 
          .S1(n108[12]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_13.INIT0 = 16'h5555;
    defparam sub_36_add_2_13.INIT1 = 16'h5555;
    defparam sub_36_add_2_13.INJECT1_0 = "NO";
    defparam sub_36_add_2_13.INJECT1_1 = "NO";
    FD1P3AY lcl_data_i6 (.D(\lcl_data_7__N_511[6] ), .SP(dac_clk_p_c_enable_321), 
            .CK(dac_clk_p_c), .Q(\lcl_data[6] )) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(139[9] 143[40])
    defparam lcl_data_i6.GSR = "DISABLED";
    FD1P3AY lcl_data_i5 (.D(\lcl_data_7__N_511[5] ), .SP(dac_clk_p_c_enable_321), 
            .CK(dac_clk_p_c), .Q(\lcl_data[5] )) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(139[9] 143[40])
    defparam lcl_data_i5.GSR = "DISABLED";
    FD1P3AY lcl_data_i4 (.D(\lcl_data_7__N_511[4] ), .SP(dac_clk_p_c_enable_321), 
            .CK(dac_clk_p_c), .Q(\lcl_data[4] )) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(139[9] 143[40])
    defparam lcl_data_i4.GSR = "DISABLED";
    FD1P3AY lcl_data_i3 (.D(\lcl_data_7__N_511[3] ), .SP(dac_clk_p_c_enable_321), 
            .CK(dac_clk_p_c), .Q(\lcl_data[3] )) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(139[9] 143[40])
    defparam lcl_data_i3.GSR = "DISABLED";
    FD1P3AY lcl_data_i2 (.D(\lcl_data_7__N_511[2] ), .SP(dac_clk_p_c_enable_321), 
            .CK(dac_clk_p_c), .Q(\lcl_data[2] )) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(139[9] 143[40])
    defparam lcl_data_i2.GSR = "DISABLED";
    FD1P3AY lcl_data_i1 (.D(\lcl_data_7__N_511[1] ), .SP(dac_clk_p_c_enable_321), 
            .CK(dac_clk_p_c), .Q(\lcl_data[1] )) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(139[9] 143[40])
    defparam lcl_data_i1.GSR = "DISABLED";
    CCU2D sub_36_add_2_11 (.A0(baud_counter[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17403), .COUT(n17404), .S0(n108[9]), .S1(n108[10]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_11.INIT0 = 16'h5555;
    defparam sub_36_add_2_11.INIT1 = 16'h5555;
    defparam sub_36_add_2_11.INJECT1_0 = "NO";
    defparam sub_36_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_36_add_2_9 (.A0(baud_counter[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17402), .COUT(n17403), .S0(n108[7]), .S1(n108[8]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_9.INIT0 = 16'h5555;
    defparam sub_36_add_2_9.INIT1 = 16'h5555;
    defparam sub_36_add_2_9.INJECT1_0 = "NO";
    defparam sub_36_add_2_9.INJECT1_1 = "NO";
    LUT4 baud_counter_23__I_10_i14_4_lut (.A(n26540), .B(n133[13]), .C(n26427), 
         .D(zero_baud_counter_N_528), .Z(baud_counter_23__N_483[13])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((C+(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(217[12] 224[43])
    defparam baud_counter_23__I_10_i14_4_lut.init = 16'ha0ac;
    LUT4 i11557_2_lut (.A(n108[13]), .B(zero_baud_counter), .Z(n133[13])) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(224[4:43])
    defparam i11557_2_lut.init = 16'heeee;
    CCU2D sub_36_add_2_7 (.A0(baud_counter[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17401), .COUT(n17402), .S0(n108[5]), .S1(n108[6]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_7.INIT0 = 16'h5555;
    defparam sub_36_add_2_7.INIT1 = 16'h5555;
    defparam sub_36_add_2_7.INJECT1_0 = "NO";
    defparam sub_36_add_2_7.INJECT1_1 = "NO";
    LUT4 baud_counter_23__I_10_i11_4_lut (.A(n26540), .B(n133[10]), .C(n26427), 
         .D(zero_baud_counter_N_528), .Z(baud_counter_23__N_483[10])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((C+(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(217[12] 224[43])
    defparam baud_counter_23__I_10_i11_4_lut.init = 16'ha0ac;
    LUT4 i11558_2_lut (.A(n108[10]), .B(zero_baud_counter), .Z(n133[10])) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(224[4:43])
    defparam i11558_2_lut.init = 16'heeee;
    LUT4 baud_counter_23__I_10_i10_4_lut (.A(n26540), .B(n133[9]), .C(n26427), 
         .D(zero_baud_counter_N_528), .Z(baud_counter_23__N_483[9])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((C+(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(217[12] 224[43])
    defparam baud_counter_23__I_10_i10_4_lut.init = 16'ha0ac;
    LUT4 i11559_2_lut (.A(n108[9]), .B(zero_baud_counter), .Z(n133[9])) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(224[4:43])
    defparam i11559_2_lut.init = 16'heeee;
    LUT4 baud_counter_23__I_10_i9_4_lut (.A(n26540), .B(n133[8]), .C(n26427), 
         .D(zero_baud_counter_N_528), .Z(baud_counter_23__N_483[8])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((C+(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(217[12] 224[43])
    defparam baud_counter_23__I_10_i9_4_lut.init = 16'ha0ac;
    LUT4 i11560_2_lut (.A(n108[8]), .B(zero_baud_counter), .Z(n133[8])) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(224[4:43])
    defparam i11560_2_lut.init = 16'heeee;
    LUT4 baud_counter_23__I_10_i4_4_lut (.A(n26540), .B(n133[3]), .C(n26427), 
         .D(zero_baud_counter_N_528), .Z(baud_counter_23__N_483[3])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((C+(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(217[12] 224[43])
    defparam baud_counter_23__I_10_i4_4_lut.init = 16'ha0ac;
    LUT4 i11561_2_lut (.A(n108[3]), .B(zero_baud_counter), .Z(n133[3])) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(224[4:43])
    defparam i11561_2_lut.init = 16'heeee;
    LUT4 baud_counter_23__I_10_i3_4_lut (.A(n26540), .B(n133[2]), .C(n26427), 
         .D(zero_baud_counter_N_528), .Z(baud_counter_23__N_483[2])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((C+(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(217[12] 224[43])
    defparam baud_counter_23__I_10_i3_4_lut.init = 16'ha0ac;
    LUT4 i11562_2_lut (.A(n108[2]), .B(zero_baud_counter), .Z(n133[2])) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(224[4:43])
    defparam i11562_2_lut.init = 16'heeee;
    LUT4 baud_counter_23__I_10_i2_4_lut (.A(n26540), .B(n133[1]), .C(n26427), 
         .D(zero_baud_counter_N_528), .Z(baud_counter_23__N_483[1])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((C+(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(217[12] 224[43])
    defparam baud_counter_23__I_10_i2_4_lut.init = 16'ha0ac;
    LUT4 i11563_2_lut (.A(n108[1]), .B(zero_baud_counter), .Z(n133[1])) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(224[4:43])
    defparam i11563_2_lut.init = 16'heeee;
    CCU2D sub_36_add_2_5 (.A0(baud_counter[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17400), .COUT(n17401), .S0(n108[3]), .S1(n108[4]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_5.INIT0 = 16'h5555;
    defparam sub_36_add_2_5.INIT1 = 16'h5555;
    defparam sub_36_add_2_5.INJECT1_0 = "NO";
    defparam sub_36_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_36_add_2_3 (.A0(baud_counter[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17399), .COUT(n17400), .S0(n108[1]), .S1(n108[2]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_3.INIT0 = 16'h5555;
    defparam sub_36_add_2_3.INIT1 = 16'h5555;
    defparam sub_36_add_2_3.INJECT1_0 = "NO";
    defparam sub_36_add_2_3.INJECT1_1 = "NO";
    LUT4 i22381_2_lut (.A(o_busy_N_536), .B(zero_baud_counter), .Z(n8876)) /* synthesis lut_function=(!(A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(97[8] 113[6])
    defparam i22381_2_lut.init = 16'h7777;
    LUT4 i732_4_lut (.A(state_c[2]), .B(state_c[3]), .C(state_c[1]), .D(state[0]), 
         .Z(o_busy_N_536)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;
    defparam i732_4_lut.init = 16'hccc8;
    LUT4 state_544_mux_6_i2_4_lut (.A(state_c[1]), .B(n26540), .C(o_busy_N_536), 
         .D(state[0]), .Z(n27[1])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(110[14:26])
    defparam state_544_mux_6_i2_4_lut.init = 16'h353a;
    CCU2D sub_36_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(baud_counter[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n17399), .S1(n108[0]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_1.INIT0 = 16'hF000;
    defparam sub_36_add_2_1.INIT1 = 16'h5555;
    defparam sub_36_add_2_1.INJECT1_0 = "NO";
    defparam sub_36_add_2_1.INJECT1_1 = "NO";
    LUT4 zero_baud_counter_I_0_51_4_lut (.A(n26540), .B(n20118), .C(n26427), 
         .D(zero_baud_counter_N_528), .Z(zero_baud_counter_N_525)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C))+!A !((C+(D))+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(217[12] 224[43])
    defparam zero_baud_counter_I_0_51_4_lut.init = 16'h5f53;
    LUT4 i1_4_lut (.A(n20526), .B(n20534), .C(n20532), .D(n20524), .Z(n20118)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(207[24:43])
    defparam i1_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_105 (.A(baud_counter[1]), .B(baud_counter[4]), .C(baud_counter[17]), 
         .D(baud_counter[5]), .Z(n20526)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(207[24:43])
    defparam i1_4_lut_adj_105.init = 16'hfffe;
    LUT4 i1_4_lut_adj_106 (.A(n20510), .B(baud_counter[0]), .C(n20520), 
         .D(baud_counter[19]), .Z(n20534)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(207[24:43])
    defparam i1_4_lut_adj_106.init = 16'hfffb;
    LUT4 i1_4_lut_adj_107 (.A(baud_counter[22]), .B(n20522), .C(n20512), 
         .D(baud_counter[12]), .Z(n20532)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(207[24:43])
    defparam i1_4_lut_adj_107.init = 16'hfffe;
    LUT4 i1_2_lut_rep_574 (.A(state[0]), .B(state_c[3]), .Z(n26534)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(110[14:26])
    defparam i1_2_lut_rep_574.init = 16'h8888;
    LUT4 i1_3_lut_rep_467_4_lut (.A(state[0]), .B(state_c[3]), .C(state_c[1]), 
         .D(state_c[2]), .Z(n26427)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(110[14:26])
    defparam i1_3_lut_rep_467_4_lut.init = 16'h8000;
    LUT4 i1_4_lut_adj_108 (.A(baud_counter[18]), .B(baud_counter[11]), .C(baud_counter[9]), 
         .D(baud_counter[20]), .Z(n20524)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(207[24:43])
    defparam i1_4_lut_adj_108.init = 16'hfffe;
    LUT4 i1_2_lut (.A(baud_counter[8]), .B(baud_counter[6]), .Z(n20510)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(207[24:43])
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i1_4_lut_adj_109 (.A(baud_counter[13]), .B(baud_counter[23]), .C(baud_counter[3]), 
         .D(baud_counter[16]), .Z(n20520)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(207[24:43])
    defparam i1_4_lut_adj_109.init = 16'hfffe;
    LUT4 i1_4_lut_adj_110 (.A(baud_counter[7]), .B(baud_counter[2]), .C(baud_counter[15]), 
         .D(baud_counter[14]), .Z(n20522)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(207[24:43])
    defparam i1_4_lut_adj_110.init = 16'hfffe;
    LUT4 i11020_2_lut (.A(n108[0]), .B(zero_baud_counter), .Z(n133[0])) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(224[4:43])
    defparam i11020_2_lut.init = 16'heeee;
    FD1S3JX r_busy_45 (.D(n8876), .CK(dac_clk_p_c), .PD(n26540), .Q(tx_busy)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(92[9] 114[5])
    defparam r_busy_45.GSR = "DISABLED";
    LUT4 i1_2_lut_adj_111 (.A(baud_counter[21]), .B(baud_counter[10]), .Z(n20512)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(207[24:43])
    defparam i1_2_lut_adj_111.init = 16'heeee;
    PFUMX i24491 (.BLUT(n26781), .ALUT(n26782), .C0(state_c[3]), .Z(n26783));
    FD1P3AX state_544__i3 (.D(n26783), .SP(zero_baud_counter), .CK(dac_clk_p_c), 
            .Q(state_c[3]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(110[14:26])
    defparam state_544__i3.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_112 (.A(state_c[1]), .B(n26534), .C(state_c[2]), 
         .D(zero_baud_counter), .Z(zero_baud_counter_N_528)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_adj_112.init = 16'h0400;
    PFUMX i24489 (.BLUT(n26778), .ALUT(n26779), .C0(state_c[2]), .Z(n26780));
    FD1P3AX state_544__i2 (.D(n26780), .SP(zero_baud_counter), .CK(dac_clk_p_c), 
            .Q(state_c[2]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(110[14:26])
    defparam state_544__i2.GSR = "DISABLED";
    FD1P3AX state_544__i1 (.D(n27[1]), .SP(zero_baud_counter), .CK(dac_clk_p_c), 
            .Q(state_c[1]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(110[14:26])
    defparam state_544__i1.GSR = "DISABLED";
    FD1P3AX state_544__i0 (.D(n17598), .SP(zero_baud_counter), .CK(dac_clk_p_c), 
            .Q(state[0]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(110[14:26])
    defparam state_544__i0.GSR = "DISABLED";
    LUT4 baud_counter_23__I_10_i1_4_lut (.A(n26540), .B(n133[0]), .C(n26427), 
         .D(zero_baud_counter_N_528), .Z(baud_counter_23__N_483[0])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((C+(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(217[12] 224[43])
    defparam baud_counter_23__I_10_i1_4_lut.init = 16'ha0ac;
    
endmodule
//
// Verilog Description of module efb_inst
//

module efb_inst (dac_clk_p_c, n26683, wb_cyc, wb_lo_data_7__N_96, wb_we, 
            \wb_addr[7] , \wb_addr[6] , \wb_addr[5] , \wb_addr[4] , 
            \wb_addr[3] , \wb_addr[2] , \wb_addr[1] , \wb_addr[0] , 
            \wb_odata[7] , \wb_odata[6] , \wb_odata[5] , \wb_odata[4] , 
            \wb_odata[3] , \wb_odata[2] , \wb_odata[1] , \wb_odata[0] , 
            pll_data_o, pll_ack, wb_lo_data, wb_lo_ack, pll_clk, pll_rst, 
            pll_stb, pll_we, pll_addr, pll_data_i, GND_net, VCC_net) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;
    input dac_clk_p_c;
    input n26683;
    input wb_cyc;
    input wb_lo_data_7__N_96;
    input wb_we;
    input \wb_addr[7] ;
    input \wb_addr[6] ;
    input \wb_addr[5] ;
    input \wb_addr[4] ;
    input \wb_addr[3] ;
    input \wb_addr[2] ;
    input \wb_addr[1] ;
    input \wb_addr[0] ;
    input \wb_odata[7] ;
    input \wb_odata[6] ;
    input \wb_odata[5] ;
    input \wb_odata[4] ;
    input \wb_odata[3] ;
    input \wb_odata[2] ;
    input \wb_odata[1] ;
    input \wb_odata[0] ;
    input [7:0]pll_data_o;
    input pll_ack;
    output [7:0]wb_lo_data;
    output wb_lo_ack;
    output pll_clk;
    output pll_rst;
    output pll_stb;
    output pll_we;
    output [4:0]pll_addr;
    output [7:0]pll_data_i;
    input GND_net;
    input VCC_net;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(29[49:58])
    
    EFB EFBInst_0 (.WBCLKI(dac_clk_p_c), .WBRSTI(n26683), .WBCYCI(wb_cyc), 
        .WBSTBI(wb_lo_data_7__N_96), .WBWEI(wb_we), .WBADRI0(\wb_addr[0] ), 
        .WBADRI1(\wb_addr[1] ), .WBADRI2(\wb_addr[2] ), .WBADRI3(\wb_addr[3] ), 
        .WBADRI4(\wb_addr[4] ), .WBADRI5(\wb_addr[5] ), .WBADRI6(\wb_addr[6] ), 
        .WBADRI7(\wb_addr[7] ), .WBDATI0(\wb_odata[0] ), .WBDATI1(\wb_odata[1] ), 
        .WBDATI2(\wb_odata[2] ), .WBDATI3(\wb_odata[3] ), .WBDATI4(\wb_odata[4] ), 
        .WBDATI5(\wb_odata[5] ), .WBDATI6(\wb_odata[6] ), .WBDATI7(\wb_odata[7] ), 
        .I2C1SCLI(GND_net), .I2C1SDAI(GND_net), .I2C2SCLI(GND_net), .I2C2SDAI(GND_net), 
        .SPISCKI(GND_net), .SPIMISOI(GND_net), .SPIMOSII(GND_net), .SPISCSN(GND_net), 
        .TCCLKI(GND_net), .TCRSTN(GND_net), .TCIC(GND_net), .UFMSN(VCC_net), 
        .PLL0DATI0(pll_data_o[0]), .PLL0DATI1(pll_data_o[1]), .PLL0DATI2(pll_data_o[2]), 
        .PLL0DATI3(pll_data_o[3]), .PLL0DATI4(pll_data_o[4]), .PLL0DATI5(pll_data_o[5]), 
        .PLL0DATI6(pll_data_o[6]), .PLL0DATI7(pll_data_o[7]), .PLL0ACKI(pll_ack), 
        .PLL1DATI0(GND_net), .PLL1DATI1(GND_net), .PLL1DATI2(GND_net), 
        .PLL1DATI3(GND_net), .PLL1DATI4(GND_net), .PLL1DATI5(GND_net), 
        .PLL1DATI6(GND_net), .PLL1DATI7(GND_net), .PLL1ACKI(GND_net), 
        .WBDATO0(wb_lo_data[0]), .WBDATO1(wb_lo_data[1]), .WBDATO2(wb_lo_data[2]), 
        .WBDATO3(wb_lo_data[3]), .WBDATO4(wb_lo_data[4]), .WBDATO5(wb_lo_data[5]), 
        .WBDATO6(wb_lo_data[6]), .WBDATO7(wb_lo_data[7]), .WBACKO(wb_lo_ack), 
        .PLLCLKO(pll_clk), .PLLRSTO(pll_rst), .PLL0STBO(pll_stb), .PLLWEO(pll_we), 
        .PLLADRO0(pll_addr[0]), .PLLADRO1(pll_addr[1]), .PLLADRO2(pll_addr[2]), 
        .PLLADRO3(pll_addr[3]), .PLLADRO4(pll_addr[4]), .PLLDATO0(pll_data_i[0]), 
        .PLLDATO1(pll_data_i[1]), .PLLDATO2(pll_data_i[2]), .PLLDATO3(pll_data_i[3]), 
        .PLLDATO4(pll_data_i[4]), .PLLDATO5(pll_data_i[5]), .PLLDATO6(pll_data_i[6]), 
        .PLLDATO7(pll_data_i[7])) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=8, LSE_LCOL=10, LSE_RCOL=3, LSE_LLINE=177, LSE_RLINE=189 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(177[10] 189[3])
    defparam EFBInst_0.EFB_I2C1 = "DISABLED";
    defparam EFBInst_0.EFB_I2C2 = "DISABLED";
    defparam EFBInst_0.EFB_SPI = "DISABLED";
    defparam EFBInst_0.EFB_TC = "DISABLED";
    defparam EFBInst_0.EFB_TC_PORTMODE = "WB";
    defparam EFBInst_0.EFB_UFM = "DISABLED";
    defparam EFBInst_0.EFB_WB_CLK_FREQ = "50.0";
    defparam EFBInst_0.DEV_DENSITY = "6900L";
    defparam EFBInst_0.UFM_INIT_PAGES = 0;
    defparam EFBInst_0.UFM_INIT_START_PAGE = 0;
    defparam EFBInst_0.UFM_INIT_ALL_ZEROS = "ENABLED";
    defparam EFBInst_0.UFM_INIT_FILE_NAME = "NONE";
    defparam EFBInst_0.UFM_INIT_FILE_FORMAT = "HEX";
    defparam EFBInst_0.I2C1_ADDRESSING = "7BIT";
    defparam EFBInst_0.I2C2_ADDRESSING = "7BIT";
    defparam EFBInst_0.I2C1_SLAVE_ADDR = "0b1000001";
    defparam EFBInst_0.I2C2_SLAVE_ADDR = "0b1000010";
    defparam EFBInst_0.I2C1_BUS_PERF = "100kHz";
    defparam EFBInst_0.I2C2_BUS_PERF = "100kHz";
    defparam EFBInst_0.I2C1_CLK_DIVIDER = 1;
    defparam EFBInst_0.I2C2_CLK_DIVIDER = 1;
    defparam EFBInst_0.I2C1_GEN_CALL = "DISABLED";
    defparam EFBInst_0.I2C2_GEN_CALL = "DISABLED";
    defparam EFBInst_0.I2C1_WAKEUP = "DISABLED";
    defparam EFBInst_0.I2C2_WAKEUP = "DISABLED";
    defparam EFBInst_0.SPI_MODE = "MASTER";
    defparam EFBInst_0.SPI_CLK_DIVIDER = 1;
    defparam EFBInst_0.SPI_LSB_FIRST = "DISABLED";
    defparam EFBInst_0.SPI_CLK_INV = "DISABLED";
    defparam EFBInst_0.SPI_PHASE_ADJ = "DISABLED";
    defparam EFBInst_0.SPI_SLAVE_HANDSHAKE = "DISABLED";
    defparam EFBInst_0.SPI_INTR_TXRDY = "DISABLED";
    defparam EFBInst_0.SPI_INTR_RXRDY = "DISABLED";
    defparam EFBInst_0.SPI_INTR_TXOVR = "DISABLED";
    defparam EFBInst_0.SPI_INTR_RXOVR = "DISABLED";
    defparam EFBInst_0.SPI_WAKEUP = "DISABLED";
    defparam EFBInst_0.TC_MODE = "CTCM";
    defparam EFBInst_0.TC_SCLK_SEL = "PCLOCK";
    defparam EFBInst_0.TC_CCLK_SEL = 1;
    defparam EFBInst_0.GSR = "ENABLED";
    defparam EFBInst_0.TC_TOP_SET = 65535;
    defparam EFBInst_0.TC_OCR_SET = 32767;
    defparam EFBInst_0.TC_OC_MODE = "TOGGLE";
    defparam EFBInst_0.TC_RESETN = "ENABLED";
    defparam EFBInst_0.TC_TOP_SEL = "OFF";
    defparam EFBInst_0.TC_OV_INT = "OFF";
    defparam EFBInst_0.TC_OCR_INT = "OFF";
    defparam EFBInst_0.TC_ICR_INT = "OFF";
    defparam EFBInst_0.TC_OVERFLOW = "DISABLED";
    defparam EFBInst_0.TC_ICAPTURE = "DISABLED";
    
endmodule
//
// Verilog Description of module TSALL
// module not written out since it is a black-box. 
//

//
// Verilog Description of module clock_phase_shifter
//

module clock_phase_shifter (q_clk_p_c, i_clk_2f_N_2250, q_clk_n_c, i_clk_p_c, 
            lo_pll_out, i_clk_n_c) /* synthesis syn_module_defined=1 */ ;
    output q_clk_p_c;
    input i_clk_2f_N_2250;
    input q_clk_n_c;
    output i_clk_p_c;
    input lo_pll_out;
    input i_clk_n_c;
    
    wire i_clk_2f_N_2250 /* synthesis is_inv_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/clock_phase_shifter.v(11[21:28])
    wire lo_pll_out /* synthesis is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(157[6:16])
    
    FD1S3AX o_clk_q_10 (.D(q_clk_n_c), .CK(i_clk_2f_N_2250), .Q(q_clk_p_c)) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=21, LSE_RCOL=2, LSE_LLINE=158, LSE_RLINE=162 */ ;   // d:/documents/git_local/fm_modulator/rtl/clock_phase_shifter.v(17[8] 19[4])
    defparam o_clk_q_10.GSR = "DISABLED";
    FD1S3AX o_clk_i_9 (.D(i_clk_n_c), .CK(lo_pll_out), .Q(i_clk_p_c)) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=21, LSE_RCOL=2, LSE_LLINE=158, LSE_RLINE=162 */ ;   // d:/documents/git_local/fm_modulator/rtl/clock_phase_shifter.v(13[8] 15[4])
    defparam o_clk_i_9.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module sys_clk
//

module sys_clk (i_ref_clk_c, dac_clk_p_c, GND_net) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;
    input i_ref_clk_c;
    output dac_clk_p_c;
    input GND_net;
    
    wire i_ref_clk_c /* synthesis is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(23[12:21])
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(29[49:58])
    
    EHXPLLJ PLLInst_0 (.CLKI(i_ref_clk_c), .CLKFB(dac_clk_p_c), .PHASESEL0(GND_net), 
            .PHASESEL1(GND_net), .PHASEDIR(GND_net), .PHASESTEP(GND_net), 
            .LOADREG(GND_net), .STDBY(GND_net), .PLLWAKESYNC(GND_net), 
            .RST(GND_net), .RESETC(GND_net), .RESETD(GND_net), .RESETM(GND_net), 
            .ENCLKOP(GND_net), .ENCLKOS(GND_net), .ENCLKOS2(GND_net), 
            .ENCLKOS3(GND_net), .PLLCLK(GND_net), .PLLRST(GND_net), .PLLSTB(GND_net), 
            .PLLWE(GND_net), .PLLDATI0(GND_net), .PLLDATI1(GND_net), .PLLDATI2(GND_net), 
            .PLLDATI3(GND_net), .PLLDATI4(GND_net), .PLLDATI5(GND_net), 
            .PLLDATI6(GND_net), .PLLDATI7(GND_net), .PLLADDR0(GND_net), 
            .PLLADDR1(GND_net), .PLLADDR2(GND_net), .PLLADDR3(GND_net), 
            .PLLADDR4(GND_net), .CLKOP(dac_clk_p_c)) /* synthesis FREQUENCY_PIN_CLKOP="72.000000", FREQUENCY_PIN_CLKI="12.000000", ICP_CURRENT="9", LPF_RESISTOR="72", syn_instantiated=1, LSE_LINE_FILE_ID=8, LSE_LCOL=10, LSE_RCOL=54, LSE_LLINE=38, LSE_RLINE=38 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(38[10:54])
    defparam PLLInst_0.CLKI_DIV = 1;
    defparam PLLInst_0.CLKFB_DIV = 6;
    defparam PLLInst_0.CLKOP_DIV = 7;
    defparam PLLInst_0.CLKOS_DIV = 1;
    defparam PLLInst_0.CLKOS2_DIV = 1;
    defparam PLLInst_0.CLKOS3_DIV = 1;
    defparam PLLInst_0.CLKOP_ENABLE = "ENABLED";
    defparam PLLInst_0.CLKOS_ENABLE = "DISABLED";
    defparam PLLInst_0.CLKOS2_ENABLE = "DISABLED";
    defparam PLLInst_0.CLKOS3_ENABLE = "DISABLED";
    defparam PLLInst_0.VCO_BYPASS_A0 = "DISABLED";
    defparam PLLInst_0.VCO_BYPASS_B0 = "DISABLED";
    defparam PLLInst_0.VCO_BYPASS_C0 = "DISABLED";
    defparam PLLInst_0.VCO_BYPASS_D0 = "DISABLED";
    defparam PLLInst_0.CLKOP_CPHASE = 6;
    defparam PLLInst_0.CLKOS_CPHASE = 0;
    defparam PLLInst_0.CLKOS2_CPHASE = 0;
    defparam PLLInst_0.CLKOS3_CPHASE = 0;
    defparam PLLInst_0.CLKOP_FPHASE = 0;
    defparam PLLInst_0.CLKOS_FPHASE = 0;
    defparam PLLInst_0.CLKOS2_FPHASE = 0;
    defparam PLLInst_0.CLKOS3_FPHASE = 0;
    defparam PLLInst_0.FEEDBK_PATH = "CLKOP";
    defparam PLLInst_0.FRACN_ENABLE = "DISABLED";
    defparam PLLInst_0.FRACN_DIV = 0;
    defparam PLLInst_0.CLKOP_TRIM_POL = "RISING";
    defparam PLLInst_0.CLKOP_TRIM_DELAY = 0;
    defparam PLLInst_0.CLKOS_TRIM_POL = "FALLING";
    defparam PLLInst_0.CLKOS_TRIM_DELAY = 0;
    defparam PLLInst_0.PLL_USE_WB = "DISABLED";
    defparam PLLInst_0.PREDIVIDER_MUXA1 = 0;
    defparam PLLInst_0.PREDIVIDER_MUXB1 = 0;
    defparam PLLInst_0.PREDIVIDER_MUXC1 = 0;
    defparam PLLInst_0.PREDIVIDER_MUXD1 = 0;
    defparam PLLInst_0.OUTDIVIDER_MUXA2 = "DIVA";
    defparam PLLInst_0.OUTDIVIDER_MUXB2 = "DIVB";
    defparam PLLInst_0.OUTDIVIDER_MUXC2 = "DIVC";
    defparam PLLInst_0.OUTDIVIDER_MUXD2 = "DIVD";
    defparam PLLInst_0.PLL_LOCK_MODE = 0;
    defparam PLLInst_0.STDBY_ENABLE = "DISABLED";
    defparam PLLInst_0.DPHASE_SOURCE = "DISABLED";
    defparam PLLInst_0.PLLRST_ENA = "DISABLED";
    defparam PLLInst_0.MRST_ENA = "DISABLED";
    defparam PLLInst_0.DCRST_ENA = "DISABLED";
    defparam PLLInst_0.DDRST_ENA = "DISABLED";
    defparam PLLInst_0.INTFB_WAKE = "DISABLED";
    
endmodule
//
// Verilog Description of module fm_generator_wb_slave
//

module fm_generator_wb_slave (dac_clk_p_c, wb_odata, n26683, wb_fm_data, 
            \wb_addr[1] , wb_fm_ack, o_dac_a_9__N_1, GND_net, \wb_addr[0] , 
            \power_counter[1] , \smpl_register[1] , n2035, n26563, n38, 
            n34, \wb_addr[8] , \wb_addr[12] , n26557, \wb_addr[15] , 
            \wb_addr[9] , o_dac_cw_b_c_c, n2, \smpl_register[16] , n26331, 
            n2_adj_1, \smpl_register[10] , n26342, n2_adj_2, \smpl_register[9] , 
            n26341, n2_adj_3, \smpl_register[29] , n26339, n2_adj_4, 
            \smpl_register[20] , n26337, n2_adj_5, \smpl_register[5] , 
            n26336, n2_adj_6, \smpl_register[18] , n26333, n2_adj_7, 
            \smpl_register[17] , n26332, o_dac_a_c_5, o_dac_b_c_15, 
            o_dac_b_c_9, n26643, o_dac_a_c_9, n20438, n20864, n20416, 
            n20402, n20422, o_dac_b_c_7, \o_sample_i[7] , \o_sample_i[14] , 
            \o_sample_i[13] , \o_sample_i[11] , \o_sample_i[10] , \o_sample_i[9] , 
            \o_sample_i[8] , n29209, o_dac_b_c_14, o_dac_b_c_13, o_dac_b_c_12, 
            o_dac_b_c_11, o_dac_b_c_10, n3537, o_dac_b_c_8) /* synthesis syn_module_defined=1 */ ;
    input dac_clk_p_c;
    input [31:0]wb_odata;
    input n26683;
    output [31:0]wb_fm_data;
    input \wb_addr[1] ;
    output wb_fm_ack;
    input o_dac_a_9__N_1;
    input GND_net;
    input \wb_addr[0] ;
    input \power_counter[1] ;
    input \smpl_register[1] ;
    output n2035;
    input n26563;
    input n38;
    input n34;
    input \wb_addr[8] ;
    input \wb_addr[12] ;
    input n26557;
    input \wb_addr[15] ;
    input \wb_addr[9] ;
    input o_dac_cw_b_c_c;
    input n2;
    input \smpl_register[16] ;
    output n26331;
    input n2_adj_1;
    input \smpl_register[10] ;
    output n26342;
    input n2_adj_2;
    input \smpl_register[9] ;
    output n26341;
    input n2_adj_3;
    input \smpl_register[29] ;
    output n26339;
    input n2_adj_4;
    input \smpl_register[20] ;
    output n26337;
    input n2_adj_5;
    input \smpl_register[5] ;
    output n26336;
    input n2_adj_6;
    input \smpl_register[18] ;
    output n26333;
    input n2_adj_7;
    input \smpl_register[17] ;
    output n26332;
    output o_dac_a_c_5;
    output o_dac_b_c_15;
    output o_dac_b_c_9;
    output n26643;
    output o_dac_a_c_9;
    input n20438;
    input n20864;
    input n20416;
    input n20402;
    input n20422;
    output o_dac_b_c_7;
    output \o_sample_i[7] ;
    output \o_sample_i[14] ;
    output \o_sample_i[13] ;
    output \o_sample_i[11] ;
    output \o_sample_i[10] ;
    output \o_sample_i[9] ;
    output \o_sample_i[8] ;
    input n29209;
    output o_dac_b_c_14;
    output o_dac_b_c_13;
    output o_dac_b_c_12;
    output o_dac_b_c_11;
    output o_dac_b_c_10;
    output n3537;
    output o_dac_b_c_8;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(29[49:58])
    wire [15:0]modulation_output /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(73[39:56])
    wire [15:0]o_sample_i /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[39:49])
    wire o_dac_b_c_15 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire o_dac_b_c_7 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire \o_sample_i[7]  /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[39:49])
    wire \o_sample_i[14]  /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[39:49])
    wire \o_sample_i[13]  /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[39:49])
    wire \o_sample_i[11]  /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[39:49])
    wire \o_sample_i[10]  /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[39:49])
    wire \o_sample_i[9]  /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[39:49])
    wire \o_sample_i[8]  /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[39:49])
    wire o_dac_b_c_14 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire o_dac_b_c_13 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire o_dac_b_c_12 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire o_dac_b_c_11 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire o_dac_b_c_10 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire n3537 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire o_dac_b_c_8 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire [31:0]\addr_space[3] ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(36[12:22])
    
    wire dac_clk_p_c_enable_143;
    wire [31:0]\addr_space[0] ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(36[12:22])
    
    wire dac_clk_p_c_enable_114;
    wire [31:0]\addr_space[1] ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(36[12:22])
    
    wire dac_clk_p_c_enable_71;
    wire [31:0]\addr_space[2] ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(36[12:22])
    
    wire dac_clk_p_c_enable_103;
    wire [30:0]carrier_center_increment_offset_ls;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(63[31:65])
    wire [30:0]n1;
    wire [31:0]o_wb_data_31__N_1337;
    wire [30:0]carrier_center_increment_offset_rs;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(63[67:101])
    wire [30:0]carrier_center_increment_offset_rs_30__N_1560;
    wire [30:0]carrier_increment;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(64[31:48])
    wire [30:0]carrier_increment_30__N_1591;
    wire [16:0]sine_lookup_width_minus_modulation_deviation_amount;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(85[27:78])
    wire [31:0]sine_lookup_width_minus_modulation_deviation_amount_16__N_1622;
    wire [16:0]modulation_deviation_amount_minus_sine_lookup_width;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(85[80:131])
    
    wire n21740, n21741, n63, n94, n22092, n64, n95, n17377, 
        n14347, n17376, n17375, n17374, n17373, n17372, n17371, 
        n17370, n17369, n17368, n17367, n21743, n21744, n17366, 
        n17365, n17364, n17363, n17361, n21746, n21747, n21749, 
        n21750, n21752, n21753, n17360, n17359, n21755, n21756, 
        n17428;
    wire [17:0]modulation_deviation_amount_minus_sine_lookup_width_16__N_1639;
    
    wire n17427, n17358, n17426, n17425, n26533, n26355, n58, 
        n89, n17424, n17423, n17357, n17356, n20073, n17355, n17354, 
        n21738, n21737, n26558, n72, n20634, n20636, n20638, n20624, 
        n178, n13449, n36_adj_2995, n13450, n40_adj_2996, n44_adj_2997, 
        n71, n9, n11, n13, n15, n13451, n7, n13448, n26409, 
        n13457, n37_adj_2998, n33_adj_2999, n41_adj_3000, n45_adj_3001, 
        n72_adj_3002, n14, n10, n12, n21735, n6, n8, n13456, 
        n38_adj_3003, n42_adj_3004, n46_adj_3005, n73, n21734, n20348, 
        n20362, n20360, n20346, n20350, n85, n26379, n26380, n21006, 
        n81, n26364, n80, n88, n26365, n21005, n21003, n21002, 
        n21000, n20999, n73_adj_3006, n104, n21926, n135, n78, 
        n101, n79, n102, n103, n134, n82, n59_adj_3007, n26553, 
        n105, n47_adj_3008, n74, n83, n60_adj_3009, n106, n48_adj_3010, 
        n75, n21858, n26399, n26366, n21857, n21855, n21854, n26400, 
        n43_adj_3011, n21852, n21851, n21849, n21848, n21846, n21845, 
        n26325, n26324, n26326, n21843, n26319, n26318, n26320, 
        n21842, n26313, n26312, n26314, n21840, n21839, n21837, 
        n21836, n21834, n26267, n39_adj_3012, n26268, n21833, n20488, 
        n20482, n20480, n21831, n21830, n8972, n8970, n21828, 
        n70, n178_adj_3015, n52_adj_3016, n25, n27, n56_adj_3017, 
        n29, n17, n19, n21, n23, n95_adj_3018, n26445, n49_adj_3019, 
        n53_adj_3020, n57_adj_3021, n30, n18, n20, n22, n24, n21827, 
        n26, n28, n96, n26556, n21825, n50_adj_3022, n54_adj_3023, 
        n97, n113, n16, n51_adj_3024, n55_adj_3025, n98, n114, 
        n21824, n99, n115, n76, n45_adj_3026, n84, n26555, n100, 
        n26363, n77, n46_adj_3027, n21822, n132, n133, n136, n21821, 
        n137, n107, n123, n21813, n108, n21812, n26398, n21804, 
        n24273, n24274, n21803, n21795, n21794, n21786, n21785, 
        n21777, n21776, n21771, n21770, n21762, n21761, n21759, 
        n21758, n26425, n24275, n26266, n26269, n26615, n117, 
        n118, n20296, n20112, n20302, n20298;
    wire [15:0]quarter_wave_sample_register_q;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(22[56:86])
    
    FD1P3AX \addr_space_3[[30__265  (.D(wb_odata[30]), .SP(dac_clk_p_c_enable_143), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[30__265 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[29__267  (.D(wb_odata[29]), .SP(dac_clk_p_c_enable_143), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[29__267 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[28__269  (.D(wb_odata[28]), .SP(dac_clk_p_c_enable_143), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[28__269 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[27__271  (.D(wb_odata[27]), .SP(dac_clk_p_c_enable_143), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[27__271 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[26__273  (.D(wb_odata[26]), .SP(dac_clk_p_c_enable_143), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[26__273 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[30__166  (.D(wb_odata[30]), .SP(dac_clk_p_c_enable_114), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[0] [30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[30__166 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[29__167  (.D(wb_odata[29]), .SP(dac_clk_p_c_enable_114), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[0] [29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[29__167 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[28__168  (.D(wb_odata[28]), .SP(dac_clk_p_c_enable_114), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[0] [28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[28__168 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[27__169  (.D(wb_odata[27]), .SP(dac_clk_p_c_enable_114), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[0] [27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[27__169 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[26__170  (.D(wb_odata[26]), .SP(dac_clk_p_c_enable_114), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[0] [26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[26__170 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[25__171  (.D(wb_odata[25]), .SP(dac_clk_p_c_enable_114), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[0] [25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[25__171 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[24__172  (.D(wb_odata[24]), .SP(dac_clk_p_c_enable_114), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[0] [24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[24__172 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[23__173  (.D(wb_odata[23]), .SP(dac_clk_p_c_enable_114), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[0] [23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[23__173 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[21__176  (.D(wb_odata[21]), .SP(dac_clk_p_c_enable_114), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[0] [21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[21__176 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[20__177  (.D(wb_odata[20]), .SP(dac_clk_p_c_enable_114), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[0] [20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[20__177 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[19__178  (.D(wb_odata[19]), .SP(dac_clk_p_c_enable_114), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[0] [19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[19__178 .GSR = "DISABLED";
    FD1P3BX \addr_space_0[[18__179  (.D(wb_odata[18]), .SP(dac_clk_p_c_enable_114), 
            .CK(dac_clk_p_c), .PD(n26683), .Q(\addr_space[0] [18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[18__179 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[17__180  (.D(wb_odata[17]), .SP(dac_clk_p_c_enable_114), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[0] [17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[17__180 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[16__181  (.D(wb_odata[16]), .SP(dac_clk_p_c_enable_114), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[0] [16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[16__181 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[15__182  (.D(wb_odata[15]), .SP(dac_clk_p_c_enable_114), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[0] [15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[15__182 .GSR = "DISABLED";
    FD1P3BX \addr_space_0[[14__183  (.D(wb_odata[14]), .SP(dac_clk_p_c_enable_114), 
            .CK(dac_clk_p_c), .PD(n26683), .Q(\addr_space[0] [14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[14__183 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[13__184  (.D(wb_odata[13]), .SP(dac_clk_p_c_enable_114), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[0] [13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[13__184 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[12__185  (.D(wb_odata[12]), .SP(dac_clk_p_c_enable_114), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[0] [12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[12__185 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[11__186  (.D(wb_odata[11]), .SP(dac_clk_p_c_enable_114), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[0] [11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[11__186 .GSR = "DISABLED";
    FD1P3BX \addr_space_0[[10__187  (.D(wb_odata[10]), .SP(dac_clk_p_c_enable_114), 
            .CK(dac_clk_p_c), .PD(n26683), .Q(\addr_space[0] [10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[10__187 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[9__188  (.D(wb_odata[9]), .SP(dac_clk_p_c_enable_114), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[0] [9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[9__188 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[8__189  (.D(wb_odata[8]), .SP(dac_clk_p_c_enable_114), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[0] [8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[8__189 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[7__190  (.D(wb_odata[7]), .SP(dac_clk_p_c_enable_114), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[0] [7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[7__190 .GSR = "DISABLED";
    FD1P3BX \addr_space_0[[6__191  (.D(wb_odata[6]), .SP(dac_clk_p_c_enable_114), 
            .CK(dac_clk_p_c), .PD(n26683), .Q(\addr_space[0] [6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[6__191 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[5__192  (.D(wb_odata[5]), .SP(dac_clk_p_c_enable_114), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[0] [5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[5__192 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[4__193  (.D(wb_odata[4]), .SP(dac_clk_p_c_enable_114), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[0] [4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[4__193 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[3__194  (.D(wb_odata[3]), .SP(dac_clk_p_c_enable_114), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[0] [3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[3__194 .GSR = "DISABLED";
    FD1P3BX \addr_space_0[[2__195  (.D(wb_odata[2]), .SP(dac_clk_p_c_enable_114), 
            .CK(dac_clk_p_c), .PD(n26683), .Q(\addr_space[0] [2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[2__195 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[1__196  (.D(wb_odata[1]), .SP(dac_clk_p_c_enable_114), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[0] [1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[1__196 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[0__197  (.D(wb_odata[0]), .SP(dac_clk_p_c_enable_114), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[0] [0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[0__197 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[31__198  (.D(wb_odata[31]), .SP(dac_clk_p_c_enable_71), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[1] [31])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[31__198 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[30__199  (.D(wb_odata[30]), .SP(dac_clk_p_c_enable_71), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[1] [30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[30__199 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[29__200  (.D(wb_odata[29]), .SP(dac_clk_p_c_enable_71), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[1] [29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[29__200 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[28__201  (.D(wb_odata[28]), .SP(dac_clk_p_c_enable_71), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[1] [28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[28__201 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[27__202  (.D(wb_odata[27]), .SP(dac_clk_p_c_enable_71), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[1] [27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[27__202 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[26__203  (.D(wb_odata[26]), .SP(dac_clk_p_c_enable_71), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[1] [26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[26__203 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[25__204  (.D(wb_odata[25]), .SP(dac_clk_p_c_enable_71), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[1] [25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[25__204 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[24__205  (.D(wb_odata[24]), .SP(dac_clk_p_c_enable_71), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[1] [24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[24__205 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[23__206  (.D(wb_odata[23]), .SP(dac_clk_p_c_enable_71), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[1] [23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[23__206 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[22__207  (.D(wb_odata[22]), .SP(dac_clk_p_c_enable_71), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[1] [22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[22__207 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[21__208  (.D(wb_odata[21]), .SP(dac_clk_p_c_enable_71), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[1] [21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[21__208 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[20__209  (.D(wb_odata[20]), .SP(dac_clk_p_c_enable_71), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[1] [20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[20__209 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[19__210  (.D(wb_odata[19]), .SP(dac_clk_p_c_enable_71), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[1] [19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[19__210 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[18__211  (.D(wb_odata[18]), .SP(dac_clk_p_c_enable_71), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[1] [18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[18__211 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[17__212  (.D(wb_odata[17]), .SP(dac_clk_p_c_enable_71), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[1] [17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[17__212 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[16__213  (.D(wb_odata[16]), .SP(dac_clk_p_c_enable_71), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[1] [16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[16__213 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[15__214  (.D(wb_odata[15]), .SP(dac_clk_p_c_enable_71), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[1] [15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[15__214 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[14__215  (.D(wb_odata[14]), .SP(dac_clk_p_c_enable_71), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[1] [14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[14__215 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[13__216  (.D(wb_odata[13]), .SP(dac_clk_p_c_enable_71), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[1] [13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[13__216 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[12__217  (.D(wb_odata[12]), .SP(dac_clk_p_c_enable_71), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[1] [12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[12__217 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[11__218  (.D(wb_odata[11]), .SP(dac_clk_p_c_enable_71), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[1] [11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[11__218 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[10__219  (.D(wb_odata[10]), .SP(dac_clk_p_c_enable_71), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[1] [10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[10__219 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[9__220  (.D(wb_odata[9]), .SP(dac_clk_p_c_enable_71), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[1] [9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[9__220 .GSR = "DISABLED";
    FD1P3BX \addr_space_1[[8__221  (.D(wb_odata[8]), .SP(dac_clk_p_c_enable_71), 
            .CK(dac_clk_p_c), .PD(n26683), .Q(\addr_space[1] [8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[8__221 .GSR = "DISABLED";
    FD1P3BX \addr_space_1[[7__222  (.D(wb_odata[7]), .SP(dac_clk_p_c_enable_71), 
            .CK(dac_clk_p_c), .PD(n26683), .Q(\addr_space[1] [7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[7__222 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[6__223  (.D(wb_odata[6]), .SP(dac_clk_p_c_enable_71), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[1] [6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[6__223 .GSR = "DISABLED";
    FD1P3BX \addr_space_1[[5__224  (.D(wb_odata[5]), .SP(dac_clk_p_c_enable_71), 
            .CK(dac_clk_p_c), .PD(n26683), .Q(\addr_space[1] [5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[5__224 .GSR = "DISABLED";
    FD1P3BX \addr_space_1[[4__225  (.D(wb_odata[4]), .SP(dac_clk_p_c_enable_71), 
            .CK(dac_clk_p_c), .PD(n26683), .Q(\addr_space[1] [4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[4__225 .GSR = "DISABLED";
    FD1P3BX \addr_space_1[[3__226  (.D(wb_odata[3]), .SP(dac_clk_p_c_enable_71), 
            .CK(dac_clk_p_c), .PD(n26683), .Q(\addr_space[1] [3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[3__226 .GSR = "DISABLED";
    FD1P3BX \addr_space_1[[2__227  (.D(wb_odata[2]), .SP(dac_clk_p_c_enable_71), 
            .CK(dac_clk_p_c), .PD(n26683), .Q(\addr_space[1] [2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[2__227 .GSR = "DISABLED";
    FD1P3BX \addr_space_1[[1__228  (.D(wb_odata[1]), .SP(dac_clk_p_c_enable_71), 
            .CK(dac_clk_p_c), .PD(n26683), .Q(\addr_space[1] [1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[1__228 .GSR = "DISABLED";
    FD1P3BX \addr_space_1[[0__229  (.D(wb_odata[0]), .SP(dac_clk_p_c_enable_71), 
            .CK(dac_clk_p_c), .PD(n26683), .Q(\addr_space[1] [0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_1[[0__229 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[31__230  (.D(wb_odata[31]), .SP(dac_clk_p_c_enable_103), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[2] [31])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[31__230 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[30__231  (.D(wb_odata[30]), .SP(dac_clk_p_c_enable_103), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[2] [30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[30__231 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[29__232  (.D(wb_odata[29]), .SP(dac_clk_p_c_enable_103), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[2] [29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[29__232 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[28__233  (.D(wb_odata[28]), .SP(dac_clk_p_c_enable_103), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[2] [28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[28__233 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[27__234  (.D(wb_odata[27]), .SP(dac_clk_p_c_enable_103), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[2] [27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[27__234 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[26__235  (.D(wb_odata[26]), .SP(dac_clk_p_c_enable_103), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[2] [26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[26__235 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[25__236  (.D(wb_odata[25]), .SP(dac_clk_p_c_enable_103), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[2] [25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[25__236 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[24__237  (.D(wb_odata[24]), .SP(dac_clk_p_c_enable_103), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[2] [24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[24__237 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[23__238  (.D(wb_odata[23]), .SP(dac_clk_p_c_enable_103), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[2] [23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[23__238 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[22__239  (.D(wb_odata[22]), .SP(dac_clk_p_c_enable_103), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[2] [22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[22__239 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[21__240  (.D(wb_odata[21]), .SP(dac_clk_p_c_enable_103), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[2] [21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[21__240 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[20__241  (.D(wb_odata[20]), .SP(dac_clk_p_c_enable_103), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[2] [20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[20__241 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[19__242  (.D(wb_odata[19]), .SP(dac_clk_p_c_enable_103), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[2] [19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[19__242 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[18__243  (.D(wb_odata[18]), .SP(dac_clk_p_c_enable_103), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[2] [18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[18__243 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[17__244  (.D(wb_odata[17]), .SP(dac_clk_p_c_enable_103), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[2] [17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[17__244 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[16__245  (.D(wb_odata[16]), .SP(dac_clk_p_c_enable_103), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[2] [16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[16__245 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[15__246  (.D(wb_odata[15]), .SP(dac_clk_p_c_enable_103), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[2] [15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[15__246 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[14__247  (.D(wb_odata[14]), .SP(dac_clk_p_c_enable_103), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[2] [14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[14__247 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[13__248  (.D(wb_odata[13]), .SP(dac_clk_p_c_enable_103), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[2] [13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[13__248 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[12__249  (.D(wb_odata[12]), .SP(dac_clk_p_c_enable_103), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[2] [12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[12__249 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[11__250  (.D(wb_odata[11]), .SP(dac_clk_p_c_enable_103), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[2] [11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[11__250 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[10__251  (.D(wb_odata[10]), .SP(dac_clk_p_c_enable_103), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[2] [10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[10__251 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[9__252  (.D(wb_odata[9]), .SP(dac_clk_p_c_enable_103), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[2] [9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[9__252 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[8__253  (.D(wb_odata[8]), .SP(dac_clk_p_c_enable_103), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[2] [8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[8__253 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[7__254  (.D(wb_odata[7]), .SP(dac_clk_p_c_enable_103), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[2] [7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[7__254 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[6__255  (.D(wb_odata[6]), .SP(dac_clk_p_c_enable_103), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[2] [6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[6__255 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[5__256  (.D(wb_odata[5]), .SP(dac_clk_p_c_enable_103), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[2] [5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[5__256 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[4__257  (.D(wb_odata[4]), .SP(dac_clk_p_c_enable_103), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[2] [4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[4__257 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[3__258  (.D(wb_odata[3]), .SP(dac_clk_p_c_enable_103), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[2] [3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[3__258 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[2__259  (.D(wb_odata[2]), .SP(dac_clk_p_c_enable_103), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[2] [2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[2__259 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[1__260  (.D(wb_odata[1]), .SP(dac_clk_p_c_enable_103), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[2] [1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[1__260 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[0__261  (.D(wb_odata[0]), .SP(dac_clk_p_c_enable_103), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[2] [0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_2[[0__261 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[25__275  (.D(wb_odata[25]), .SP(dac_clk_p_c_enable_143), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[25__275 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[24__277  (.D(wb_odata[24]), .SP(dac_clk_p_c_enable_143), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[24__277 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[23__279  (.D(wb_odata[23]), .SP(dac_clk_p_c_enable_143), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[23__279 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[22__281  (.D(wb_odata[22]), .SP(dac_clk_p_c_enable_143), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[22__281 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[21__283  (.D(wb_odata[21]), .SP(dac_clk_p_c_enable_143), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[21__283 .GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i0 (.D(n1[0]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(carrier_center_increment_offset_ls[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_center_increment_offset_ls__i0.GSR = "DISABLED";
    FD1S3AX o_wb_data_i0 (.D(o_wb_data_31__N_1337[0]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i0.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_rs_i1 (.D(carrier_center_increment_offset_rs_30__N_1560[0]), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(carrier_center_increment_offset_rs[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_center_increment_offset_rs_i1.GSR = "DISABLED";
    FD1P3AX \addr_space_3[[20__285  (.D(wb_odata[20]), .SP(dac_clk_p_c_enable_143), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[20__285 .GSR = "DISABLED";
    FD1S3DX carrier_increment_i0 (.D(carrier_increment_30__N_1591[0]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(carrier_increment[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_increment_i0.GSR = "DISABLED";
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i0 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[0]), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(sine_lookup_width_minus_modulation_deviation_amount[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i0.GSR = "DISABLED";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i0 (.D(\addr_space[2] [0]), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(modulation_deviation_amount_minus_sine_lookup_width[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i0.GSR = "DISABLED";
    FD1P3DX \addr_space_0[[31__165  (.D(wb_odata[31]), .SP(dac_clk_p_c_enable_114), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(\addr_space[0] [31])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[31__165 .GSR = "DISABLED";
    FD1P3BX \addr_space_0[[22__175  (.D(wb_odata[22]), .SP(dac_clk_p_c_enable_114), 
            .CK(dac_clk_p_c), .PD(n26683), .Q(\addr_space[0] [22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_0[[22__175 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[19__287  (.D(wb_odata[19]), .SP(dac_clk_p_c_enable_143), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[19__287 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[18__289  (.D(wb_odata[18]), .SP(dac_clk_p_c_enable_143), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[18__289 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[17__291  (.D(wb_odata[17]), .SP(dac_clk_p_c_enable_143), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[17__291 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[16__293  (.D(wb_odata[16]), .SP(dac_clk_p_c_enable_143), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[16__293 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[15__295  (.D(wb_odata[15]), .SP(dac_clk_p_c_enable_143), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[15__295 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[14__297  (.D(wb_odata[14]), .SP(dac_clk_p_c_enable_143), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[14__297 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[13__299  (.D(wb_odata[13]), .SP(dac_clk_p_c_enable_143), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[13__299 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[12__301  (.D(wb_odata[12]), .SP(dac_clk_p_c_enable_143), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[12__301 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[11__303  (.D(wb_odata[11]), .SP(dac_clk_p_c_enable_143), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[11__303 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[10__305  (.D(wb_odata[10]), .SP(dac_clk_p_c_enable_143), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[10__305 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[9__307  (.D(wb_odata[9]), .SP(dac_clk_p_c_enable_143), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[9__307 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[8__309  (.D(wb_odata[8]), .SP(dac_clk_p_c_enable_143), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[8__309 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[7__311  (.D(wb_odata[7]), .SP(dac_clk_p_c_enable_143), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[7__311 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[6__313  (.D(wb_odata[6]), .SP(dac_clk_p_c_enable_143), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[6__313 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[5__315  (.D(wb_odata[5]), .SP(dac_clk_p_c_enable_143), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[5__315 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[4__317  (.D(wb_odata[4]), .SP(dac_clk_p_c_enable_143), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[4__317 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[3__319  (.D(wb_odata[3]), .SP(dac_clk_p_c_enable_143), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[3__319 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[2__321  (.D(wb_odata[2]), .SP(dac_clk_p_c_enable_143), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[2__321 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[1__323  (.D(wb_odata[1]), .SP(dac_clk_p_c_enable_143), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[1__323 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[0__325  (.D(wb_odata[0]), .SP(dac_clk_p_c_enable_143), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[0__325 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[31__263  (.D(wb_odata[31]), .SP(dac_clk_p_c_enable_143), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [31])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[11] 47[5])
    defparam \addr_space_3[[31__263 .GSR = "DISABLED";
    PFUMX i19422 (.BLUT(n21740), .ALUT(n21741), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[30]));
    FD1S3IX o_wb_ack_327 (.D(o_dac_a_9__N_1), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(wb_fm_ack)) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(54[8] 59[4])
    defparam o_wb_ack_327.GSR = "DISABLED";
    PFUMX i6621 (.BLUT(n63), .ALUT(n94), .C0(n22092), .Z(carrier_center_increment_offset_rs_30__N_1560[0]));
    PFUMX i6623 (.BLUT(n64), .ALUT(n95), .C0(n22092), .Z(carrier_center_increment_offset_rs_30__N_1560[1]));
    CCU2D add_379_31 (.A0(\addr_space[0] [29]), .B0(n14347), .C0(carrier_center_increment_offset_rs[30]), 
          .D0(carrier_center_increment_offset_ls[29]), .A1(\addr_space[0] [30]), 
          .B1(n14347), .C1(carrier_center_increment_offset_rs[30]), .D1(carrier_center_increment_offset_ls[30]), 
          .CIN(n17377), .S0(carrier_increment_30__N_1591[29]), .S1(carrier_increment_30__N_1591[30]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(103[4:87])
    defparam add_379_31.INIT0 = 16'h569a;
    defparam add_379_31.INIT1 = 16'h569a;
    defparam add_379_31.INJECT1_0 = "NO";
    defparam add_379_31.INJECT1_1 = "NO";
    CCU2D add_379_29 (.A0(\addr_space[0] [27]), .B0(n14347), .C0(carrier_center_increment_offset_rs[30]), 
          .D0(carrier_center_increment_offset_ls[27]), .A1(\addr_space[0] [28]), 
          .B1(n14347), .C1(carrier_center_increment_offset_rs[30]), .D1(carrier_center_increment_offset_ls[28]), 
          .CIN(n17376), .COUT(n17377), .S0(carrier_increment_30__N_1591[27]), 
          .S1(carrier_increment_30__N_1591[28]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(103[4:87])
    defparam add_379_29.INIT0 = 16'h569a;
    defparam add_379_29.INIT1 = 16'h569a;
    defparam add_379_29.INJECT1_0 = "NO";
    defparam add_379_29.INJECT1_1 = "NO";
    CCU2D add_379_27 (.A0(\addr_space[0] [25]), .B0(n14347), .C0(carrier_center_increment_offset_rs[30]), 
          .D0(carrier_center_increment_offset_ls[25]), .A1(\addr_space[0] [26]), 
          .B1(n14347), .C1(carrier_center_increment_offset_rs[30]), .D1(carrier_center_increment_offset_ls[26]), 
          .CIN(n17375), .COUT(n17376), .S0(carrier_increment_30__N_1591[25]), 
          .S1(carrier_increment_30__N_1591[26]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(103[4:87])
    defparam add_379_27.INIT0 = 16'h569a;
    defparam add_379_27.INIT1 = 16'h569a;
    defparam add_379_27.INJECT1_0 = "NO";
    defparam add_379_27.INJECT1_1 = "NO";
    CCU2D add_379_25 (.A0(\addr_space[0] [23]), .B0(n14347), .C0(carrier_center_increment_offset_rs[30]), 
          .D0(carrier_center_increment_offset_ls[23]), .A1(\addr_space[0] [24]), 
          .B1(n14347), .C1(carrier_center_increment_offset_rs[30]), .D1(carrier_center_increment_offset_ls[24]), 
          .CIN(n17374), .COUT(n17375), .S0(carrier_increment_30__N_1591[23]), 
          .S1(carrier_increment_30__N_1591[24]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(103[4:87])
    defparam add_379_25.INIT0 = 16'h569a;
    defparam add_379_25.INIT1 = 16'h569a;
    defparam add_379_25.INJECT1_0 = "NO";
    defparam add_379_25.INJECT1_1 = "NO";
    CCU2D add_379_23 (.A0(\addr_space[0] [21]), .B0(n14347), .C0(carrier_center_increment_offset_rs[30]), 
          .D0(carrier_center_increment_offset_ls[21]), .A1(\addr_space[0] [22]), 
          .B1(n14347), .C1(carrier_center_increment_offset_rs[30]), .D1(carrier_center_increment_offset_ls[22]), 
          .CIN(n17373), .COUT(n17374), .S0(carrier_increment_30__N_1591[21]), 
          .S1(carrier_increment_30__N_1591[22]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(103[4:87])
    defparam add_379_23.INIT0 = 16'h569a;
    defparam add_379_23.INIT1 = 16'h569a;
    defparam add_379_23.INJECT1_0 = "NO";
    defparam add_379_23.INJECT1_1 = "NO";
    CCU2D add_379_21 (.A0(\addr_space[0] [19]), .B0(n14347), .C0(carrier_center_increment_offset_rs[30]), 
          .D0(carrier_center_increment_offset_ls[19]), .A1(\addr_space[0] [20]), 
          .B1(n14347), .C1(carrier_center_increment_offset_rs[30]), .D1(carrier_center_increment_offset_ls[20]), 
          .CIN(n17372), .COUT(n17373), .S0(carrier_increment_30__N_1591[19]), 
          .S1(carrier_increment_30__N_1591[20]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(103[4:87])
    defparam add_379_21.INIT0 = 16'h569a;
    defparam add_379_21.INIT1 = 16'h569a;
    defparam add_379_21.INJECT1_0 = "NO";
    defparam add_379_21.INJECT1_1 = "NO";
    CCU2D add_379_19 (.A0(\addr_space[0] [17]), .B0(n14347), .C0(carrier_center_increment_offset_rs[30]), 
          .D0(carrier_center_increment_offset_ls[17]), .A1(\addr_space[0] [18]), 
          .B1(n14347), .C1(carrier_center_increment_offset_rs[30]), .D1(carrier_center_increment_offset_ls[18]), 
          .CIN(n17371), .COUT(n17372), .S0(carrier_increment_30__N_1591[17]), 
          .S1(carrier_increment_30__N_1591[18]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(103[4:87])
    defparam add_379_19.INIT0 = 16'h569a;
    defparam add_379_19.INIT1 = 16'h569a;
    defparam add_379_19.INJECT1_0 = "NO";
    defparam add_379_19.INJECT1_1 = "NO";
    CCU2D add_379_17 (.A0(\addr_space[0] [15]), .B0(n14347), .C0(carrier_center_increment_offset_rs[30]), 
          .D0(carrier_center_increment_offset_ls[15]), .A1(\addr_space[0] [16]), 
          .B1(n14347), .C1(carrier_center_increment_offset_rs[30]), .D1(carrier_center_increment_offset_ls[16]), 
          .CIN(n17370), .COUT(n17371), .S0(carrier_increment_30__N_1591[15]), 
          .S1(carrier_increment_30__N_1591[16]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(103[4:87])
    defparam add_379_17.INIT0 = 16'h569a;
    defparam add_379_17.INIT1 = 16'h569a;
    defparam add_379_17.INJECT1_0 = "NO";
    defparam add_379_17.INJECT1_1 = "NO";
    CCU2D add_379_15 (.A0(\addr_space[0] [13]), .B0(n14347), .C0(carrier_center_increment_offset_rs[13]), 
          .D0(carrier_center_increment_offset_ls[13]), .A1(\addr_space[0] [14]), 
          .B1(n14347), .C1(carrier_center_increment_offset_rs[14]), .D1(carrier_center_increment_offset_ls[14]), 
          .CIN(n17369), .COUT(n17370), .S0(carrier_increment_30__N_1591[13]), 
          .S1(carrier_increment_30__N_1591[14]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(103[4:87])
    defparam add_379_15.INIT0 = 16'h569a;
    defparam add_379_15.INIT1 = 16'h569a;
    defparam add_379_15.INJECT1_0 = "NO";
    defparam add_379_15.INJECT1_1 = "NO";
    CCU2D add_379_13 (.A0(\addr_space[0] [11]), .B0(n14347), .C0(carrier_center_increment_offset_rs[11]), 
          .D0(carrier_center_increment_offset_ls[11]), .A1(\addr_space[0] [12]), 
          .B1(n14347), .C1(carrier_center_increment_offset_rs[12]), .D1(carrier_center_increment_offset_ls[12]), 
          .CIN(n17368), .COUT(n17369), .S0(carrier_increment_30__N_1591[11]), 
          .S1(carrier_increment_30__N_1591[12]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(103[4:87])
    defparam add_379_13.INIT0 = 16'h569a;
    defparam add_379_13.INIT1 = 16'h569a;
    defparam add_379_13.INJECT1_0 = "NO";
    defparam add_379_13.INJECT1_1 = "NO";
    CCU2D add_379_11 (.A0(\addr_space[0] [9]), .B0(n14347), .C0(carrier_center_increment_offset_rs[9]), 
          .D0(carrier_center_increment_offset_ls[9]), .A1(\addr_space[0] [10]), 
          .B1(n14347), .C1(carrier_center_increment_offset_rs[10]), .D1(carrier_center_increment_offset_ls[10]), 
          .CIN(n17367), .COUT(n17368), .S0(carrier_increment_30__N_1591[9]), 
          .S1(carrier_increment_30__N_1591[10]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(103[4:87])
    defparam add_379_11.INIT0 = 16'h569a;
    defparam add_379_11.INIT1 = 16'h569a;
    defparam add_379_11.INJECT1_0 = "NO";
    defparam add_379_11.INJECT1_1 = "NO";
    PFUMX i19425 (.BLUT(n21743), .ALUT(n21744), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[29]));
    CCU2D add_379_9 (.A0(\addr_space[0] [7]), .B0(n14347), .C0(carrier_center_increment_offset_rs[7]), 
          .D0(carrier_center_increment_offset_ls[7]), .A1(\addr_space[0] [8]), 
          .B1(n14347), .C1(carrier_center_increment_offset_rs[8]), .D1(carrier_center_increment_offset_ls[8]), 
          .CIN(n17366), .COUT(n17367), .S0(carrier_increment_30__N_1591[7]), 
          .S1(carrier_increment_30__N_1591[8]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(103[4:87])
    defparam add_379_9.INIT0 = 16'h569a;
    defparam add_379_9.INIT1 = 16'h569a;
    defparam add_379_9.INJECT1_0 = "NO";
    defparam add_379_9.INJECT1_1 = "NO";
    CCU2D add_379_7 (.A0(\addr_space[0] [5]), .B0(n14347), .C0(carrier_center_increment_offset_rs[5]), 
          .D0(carrier_center_increment_offset_ls[5]), .A1(\addr_space[0] [6]), 
          .B1(n14347), .C1(carrier_center_increment_offset_rs[6]), .D1(carrier_center_increment_offset_ls[6]), 
          .CIN(n17365), .COUT(n17366), .S0(carrier_increment_30__N_1591[5]), 
          .S1(carrier_increment_30__N_1591[6]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(103[4:87])
    defparam add_379_7.INIT0 = 16'h569a;
    defparam add_379_7.INIT1 = 16'h569a;
    defparam add_379_7.INJECT1_0 = "NO";
    defparam add_379_7.INJECT1_1 = "NO";
    CCU2D add_379_5 (.A0(\addr_space[0] [3]), .B0(n14347), .C0(carrier_center_increment_offset_rs[3]), 
          .D0(carrier_center_increment_offset_ls[3]), .A1(\addr_space[0] [4]), 
          .B1(n14347), .C1(carrier_center_increment_offset_rs[4]), .D1(carrier_center_increment_offset_ls[4]), 
          .CIN(n17364), .COUT(n17365), .S0(carrier_increment_30__N_1591[3]), 
          .S1(carrier_increment_30__N_1591[4]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(103[4:87])
    defparam add_379_5.INIT0 = 16'h569a;
    defparam add_379_5.INIT1 = 16'h569a;
    defparam add_379_5.INJECT1_0 = "NO";
    defparam add_379_5.INJECT1_1 = "NO";
    CCU2D add_379_3 (.A0(\addr_space[0] [1]), .B0(n14347), .C0(carrier_center_increment_offset_rs[1]), 
          .D0(carrier_center_increment_offset_ls[1]), .A1(\addr_space[0] [2]), 
          .B1(n14347), .C1(carrier_center_increment_offset_rs[2]), .D1(carrier_center_increment_offset_ls[2]), 
          .CIN(n17363), .COUT(n17364), .S0(carrier_increment_30__N_1591[1]), 
          .S1(carrier_increment_30__N_1591[2]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(103[4:87])
    defparam add_379_3.INIT0 = 16'h569a;
    defparam add_379_3.INIT1 = 16'h569a;
    defparam add_379_3.INJECT1_0 = "NO";
    defparam add_379_3.INJECT1_1 = "NO";
    CCU2D add_379_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\addr_space[0] [0]), .B1(n14347), .C1(carrier_center_increment_offset_rs[0]), 
          .D1(carrier_center_increment_offset_ls[0]), .COUT(n17363), .S1(carrier_increment_30__N_1591[0]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(103[4:87])
    defparam add_379_1.INIT0 = 16'hF000;
    defparam add_379_1.INIT1 = 16'h569a;
    defparam add_379_1.INJECT1_0 = "NO";
    defparam add_379_1.INJECT1_1 = "NO";
    CCU2D sub_391_add_2_17 (.A0(\addr_space[2] [15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\addr_space[2] [16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17361), .S0(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[15]), 
          .S1(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[16]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(96[58:109])
    defparam sub_391_add_2_17.INIT0 = 16'hf555;
    defparam sub_391_add_2_17.INIT1 = 16'hf555;
    defparam sub_391_add_2_17.INJECT1_0 = "NO";
    defparam sub_391_add_2_17.INJECT1_1 = "NO";
    PFUMX i19428 (.BLUT(n21746), .ALUT(n21747), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[28]));
    PFUMX i19431 (.BLUT(n21749), .ALUT(n21750), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[27]));
    PFUMX i19434 (.BLUT(n21752), .ALUT(n21753), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[26]));
    LUT4 mux_388_Mux_1_i3_4_lut_4_lut_4_lut (.A(\wb_addr[0] ), .B(\wb_addr[1] ), 
         .C(\power_counter[1] ), .D(\smpl_register[1] ), .Z(n2035)) /* synthesis lut_function=(A (B (C)+!B (D))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(45[4:25])
    defparam mux_388_Mux_1_i3_4_lut_4_lut_4_lut.init = 16'hb391;
    LUT4 sub_391_inv_0_i1_1_lut (.A(\addr_space[2] [0]), .Z(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[0])) /* synthesis lut_function=(!(A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(96[58:109])
    defparam sub_391_inv_0_i1_1_lut.init = 16'h5555;
    CCU2D sub_391_add_2_15 (.A0(\addr_space[2] [13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\addr_space[2] [14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17360), .COUT(n17361), .S0(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[13]), 
          .S1(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[14]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(96[58:109])
    defparam sub_391_add_2_15.INIT0 = 16'hf555;
    defparam sub_391_add_2_15.INIT1 = 16'hf555;
    defparam sub_391_add_2_15.INJECT1_0 = "NO";
    defparam sub_391_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_391_add_2_13 (.A0(\addr_space[2] [11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\addr_space[2] [12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17359), .COUT(n17360), .S0(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[11]), 
          .S1(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[12]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(96[58:109])
    defparam sub_391_add_2_13.INIT0 = 16'hf555;
    defparam sub_391_add_2_13.INIT1 = 16'hf555;
    defparam sub_391_add_2_13.INJECT1_0 = "NO";
    defparam sub_391_add_2_13.INJECT1_1 = "NO";
    PFUMX i19437 (.BLUT(n21755), .ALUT(n21756), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[25]));
    CCU2D sub_108_add_2_13 (.A0(\addr_space[2] [15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\addr_space[2] [16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17428), .S0(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[15]), 
          .S1(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[16]));
    defparam sub_108_add_2_13.INIT0 = 16'h5555;
    defparam sub_108_add_2_13.INIT1 = 16'h5555;
    defparam sub_108_add_2_13.INJECT1_0 = "NO";
    defparam sub_108_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_108_add_2_11 (.A0(\addr_space[2] [13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\addr_space[2] [14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17427), .COUT(n17428), .S0(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[13]), 
          .S1(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[14]));
    defparam sub_108_add_2_11.INIT0 = 16'h5555;
    defparam sub_108_add_2_11.INIT1 = 16'h5555;
    defparam sub_108_add_2_11.INJECT1_0 = "NO";
    defparam sub_108_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_391_add_2_11 (.A0(\addr_space[2] [9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\addr_space[2] [10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17358), .COUT(n17359), .S0(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[9]), 
          .S1(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[10]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(96[58:109])
    defparam sub_391_add_2_11.INIT0 = 16'hf555;
    defparam sub_391_add_2_11.INIT1 = 16'hf555;
    defparam sub_391_add_2_11.INJECT1_0 = "NO";
    defparam sub_391_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_108_add_2_9 (.A0(\addr_space[2] [11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\addr_space[2] [12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17426), .COUT(n17427), .S0(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[11]), 
          .S1(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[12]));
    defparam sub_108_add_2_9.INIT0 = 16'h5555;
    defparam sub_108_add_2_9.INIT1 = 16'h5555;
    defparam sub_108_add_2_9.INJECT1_0 = "NO";
    defparam sub_108_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_108_add_2_7 (.A0(\addr_space[2] [9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\addr_space[2] [10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17425), .COUT(n17426), .S0(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[9]), 
          .S1(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[10]));
    defparam sub_108_add_2_7.INIT0 = 16'h5555;
    defparam sub_108_add_2_7.INIT1 = 16'h5555;
    defparam sub_108_add_2_7.INJECT1_0 = "NO";
    defparam sub_108_add_2_7.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_395_3_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .B(n26533), .C(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .D(modulation_deviation_amount_minus_sine_lookup_width[2]), .Z(n26355)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam i1_2_lut_rep_395_3_lut_4_lut.init = 16'h0004;
    LUT4 i10922_3_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .B(n26533), .C(modulation_deviation_amount_minus_sine_lookup_width[2]), 
         .D(n58), .Z(n89)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam i10922_3_lut_4_lut.init = 16'h4f40;
    CCU2D sub_108_add_2_5 (.A0(\addr_space[2] [7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\addr_space[2] [8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17424), .COUT(n17425), .S0(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[7]), 
          .S1(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[8]));
    defparam sub_108_add_2_5.INIT0 = 16'h5555;
    defparam sub_108_add_2_5.INIT1 = 16'h5555;
    defparam sub_108_add_2_5.INJECT1_0 = "NO";
    defparam sub_108_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_108_add_2_3 (.A0(\addr_space[2] [5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\addr_space[2] [6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17423), .COUT(n17424), .S0(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[5]), 
          .S1(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[6]));
    defparam sub_108_add_2_3.INIT0 = 16'h5555;
    defparam sub_108_add_2_3.INIT1 = 16'h5555;
    defparam sub_108_add_2_3.INJECT1_0 = "NO";
    defparam sub_108_add_2_3.INJECT1_1 = "NO";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i16 (.D(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[16]), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(modulation_deviation_amount_minus_sine_lookup_width[16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i16.GSR = "DISABLED";
    CCU2D sub_108_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\addr_space[2] [4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n17423), .S1(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[4]));
    defparam sub_108_add_2_1.INIT0 = 16'hF000;
    defparam sub_108_add_2_1.INIT1 = 16'h5555;
    defparam sub_108_add_2_1.INJECT1_0 = "NO";
    defparam sub_108_add_2_1.INJECT1_1 = "NO";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i15 (.D(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[15]), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(modulation_deviation_amount_minus_sine_lookup_width[15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i15.GSR = "DISABLED";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i14 (.D(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[14]), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(modulation_deviation_amount_minus_sine_lookup_width[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i14.GSR = "DISABLED";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i13 (.D(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[13]), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(modulation_deviation_amount_minus_sine_lookup_width[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i13.GSR = "DISABLED";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i12 (.D(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[12]), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(modulation_deviation_amount_minus_sine_lookup_width[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i12.GSR = "DISABLED";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i11 (.D(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[11]), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(modulation_deviation_amount_minus_sine_lookup_width[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i11.GSR = "DISABLED";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i10 (.D(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[10]), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(modulation_deviation_amount_minus_sine_lookup_width[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i10.GSR = "DISABLED";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i9 (.D(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[9]), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(modulation_deviation_amount_minus_sine_lookup_width[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i9.GSR = "DISABLED";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i8 (.D(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[8]), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(modulation_deviation_amount_minus_sine_lookup_width[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i8.GSR = "DISABLED";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i7 (.D(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[7]), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(modulation_deviation_amount_minus_sine_lookup_width[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i7.GSR = "DISABLED";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i6 (.D(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[6]), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(modulation_deviation_amount_minus_sine_lookup_width[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i6.GSR = "DISABLED";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i5 (.D(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[5]), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(modulation_deviation_amount_minus_sine_lookup_width[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i5.GSR = "DISABLED";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i4 (.D(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[4]), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(modulation_deviation_amount_minus_sine_lookup_width[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i4.GSR = "DISABLED";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i3 (.D(\addr_space[2] [3]), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(modulation_deviation_amount_minus_sine_lookup_width[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i3.GSR = "DISABLED";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i2 (.D(\addr_space[2] [2]), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(modulation_deviation_amount_minus_sine_lookup_width[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i2.GSR = "DISABLED";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i1 (.D(\addr_space[2] [1]), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(modulation_deviation_amount_minus_sine_lookup_width[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i1.GSR = "DISABLED";
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i16 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[16]), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(sine_lookup_width_minus_modulation_deviation_amount[16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i16.GSR = "DISABLED";
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i15 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[15]), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(sine_lookup_width_minus_modulation_deviation_amount[15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i15.GSR = "DISABLED";
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i14 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[14]), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(sine_lookup_width_minus_modulation_deviation_amount[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i14.GSR = "DISABLED";
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i13 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[13]), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(sine_lookup_width_minus_modulation_deviation_amount[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i13.GSR = "DISABLED";
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i12 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[12]), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(sine_lookup_width_minus_modulation_deviation_amount[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i12.GSR = "DISABLED";
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i11 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[11]), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(sine_lookup_width_minus_modulation_deviation_amount[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i11.GSR = "DISABLED";
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i10 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[10]), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(sine_lookup_width_minus_modulation_deviation_amount[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i10.GSR = "DISABLED";
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i9 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[9]), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(sine_lookup_width_minus_modulation_deviation_amount[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i9.GSR = "DISABLED";
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i8 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[8]), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(sine_lookup_width_minus_modulation_deviation_amount[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i8.GSR = "DISABLED";
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i7 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[7]), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(sine_lookup_width_minus_modulation_deviation_amount[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i7.GSR = "DISABLED";
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i6 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[6]), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(sine_lookup_width_minus_modulation_deviation_amount[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i6.GSR = "DISABLED";
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i5 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[5]), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(sine_lookup_width_minus_modulation_deviation_amount[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i5.GSR = "DISABLED";
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i4 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[4]), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(sine_lookup_width_minus_modulation_deviation_amount[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i4.GSR = "DISABLED";
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i3 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[3]), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(sine_lookup_width_minus_modulation_deviation_amount[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i3.GSR = "DISABLED";
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i2 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[2]), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(sine_lookup_width_minus_modulation_deviation_amount[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i2.GSR = "DISABLED";
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i1 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[1]), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(sine_lookup_width_minus_modulation_deviation_amount[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i1.GSR = "DISABLED";
    FD1S3DX carrier_increment_i30 (.D(carrier_increment_30__N_1591[30]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(carrier_increment[30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_increment_i30.GSR = "DISABLED";
    FD1S3DX carrier_increment_i29 (.D(carrier_increment_30__N_1591[29]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(carrier_increment[29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_increment_i29.GSR = "DISABLED";
    FD1S3DX carrier_increment_i28 (.D(carrier_increment_30__N_1591[28]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(carrier_increment[28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_increment_i28.GSR = "DISABLED";
    FD1S3DX carrier_increment_i27 (.D(carrier_increment_30__N_1591[27]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(carrier_increment[27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_increment_i27.GSR = "DISABLED";
    CCU2D sub_391_add_2_9 (.A0(\addr_space[2] [7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\addr_space[2] [8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17357), .COUT(n17358), .S0(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[7]), 
          .S1(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[8]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(96[58:109])
    defparam sub_391_add_2_9.INIT0 = 16'hf555;
    defparam sub_391_add_2_9.INIT1 = 16'hf555;
    defparam sub_391_add_2_9.INJECT1_0 = "NO";
    defparam sub_391_add_2_9.INJECT1_1 = "NO";
    FD1S3DX carrier_increment_i26 (.D(carrier_increment_30__N_1591[26]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(carrier_increment[26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_increment_i26.GSR = "DISABLED";
    FD1S3DX carrier_increment_i25 (.D(carrier_increment_30__N_1591[25]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(carrier_increment[25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_increment_i25.GSR = "DISABLED";
    FD1S3DX carrier_increment_i24 (.D(carrier_increment_30__N_1591[24]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(carrier_increment[24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_increment_i24.GSR = "DISABLED";
    CCU2D sub_391_add_2_7 (.A0(\addr_space[2] [5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\addr_space[2] [6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17356), .COUT(n17357), .S0(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[5]), 
          .S1(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[6]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(96[58:109])
    defparam sub_391_add_2_7.INIT0 = 16'hf555;
    defparam sub_391_add_2_7.INIT1 = 16'hf555;
    defparam sub_391_add_2_7.INJECT1_0 = "NO";
    defparam sub_391_add_2_7.INJECT1_1 = "NO";
    FD1S3DX carrier_increment_i23 (.D(carrier_increment_30__N_1591[23]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(carrier_increment[23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_increment_i23.GSR = "DISABLED";
    FD1S3DX carrier_increment_i22 (.D(carrier_increment_30__N_1591[22]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(carrier_increment[22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_increment_i22.GSR = "DISABLED";
    FD1S3DX carrier_increment_i21 (.D(carrier_increment_30__N_1591[21]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(carrier_increment[21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_increment_i21.GSR = "DISABLED";
    FD1S3DX carrier_increment_i20 (.D(carrier_increment_30__N_1591[20]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(carrier_increment[20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_increment_i20.GSR = "DISABLED";
    FD1S3DX carrier_increment_i19 (.D(carrier_increment_30__N_1591[19]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(carrier_increment[19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_increment_i19.GSR = "DISABLED";
    FD1S3DX carrier_increment_i18 (.D(carrier_increment_30__N_1591[18]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(carrier_increment[18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_increment_i18.GSR = "DISABLED";
    FD1S3DX carrier_increment_i17 (.D(carrier_increment_30__N_1591[17]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(carrier_increment[17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_increment_i17.GSR = "DISABLED";
    FD1S3DX carrier_increment_i16 (.D(carrier_increment_30__N_1591[16]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(carrier_increment[16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_increment_i16.GSR = "DISABLED";
    FD1S3DX carrier_increment_i15 (.D(carrier_increment_30__N_1591[15]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(carrier_increment[15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_increment_i15.GSR = "DISABLED";
    FD1S3DX carrier_increment_i14 (.D(carrier_increment_30__N_1591[14]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(carrier_increment[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_increment_i14.GSR = "DISABLED";
    FD1S3DX carrier_increment_i13 (.D(carrier_increment_30__N_1591[13]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(carrier_increment[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_increment_i13.GSR = "DISABLED";
    FD1S3DX carrier_increment_i12 (.D(carrier_increment_30__N_1591[12]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(carrier_increment[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_increment_i12.GSR = "DISABLED";
    FD1S3DX carrier_increment_i11 (.D(carrier_increment_30__N_1591[11]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(carrier_increment[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_increment_i11.GSR = "DISABLED";
    FD1S3DX carrier_increment_i10 (.D(carrier_increment_30__N_1591[10]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(carrier_increment[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_increment_i10.GSR = "DISABLED";
    FD1S3DX carrier_increment_i9 (.D(carrier_increment_30__N_1591[9]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(carrier_increment[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_increment_i9.GSR = "DISABLED";
    FD1S3DX carrier_increment_i8 (.D(carrier_increment_30__N_1591[8]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(carrier_increment[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_increment_i8.GSR = "DISABLED";
    FD1S3DX carrier_increment_i7 (.D(carrier_increment_30__N_1591[7]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(carrier_increment[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_increment_i7.GSR = "DISABLED";
    FD1S3DX carrier_increment_i6 (.D(carrier_increment_30__N_1591[6]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(carrier_increment[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_increment_i6.GSR = "DISABLED";
    FD1S3DX carrier_increment_i5 (.D(carrier_increment_30__N_1591[5]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(carrier_increment[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_increment_i5.GSR = "DISABLED";
    FD1S3DX carrier_increment_i4 (.D(carrier_increment_30__N_1591[4]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(carrier_increment[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_increment_i4.GSR = "DISABLED";
    FD1S3DX carrier_increment_i3 (.D(carrier_increment_30__N_1591[3]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(carrier_increment[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_increment_i3.GSR = "DISABLED";
    FD1S3DX carrier_increment_i2 (.D(carrier_increment_30__N_1591[2]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(carrier_increment[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_increment_i2.GSR = "DISABLED";
    FD1S3DX carrier_increment_i1 (.D(carrier_increment_30__N_1591[1]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(carrier_increment[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_increment_i1.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_rs_i16 (.D(modulation_output[15]), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(carrier_center_increment_offset_rs[30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_center_increment_offset_rs_i16.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_rs_i15 (.D(carrier_center_increment_offset_rs_30__N_1560[14]), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(carrier_center_increment_offset_rs[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_center_increment_offset_rs_i15.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_rs_i14 (.D(carrier_center_increment_offset_rs_30__N_1560[13]), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(carrier_center_increment_offset_rs[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_center_increment_offset_rs_i14.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_rs_i13 (.D(carrier_center_increment_offset_rs_30__N_1560[12]), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(carrier_center_increment_offset_rs[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_center_increment_offset_rs_i13.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_rs_i12 (.D(carrier_center_increment_offset_rs_30__N_1560[11]), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(carrier_center_increment_offset_rs[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_center_increment_offset_rs_i12.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_rs_i11 (.D(carrier_center_increment_offset_rs_30__N_1560[10]), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(carrier_center_increment_offset_rs[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_center_increment_offset_rs_i11.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_rs_i10 (.D(carrier_center_increment_offset_rs_30__N_1560[9]), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(carrier_center_increment_offset_rs[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_center_increment_offset_rs_i10.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_rs_i9 (.D(carrier_center_increment_offset_rs_30__N_1560[8]), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(carrier_center_increment_offset_rs[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_center_increment_offset_rs_i9.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_rs_i8 (.D(carrier_center_increment_offset_rs_30__N_1560[7]), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(carrier_center_increment_offset_rs[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_center_increment_offset_rs_i8.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_rs_i7 (.D(carrier_center_increment_offset_rs_30__N_1560[6]), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(carrier_center_increment_offset_rs[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_center_increment_offset_rs_i7.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_rs_i6 (.D(carrier_center_increment_offset_rs_30__N_1560[5]), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(carrier_center_increment_offset_rs[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_center_increment_offset_rs_i6.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_rs_i5 (.D(carrier_center_increment_offset_rs_30__N_1560[4]), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(carrier_center_increment_offset_rs[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_center_increment_offset_rs_i5.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_rs_i4 (.D(carrier_center_increment_offset_rs_30__N_1560[3]), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(carrier_center_increment_offset_rs[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_center_increment_offset_rs_i4.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_rs_i3 (.D(carrier_center_increment_offset_rs_30__N_1560[2]), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(carrier_center_increment_offset_rs[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_center_increment_offset_rs_i3.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_rs_i2 (.D(carrier_center_increment_offset_rs_30__N_1560[1]), 
            .CK(dac_clk_p_c), .CD(n26683), .Q(carrier_center_increment_offset_rs[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_center_increment_offset_rs_i2.GSR = "DISABLED";
    FD1S3AX o_wb_data_i31 (.D(o_wb_data_31__N_1337[31]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[31])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i31.GSR = "DISABLED";
    FD1S3AX o_wb_data_i30 (.D(o_wb_data_31__N_1337[30]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i30.GSR = "DISABLED";
    FD1S3AX o_wb_data_i29 (.D(o_wb_data_31__N_1337[29]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i29.GSR = "DISABLED";
    FD1S3AX o_wb_data_i28 (.D(o_wb_data_31__N_1337[28]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i28.GSR = "DISABLED";
    FD1S3AX o_wb_data_i27 (.D(o_wb_data_31__N_1337[27]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i27.GSR = "DISABLED";
    FD1S3AX o_wb_data_i26 (.D(o_wb_data_31__N_1337[26]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i26.GSR = "DISABLED";
    FD1S3AX o_wb_data_i25 (.D(o_wb_data_31__N_1337[25]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i25.GSR = "DISABLED";
    FD1S3AX o_wb_data_i24 (.D(o_wb_data_31__N_1337[24]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i24.GSR = "DISABLED";
    FD1S3AX o_wb_data_i23 (.D(o_wb_data_31__N_1337[23]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i23.GSR = "DISABLED";
    FD1S3AX o_wb_data_i22 (.D(o_wb_data_31__N_1337[22]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i22.GSR = "DISABLED";
    FD1S3AX o_wb_data_i21 (.D(o_wb_data_31__N_1337[21]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i21.GSR = "DISABLED";
    FD1S3AX o_wb_data_i20 (.D(o_wb_data_31__N_1337[20]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i20.GSR = "DISABLED";
    FD1S3AX o_wb_data_i19 (.D(o_wb_data_31__N_1337[19]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i19.GSR = "DISABLED";
    FD1S3AX o_wb_data_i18 (.D(o_wb_data_31__N_1337[18]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i18.GSR = "DISABLED";
    FD1S3AX o_wb_data_i17 (.D(o_wb_data_31__N_1337[17]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i17.GSR = "DISABLED";
    FD1S3AX o_wb_data_i16 (.D(o_wb_data_31__N_1337[16]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i16.GSR = "DISABLED";
    FD1S3AX o_wb_data_i15 (.D(o_wb_data_31__N_1337[15]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i15.GSR = "DISABLED";
    FD1S3AX o_wb_data_i14 (.D(o_wb_data_31__N_1337[14]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i14.GSR = "DISABLED";
    FD1S3AX o_wb_data_i13 (.D(o_wb_data_31__N_1337[13]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i13.GSR = "DISABLED";
    FD1S3AX o_wb_data_i12 (.D(o_wb_data_31__N_1337[12]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i12.GSR = "DISABLED";
    FD1S3AX o_wb_data_i11 (.D(o_wb_data_31__N_1337[11]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i11.GSR = "DISABLED";
    FD1S3AX o_wb_data_i10 (.D(o_wb_data_31__N_1337[10]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i10.GSR = "DISABLED";
    FD1S3AX o_wb_data_i9 (.D(o_wb_data_31__N_1337[9]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i9.GSR = "DISABLED";
    FD1S3AX o_wb_data_i8 (.D(o_wb_data_31__N_1337[8]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i8.GSR = "DISABLED";
    FD1S3AX o_wb_data_i7 (.D(o_wb_data_31__N_1337[7]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i7.GSR = "DISABLED";
    FD1S3AX o_wb_data_i6 (.D(o_wb_data_31__N_1337[6]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i6.GSR = "DISABLED";
    FD1S3AX o_wb_data_i5 (.D(o_wb_data_31__N_1337[5]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i5.GSR = "DISABLED";
    FD1S3AX o_wb_data_i4 (.D(o_wb_data_31__N_1337[4]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i4.GSR = "DISABLED";
    FD1S3AX o_wb_data_i3 (.D(o_wb_data_31__N_1337[3]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i3.GSR = "DISABLED";
    FD1S3AX o_wb_data_i2 (.D(o_wb_data_31__N_1337[2]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i2.GSR = "DISABLED";
    FD1S3AX o_wb_data_i1 (.D(o_wb_data_31__N_1337[1]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(50[8] 52[4])
    defparam o_wb_data_i1.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i30 (.D(n1[30]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(carrier_center_increment_offset_ls[30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_center_increment_offset_ls__i30.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i29 (.D(n1[29]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(carrier_center_increment_offset_ls[29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_center_increment_offset_ls__i29.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i28 (.D(n1[28]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(carrier_center_increment_offset_ls[28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_center_increment_offset_ls__i28.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i27 (.D(n1[27]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(carrier_center_increment_offset_ls[27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_center_increment_offset_ls__i27.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i26 (.D(n1[26]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(carrier_center_increment_offset_ls[26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_center_increment_offset_ls__i26.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i25 (.D(n1[25]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(carrier_center_increment_offset_ls[25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_center_increment_offset_ls__i25.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i24 (.D(n1[24]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(carrier_center_increment_offset_ls[24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_center_increment_offset_ls__i24.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i23 (.D(n1[23]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(carrier_center_increment_offset_ls[23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_center_increment_offset_ls__i23.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i22 (.D(n1[22]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(carrier_center_increment_offset_ls[22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_center_increment_offset_ls__i22.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i21 (.D(n1[21]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(carrier_center_increment_offset_ls[21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_center_increment_offset_ls__i21.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i20 (.D(n1[20]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(carrier_center_increment_offset_ls[20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_center_increment_offset_ls__i20.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i19 (.D(n1[19]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(carrier_center_increment_offset_ls[19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_center_increment_offset_ls__i19.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i18 (.D(n1[18]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(carrier_center_increment_offset_ls[18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_center_increment_offset_ls__i18.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i17 (.D(n1[17]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(carrier_center_increment_offset_ls[17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_center_increment_offset_ls__i17.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i16 (.D(n1[16]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(carrier_center_increment_offset_ls[16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_center_increment_offset_ls__i16.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i15 (.D(n1[15]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(carrier_center_increment_offset_ls[15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_center_increment_offset_ls__i15.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i14 (.D(n1[14]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(carrier_center_increment_offset_ls[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_center_increment_offset_ls__i14.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i13 (.D(n1[13]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(carrier_center_increment_offset_ls[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_center_increment_offset_ls__i13.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i12 (.D(n1[12]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(carrier_center_increment_offset_ls[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_center_increment_offset_ls__i12.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i11 (.D(n1[11]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(carrier_center_increment_offset_ls[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_center_increment_offset_ls__i11.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i10 (.D(n1[10]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(carrier_center_increment_offset_ls[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_center_increment_offset_ls__i10.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i9 (.D(n1[9]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(carrier_center_increment_offset_ls[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_center_increment_offset_ls__i9.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i8 (.D(n1[8]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(carrier_center_increment_offset_ls[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_center_increment_offset_ls__i8.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i7 (.D(n1[7]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(carrier_center_increment_offset_ls[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_center_increment_offset_ls__i7.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i6 (.D(n1[6]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(carrier_center_increment_offset_ls[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_center_increment_offset_ls__i6.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i5 (.D(n1[5]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(carrier_center_increment_offset_ls[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_center_increment_offset_ls__i5.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i4 (.D(n1[4]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(carrier_center_increment_offset_ls[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_center_increment_offset_ls__i4.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i3 (.D(n1[3]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(carrier_center_increment_offset_ls[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_center_increment_offset_ls__i3.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i2 (.D(n1[2]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(carrier_center_increment_offset_ls[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_center_increment_offset_ls__i2.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i1 (.D(n20073), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(carrier_center_increment_offset_ls[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam carrier_center_increment_offset_ls__i1.GSR = "DISABLED";
    CCU2D sub_391_add_2_5 (.A0(\addr_space[2] [3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\addr_space[2] [4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17355), .COUT(n17356), .S0(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[3]), 
          .S1(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[4]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(96[58:109])
    defparam sub_391_add_2_5.INIT0 = 16'hf555;
    defparam sub_391_add_2_5.INIT1 = 16'h0aaa;
    defparam sub_391_add_2_5.INJECT1_0 = "NO";
    defparam sub_391_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_391_add_2_3 (.A0(\addr_space[2] [1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\addr_space[2] [2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17354), .COUT(n17355), .S0(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[1]), 
          .S1(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[2]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(96[58:109])
    defparam sub_391_add_2_3.INIT0 = 16'hf555;
    defparam sub_391_add_2_3.INIT1 = 16'hf555;
    defparam sub_391_add_2_3.INJECT1_0 = "NO";
    defparam sub_391_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_391_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\addr_space[2] [0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n17354));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(96[58:109])
    defparam sub_391_add_2_1.INIT0 = 16'h0000;
    defparam sub_391_add_2_1.INIT1 = 16'h0aaa;
    defparam sub_391_add_2_1.INJECT1_0 = "NO";
    defparam sub_391_add_2_1.INJECT1_1 = "NO";
    LUT4 i19418_3_lut (.A(\addr_space[2] [31]), .B(\addr_space[3] [31]), 
         .C(\wb_addr[0] ), .Z(n21738)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19418_3_lut.init = 16'hcaca;
    LUT4 i19417_3_lut (.A(\addr_space[0] [31]), .B(\addr_space[1] [31]), 
         .C(\wb_addr[0] ), .Z(n21737)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19417_3_lut.init = 16'hcaca;
    LUT4 i19420_3_lut (.A(\addr_space[0] [30]), .B(\addr_space[1] [30]), 
         .C(\wb_addr[0] ), .Z(n21740)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19420_3_lut.init = 16'hcaca;
    LUT4 i6546_3_lut_4_lut (.A(n26558), .B(modulation_deviation_amount_minus_sine_lookup_width[2]), 
         .C(modulation_output[14]), .D(modulation_output[15]), .Z(n72)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam i6546_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_4_lut (.A(n20634), .B(n20636), .C(n20638), .D(n20624), .Z(n178)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam i1_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut (.A(sine_lookup_width_minus_modulation_deviation_amount[14]), 
         .B(sine_lookup_width_minus_modulation_deviation_amount[5]), .Z(n20634)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i1_4_lut_adj_87 (.A(sine_lookup_width_minus_modulation_deviation_amount[6]), 
         .B(sine_lookup_width_minus_modulation_deviation_amount[15]), .C(sine_lookup_width_minus_modulation_deviation_amount[16]), 
         .D(sine_lookup_width_minus_modulation_deviation_amount[9]), .Z(n20636)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam i1_4_lut_adj_87.init = 16'hfffe;
    LUT4 i1_4_lut_adj_88 (.A(sine_lookup_width_minus_modulation_deviation_amount[12]), 
         .B(sine_lookup_width_minus_modulation_deviation_amount[8]), .C(sine_lookup_width_minus_modulation_deviation_amount[11]), 
         .D(sine_lookup_width_minus_modulation_deviation_amount[13]), .Z(n20638)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam i1_4_lut_adj_88.init = 16'hfffe;
    LUT4 i10909_3_lut (.A(n13449), .B(n36_adj_2995), .C(sine_lookup_width_minus_modulation_deviation_amount[2]), 
         .Z(n13450)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(85[27:78])
    defparam i10909_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i71_3_lut (.A(n40_adj_2996), .B(n44_adj_2997), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[2]), .Z(n71)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_i71_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i40_3_lut (.A(n9), .B(n11), .C(sine_lookup_width_minus_modulation_deviation_amount[1]), 
         .Z(n40_adj_2996)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_i40_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i44_3_lut (.A(n13), .B(n15), .C(sine_lookup_width_minus_modulation_deviation_amount[1]), 
         .Z(n44_adj_2997)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_i44_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i15_3_lut (.A(modulation_output[14]), .B(modulation_output[15]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[0]), .Z(n15)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_i15_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i13_3_lut (.A(modulation_output[12]), .B(modulation_output[13]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[0]), .Z(n13)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_i13_3_lut.init = 16'hcaca;
    LUT4 i10908_3_lut (.A(modulation_output[2]), .B(modulation_output[3]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[0]), .Z(n13449)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(85[27:78])
    defparam i10908_3_lut.init = 16'hcaca;
    LUT4 i10912_3_lut (.A(n13451), .B(n7), .C(sine_lookup_width_minus_modulation_deviation_amount[1]), 
         .Z(n36_adj_2995)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(85[27:78])
    defparam i10912_3_lut.init = 16'hcaca;
    LUT4 i10910_3_lut (.A(modulation_output[4]), .B(modulation_output[5]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[0]), .Z(n13451)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(85[27:78])
    defparam i10910_3_lut.init = 16'hcaca;
    LUT4 i10911_3_lut (.A(modulation_output[6]), .B(modulation_output[7]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[0]), .Z(n7)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(85[27:78])
    defparam i10911_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i9_3_lut (.A(modulation_output[8]), .B(modulation_output[9]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[0]), .Z(n9)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_i9_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i11_3_lut (.A(modulation_output[10]), .B(modulation_output[11]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[0]), .Z(n11)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_i11_3_lut.init = 16'hcaca;
    LUT4 i10907_3_lut (.A(modulation_output[0]), .B(modulation_output[1]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[0]), .Z(n13448)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(85[27:78])
    defparam i10907_3_lut.init = 16'hcaca;
    LUT4 i22414_4_lut (.A(n26409), .B(sine_lookup_width_minus_modulation_deviation_amount[3]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[2]), .D(sine_lookup_width_minus_modulation_deviation_amount[1]), 
         .Z(n22092)) /* synthesis lut_function=(A+!(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam i22414_4_lut.init = 16'haaab;
    LUT4 i10917_3_lut (.A(n13457), .B(n37_adj_2998), .C(sine_lookup_width_minus_modulation_deviation_amount[2]), 
         .Z(n33_adj_2999)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(85[27:78])
    defparam i10917_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i72_3_lut (.A(n41_adj_3000), .B(n45_adj_3001), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[2]), .Z(n72_adj_3002)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_i72_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i45_3_lut (.A(n14), .B(modulation_output[15]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[1]), .Z(n45_adj_3001)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_i45_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i14_3_lut (.A(modulation_output[13]), .B(modulation_output[14]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[0]), .Z(n14)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_i14_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i41_3_lut (.A(n10), .B(n12), .C(sine_lookup_width_minus_modulation_deviation_amount[1]), 
         .Z(n41_adj_3000)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_i41_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i10_3_lut (.A(modulation_output[9]), .B(modulation_output[10]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[0]), .Z(n10)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_i10_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i12_3_lut (.A(modulation_output[11]), .B(modulation_output[12]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[0]), .Z(n12)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_i12_3_lut.init = 16'hcaca;
    LUT4 i10916_3_lut (.A(modulation_output[3]), .B(modulation_output[4]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[0]), .Z(n13457)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(85[27:78])
    defparam i10916_3_lut.init = 16'hcaca;
    LUT4 i19415_3_lut (.A(\addr_space[2] [0]), .B(\addr_space[3] [0]), .C(\wb_addr[0] ), 
         .Z(n21735)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19415_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_89 (.A(sine_lookup_width_minus_modulation_deviation_amount[7]), 
         .B(sine_lookup_width_minus_modulation_deviation_amount[10]), .Z(n20624)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam i1_2_lut_adj_89.init = 16'heeee;
    LUT4 modulation_output_15__I_0_i37_3_lut (.A(n6), .B(n8), .C(sine_lookup_width_minus_modulation_deviation_amount[1]), 
         .Z(n37_adj_2998)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_i37_3_lut.init = 16'hcaca;
    LUT4 i10918_3_lut (.A(modulation_output[5]), .B(modulation_output[6]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[0]), .Z(n6)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(85[27:78])
    defparam i10918_3_lut.init = 16'hcaca;
    LUT4 i10924_3_lut (.A(modulation_output[7]), .B(modulation_output[8]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[0]), .Z(n8)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(85[27:78])
    defparam i10924_3_lut.init = 16'hcaca;
    LUT4 i10915_3_lut (.A(modulation_output[1]), .B(modulation_output[2]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[0]), .Z(n13456)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(85[27:78])
    defparam i10915_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i38_3_lut (.A(n7), .B(n9), .C(sine_lookup_width_minus_modulation_deviation_amount[1]), 
         .Z(n38_adj_3003)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_i38_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i73_3_lut (.A(n42_adj_3004), .B(n46_adj_3005), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[2]), .Z(n73)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_i73_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i42_3_lut (.A(n11), .B(n13), .C(sine_lookup_width_minus_modulation_deviation_amount[1]), 
         .Z(n42_adj_3004)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_i42_3_lut.init = 16'hcaca;
    LUT4 i19414_3_lut (.A(\addr_space[0] [0]), .B(\addr_space[1] [0]), .C(\wb_addr[0] ), 
         .Z(n21734)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19414_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_90 (.A(n20348), .B(n20362), .C(n20360), .D(\addr_space[2] [4]), 
         .Z(n14347)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_90.init = 16'hfffe;
    LUT4 i1_2_lut_adj_91 (.A(\addr_space[2] [12]), .B(\addr_space[2] [13]), 
         .Z(n20348)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_91.init = 16'heeee;
    LUT4 i1_4_lut_adj_92 (.A(\addr_space[2] [16]), .B(n20346), .C(n20350), 
         .D(\addr_space[2] [8]), .Z(n20362)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_92.init = 16'hfffe;
    LUT4 i1_4_lut_adj_93 (.A(\addr_space[2] [6]), .B(\addr_space[2] [9]), 
         .C(\addr_space[2] [15]), .D(\addr_space[2] [7]), .Z(n20360)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_93.init = 16'hfffe;
    LUT4 i1_2_lut_adj_94 (.A(\addr_space[2] [5]), .B(\addr_space[2] [14]), 
         .Z(n20346)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_94.init = 16'heeee;
    LUT4 i1_2_lut_adj_95 (.A(\addr_space[2] [11]), .B(\addr_space[2] [10]), 
         .Z(n20350)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_95.init = 16'heeee;
    LUT4 i11874_2_lut_4_lut (.A(n85), .B(n26379), .C(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .D(n26380), .Z(n1[8])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(85[80:131])
    defparam i11874_2_lut_4_lut.init = 16'h00ca;
    LUT4 i18686_3_lut (.A(\addr_space[2] [1]), .B(\addr_space[3] [1]), .C(\wb_addr[0] ), 
         .Z(n21006)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18686_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_336_i112_3_lut_rep_404 (.A(n81), .B(n89), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[3]), .Z(n26364)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam modulation_output_15__I_0_336_i112_3_lut_rep_404.init = 16'hcaca;
    LUT4 i11878_2_lut_4_lut (.A(n81), .B(n89), .C(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .D(n26380), .Z(n1[12])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam i11878_2_lut_4_lut.init = 16'h00ca;
    LUT4 modulation_output_15__I_0_336_i111_3_lut_rep_405 (.A(n80), .B(n88), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[3]), .Z(n26365)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam modulation_output_15__I_0_336_i111_3_lut_rep_405.init = 16'hcaca;
    LUT4 i18685_3_lut (.A(\addr_space[0] [1]), .B(\addr_space[1] [1]), .C(\wb_addr[0] ), 
         .Z(n21005)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18685_3_lut.init = 16'hcaca;
    LUT4 i18683_3_lut (.A(\addr_space[2] [2]), .B(\addr_space[3] [2]), .C(\wb_addr[0] ), 
         .Z(n21003)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18683_3_lut.init = 16'hcaca;
    LUT4 i18682_3_lut (.A(\addr_space[0] [2]), .B(\addr_space[1] [2]), .C(\wb_addr[0] ), 
         .Z(n21002)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18682_3_lut.init = 16'hcaca;
    LUT4 i18680_3_lut (.A(\addr_space[2] [3]), .B(\addr_space[3] [3]), .C(\wb_addr[0] ), 
         .Z(n21000)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18680_3_lut.init = 16'hcaca;
    LUT4 i18679_3_lut (.A(\addr_space[0] [3]), .B(\addr_space[1] [3]), .C(\wb_addr[0] ), 
         .Z(n20999)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18679_3_lut.init = 16'hcaca;
    PFUMX modulation_output_15__I_0_336_i135 (.BLUT(n73_adj_3006), .ALUT(n104), 
          .C0(n21926), .Z(n135)) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;
    LUT4 modulation_output_15__I_0_336_i101_3_lut (.A(modulation_output[15]), 
         .B(n78), .C(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .Z(n101)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam modulation_output_15__I_0_336_i101_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_336_i102_3_lut (.A(modulation_output[15]), 
         .B(n79), .C(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .Z(n102)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam modulation_output_15__I_0_336_i102_3_lut.init = 16'hcaca;
    PFUMX modulation_output_15__I_0_336_i134 (.BLUT(n72), .ALUT(n103), .C0(n21926), 
          .Z(n134)) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;
    LUT4 modulation_output_15__I_0_336_i105_4_lut (.A(n82), .B(n59_adj_3007), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[4]), .D(n26553), 
         .Z(n105)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam modulation_output_15__I_0_336_i105_4_lut.init = 16'hca0a;
    LUT4 modulation_output_15__I_0_336_i74_3_lut (.A(modulation_output[15]), 
         .B(n47_adj_3008), .C(modulation_deviation_amount_minus_sine_lookup_width[2]), 
         .Z(n74)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam modulation_output_15__I_0_336_i74_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_336_i106_4_lut (.A(n83), .B(n60_adj_3009), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[4]), .D(n26553), 
         .Z(n106)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam modulation_output_15__I_0_336_i106_4_lut.init = 16'hca0a;
    LUT4 modulation_output_15__I_0_336_i75_3_lut (.A(modulation_output[15]), 
         .B(n48_adj_3010), .C(modulation_deviation_amount_minus_sine_lookup_width[2]), 
         .Z(n75)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam modulation_output_15__I_0_336_i75_3_lut.init = 16'hcaca;
    LUT4 i19538_3_lut (.A(\addr_space[2] [4]), .B(\addr_space[3] [4]), .C(\wb_addr[0] ), 
         .Z(n21858)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19538_3_lut.init = 16'hcaca;
    LUT4 i11879_2_lut_4_lut (.A(n80), .B(n88), .C(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .D(n26380), .Z(n1[13])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam i11879_2_lut_4_lut.init = 16'h00ca;
    LUT4 modulation_output_15__I_0_336_i110_3_lut_rep_406 (.A(n79), .B(n26399), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[3]), .Z(n26366)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam modulation_output_15__I_0_336_i110_3_lut_rep_406.init = 16'hcaca;
    LUT4 i19537_3_lut (.A(\addr_space[0] [4]), .B(\addr_space[1] [4]), .C(\wb_addr[0] ), 
         .Z(n21857)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19537_3_lut.init = 16'hcaca;
    LUT4 i11880_2_lut_4_lut (.A(n79), .B(n26399), .C(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .D(n26380), .Z(n1[14])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam i11880_2_lut_4_lut.init = 16'h00ca;
    LUT4 i19535_3_lut (.A(\addr_space[2] [5]), .B(\addr_space[3] [5]), .C(\wb_addr[0] ), 
         .Z(n21855)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19535_3_lut.init = 16'hcaca;
    LUT4 i19534_3_lut (.A(\addr_space[0] [5]), .B(\addr_space[1] [5]), .C(\wb_addr[0] ), 
         .Z(n21854)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19534_3_lut.init = 16'hcaca;
    LUT4 i6645_3_lut_4_lut (.A(sine_lookup_width_minus_modulation_deviation_amount[2]), 
         .B(n26400), .C(modulation_output[15]), .D(n44_adj_2997), .Z(carrier_center_increment_offset_rs_30__N_1560[12])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam i6645_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i6643_3_lut_4_lut (.A(sine_lookup_width_minus_modulation_deviation_amount[2]), 
         .B(n26400), .C(modulation_output[15]), .D(n43_adj_3011), .Z(carrier_center_increment_offset_rs_30__N_1560[11])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam i6643_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i19532_3_lut (.A(\addr_space[2] [6]), .B(\addr_space[3] [6]), .C(\wb_addr[0] ), 
         .Z(n21852)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19532_3_lut.init = 16'hcaca;
    LUT4 i19531_3_lut (.A(\addr_space[0] [6]), .B(\addr_space[1] [6]), .C(\wb_addr[0] ), 
         .Z(n21851)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19531_3_lut.init = 16'hcaca;
    LUT4 i19529_3_lut (.A(\addr_space[2] [7]), .B(\addr_space[3] [7]), .C(\wb_addr[0] ), 
         .Z(n21849)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19529_3_lut.init = 16'hcaca;
    LUT4 i19528_3_lut (.A(\addr_space[0] [7]), .B(\addr_space[1] [7]), .C(\wb_addr[0] ), 
         .Z(n21848)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19528_3_lut.init = 16'hcaca;
    LUT4 i19526_3_lut (.A(\addr_space[2] [8]), .B(\addr_space[3] [8]), .C(\wb_addr[0] ), 
         .Z(n21846)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19526_3_lut.init = 16'hcaca;
    LUT4 i19525_3_lut (.A(\addr_space[0] [8]), .B(\addr_space[1] [8]), .C(\wb_addr[0] ), 
         .Z(n21845)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19525_3_lut.init = 16'hcaca;
    PFUMX i24464 (.BLUT(n26325), .ALUT(n26324), .C0(sine_lookup_width_minus_modulation_deviation_amount[3]), 
          .Z(n26326));
    LUT4 i19523_3_lut (.A(\addr_space[2] [9]), .B(\addr_space[3] [9]), .C(\wb_addr[0] ), 
         .Z(n21843)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19523_3_lut.init = 16'hcaca;
    PFUMX i24462 (.BLUT(n26319), .ALUT(n26318), .C0(sine_lookup_width_minus_modulation_deviation_amount[3]), 
          .Z(n26320));
    LUT4 i19522_3_lut (.A(\addr_space[0] [9]), .B(\addr_space[1] [9]), .C(\wb_addr[0] ), 
         .Z(n21842)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19522_3_lut.init = 16'hcaca;
    PFUMX i24459 (.BLUT(n26313), .ALUT(n26312), .C0(sine_lookup_width_minus_modulation_deviation_amount[3]), 
          .Z(n26314));
    LUT4 i19520_3_lut (.A(\addr_space[2] [10]), .B(\addr_space[3] [10]), 
         .C(\wb_addr[0] ), .Z(n21840)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19520_3_lut.init = 16'hcaca;
    LUT4 i19519_3_lut (.A(\addr_space[0] [10]), .B(\addr_space[1] [10]), 
         .C(\wb_addr[0] ), .Z(n21839)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19519_3_lut.init = 16'hcaca;
    LUT4 i19517_3_lut (.A(\addr_space[2] [11]), .B(\addr_space[3] [11]), 
         .C(\wb_addr[0] ), .Z(n21837)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19517_3_lut.init = 16'hcaca;
    LUT4 i19516_3_lut (.A(\addr_space[0] [11]), .B(\addr_space[1] [11]), 
         .C(\wb_addr[0] ), .Z(n21836)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19516_3_lut.init = 16'hcaca;
    LUT4 i19514_3_lut (.A(\addr_space[2] [12]), .B(\addr_space[3] [12]), 
         .C(\wb_addr[0] ), .Z(n21834)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19514_3_lut.init = 16'hcaca;
    PFUMX i24418 (.BLUT(n26267), .ALUT(n39_adj_3012), .C0(sine_lookup_width_minus_modulation_deviation_amount[2]), 
          .Z(n26268));
    LUT4 i19513_3_lut (.A(\addr_space[0] [12]), .B(\addr_space[1] [12]), 
         .C(\wb_addr[0] ), .Z(n21833)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19513_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_96 (.A(n26563), .B(n38), .C(n34), .D(n20488), 
         .Z(dac_clk_p_c_enable_143)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut_adj_96.init = 16'h0100;
    LUT4 i1_4_lut_adj_97 (.A(n20482), .B(\wb_addr[8] ), .C(\wb_addr[12] ), 
         .D(n20480), .Z(n20488)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_4_lut_adj_97.init = 16'h0200;
    LUT4 i19511_3_lut (.A(\addr_space[2] [13]), .B(\addr_space[3] [13]), 
         .C(\wb_addr[0] ), .Z(n21831)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19511_3_lut.init = 16'hcaca;
    LUT4 i19510_3_lut (.A(\addr_space[0] [13]), .B(\addr_space[1] [13]), 
         .C(\wb_addr[0] ), .Z(n21830)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19510_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_98 (.A(n26557), .B(\wb_addr[15] ), .C(\wb_addr[9] ), 
         .D(o_dac_cw_b_c_c), .Z(n20482)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_98.init = 16'h8000;
    LUT4 i1_2_lut_adj_99 (.A(\wb_addr[0] ), .B(\wb_addr[1] ), .Z(n20480)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_99.init = 16'h8888;
    LUT4 i6649_4_lut (.A(modulation_output[14]), .B(modulation_output[15]), 
         .C(n8972), .D(n26400), .Z(carrier_center_increment_offset_rs_30__N_1560[14])) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam i6649_4_lut.init = 16'hccca;
    LUT4 i6647_4_lut (.A(n14), .B(modulation_output[15]), .C(n8970), .D(n26400), 
         .Z(carrier_center_increment_offset_rs_30__N_1560[13])) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam i6647_4_lut.init = 16'hccca;
    LUT4 i6589_2_lut (.A(sine_lookup_width_minus_modulation_deviation_amount[1]), 
         .B(sine_lookup_width_minus_modulation_deviation_amount[2]), .Z(n8970)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam i6589_2_lut.init = 16'heeee;
    LUT4 modulation_output_15__I_0_i43_3_lut (.A(n12), .B(n14), .C(sine_lookup_width_minus_modulation_deviation_amount[1]), 
         .Z(n43_adj_3011)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_i43_3_lut.init = 16'hcaca;
    LUT4 i6641_3_lut (.A(n73), .B(modulation_output[15]), .C(n26400), 
         .Z(carrier_center_increment_offset_rs_30__N_1560[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam i6641_3_lut.init = 16'hcaca;
    LUT4 i6639_3_lut (.A(n72_adj_3002), .B(modulation_output[15]), .C(n26400), 
         .Z(carrier_center_increment_offset_rs_30__N_1560[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam i6639_3_lut.init = 16'hcaca;
    LUT4 i6637_3_lut (.A(n71), .B(modulation_output[15]), .C(n26400), 
         .Z(carrier_center_increment_offset_rs_30__N_1560[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam i6637_3_lut.init = 16'hcaca;
    LUT4 i19508_3_lut (.A(\addr_space[2] [14]), .B(\addr_space[3] [14]), 
         .C(\wb_addr[0] ), .Z(n21828)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19508_3_lut.init = 16'hcaca;
    LUT4 i6635_3_lut (.A(n70), .B(modulation_output[15]), .C(n26400), 
         .Z(carrier_center_increment_offset_rs_30__N_1560[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam i6635_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i70_3_lut (.A(n39_adj_3012), .B(n43_adj_3011), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[2]), .Z(n70)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_i70_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i39_3_lut (.A(n8), .B(n10), .C(sine_lookup_width_minus_modulation_deviation_amount[1]), 
         .Z(n39_adj_3012)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_i39_3_lut.init = 16'hcaca;
    LUT4 i11075_4_lut (.A(modulation_output[15]), .B(n178_adj_3015), .C(n26366), 
         .D(modulation_deviation_amount_minus_sine_lookup_width[4]), .Z(n1[30])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam i11075_4_lut.init = 16'h3022;
    LUT4 modulation_output_15__I_0_336_i79_3_lut (.A(n48_adj_3010), .B(n52_adj_3016), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[2]), .Z(n79)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam modulation_output_15__I_0_336_i79_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_336_i56_3_lut (.A(n25), .B(n27), .C(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .Z(n56_adj_3017)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam modulation_output_15__I_0_336_i56_3_lut.init = 16'hcaca;
    LUT4 i10925_3_lut (.A(modulation_output[2]), .B(modulation_output[1]), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[0]), .Z(n29)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(85[80:131])
    defparam i10925_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_336_i48_3_lut (.A(n17), .B(n19), .C(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .Z(n48_adj_3010)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam modulation_output_15__I_0_336_i48_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_336_i52_3_lut (.A(n21), .B(n23), .C(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .Z(n52_adj_3016)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam modulation_output_15__I_0_336_i52_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_336_i21_3_lut (.A(modulation_output[10]), 
         .B(modulation_output[9]), .C(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .Z(n21)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam modulation_output_15__I_0_336_i21_3_lut.init = 16'hcaca;
    LUT4 i10923_3_lut (.A(modulation_output[8]), .B(modulation_output[7]), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[0]), .Z(n23)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(85[80:131])
    defparam i10923_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_336_i17_3_lut (.A(modulation_output[14]), 
         .B(modulation_output[13]), .C(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .Z(n17)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam modulation_output_15__I_0_336_i17_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_336_i19_3_lut (.A(modulation_output[12]), 
         .B(modulation_output[11]), .C(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .Z(n19)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam modulation_output_15__I_0_336_i19_3_lut.init = 16'hcaca;
    LUT4 i10926_3_lut (.A(modulation_output[6]), .B(modulation_output[5]), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[0]), .Z(n25)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(85[80:131])
    defparam i10926_3_lut.init = 16'hcaca;
    LUT4 i10931_3_lut (.A(modulation_output[4]), .B(modulation_output[3]), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[0]), .Z(n27)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(85[80:131])
    defparam i10931_3_lut.init = 16'hcaca;
    LUT4 i11076_4_lut (.A(n95_adj_3018), .B(n178_adj_3015), .C(n26365), 
         .D(modulation_deviation_amount_minus_sine_lookup_width[4]), .Z(n1[29])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam i11076_4_lut.init = 16'h3022;
    LUT4 i6554_4_lut (.A(modulation_output[15]), .B(modulation_output[14]), 
         .C(n26445), .D(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .Z(n95_adj_3018)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C (D)))) */ ;
    defparam i6554_4_lut.init = 16'hcaaa;
    LUT4 modulation_output_15__I_0_336_i80_3_lut (.A(n49_adj_3019), .B(n53_adj_3020), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[2]), .Z(n80)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam modulation_output_15__I_0_336_i80_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_336_i88_4_lut (.A(n57_adj_3021), .B(n30), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[2]), .D(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .Z(n88)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam modulation_output_15__I_0_336_i88_4_lut.init = 16'h0aca;
    LUT4 modulation_output_15__I_0_336_i49_3_lut (.A(n18), .B(n20), .C(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .Z(n49_adj_3019)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam modulation_output_15__I_0_336_i49_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_336_i53_3_lut (.A(n22), .B(n24), .C(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .Z(n53_adj_3020)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam modulation_output_15__I_0_336_i53_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_336_i22_3_lut (.A(modulation_output[9]), 
         .B(modulation_output[8]), .C(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .Z(n22)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam modulation_output_15__I_0_336_i22_3_lut.init = 16'hcaca;
    LUT4 i10928_3_lut (.A(modulation_output[7]), .B(modulation_output[6]), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[0]), .Z(n24)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(85[80:131])
    defparam i10928_3_lut.init = 16'hcaca;
    LUT4 i19507_3_lut (.A(\addr_space[0] [14]), .B(\addr_space[1] [14]), 
         .C(\wb_addr[0] ), .Z(n21827)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19507_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_336_i18_3_lut (.A(modulation_output[13]), 
         .B(modulation_output[12]), .C(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .Z(n18)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam modulation_output_15__I_0_336_i18_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_336_i20_3_lut (.A(modulation_output[11]), 
         .B(modulation_output[10]), .C(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .Z(n20)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam modulation_output_15__I_0_336_i20_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_336_i57_3_lut (.A(n26), .B(n28), .C(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .Z(n57_adj_3021)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam modulation_output_15__I_0_336_i57_3_lut.init = 16'hcaca;
    LUT4 i10927_3_lut (.A(modulation_output[1]), .B(modulation_output[0]), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[0]), .Z(n30)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(85[80:131])
    defparam i10927_3_lut.init = 16'hcaca;
    LUT4 i10929_3_lut (.A(modulation_output[5]), .B(modulation_output[4]), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[0]), .Z(n26)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(85[80:131])
    defparam i10929_3_lut.init = 16'hcaca;
    LUT4 i10930_3_lut (.A(modulation_output[3]), .B(modulation_output[2]), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[0]), .Z(n28)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(85[80:131])
    defparam i10930_3_lut.init = 16'hcaca;
    LUT4 i11077_4_lut (.A(n96), .B(n178_adj_3015), .C(n26364), .D(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .Z(n1[28])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam i11077_4_lut.init = 16'h3022;
    LUT4 i6556_4_lut (.A(modulation_output[15]), .B(n17), .C(n26556), 
         .D(modulation_deviation_amount_minus_sine_lookup_width[3]), .Z(n96)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C (D)))) */ ;
    defparam i6556_4_lut.init = 16'hcaaa;
    LUT4 i19505_3_lut (.A(\addr_space[2] [15]), .B(\addr_space[3] [15]), 
         .C(\wb_addr[0] ), .Z(n21825)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19505_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_336_i81_3_lut (.A(n50_adj_3022), .B(n54_adj_3023), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[2]), .Z(n81)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam modulation_output_15__I_0_336_i81_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_336_i50_3_lut (.A(n19), .B(n21), .C(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .Z(n50_adj_3022)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam modulation_output_15__I_0_336_i50_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_336_i54_3_lut (.A(n23), .B(n25), .C(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .Z(n54_adj_3023)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam modulation_output_15__I_0_336_i54_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_336_i58_3_lut (.A(n27), .B(n29), .C(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .Z(n58)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam modulation_output_15__I_0_336_i58_3_lut.init = 16'hcaca;
    LUT4 i11078_4_lut (.A(n97), .B(n178_adj_3015), .C(n113), .D(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .Z(n1[27])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam i11078_4_lut.init = 16'h3022;
    LUT4 modulation_output_15__I_0_336_i47_3_lut (.A(n16), .B(n18), .C(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .Z(n47_adj_3008)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam modulation_output_15__I_0_336_i47_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_336_i16_3_lut (.A(modulation_output[15]), 
         .B(modulation_output[14]), .C(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .Z(n16)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam modulation_output_15__I_0_336_i16_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_336_i113_4_lut (.A(n82), .B(n59_adj_3007), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[3]), .D(modulation_deviation_amount_minus_sine_lookup_width[2]), 
         .Z(n113)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam modulation_output_15__I_0_336_i113_4_lut.init = 16'h0aca;
    LUT4 modulation_output_15__I_0_336_i82_3_lut (.A(n51_adj_3024), .B(n55_adj_3025), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[2]), .Z(n82)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam modulation_output_15__I_0_336_i82_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_336_i59_3_lut (.A(n28), .B(n30), .C(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .Z(n59_adj_3007)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam modulation_output_15__I_0_336_i59_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_336_i51_3_lut (.A(n20), .B(n22), .C(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .Z(n51_adj_3024)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam modulation_output_15__I_0_336_i51_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_336_i55_3_lut (.A(n24), .B(n26), .C(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .Z(n55_adj_3025)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam modulation_output_15__I_0_336_i55_3_lut.init = 16'hcaca;
    LUT4 i11079_4_lut (.A(n98), .B(n178_adj_3015), .C(n114), .D(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .Z(n1[26])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam i11079_4_lut.init = 16'h3022;
    LUT4 i19504_3_lut (.A(\addr_space[0] [15]), .B(\addr_space[1] [15]), 
         .C(\wb_addr[0] ), .Z(n21824)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19504_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_336_i114_4_lut (.A(n83), .B(n60_adj_3009), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[3]), .D(modulation_deviation_amount_minus_sine_lookup_width[2]), 
         .Z(n114)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam modulation_output_15__I_0_336_i114_4_lut.init = 16'h0aca;
    LUT4 modulation_output_15__I_0_336_i83_3_lut (.A(n52_adj_3016), .B(n56_adj_3017), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[2]), .Z(n83)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam modulation_output_15__I_0_336_i83_3_lut.init = 16'hcaca;
    LUT4 i11080_4_lut (.A(n99), .B(n178_adj_3015), .C(n115), .D(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .Z(n1[25])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam i11080_4_lut.init = 16'h3022;
    LUT4 modulation_output_15__I_0_336_i99_3_lut (.A(modulation_output[15]), 
         .B(n76), .C(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .Z(n99)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam modulation_output_15__I_0_336_i99_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_336_i76_3_lut (.A(n45_adj_3026), .B(n49_adj_3019), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[2]), .Z(n76)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam modulation_output_15__I_0_336_i76_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_336_i115_4_lut (.A(n84), .B(n30), .C(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .D(n26555), .Z(n115)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam modulation_output_15__I_0_336_i115_4_lut.init = 16'h0aca;
    LUT4 modulation_output_15__I_0_336_i84_3_lut (.A(n53_adj_3020), .B(n57_adj_3021), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[2]), .Z(n84)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam modulation_output_15__I_0_336_i84_3_lut.init = 16'hcaca;
    LUT4 i11081_4_lut (.A(n100), .B(n178_adj_3015), .C(n26363), .D(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .Z(n1[24])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam i11081_4_lut.init = 16'h3022;
    LUT4 modulation_output_15__I_0_336_i100_3_lut (.A(modulation_output[15]), 
         .B(n77), .C(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .Z(n100)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam modulation_output_15__I_0_336_i100_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_336_i77_3_lut (.A(n46_adj_3027), .B(n50_adj_3022), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[2]), .Z(n77)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam modulation_output_15__I_0_336_i77_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_336_i46_3_lut (.A(modulation_output[15]), 
         .B(n17), .C(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .Z(n46_adj_3027)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam modulation_output_15__I_0_336_i46_3_lut.init = 16'hcaca;
    LUT4 i19502_3_lut (.A(\addr_space[2] [16]), .B(\addr_space[3] [16]), 
         .C(\wb_addr[0] ), .Z(n21822)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19502_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_336_i85_3_lut (.A(n54_adj_3023), .B(n58), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[2]), .Z(n85)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam modulation_output_15__I_0_336_i85_3_lut.init = 16'hcaca;
    LUT4 i11082_2_lut (.A(n132), .B(n178_adj_3015), .Z(n1[23])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam i11082_2_lut.init = 16'h2222;
    LUT4 i11084_2_lut (.A(n133), .B(n178_adj_3015), .Z(n1[22])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam i11084_2_lut.init = 16'h2222;
    LUT4 i11085_2_lut (.A(n134), .B(n178_adj_3015), .Z(n1[21])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam i11085_2_lut.init = 16'h2222;
    LUT4 i11086_2_lut (.A(n135), .B(n178_adj_3015), .Z(n1[20])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam i11086_2_lut.init = 16'h2222;
    LUT4 i11087_2_lut (.A(n136), .B(n178_adj_3015), .Z(n1[19])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam i11087_2_lut.init = 16'h2222;
    LUT4 i19501_3_lut (.A(\addr_space[0] [16]), .B(\addr_space[1] [16]), 
         .C(\wb_addr[0] ), .Z(n21821)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19501_3_lut.init = 16'hcaca;
    LUT4 i11088_2_lut (.A(n137), .B(n178_adj_3015), .Z(n1[18])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam i11088_2_lut.init = 16'h2222;
    LUT4 i11089_4_lut (.A(n107), .B(n178_adj_3015), .C(n123), .D(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .Z(n1[17])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam i11089_4_lut.init = 16'h3022;
    LUT4 i19493_3_lut (.A(\addr_space[2] [17]), .B(\addr_space[3] [17]), 
         .C(\wb_addr[0] ), .Z(n21813)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19493_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_336_i107_3_lut (.A(n76), .B(n84), .C(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .Z(n107)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam modulation_output_15__I_0_336_i107_3_lut.init = 16'hcaca;
    LUT4 i11090_4_lut (.A(n108), .B(n178_adj_3015), .C(n26355), .D(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .Z(n1[16])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam i11090_4_lut.init = 16'h3022;
    LUT4 modulation_output_15__I_0_336_i108_3_lut (.A(n77), .B(n85), .C(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .Z(n108)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam modulation_output_15__I_0_336_i108_3_lut.init = 16'hcaca;
    LUT4 i19492_3_lut (.A(\addr_space[0] [17]), .B(\addr_space[1] [17]), 
         .C(\wb_addr[0] ), .Z(n21812)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19492_3_lut.init = 16'hcaca;
    LUT4 i11882_4_lut (.A(n78), .B(n26380), .C(n26398), .D(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .Z(n1[15])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam i11882_4_lut.init = 16'h3022;
    LUT4 modulation_output_15__I_0_336_i78_3_lut (.A(n47_adj_3008), .B(n51_adj_3024), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[2]), .Z(n78)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam modulation_output_15__I_0_336_i78_3_lut.init = 16'hcaca;
    LUT4 i19484_3_lut (.A(\addr_space[2] [18]), .B(\addr_space[3] [18]), 
         .C(\wb_addr[0] ), .Z(n21804)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19484_3_lut.init = 16'hcaca;
    PFUMX i22702 (.BLUT(n24273), .ALUT(n38_adj_3003), .C0(sine_lookup_width_minus_modulation_deviation_amount[2]), 
          .Z(n24274));
    LUT4 i19483_3_lut (.A(\addr_space[0] [18]), .B(\addr_space[1] [18]), 
         .C(\wb_addr[0] ), .Z(n21803)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19483_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_336_i86_3_lut_rep_438 (.A(n55_adj_3025), 
         .B(n59_adj_3007), .C(modulation_deviation_amount_minus_sine_lookup_width[2]), 
         .Z(n26398)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam modulation_output_15__I_0_336_i86_3_lut_rep_438.init = 16'hcaca;
    LUT4 i19475_3_lut (.A(\addr_space[2] [19]), .B(\addr_space[3] [19]), 
         .C(\wb_addr[0] ), .Z(n21795)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19475_3_lut.init = 16'hcaca;
    LUT4 i19474_3_lut (.A(\addr_space[0] [19]), .B(\addr_space[1] [19]), 
         .C(\wb_addr[0] ), .Z(n21794)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19474_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_336_i87_3_lut_rep_439 (.A(n56_adj_3017), 
         .B(n60_adj_3009), .C(modulation_deviation_amount_minus_sine_lookup_width[2]), 
         .Z(n26399)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam modulation_output_15__I_0_336_i87_3_lut_rep_439.init = 16'hcaca;
    LUT4 i19466_3_lut (.A(\addr_space[2] [20]), .B(\addr_space[3] [20]), 
         .C(\wb_addr[0] ), .Z(n21786)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19466_3_lut.init = 16'hcaca;
    LUT4 i19465_3_lut (.A(\addr_space[0] [20]), .B(\addr_space[1] [20]), 
         .C(\wb_addr[0] ), .Z(n21785)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19465_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_rep_440 (.A(sine_lookup_width_minus_modulation_deviation_amount[3]), 
         .B(n178), .C(sine_lookup_width_minus_modulation_deviation_amount[4]), 
         .Z(n26400)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam i1_3_lut_rep_440.init = 16'hfefe;
    LUT4 i19457_3_lut (.A(\addr_space[2] [21]), .B(\addr_space[3] [21]), 
         .C(\wb_addr[0] ), .Z(n21777)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19457_3_lut.init = 16'hcaca;
    LUT4 i19456_3_lut (.A(\addr_space[0] [21]), .B(\addr_space[1] [21]), 
         .C(\wb_addr[0] ), .Z(n21776)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19456_3_lut.init = 16'hcaca;
    LUT4 i19451_3_lut (.A(\addr_space[2] [22]), .B(\addr_space[3] [22]), 
         .C(\wb_addr[0] ), .Z(n21771)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19451_3_lut.init = 16'hcaca;
    LUT4 i19450_3_lut (.A(\addr_space[0] [22]), .B(\addr_space[1] [22]), 
         .C(\wb_addr[0] ), .Z(n21770)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19450_3_lut.init = 16'hcaca;
    LUT4 i19442_3_lut (.A(\addr_space[2] [23]), .B(\addr_space[3] [23]), 
         .C(\wb_addr[0] ), .Z(n21762)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19442_3_lut.init = 16'hcaca;
    LUT4 i19441_3_lut (.A(\addr_space[0] [23]), .B(\addr_space[1] [23]), 
         .C(\wb_addr[0] ), .Z(n21761)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19441_3_lut.init = 16'hcaca;
    LUT4 i19439_3_lut (.A(\addr_space[2] [24]), .B(\addr_space[3] [24]), 
         .C(\wb_addr[0] ), .Z(n21759)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19439_3_lut.init = 16'hcaca;
    LUT4 i19438_3_lut (.A(\addr_space[0] [24]), .B(\addr_space[1] [24]), 
         .C(\wb_addr[0] ), .Z(n21758)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19438_3_lut.init = 16'hcaca;
    LUT4 i22471_2_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[3]), .Z(n21926)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam i22471_2_lut.init = 16'heeee;
    LUT4 n38_bdd_3_lut_23493 (.A(n13449), .B(n13451), .C(sine_lookup_width_minus_modulation_deviation_amount[1]), 
         .Z(n24273)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n38_bdd_3_lut_23493.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[2]), 
         .B(n26425), .C(n26380), .D(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .Z(n1[0])) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0004;
    LUT4 i10914_3_lut_rep_403_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[2]), 
         .B(n26425), .C(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .D(n85), .Z(n26363)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam i10914_3_lut_rep_403_4_lut.init = 16'h4f40;
    LUT4 n24274_bdd_3_lut (.A(n24274), .B(n73), .C(sine_lookup_width_minus_modulation_deviation_amount[3]), 
         .Z(n24275)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n24274_bdd_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_420 (.A(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .B(n178_adj_3015), .Z(n26380)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam i1_2_lut_rep_420.init = 16'heeee;
    LUT4 i11888_2_lut_3_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .B(n178_adj_3015), .C(n88), .D(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .Z(n1[5])) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam i11888_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 i11881_2_lut_3_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .B(n178_adj_3015), .C(n26398), .D(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .Z(n1[7])) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam i11881_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 i11909_2_lut_3_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .B(n178_adj_3015), .C(n60_adj_3009), .D(n26553), .Z(n1[2])) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam i11909_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 i11883_2_lut_3_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .B(n178_adj_3015), .C(n26399), .D(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .Z(n1[6])) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam i11883_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 i11666_2_lut_3_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .B(n178_adj_3015), .C(n59_adj_3007), .D(n26553), .Z(n1[3])) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam i11666_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 i11664_2_lut_3_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .B(n178_adj_3015), .C(n89), .D(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .Z(n1[4])) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam i11664_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 i11877_2_lut_3_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .B(n178_adj_3015), .C(n113), .Z(n1[11])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam i11877_2_lut_3_lut.init = 16'h1010;
    LUT4 n39_bdd_3_lut_25269 (.A(n13457), .B(n6), .C(sine_lookup_width_minus_modulation_deviation_amount[1]), 
         .Z(n26267)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n39_bdd_3_lut_25269.init = 16'hcaca;
    LUT4 n39_bdd_3_lut_24417 (.A(n43_adj_3011), .B(modulation_output[15]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[2]), .Z(n26266)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n39_bdd_3_lut_24417.init = 16'hcaca;
    LUT4 i11876_2_lut_3_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .B(n178_adj_3015), .C(n114), .Z(n1[10])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam i11876_2_lut_3_lut.init = 16'h1010;
    PFUMX i19440 (.BLUT(n21758), .ALUT(n21759), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[24]));
    LUT4 i11875_2_lut_3_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .B(n178_adj_3015), .C(n115), .Z(n1[9])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam i11875_2_lut_3_lut.init = 16'h1010;
    PFUMX i19443 (.BLUT(n21761), .ALUT(n21762), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[23]));
    LUT4 n26268_bdd_3_lut (.A(n26268), .B(n26266), .C(sine_lookup_width_minus_modulation_deviation_amount[3]), 
         .Z(n26269)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n26268_bdd_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .B(n178_adj_3015), .C(n123), .Z(n20073)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam i1_2_lut_3_lut.init = 16'h1010;
    LUT4 n36_bdd_3_lut_24629 (.A(n36_adj_2995), .B(n40_adj_2996), .C(sine_lookup_width_minus_modulation_deviation_amount[2]), 
         .Z(n26313)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n36_bdd_3_lut_24629.init = 16'hcaca;
    LUT4 n36_bdd_3_lut_24458 (.A(n44_adj_2997), .B(modulation_output[15]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[2]), .Z(n26312)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n36_bdd_3_lut_24458.init = 16'hcaca;
    LUT4 n37_bdd_3_lut_24632 (.A(n37_adj_2998), .B(n41_adj_3000), .C(sine_lookup_width_minus_modulation_deviation_amount[2]), 
         .Z(n26319)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n37_bdd_3_lut_24632.init = 16'hcaca;
    LUT4 n37_bdd_4_lut (.A(n14), .B(modulation_output[15]), .C(sine_lookup_width_minus_modulation_deviation_amount[2]), 
         .D(sine_lookup_width_minus_modulation_deviation_amount[1]), .Z(n26318)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;
    defparam n37_bdd_4_lut.init = 16'hccca;
    LUT4 n38_bdd_3_lut_24648 (.A(n38_adj_3003), .B(n42_adj_3004), .C(sine_lookup_width_minus_modulation_deviation_amount[2]), 
         .Z(n26325)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n38_bdd_3_lut_24648.init = 16'hcaca;
    LUT4 n38_bdd_4_lut (.A(modulation_output[14]), .B(modulation_output[15]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[2]), .D(n26615), 
         .Z(n26324)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;
    defparam n38_bdd_4_lut.init = 16'hccca;
    PFUMX i19452 (.BLUT(n21770), .ALUT(n21771), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[22]));
    PFUMX i19458 (.BLUT(n21776), .ALUT(n21777), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[21]));
    PFUMX i19467 (.BLUT(n21785), .ALUT(n21786), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[20]));
    PFUMX i19476 (.BLUT(n21794), .ALUT(n21795), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[19]));
    PFUMX i19485 (.BLUT(n21803), .ALUT(n21804), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[18]));
    PFUMX i19494 (.BLUT(n21812), .ALUT(n21813), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[17]));
    PFUMX i19503 (.BLUT(n21821), .ALUT(n21822), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[16]));
    LUT4 i11054_2_lut_4_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[2]), .C(n59_adj_3007), 
         .D(n55_adj_3025), .Z(n117)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam i11054_2_lut_4_lut_4_lut.init = 16'h5140;
    LUT4 modulation_output_15__I_0_336_i104_4_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[4]), .C(n89), 
         .D(n81), .Z(n104)) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C)+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam modulation_output_15__I_0_336_i104_4_lut_4_lut.init = 16'h7340;
    PFUMX i19506 (.BLUT(n21824), .ALUT(n21825), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[15]));
    LUT4 i11055_2_lut_4_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[2]), .C(n60_adj_3009), 
         .D(n56_adj_3017), .Z(n118)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam i11055_2_lut_4_lut_4_lut.init = 16'h5140;
    LUT4 modulation_output_15__I_0_336_i103_4_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[4]), .C(n88), 
         .D(n80), .Z(n103)) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C)+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam modulation_output_15__I_0_336_i103_4_lut_4_lut.init = 16'h7340;
    PFUMX i19509 (.BLUT(n21827), .ALUT(n21828), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[14]));
    LUT4 smpl_register_16__bdd_4_lut_4_lut (.A(\wb_addr[0] ), .B(\wb_addr[1] ), 
         .C(n2), .D(\smpl_register[16] ), .Z(n26331)) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(45[4:25])
    defparam smpl_register_16__bdd_4_lut_4_lut.init = 16'hf3d1;
    PFUMX i19512 (.BLUT(n21830), .ALUT(n21831), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[13]));
    LUT4 smpl_register_10__bdd_4_lut_4_lut (.A(\wb_addr[0] ), .B(\wb_addr[1] ), 
         .C(n2_adj_1), .D(\smpl_register[10] ), .Z(n26342)) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(45[4:25])
    defparam smpl_register_10__bdd_4_lut_4_lut.init = 16'hf3d1;
    LUT4 smpl_register_9__bdd_4_lut_4_lut (.A(\wb_addr[0] ), .B(\wb_addr[1] ), 
         .C(n2_adj_2), .D(\smpl_register[9] ), .Z(n26341)) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(45[4:25])
    defparam smpl_register_9__bdd_4_lut_4_lut.init = 16'hf3d1;
    PFUMX i19515 (.BLUT(n21833), .ALUT(n21834), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[12]));
    LUT4 smpl_register_29__bdd_4_lut_4_lut (.A(\wb_addr[0] ), .B(\wb_addr[1] ), 
         .C(n2_adj_3), .D(\smpl_register[29] ), .Z(n26339)) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(45[4:25])
    defparam smpl_register_29__bdd_4_lut_4_lut.init = 16'hf3d1;
    LUT4 smpl_register_20__bdd_4_lut_4_lut (.A(\wb_addr[0] ), .B(\wb_addr[1] ), 
         .C(n2_adj_4), .D(\smpl_register[20] ), .Z(n26337)) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(45[4:25])
    defparam smpl_register_20__bdd_4_lut_4_lut.init = 16'hf3d1;
    LUT4 smpl_register_5__bdd_4_lut_4_lut (.A(\wb_addr[0] ), .B(\wb_addr[1] ), 
         .C(n2_adj_5), .D(\smpl_register[5] ), .Z(n26336)) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(45[4:25])
    defparam smpl_register_5__bdd_4_lut_4_lut.init = 16'hf3d1;
    LUT4 i22507_2_lut_rep_593 (.A(modulation_deviation_amount_minus_sine_lookup_width[2]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[3]), .Z(n26553)) /* synthesis lut_function=(!(A+(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam i22507_2_lut_rep_593.init = 16'h1111;
    LUT4 i6549_2_lut_rep_595 (.A(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[2]), .Z(n26555)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam i6549_2_lut_rep_595.init = 16'heeee;
    LUT4 i11917_3_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[2]), .C(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .D(n30), .Z(n123)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam i11917_3_lut_4_lut.init = 16'h0100;
    LUT4 i6558_3_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[2]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[3]), .C(n47_adj_3008), 
         .D(modulation_output[15]), .Z(n97)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam i6558_3_lut_4_lut.init = 16'hf780;
    LUT4 i6560_3_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[2]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[3]), .C(n48_adj_3010), 
         .D(modulation_output[15]), .Z(n98)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam i6560_3_lut_4_lut.init = 16'hf780;
    LUT4 i6547_2_lut_rep_596 (.A(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[2]), .Z(n26556)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam i6547_2_lut_rep_596.init = 16'h8888;
    LUT4 i6548_3_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[2]), .C(n17), 
         .D(modulation_output[15]), .Z(n73_adj_3006)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam i6548_3_lut_4_lut.init = 16'hf780;
    LUT4 i6539_2_lut_rep_598 (.A(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[1]), .Z(n26558)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam i6539_2_lut_rep_598.init = 16'h8888;
    LUT4 i6545_2_lut_rep_485_3_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[1]), .C(modulation_deviation_amount_minus_sine_lookup_width[2]), 
         .Z(n26445)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam i6545_2_lut_rep_485_3_lut.init = 16'h8080;
    LUT4 i6540_3_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[1]), .C(modulation_output[14]), 
         .D(modulation_output[15]), .Z(n45_adj_3026)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam i6540_3_lut_4_lut.init = 16'hf780;
    LUT4 smpl_register_18__bdd_4_lut_4_lut (.A(\wb_addr[0] ), .B(\wb_addr[1] ), 
         .C(n2_adj_6), .D(\smpl_register[18] ), .Z(n26333)) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(45[4:25])
    defparam smpl_register_18__bdd_4_lut_4_lut.init = 16'hf3d1;
    PFUMX i19518 (.BLUT(n21836), .ALUT(n21837), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[11]));
    LUT4 smpl_register_17__bdd_4_lut_4_lut (.A(\wb_addr[0] ), .B(\wb_addr[1] ), 
         .C(n2_adj_7), .D(\smpl_register[17] ), .Z(n26332)) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(45[4:25])
    defparam smpl_register_17__bdd_4_lut_4_lut.init = 16'hf3d1;
    LUT4 i11539_2_lut (.A(o_sample_i[12]), .B(o_dac_cw_b_c_c), .Z(o_dac_a_c_5)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(29[18:124])
    defparam i11539_2_lut.init = 16'heeee;
    LUT4 i791_1_lut (.A(o_dac_b_c_15), .Z(o_dac_b_c_9)) /* synthesis lut_function=(!(A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(28[31:66])
    defparam i791_1_lut.init = 16'h5555;
    PFUMX i19521 (.BLUT(n21839), .ALUT(n21840), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[10]));
    PFUMX i19524 (.BLUT(n21842), .ALUT(n21843), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[9]));
    PFUMX i19527 (.BLUT(n21845), .ALUT(n21846), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[8]));
    LUT4 i19436_3_lut (.A(\addr_space[2] [25]), .B(\addr_space[3] [25]), 
         .C(\wb_addr[0] ), .Z(n21756)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19436_3_lut.init = 16'hcaca;
    LUT4 i19435_3_lut (.A(\addr_space[0] [25]), .B(\addr_space[1] [25]), 
         .C(\wb_addr[0] ), .Z(n21755)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19435_3_lut.init = 16'hcaca;
    LUT4 i19433_3_lut (.A(\addr_space[2] [26]), .B(\addr_space[3] [26]), 
         .C(\wb_addr[0] ), .Z(n21753)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19433_3_lut.init = 16'hcaca;
    PFUMX i19530 (.BLUT(n21848), .ALUT(n21849), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[7]));
    PFUMX i19533 (.BLUT(n21851), .ALUT(n21852), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[6]));
    LUT4 i19432_3_lut (.A(\addr_space[0] [26]), .B(\addr_space[1] [26]), 
         .C(\wb_addr[0] ), .Z(n21752)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19432_3_lut.init = 16'hcaca;
    LUT4 i12208_2_lut_rep_683 (.A(o_sample_i[15]), .B(o_dac_cw_b_c_c), .Z(n26643)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i12208_2_lut_rep_683.init = 16'heeee;
    LUT4 i12209_1_lut_2_lut (.A(o_sample_i[15]), .B(o_dac_cw_b_c_c), .Z(o_dac_a_c_9)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i12209_1_lut_2_lut.init = 16'h1111;
    PFUMX i19536 (.BLUT(n21854), .ALUT(n21855), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[5]));
    LUT4 i19430_3_lut (.A(\addr_space[2] [27]), .B(\addr_space[3] [27]), 
         .C(\wb_addr[0] ), .Z(n21750)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19430_3_lut.init = 16'hcaca;
    PFUMX i19539 (.BLUT(n21857), .ALUT(n21858), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[4]));
    LUT4 i19429_3_lut (.A(\addr_space[0] [27]), .B(\addr_space[1] [27]), 
         .C(\wb_addr[0] ), .Z(n21749)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19429_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_100 (.A(n20296), .B(n20112), .C(n20302), .D(n20298), 
         .Z(n178_adj_3015)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam i1_4_lut_adj_100.init = 16'hfffe;
    PFUMX modulation_output_15__I_0_336_i137 (.BLUT(n75), .ALUT(n106), .C0(n21926), 
          .Z(n137)) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;
    PFUMX modulation_output_15__I_0_336_i136 (.BLUT(n74), .ALUT(n105), .C0(n21926), 
          .Z(n136)) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;
    PFUMX modulation_output_15__I_0_336_i133 (.BLUT(n102), .ALUT(n118), 
          .C0(modulation_deviation_amount_minus_sine_lookup_width[4]), .Z(n133)) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;
    PFUMX modulation_output_15__I_0_336_i132 (.BLUT(n101), .ALUT(n117), 
          .C0(modulation_deviation_amount_minus_sine_lookup_width[4]), .Z(n132)) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=120, LSE_RLINE=132 */ ;
    LUT4 i19427_3_lut (.A(\addr_space[2] [28]), .B(\addr_space[3] [28]), 
         .C(\wb_addr[0] ), .Z(n21747)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19427_3_lut.init = 16'hcaca;
    PFUMX i18681 (.BLUT(n20999), .ALUT(n21000), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[3]));
    LUT4 i1_2_lut_adj_101 (.A(modulation_deviation_amount_minus_sine_lookup_width[7]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[8]), .Z(n20296)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam i1_2_lut_adj_101.init = 16'heeee;
    LUT4 i1_4_lut_adj_102 (.A(modulation_deviation_amount_minus_sine_lookup_width[5]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[13]), .C(modulation_deviation_amount_minus_sine_lookup_width[15]), 
         .D(modulation_deviation_amount_minus_sine_lookup_width[10]), .Z(n20112)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam i1_4_lut_adj_102.init = 16'hfffe;
    LUT4 i19426_3_lut (.A(\addr_space[0] [28]), .B(\addr_space[1] [28]), 
         .C(\wb_addr[0] ), .Z(n21746)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19426_3_lut.init = 16'hcaca;
    PFUMX i18684 (.BLUT(n21002), .ALUT(n21003), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[2]));
    LUT4 i19424_3_lut (.A(\addr_space[2] [29]), .B(\addr_space[3] [29]), 
         .C(\wb_addr[0] ), .Z(n21744)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19424_3_lut.init = 16'hcaca;
    PFUMX i18687 (.BLUT(n21005), .ALUT(n21006), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[1]));
    LUT4 i1_4_lut_adj_103 (.A(modulation_deviation_amount_minus_sine_lookup_width[6]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[9]), .C(modulation_deviation_amount_minus_sine_lookup_width[11]), 
         .D(modulation_deviation_amount_minus_sine_lookup_width[14]), .Z(n20302)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam i1_4_lut_adj_103.init = 16'hfffe;
    PFUMX i19416 (.BLUT(n21734), .ALUT(n21735), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[0]));
    LUT4 i6630_2_lut_rep_449 (.A(sine_lookup_width_minus_modulation_deviation_amount[4]), 
         .B(n178), .Z(n26409)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam i6630_2_lut_rep_449.init = 16'heeee;
    LUT4 i19423_3_lut (.A(\addr_space[0] [29]), .B(\addr_space[1] [29]), 
         .C(\wb_addr[0] ), .Z(n21743)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19423_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_573 (.A(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .B(modulation_output[0]), .Z(n26533)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam i1_2_lut_rep_573.init = 16'h4444;
    LUT4 n26269_bdd_3_lut_4_lut (.A(sine_lookup_width_minus_modulation_deviation_amount[4]), 
         .B(n178), .C(modulation_output[15]), .D(n26269), .Z(carrier_center_increment_offset_rs_30__N_1560[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam n26269_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n26320_bdd_3_lut_4_lut (.A(sine_lookup_width_minus_modulation_deviation_amount[4]), 
         .B(n178), .C(modulation_output[15]), .D(n26320), .Z(carrier_center_increment_offset_rs_30__N_1560[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam n26320_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_rep_465_3_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .B(modulation_output[0]), .C(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .Z(n26425)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam i1_2_lut_rep_465_3_lut.init = 16'h0404;
    LUT4 i6587_2_lut_rep_655 (.A(sine_lookup_width_minus_modulation_deviation_amount[0]), 
         .B(sine_lookup_width_minus_modulation_deviation_amount[1]), .Z(n26615)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam i6587_2_lut_rep_655.init = 16'heeee;
    LUT4 i1_2_lut_rep_419_3_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .B(modulation_output[0]), .C(modulation_deviation_amount_minus_sine_lookup_width[2]), 
         .D(modulation_deviation_amount_minus_sine_lookup_width[1]), .Z(n26379)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam i1_2_lut_rep_419_3_lut_4_lut.init = 16'h0004;
    LUT4 n26314_bdd_3_lut_4_lut (.A(sine_lookup_width_minus_modulation_deviation_amount[4]), 
         .B(n178), .C(modulation_output[15]), .D(n26314), .Z(carrier_center_increment_offset_rs_30__N_1560[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam n26314_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i6591_2_lut_3_lut (.A(sine_lookup_width_minus_modulation_deviation_amount[0]), 
         .B(sine_lookup_width_minus_modulation_deviation_amount[1]), .C(sine_lookup_width_minus_modulation_deviation_amount[2]), 
         .Z(n8972)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam i6591_2_lut_3_lut.init = 16'hfefe;
    LUT4 i6588_3_lut_4_lut (.A(sine_lookup_width_minus_modulation_deviation_amount[0]), 
         .B(sine_lookup_width_minus_modulation_deviation_amount[1]), .C(modulation_output[15]), 
         .D(modulation_output[14]), .Z(n46_adj_3005)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam i6588_3_lut_4_lut.init = 16'hf1e0;
    LUT4 modulation_output_15__I_0_336_i60_3_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .B(modulation_output[0]), .C(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .D(n29), .Z(n60_adj_3009)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(95[11] 105[5])
    defparam modulation_output_15__I_0_336_i60_3_lut_4_lut.init = 16'h4f40;
    LUT4 i22487_4_lut (.A(n20438), .B(n26557), .C(n38), .D(\wb_addr[15] ), 
         .Z(dac_clk_p_c_enable_114)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(44[3] 46[6])
    defparam i22487_4_lut.init = 16'h0400;
    LUT4 i19421_3_lut (.A(\addr_space[2] [30]), .B(\addr_space[3] [30]), 
         .C(\wb_addr[0] ), .Z(n21741)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19421_3_lut.init = 16'hcaca;
    LUT4 n26326_bdd_3_lut_4_lut (.A(sine_lookup_width_minus_modulation_deviation_amount[4]), 
         .B(n178), .C(modulation_output[15]), .D(n26326), .Z(carrier_center_increment_offset_rs_30__N_1560[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam n26326_bdd_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i19419 (.BLUT(n21737), .ALUT(n21738), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[31]));
    LUT4 n24275_bdd_3_lut_4_lut (.A(sine_lookup_width_minus_modulation_deviation_amount[4]), 
         .B(n178), .C(modulation_output[15]), .D(n24275), .Z(carrier_center_increment_offset_rs_30__N_1560[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam n24275_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 modulation_output_15__I_0_i94_3_lut_4_lut (.A(sine_lookup_width_minus_modulation_deviation_amount[4]), 
         .B(n178), .C(modulation_output[15]), .D(n13448), .Z(n94)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_i94_3_lut_4_lut.init = 16'hf1e0;
    LUT4 modulation_output_15__I_0_i95_3_lut_4_lut (.A(sine_lookup_width_minus_modulation_deviation_amount[4]), 
         .B(n178), .C(modulation_output[15]), .D(n13456), .Z(n95)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_i95_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i1_2_lut_adj_104 (.A(modulation_deviation_amount_minus_sine_lookup_width[12]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[16]), .Z(n20298)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(98[41:116])
    defparam i1_2_lut_adj_104.init = 16'heeee;
    LUT4 modulation_output_15__I_0_i64_3_lut (.A(n33_adj_2999), .B(n72_adj_3002), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[3]), .Z(n64)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(99[41:116])
    defparam modulation_output_15__I_0_i64_3_lut.init = 16'hcaca;
    LUT4 i22480_4_lut (.A(n20864), .B(n20416), .C(n20402), .D(n38), 
         .Z(dac_clk_p_c_enable_71)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(44[3] 46[6])
    defparam i22480_4_lut.init = 16'h0002;
    LUT4 i22478_4_lut (.A(n26557), .B(n20422), .C(n38), .D(\wb_addr[1] ), 
         .Z(dac_clk_p_c_enable_103)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(44[3] 46[6])
    defparam i22478_4_lut.init = 16'h0200;
    LUT4 i10913_3_lut (.A(n13450), .B(n71), .C(sine_lookup_width_minus_modulation_deviation_amount[3]), 
         .Z(n63)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(85[27:78])
    defparam i10913_3_lut.init = 16'hcaca;
    dds modulation (.dac_clk_p_c(dac_clk_p_c), .n26683(n26683), .\addr_space[1][0] (\addr_space[1] [0]), 
        .\addr_space[1][30] (\addr_space[1] [30]), .\addr_space[1][29] (\addr_space[1] [29]), 
        .\addr_space[1][28] (\addr_space[1] [28]), .\addr_space[1][27] (\addr_space[1] [27]), 
        .\addr_space[1][26] (\addr_space[1] [26]), .\addr_space[1][25] (\addr_space[1] [25]), 
        .\addr_space[1][24] (\addr_space[1] [24]), .\addr_space[1][23] (\addr_space[1] [23]), 
        .\addr_space[1][22] (\addr_space[1] [22]), .\addr_space[1][21] (\addr_space[1] [21]), 
        .\addr_space[1][20] (\addr_space[1] [20]), .\addr_space[1][19] (\addr_space[1] [19]), 
        .\addr_space[1][18] (\addr_space[1] [18]), .\addr_space[1][17] (\addr_space[1] [17]), 
        .\addr_space[1][16] (\addr_space[1] [16]), .\addr_space[1][15] (\addr_space[1] [15]), 
        .\addr_space[1][14] (\addr_space[1] [14]), .\addr_space[1][13] (\addr_space[1] [13]), 
        .\addr_space[1][12] (\addr_space[1] [12]), .\addr_space[1][11] (\addr_space[1] [11]), 
        .\addr_space[1][10] (\addr_space[1] [10]), .\addr_space[1][9] (\addr_space[1] [9]), 
        .\addr_space[1][8] (\addr_space[1] [8]), .\addr_space[1][7] (\addr_space[1] [7]), 
        .\addr_space[1][6] (\addr_space[1] [6]), .\addr_space[1][5] (\addr_space[1] [5]), 
        .\addr_space[1][4] (\addr_space[1] [4]), .\addr_space[1][3] (\addr_space[1] [3]), 
        .\addr_space[1][2] (\addr_space[1] [2]), .\addr_space[1][1] (\addr_space[1] [1]), 
        .modulation_output({modulation_output}), .o_dac_cw_b_c_c(o_dac_cw_b_c_c), 
        .\quarter_wave_sample_register_q[15] (quarter_wave_sample_register_q[15]), 
        .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(83[4:161])
    dds_U2 carrier (.dac_clk_p_c(dac_clk_p_c), .n26683(n26683), .carrier_increment({carrier_increment}), 
           .o_dac_cw_b_c_c(o_dac_cw_b_c_c), .o_dac_b_c_7(o_dac_b_c_7), .\o_sample_i[7] (\o_sample_i[7] ), 
           .\o_sample_i[15] (o_sample_i[15]), .\o_sample_i[14] (\o_sample_i[14] ), 
           .\o_sample_i[13] (\o_sample_i[13] ), .\o_sample_i[12] (o_sample_i[12]), 
           .\o_sample_i[11] (\o_sample_i[11] ), .\o_sample_i[10] (\o_sample_i[10] ), 
           .\o_sample_i[9] (\o_sample_i[9] ), .\o_sample_i[8] (\o_sample_i[8] ), 
           .\quarter_wave_sample_register_q[15] (quarter_wave_sample_register_q[15]), 
           .n29209(n29209), .o_dac_b_c_15(o_dac_b_c_15), .o_dac_b_c_14(o_dac_b_c_14), 
           .o_dac_b_c_13(o_dac_b_c_13), .o_dac_b_c_12(o_dac_b_c_12), .o_dac_b_c_11(o_dac_b_c_11), 
           .o_dac_b_c_10(o_dac_b_c_10), .n3537(n3537), .o_dac_b_c_8(o_dac_b_c_8), 
           .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(78[4:158])
    
endmodule
//
// Verilog Description of module dds
//

module dds (dac_clk_p_c, n26683, \addr_space[1][0] , \addr_space[1][30] , 
            \addr_space[1][29] , \addr_space[1][28] , \addr_space[1][27] , 
            \addr_space[1][26] , \addr_space[1][25] , \addr_space[1][24] , 
            \addr_space[1][23] , \addr_space[1][22] , \addr_space[1][21] , 
            \addr_space[1][20] , \addr_space[1][19] , \addr_space[1][18] , 
            \addr_space[1][17] , \addr_space[1][16] , \addr_space[1][15] , 
            \addr_space[1][14] , \addr_space[1][13] , \addr_space[1][12] , 
            \addr_space[1][11] , \addr_space[1][10] , \addr_space[1][9] , 
            \addr_space[1][8] , \addr_space[1][7] , \addr_space[1][6] , 
            \addr_space[1][5] , \addr_space[1][4] , \addr_space[1][3] , 
            \addr_space[1][2] , \addr_space[1][1] , modulation_output, 
            o_dac_cw_b_c_c, \quarter_wave_sample_register_q[15] , GND_net) /* synthesis syn_module_defined=1 */ ;
    input dac_clk_p_c;
    input n26683;
    input \addr_space[1][0] ;
    input \addr_space[1][30] ;
    input \addr_space[1][29] ;
    input \addr_space[1][28] ;
    input \addr_space[1][27] ;
    input \addr_space[1][26] ;
    input \addr_space[1][25] ;
    input \addr_space[1][24] ;
    input \addr_space[1][23] ;
    input \addr_space[1][22] ;
    input \addr_space[1][21] ;
    input \addr_space[1][20] ;
    input \addr_space[1][19] ;
    input \addr_space[1][18] ;
    input \addr_space[1][17] ;
    input \addr_space[1][16] ;
    input \addr_space[1][15] ;
    input \addr_space[1][14] ;
    input \addr_space[1][13] ;
    input \addr_space[1][12] ;
    input \addr_space[1][11] ;
    input \addr_space[1][10] ;
    input \addr_space[1][9] ;
    input \addr_space[1][8] ;
    input \addr_space[1][7] ;
    input \addr_space[1][6] ;
    input \addr_space[1][5] ;
    input \addr_space[1][4] ;
    input \addr_space[1][3] ;
    input \addr_space[1][2] ;
    input \addr_space[1][1] ;
    output [15:0]modulation_output;
    input o_dac_cw_b_c_c;
    input \quarter_wave_sample_register_q[15] ;
    input GND_net;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(29[49:58])
    wire [15:0]modulation_output_c /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(73[39:56])
    wire [30:0]increment;   // d:/documents/git_local/fm_modulator/rtl/dds.v(14[31:40])
    wire [11:0]o_phase;   // d:/documents/git_local/fm_modulator/rtl/dds.v(18[26:33])
    
    FD1S3DX increment_i0 (.D(\addr_space[1][0] ), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(increment[0])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=83, LSE_RLINE=83 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i0.GSR = "DISABLED";
    FD1S3DX increment_i30 (.D(\addr_space[1][30] ), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(increment[30])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=83, LSE_RLINE=83 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i30.GSR = "DISABLED";
    FD1S3DX increment_i29 (.D(\addr_space[1][29] ), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(increment[29])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=83, LSE_RLINE=83 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i29.GSR = "DISABLED";
    FD1S3DX increment_i28 (.D(\addr_space[1][28] ), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(increment[28])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=83, LSE_RLINE=83 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i28.GSR = "DISABLED";
    FD1S3DX increment_i27 (.D(\addr_space[1][27] ), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(increment[27])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=83, LSE_RLINE=83 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i27.GSR = "DISABLED";
    FD1S3DX increment_i26 (.D(\addr_space[1][26] ), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(increment[26])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=83, LSE_RLINE=83 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i26.GSR = "DISABLED";
    FD1S3DX increment_i25 (.D(\addr_space[1][25] ), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(increment[25])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=83, LSE_RLINE=83 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i25.GSR = "DISABLED";
    FD1S3DX increment_i24 (.D(\addr_space[1][24] ), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(increment[24])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=83, LSE_RLINE=83 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i24.GSR = "DISABLED";
    FD1S3DX increment_i23 (.D(\addr_space[1][23] ), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(increment[23])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=83, LSE_RLINE=83 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i23.GSR = "DISABLED";
    FD1S3DX increment_i22 (.D(\addr_space[1][22] ), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(increment[22])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=83, LSE_RLINE=83 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i22.GSR = "DISABLED";
    FD1S3DX increment_i21 (.D(\addr_space[1][21] ), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(increment[21])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=83, LSE_RLINE=83 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i21.GSR = "DISABLED";
    FD1S3DX increment_i20 (.D(\addr_space[1][20] ), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(increment[20])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=83, LSE_RLINE=83 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i20.GSR = "DISABLED";
    FD1S3DX increment_i19 (.D(\addr_space[1][19] ), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(increment[19])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=83, LSE_RLINE=83 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i19.GSR = "DISABLED";
    FD1S3DX increment_i18 (.D(\addr_space[1][18] ), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(increment[18])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=83, LSE_RLINE=83 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i18.GSR = "DISABLED";
    FD1S3DX increment_i17 (.D(\addr_space[1][17] ), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(increment[17])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=83, LSE_RLINE=83 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i17.GSR = "DISABLED";
    FD1S3DX increment_i16 (.D(\addr_space[1][16] ), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(increment[16])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=83, LSE_RLINE=83 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i16.GSR = "DISABLED";
    FD1S3DX increment_i15 (.D(\addr_space[1][15] ), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(increment[15])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=83, LSE_RLINE=83 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i15.GSR = "DISABLED";
    FD1S3DX increment_i14 (.D(\addr_space[1][14] ), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(increment[14])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=83, LSE_RLINE=83 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i14.GSR = "DISABLED";
    FD1S3DX increment_i13 (.D(\addr_space[1][13] ), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(increment[13])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=83, LSE_RLINE=83 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i13.GSR = "DISABLED";
    FD1S3DX increment_i12 (.D(\addr_space[1][12] ), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(increment[12])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=83, LSE_RLINE=83 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i12.GSR = "DISABLED";
    FD1S3DX increment_i11 (.D(\addr_space[1][11] ), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(increment[11])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=83, LSE_RLINE=83 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i11.GSR = "DISABLED";
    FD1S3DX increment_i10 (.D(\addr_space[1][10] ), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(increment[10])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=83, LSE_RLINE=83 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i10.GSR = "DISABLED";
    FD1S3DX increment_i9 (.D(\addr_space[1][9] ), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(increment[9])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=83, LSE_RLINE=83 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i9.GSR = "DISABLED";
    FD1S3DX increment_i8 (.D(\addr_space[1][8] ), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(increment[8])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=83, LSE_RLINE=83 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i8.GSR = "DISABLED";
    FD1S3DX increment_i7 (.D(\addr_space[1][7] ), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(increment[7])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=83, LSE_RLINE=83 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i7.GSR = "DISABLED";
    FD1S3DX increment_i6 (.D(\addr_space[1][6] ), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(increment[6])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=83, LSE_RLINE=83 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i6.GSR = "DISABLED";
    FD1S3DX increment_i5 (.D(\addr_space[1][5] ), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(increment[5])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=83, LSE_RLINE=83 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i5.GSR = "DISABLED";
    FD1S3DX increment_i4 (.D(\addr_space[1][4] ), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(increment[4])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=83, LSE_RLINE=83 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i4.GSR = "DISABLED";
    FD1S3DX increment_i3 (.D(\addr_space[1][3] ), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(increment[3])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=83, LSE_RLINE=83 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i3.GSR = "DISABLED";
    FD1S3DX increment_i2 (.D(\addr_space[1][2] ), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(increment[2])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=83, LSE_RLINE=83 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i2.GSR = "DISABLED";
    FD1S3DX increment_i1 (.D(\addr_space[1][1] ), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(increment[1])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=83, LSE_RLINE=83 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i1.GSR = "DISABLED";
    quarter_wave_sine_lookup qtr_inst (.dac_clk_p_c(dac_clk_p_c), .n26683(n26683), 
            .modulation_output({modulation_output}), .o_dac_cw_b_c_c(o_dac_cw_b_c_c), 
            .o_phase({o_phase}), .\quarter_wave_sample_register_q[15] (\quarter_wave_sample_register_q[15] ), 
            .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(21[70:134])
    \nco(OW=12)  nco_inst (.dac_clk_p_c(dac_clk_p_c), .n26683(n26683), .increment({increment}), 
            .o_phase({o_phase}), .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(20[49:100])
    
endmodule
//
// Verilog Description of module quarter_wave_sine_lookup
//

module quarter_wave_sine_lookup (dac_clk_p_c, n26683, modulation_output, 
            o_dac_cw_b_c_c, o_phase, \quarter_wave_sample_register_q[15] , 
            GND_net) /* synthesis syn_module_defined=1 */ ;
    input dac_clk_p_c;
    input n26683;
    output [15:0]modulation_output;
    input o_dac_cw_b_c_c;
    input [11:0]o_phase;
    input \quarter_wave_sample_register_q[15] ;
    input GND_net;
    
    wire [15:0]\o_val_pipeline_i[0]  /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(15[24:40])
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(29[49:58])
    wire [15:0]modulation_output_c /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(73[39:56])
    wire [15:0]n1086;
    
    wire n26775, n26776;
    wire [9:0]index_i;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(31[17:24])
    
    wire n26777, n26669, n26681, n526;
    wire [15:0]quarter_wave_sample_register_i;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(22[24:54])
    wire [15:0]o_val_pipeline_i_0__15__N_2158;
    wire [1:0]phase_negation_i;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(23[12:28])
    
    wire n22889, n22890, n22891, n875, n21468, n332, n25382, n22223, 
        n22224, n22231, n541, n23076;
    wire [11:0]phase_i;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(11[17:24])
    wire [9:0]index_i_9__N_2107;
    wire [14:0]quarter_wave_sample_register_i_15__N_2127;
    
    wire n23036, n23037, n23041, n22748, n22749, n22753, n506, 
        n23104, n23105, n23106, n22577, n22578, n22581, n26765, 
        n26766, n26767, n25220, n21291, n21292, n22579, n22580, 
        n22582, n28347, n26798, n22740, n26498, n26600, n254, 
        n124, n24963, n542, n573, n22734, n21765, n26625, n29179, 
        n986, n22232, n22235, n22584, n22585, n22588, n22233, 
        n22234, n22236, n22586, n22587, n22589, n22786, n22787, 
        n22791, n21407, n21408, n476, n26659, n29169, n15, n26371, 
        n20226, n26499, n254_adj_2787, n22591, n22592, n22595, n22593, 
        n22594, n22596, n21425, n21426, n21427, n21452, n26468, 
        n700, n21224, n26858, n26859, n62, n21440, n21441, n21442, 
        n23003, n23004, n23009, n26418, n701, n23024, n23025, 
        n23035, n23026, n23027, n23032, n23033, n23039, n22098, 
        n22099, n22104, n22100, n22101, n22105, n25001, n24998, 
        n25002, n22598, n22599, n22602, n22661, n22662, n22668, 
        n22144, n22145, n22146, n22600, n22601, n22603, n22172, 
        n22173, n22179, n22174, n22175, n22180, n924, n956, n22176, 
        n22177, n22181, n382, n509, n22186, n26758, n26759, n26760, 
        n21194, n21195, n21196, n22227, n22228, n22229, n22230, 
        n22776, n22777, n22780, n22781, n22788, n22782, n22783, 
        n22789, n26621, n25665, n21465, n26467, n20076, n26638, 
        n892, n19585, n12053, n11820, n11823, n364, n443, n22188, 
        n21476, n21477, n21478, n21479, n21480, n21481, n26661, 
        n397, n762, n22168, n25681, n428, n21488, n21489, n21490, 
        n26509, n24371, n604, n14972, n252, n860, n62_adj_2788, 
        n890, n26361, n955, n364_adj_2789, n22517, n26441, n189, 
        n26510, n26416, n637, n22887, n22888, n844, n26508, n316, 
        n22515, n9197, n765, n317, n93, n24426, n21267, n21498, 
        n22885, n22886, n747, n26469, n26666, n29165, n506_adj_2790, 
        n25219, n762_adj_2791, n26752, n26753, n26754, n890_adj_2792, 
        n891, n25149, n25146, n21491, n21492, n21493, n21128, 
        n475, n26348, n252_adj_2793, n26402, n22141, n19592, n26489, 
        n24341, n22877, n22878, n22883, n22884, n21494, n21495, 
        n21496, n22879, n27969, n25254, n22882, n379, n443_adj_2794, 
        n21515, n109, n21497, n21499, n460, n26391, n251, n924_adj_2795, 
        n24343, n24344, n21503, n21504, n21505, n412, n21129, 
        n21486, n26629, n29199, n25251, n21125, n21126, n21127, 
        n26624, n684, n24968, n24964, n24969, n890_adj_2796, n716, 
        n21130, n445, n699, n101, n511, n26826, n26827, n26828, 
        n21509, n21510, n21511, n26596, n763, n24191, n22518, 
        n22519, n21512, n21513, n21514, n24368, n844_adj_2797, n860_adj_2798, 
        n46, n21246, n796, n24789, n26641, n526_adj_2799, n542_adj_2800, 
        n142, n29191, n635, n21264, n29166, n21461, n21143, n21144, 
        n21145, n22525, n22526, n26785, n21516, n21517, n29193, 
        n27967, n653, n141, n21042, n26677, n397_adj_2801, n26784, 
        n26675, n26676, n25412, n26633, n188, n17546, n17547, 
        n17548, n25151, n22583, n22096, n26630, n26664, n25436, 
        n173, n189_adj_2802, n21438, n21134, n21135, n21136, n29168, 
        n14954, n1022, n19553, n491, n508, n26086, n124_adj_2803, 
        n22864, n620, n13842, n21282, n21137, n21138, n21139, 
        n26791, n26551, n475_adj_2804, n491_adj_2805, n26790, n491_adj_2806, 
        n506_adj_2807, n21276, n645, n21039, n21038, n173_adj_2808, 
        n22991, n22992, n22993, n22994, n22995, n22996, n23005, 
        n22997, n22998, n23006, n732, n763_adj_2809, n22185, n22189, 
        n22183, n22178, n22182, n891_adj_2810, n26627, n731, n26673, 
        n23014, n23015, n23030, n23018, n23019, n23020, n23021, 
        n26620, n26617, n24796, n23028, n23029, n21247, n21250, 
        n22094, n190, n25693, n22604, n21271, n22225, n325, n890_adj_2811, 
        n21259, n21262, n22097, n348, n26560, n700_adj_2812, n574, 
        n21265, n21268, n764, n24373, n21164, n1001, n22643, n22644, 
        n22659, n22645, n22646, n22660, n22647, n22648, n22649, 
        n22650, n22651, n22652, n22663, n22102, n22103, n22106, 
        n22655, n22656, n22665, n124_adj_2813, n21249, n221, n24877, 
        n24878, n22140, n22142, n22143, n22790, n22793, n22792, 
        n574_adj_2814, n21197, n26672, n21483, n22156, n22157, n22171, 
        n22158, n22159, n22160, n22161, n22162, n22163, n22164, 
        n22165, n23092, n23093, n23100, n23094, n23095, n23101, 
        n23096, n23097, n23102, n23098, n23099, n23103, n30, n23040, 
        n23043, n23038, n23042, n24199, n24192, n24200, n318, 
        n381, n22726, n22727, n22742, n22728, n22729, n22743, 
        n26679, n21764, n22730, n22731, n22744, n620_adj_2815, n635_adj_2816, 
        n636, n22735, n22746, n22590, n22597, n27963, n22736, 
        n22737, n22747, n22738, n22739, n22741, n27964, n21274, 
        n21277, n22226, n21280, n21283, n21286, n21289, n892_adj_2817, 
        n26616, n21159, n797, n828, n22764, n22765, n22766, n22767, 
        n285, n27966, n22768, n22769, n22770, n22771, n22772, 
        n22773, n22784, n460_adj_2818, n21474, n891_adj_2819, n26575, 
        n286, n22778, n22779, n859, n860_adj_2820, n684_adj_2821, 
        n21446, n26764, n21448, n908, n924_adj_2822, n541_adj_2823, 
        n891_adj_2824, n668, n669, n26639, n11926, n21434, n21435, 
        n21436, n476_adj_2825, n397_adj_2826, n26577, n413, n747_adj_2827, 
        n763_adj_2828, n93_adj_2829, n14747, n286_adj_2830, n14970, 
        n142_adj_2831, n26413, n158, n526_adj_2832, n125, n781, 
        n31, n93_adj_2833, n22863, n21149, n21150, n21151, n25668, 
        n557, n572, n23077, n26797, n25677, n732_adj_2834, n589, 
        n23078, n125_adj_2835, n28204, n252_adj_2836, n28202, n588, 
        n25679, n28205, n26796, n21040, n26611, n25689, n1002, 
        n24792, n860_adj_2837, n908_adj_2838, n21279, n28346, n475_adj_2839, 
        n21416, n21417, n21418, n70, n653_adj_2840, n684_adj_2841, 
        n21281, n21413, n21414, n21415, n684_adj_2842, n700_adj_2843, 
        n668_adj_2844, n669_adj_2845, n26814, n26815, n26816, n221_adj_2846, 
        n21245, n26474, n46_adj_2847, n22862, n19598, n1018, n620_adj_2848, 
        n635_adj_2849, n23079, n700_adj_2850, n270, n15_adj_2851, 
        n286_adj_2852, n26459, n61, n26576, n94, n460_adj_2853, 
        n892_adj_2854, n21248, n716_adj_2855, n731_adj_2856, n732_adj_2857, 
        n653_adj_2858, n475_adj_2859, n669_adj_2860, n124_adj_2861, 
        n24425, n604_adj_2862, n605, n653_adj_2863, n668_adj_2864, 
        n23080, n26769, n21466, n285_adj_2865, n22514, n699_adj_2866, 
        n23081, n21462, n21463, n573_adj_2867, n557_adj_2868, n573_adj_2869, 
        n22149, n397_adj_2870, n954, n413_adj_2871, n316_adj_2872, 
        n317_adj_2873, n270_adj_2874, n286_adj_2875, n21152, n21153, 
        n21154, n13969, n158_adj_2876, n26660, n26640, n62_adj_2877, 
        n21257, n21258, n716_adj_2878, n23082, n21161, n11912, n731_adj_2879, 
        n732_adj_2880, n26454, n31_adj_2881, n21260, n21261, n21263, 
        n747_adj_2882, n762_adj_2883, n23083, n21266, n21269, n21270, 
        n21155, n21156, n21157, n28801, n781_adj_2884, n23084, n24345, 
        n25814, n22664, n25815, n25817, n25818, n25816, n28800, 
        n28802, n28803, n28804, n28805, n812, n23085, n28806, 
        n28807, n875_adj_2885, n23087, n923, n23088, n28207, n25845, 
        n26351, n25841, n939, n954_adj_2886, n23089, n971, n986_adj_2887, 
        n23090, n875_adj_2888, n379_adj_2889, n891_adj_2890, n1002_adj_2891, 
        n1017, n23091, n859_adj_2892, n860_adj_2893, n21272, n21273, 
        n21162, n21163, n21275, n21158, n21160, n21278, n157, 
        n26480, n636_adj_2894, n24809, n26586, n24810, n21284, n21285, 
        n26665, n26682, n444, n17549, n17550, n17551, n507, n21287, 
        n21288, n460_adj_2895, n476_adj_2896, n26670, n24807, n24808, 
        n747_adj_2897, n251_adj_2898, n413_adj_2899, n26613, n24788, 
        n763_adj_2900, n24805, n24802, n24806, n17580, n17581, n17582, 
        n21437, n109_adj_2901, n125_adj_2902, n653_adj_2903, n635_adj_2904, 
        n94_adj_2905, n491_adj_2906, n24997, n30_adj_2907, n31_adj_2908, 
        n443_adj_2909, n158_adj_2910, n189_adj_2911, n316_adj_2912, 
        n412_adj_2913, n924_adj_2914, n25884, n859_adj_2915, n860_adj_2916, 
        n25885, n25890, n14741, n21506, n21507, n21508, n26406, 
        n26405, n26642, n404, n26662, n24804, n173_adj_2917, n26105, 
        n26102, n26104, n26103, n348_adj_2918, n349, n21482, n21484, 
        n22861, n11938, n11939, n93_adj_2919, n94_adj_2920, n22865, 
        n22866, n26680, n21402, n14379, n636_adj_2921, n24193, n26344, 
        n24801, n21141, n987, n22871, n22872, n26101, n301, n890_adj_2922, 
        n891_adj_2923, n22873, n22874, n812_adj_2924, n13872, n828_adj_2925, 
        n26360, n797_adj_2926, n668_adj_2927, n669_adj_2928, n24800, 
        n22988, n25942, n14872, n26345, n22989, n25941, n22875, 
        n22876, n24794, n22984, n25944, n526_adj_2929, n542_adj_2930, 
        n26085, n731_adj_2931, n11082, n252_adj_2932, n25383, n22986, 
        n24799, n24797, n24798, n26626, n26628, n15_adj_2933, n24795, 
        n24791, n26396, n24342, n24793, n24790, n26614, n475_adj_2934, 
        n333, n348_adj_2935, n15_adj_2936, n30_adj_2937, n26678, n21443, 
        n397_adj_2938, n142_adj_2939, n22516, n22521, n22522, n22523, 
        n22524, n716_adj_2940, n14714, n157_adj_2941, n93_adj_2942, 
        n700_adj_2943, n526_adj_2944, n21458, n985, n26507, n766, 
        n21165, n20368, n11838, n24196, n26377, n11839, n364_adj_2945, 
        n30_adj_2946, n24428, n24197, n413_adj_2947, n491_adj_2948, 
        n26674, n26656, n11888, n25945, n25943, n25946, n573_adj_2949, 
        n605_adj_2950, n23000, n700_adj_2951, n732_adj_2952, n1021, 
        n21475, n23016, n62_adj_2953, n317_adj_2954, n21487, n26658, 
        n85, n108, n684_adj_2955, n21147, n21146, n21148, n24872, 
        n23023, n26786, n24876, n844_adj_2956, n23086, n24879, n21520, 
        n20077, n26654, n21523, n14378, n21401, n21403, n908_adj_2957, 
        n924_adj_2958, n605_adj_2959, n573_adj_2960, n26612, n26663, 
        n26667, n348_adj_2961, n22653, n21938, n348_adj_2962, n21766, 
        n22654, n797_adj_2963, n828_adj_2964, n21521, n21522, n25843, 
        n23031, n25417, n23034, n25438, n25842, n22785, n22774, 
        n22775, n882, n890_adj_2965, n26552, n21518, n11000, n21519, 
        n221_adj_2966, n24430, n11840, n26792, n796_adj_2967, n684_adj_2968, 
        n700_adj_2969, n21454, n349_adj_2970, n21457, n21460, n507_adj_2971, 
        n21469, n763_adj_2972, n25676, n22167, n21397, n23012, n23010, 
        n221_adj_2973, n252_adj_2974, n24965, n21400, n349_adj_2975, 
        n25148, n25433, n25413, n828_adj_2976, n17398, n17397, n25252, 
        n812_adj_2977, n21421, n25692, n25690, n25691, n17396, n25680, 
        n25678, n28206, n28203, n572_adj_2978, n716_adj_2979, n25669, 
        n25666, n25670, n25667, n11930, n21396, n26368, n62_adj_2980, 
        n21459, n94_adj_2981, n21485, n21430, n21395, n26417, n301_adj_2982, 
        n349_adj_2983, n21433, n21399, n444_adj_2984, n507_adj_2985, 
        n21439, n25218, n900, n21445, n21398, n27968, n27965, 
        n17395, n26773, n21467, n491_adj_2986, n12052, n22053, n205, 
        n24198, n348_adj_2987, n21456, n444_adj_2988, n21455, n22107, 
        n21453, n572_adj_2989, n25434, n21444, n22190, n491_adj_2990, 
        n25249, n17394, n638, n157_adj_2991, n21419, n25415, n21432, 
        n21431, n21429, n21428, n142_adj_2992, n25437, n25435, n21501, 
        n24429, n24427, n19900, n333_adj_2993, n25416, n25414, n21420, 
        n24372, n25253, n25250, n17393, n17392, n17391, n25150, 
        n25147;
    
    FD1S3DX o_val_pipeline_i_1__i32 (.D(n1086[15]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(\o_val_pipeline_i[0] [15])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i32.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i31 (.D(n1086[14]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(\o_val_pipeline_i[0] [14])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i31.GSR = "DISABLED";
    PFUMX i24487 (.BLUT(n26775), .ALUT(n26776), .C0(index_i[1]), .Z(n26777));
    FD1S3DX o_val_pipeline_i_1__i30 (.D(n1086[13]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(\o_val_pipeline_i[0] [13])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i30.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i29 (.D(n1086[12]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(\o_val_pipeline_i[0] [12])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i29.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i28 (.D(n1086[11]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(\o_val_pipeline_i[0] [11])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i28.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i27 (.D(n1086[10]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(\o_val_pipeline_i[0] [10])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i27.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i26 (.D(n1086[9]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(\o_val_pipeline_i[0] [9])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i26.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i25 (.D(n1086[8]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(\o_val_pipeline_i[0] [8])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i25.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i24 (.D(n1086[7]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(\o_val_pipeline_i[0] [7])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i24.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i23 (.D(n1086[6]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(\o_val_pipeline_i[0] [6])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i23.GSR = "DISABLED";
    LUT4 mux_193_Mux_0_i526_3_lut (.A(n26669), .B(n26681), .C(index_i[3]), 
         .Z(n526)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i526_3_lut.init = 16'hcaca;
    LUT4 mux_190_i14_3_lut (.A(quarter_wave_sample_register_i[13]), .B(o_val_pipeline_i_0__15__N_2158[13]), 
         .C(phase_negation_i[1]), .Z(n1086[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam mux_190_i14_3_lut.init = 16'hcaca;
    PFUMX i20552 (.BLUT(n22889), .ALUT(n22890), .C0(index_i[8]), .Z(n22891));
    LUT4 i9489_3_lut_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n875)) /* synthesis lut_function=(A (C (D))+!A !(B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9489_3_lut_3_lut_4_lut_4_lut.init = 16'hb555;
    FD1S3DX o_val_pipeline_i_1__i22 (.D(n1086[5]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(\o_val_pipeline_i[0] [5])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i22.GSR = "DISABLED";
    LUT4 i19148_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n21468)) /* synthesis lut_function=(A (C+(D))+!A !(B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19148_3_lut_4_lut_4_lut.init = 16'haba5;
    LUT4 mux_193_Mux_6_i332_3_lut_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n332)) /* synthesis lut_function=(!(A (C)+!A !((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_6_i332_3_lut_3_lut_3_lut.init = 16'h5b5b;
    LUT4 i23291_then_3_lut (.A(index_i[0]), .B(index_i[4]), .C(index_i[3]), 
         .Z(n26776)) /* synthesis lut_function=(A (B)+!A (B (C)+!B !(C))) */ ;
    defparam i23291_then_3_lut.init = 16'hc9c9;
    FD1S3DX o_val_pipeline_i_1__i21 (.D(n1086[4]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(\o_val_pipeline_i[0] [4])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i21.GSR = "DISABLED";
    LUT4 n72_bdd_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n25382)) /* synthesis lut_function=(!(A (D)+!A !(B (D)+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n72_bdd_4_lut_4_lut_4_lut.init = 16'h54bb;
    LUT4 i19892_3_lut (.A(n22223), .B(n22224), .C(index_i[7]), .Z(n22231)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19892_3_lut.init = 16'hcaca;
    PFUMX i20737 (.BLUT(n526), .ALUT(n541), .C0(index_i[4]), .Z(n23076));
    FD1S3DX o_val_pipeline_i_1__i20 (.D(n1086[3]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(\o_val_pipeline_i[0] [3])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i20.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i19 (.D(n1086[2]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(\o_val_pipeline_i[0] [2])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i19.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i18 (.D(n1086[1]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(\o_val_pipeline_i[0] [1])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i18.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i17 (.D(n1086[0]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(\o_val_pipeline_i[0] [0])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i17.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i16 (.D(\o_val_pipeline_i[0] [15]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(modulation_output[15])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i16.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i15 (.D(\o_val_pipeline_i[0] [14]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(modulation_output[14])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i15.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i14 (.D(\o_val_pipeline_i[0] [13]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(modulation_output[13])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i14.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i13 (.D(\o_val_pipeline_i[0] [12]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(modulation_output[12])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i13.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i12 (.D(\o_val_pipeline_i[0] [11]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(modulation_output[11])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i12.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i11 (.D(\o_val_pipeline_i[0] [10]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(modulation_output[10])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i11.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i10 (.D(\o_val_pipeline_i[0] [9]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(modulation_output[9])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i10.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i9 (.D(\o_val_pipeline_i[0] [8]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(modulation_output[8])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i9.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i8 (.D(\o_val_pipeline_i[0] [7]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(modulation_output[7])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i8.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i7 (.D(\o_val_pipeline_i[0] [6]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(modulation_output[6])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i7.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i6 (.D(\o_val_pipeline_i[0] [5]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(modulation_output[5])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i6.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i0 (.D(o_phase[0]), .SP(o_dac_cw_b_c_c), .CK(dac_clk_p_c), 
            .Q(phase_i[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i0.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i5 (.D(\o_val_pipeline_i[0] [4]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(modulation_output[4])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i5.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i4 (.D(\o_val_pipeline_i[0] [3]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(modulation_output[3])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i4.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i3 (.D(\o_val_pipeline_i[0] [2]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(modulation_output[2])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i3.GSR = "DISABLED";
    FD1S3DX phase_negation_i_i0 (.D(phase_i[11]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(phase_negation_i[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_negation_i_i0.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i2 (.D(\o_val_pipeline_i[0] [1]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(modulation_output[1])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i2.GSR = "DISABLED";
    FD1S3DX index_i_i0 (.D(index_i_9__N_2107[0]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(index_i[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_i_i0.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i1 (.D(\o_val_pipeline_i[0] [0]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(modulation_output[0])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i1.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i0 (.D(quarter_wave_sample_register_i_15__N_2127[0]), 
            .CK(dac_clk_p_c), .PD(n26683), .Q(quarter_wave_sample_register_i[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i0.GSR = "DISABLED";
    FD1S3DX index_i_i9 (.D(index_i_9__N_2107[9]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(index_i[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_i_i9.GSR = "DISABLED";
    L6MUX21 i20702 (.D0(n23036), .D1(n23037), .SD(index_i[7]), .Z(n23041));
    FD1S3DX index_i_i8 (.D(index_i_9__N_2107[8]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(index_i[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_i_i8.GSR = "DISABLED";
    FD1S3DX index_i_i7 (.D(index_i_9__N_2107[7]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(index_i[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_i_i7.GSR = "DISABLED";
    FD1S3DX index_i_i6 (.D(index_i_9__N_2107[6]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(index_i[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_i_i6.GSR = "DISABLED";
    FD1S3DX index_i_i5 (.D(index_i_9__N_2107[5]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(index_i[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_i_i5.GSR = "DISABLED";
    FD1S3DX index_i_i4 (.D(index_i_9__N_2107[4]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(index_i[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_i_i4.GSR = "DISABLED";
    FD1S3DX index_i_i3 (.D(index_i_9__N_2107[3]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(index_i[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_i_i3.GSR = "DISABLED";
    FD1S3DX index_i_i2 (.D(index_i_9__N_2107[2]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(index_i[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_i_i2.GSR = "DISABLED";
    FD1S3DX index_i_i1 (.D(index_i_9__N_2107[1]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(index_i[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_i_i1.GSR = "DISABLED";
    LUT4 i23291_else_3_lut (.A(index_i[2]), .B(index_i[0]), .C(index_i[4]), 
         .D(index_i[3]), .Z(n26775)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)+!C !(D)))+!A (B (C+!(D))+!B !(C)))) */ ;
    defparam i23291_else_3_lut.init = 16'h1e38;
    FD1S3DX phase_negation_i_i1 (.D(phase_negation_i[0]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(phase_negation_i[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_negation_i_i1.GSR = "DISABLED";
    LUT4 i20414_3_lut (.A(n22748), .B(n22749), .C(index_i[7]), .Z(n22753)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20414_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_8_i506_3_lut_4_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n506)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_8_i506_3_lut_4_lut_3_lut_4_lut.init = 16'h0ef0;
    PFUMX i20767 (.BLUT(n23104), .ALUT(n23105), .C0(index_i[8]), .Z(n23106));
    PFUMX i20242 (.BLUT(n22577), .ALUT(n22578), .C0(index_i[4]), .Z(n22581));
    PFUMX i24481 (.BLUT(n26765), .ALUT(n26766), .C0(index_i[2]), .Z(n26767));
    FD1P3AX phase_i_i0_i11 (.D(o_phase[11]), .SP(o_dac_cw_b_c_c), .CK(dac_clk_p_c), 
            .Q(phase_i[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i11.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i10 (.D(o_phase[10]), .SP(o_dac_cw_b_c_c), .CK(dac_clk_p_c), 
            .Q(phase_i[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i10.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i9 (.D(o_phase[9]), .SP(o_dac_cw_b_c_c), .CK(dac_clk_p_c), 
            .Q(phase_i[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i9.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i8 (.D(o_phase[8]), .SP(o_dac_cw_b_c_c), .CK(dac_clk_p_c), 
            .Q(phase_i[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i8.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i7 (.D(o_phase[7]), .SP(o_dac_cw_b_c_c), .CK(dac_clk_p_c), 
            .Q(phase_i[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i7.GSR = "DISABLED";
    LUT4 i21850_3_lut (.A(n25220), .B(n21291), .C(index_i[5]), .Z(n21292)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21850_3_lut.init = 16'hcaca;
    PFUMX i20243 (.BLUT(n22579), .ALUT(n22580), .C0(index_i[4]), .Z(n22582));
    LUT4 i23322_else_4_lut (.A(index_i[0]), .B(index_i[4]), .C(index_i[1]), 
         .D(index_i[3]), .Z(n26765)) /* synthesis lut_function=(!(A (B (C)+!B !(C (D)+!C !(D)))+!A (B ((D)+!C)+!B !((D)+!C)))) */ ;
    defparam i23322_else_4_lut.init = 16'h394b;
    FD1P3AX phase_i_i0_i6 (.D(o_phase[6]), .SP(o_dac_cw_b_c_c), .CK(dac_clk_p_c), 
            .Q(phase_i[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i6.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i5 (.D(o_phase[5]), .SP(o_dac_cw_b_c_c), .CK(dac_clk_p_c), 
            .Q(phase_i[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i5.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i4 (.D(o_phase[4]), .SP(o_dac_cw_b_c_c), .CK(dac_clk_p_c), 
            .Q(phase_i[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i4.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i3 (.D(o_phase[3]), .SP(o_dac_cw_b_c_c), .CK(dac_clk_p_c), 
            .Q(phase_i[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i3.GSR = "DISABLED";
    LUT4 i21857_3_lut (.A(n28347), .B(n26798), .C(index_i[5]), .Z(n22740)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21857_3_lut.init = 16'hcaca;
    LUT4 i11185_2_lut_3_lut_4_lut (.A(n26498), .B(n26600), .C(index_i[6]), 
         .D(index_i[5]), .Z(n254)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i11185_2_lut_3_lut_4_lut.init = 16'hfef0;
    FD1P3AX phase_i_i0_i2 (.D(o_phase[2]), .SP(o_dac_cw_b_c_c), .CK(dac_clk_p_c), 
            .Q(phase_i[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i2.GSR = "DISABLED";
    LUT4 n476_bdd_3_lut_23320_3_lut (.A(index_i[1]), .B(index_i[4]), .C(n124), 
         .Z(n24963)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n476_bdd_3_lut_23320_3_lut.init = 16'hd1d1;
    FD1P3AX phase_i_i0_i1 (.D(o_phase[1]), .SP(o_dac_cw_b_c_c), .CK(dac_clk_p_c), 
            .Q(phase_i[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i1.GSR = "DISABLED";
    LUT4 i21867_3_lut (.A(n542), .B(n573), .C(index_i[5]), .Z(n22734)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21867_3_lut.init = 16'hcaca;
    LUT4 i19445_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21765)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A (B (C (D)+!C !(D))+!B (D))) */ ;
    defparam i19445_3_lut_4_lut.init = 16'hd926;
    LUT4 mux_193_Mux_1_i986_3_lut (.A(n26625), .B(n29179), .C(index_i[3]), 
         .Z(n986)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_1_i986_3_lut.init = 16'hcaca;
    PFUMX i19896 (.BLUT(n22231), .ALUT(n22232), .C0(index_i[8]), .Z(n22235));
    PFUMX i20249 (.BLUT(n22584), .ALUT(n22585), .C0(index_i[4]), .Z(n22588));
    L6MUX21 i19897 (.D0(n22233), .D1(n22234), .SD(index_i[8]), .Z(n22236));
    PFUMX i20250 (.BLUT(n22586), .ALUT(n22587), .C0(index_i[4]), .Z(n22589));
    L6MUX21 i20452 (.D0(n22786), .D1(n22787), .SD(index_i[7]), .Z(n22791));
    PFUMX i19089 (.BLUT(n21407), .ALUT(n21408), .C0(index_i[4]), .Z(n476));
    LUT4 mux_193_Mux_5_i15_3_lut (.A(n26659), .B(n29169), .C(index_i[3]), 
         .Z(n15)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_5_i15_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_12_i254_4_lut (.A(n26371), .B(n20226), .C(index_i[6]), 
         .D(n26499), .Z(n254_adj_2787)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_12_i254_4_lut.init = 16'hca0a;
    PFUMX i20256 (.BLUT(n22591), .ALUT(n22592), .C0(index_i[4]), .Z(n22595));
    PFUMX i20257 (.BLUT(n22593), .ALUT(n22594), .C0(index_i[4]), .Z(n22596));
    PFUMX i19107 (.BLUT(n21425), .ALUT(n21426), .C0(index_i[4]), .Z(n21427));
    LUT4 i19132_3_lut_3_lut_4_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n21452)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19132_3_lut_3_lut_4_lut_3_lut_4_lut.init = 16'h11ef;
    LUT4 i18904_3_lut_3_lut_4_lut (.A(n26468), .B(index_i[4]), .C(n700), 
         .D(index_i[5]), .Z(n21224)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18904_3_lut_3_lut_4_lut.init = 16'hf011;
    PFUMX i24541 (.BLUT(n26858), .ALUT(n26859), .C0(index_i[3]), .Z(n62));
    PFUMX i19122 (.BLUT(n21440), .ALUT(n21441), .C0(index_i[4]), .Z(n21442));
    L6MUX21 i20670 (.D0(n23003), .D1(n23004), .SD(index_i[7]), .Z(n23009));
    LUT4 mux_193_Mux_10_i701_4_lut_4_lut (.A(n26468), .B(index_i[4]), .C(index_i[5]), 
         .D(n26418), .Z(n701)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B (C (D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_10_i701_4_lut_4_lut.init = 16'h3efe;
    L6MUX21 i20696 (.D0(n23024), .D1(n23025), .SD(index_i[6]), .Z(n23035));
    L6MUX21 i20697 (.D0(n23026), .D1(n23027), .SD(index_i[6]), .Z(n23036));
    L6MUX21 i20700 (.D0(n23032), .D1(n23033), .SD(index_i[7]), .Z(n23039));
    L6MUX21 i19765 (.D0(n22098), .D1(n22099), .SD(index_i[7]), .Z(n22104));
    PFUMX i19766 (.BLUT(n22100), .ALUT(n22101), .C0(index_i[7]), .Z(n22105));
    PFUMX i23324 (.BLUT(n25001), .ALUT(n24998), .C0(index_i[6]), .Z(n25002));
    PFUMX i20263 (.BLUT(n22598), .ALUT(n22599), .C0(index_i[4]), .Z(n22602));
    L6MUX21 i20329 (.D0(n22661), .D1(n22662), .SD(index_i[7]), .Z(n22668));
    L6MUX21 i19807 (.D0(n22144), .D1(n22145), .SD(index_i[7]), .Z(n22146));
    PFUMX i20264 (.BLUT(n22600), .ALUT(n22601), .C0(index_i[4]), .Z(n22603));
    L6MUX21 i19840 (.D0(n22172), .D1(n22173), .SD(index_i[7]), .Z(n22179));
    L6MUX21 i19841 (.D0(n22174), .D1(n22175), .SD(index_i[7]), .Z(n22180));
    LUT4 mux_193_Mux_7_i956_3_lut_3_lut_4_lut (.A(n26468), .B(index_i[4]), 
         .C(n924), .D(index_i[5]), .Z(n956)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_7_i956_3_lut_3_lut_4_lut.init = 16'h11f0;
    PFUMX i19842 (.BLUT(n22176), .ALUT(n22177), .C0(index_i[7]), .Z(n22181));
    L6MUX21 i19847 (.D0(n382), .D1(n509), .SD(index_i[7]), .Z(n22186));
    PFUMX i24477 (.BLUT(n26758), .ALUT(n26759), .C0(index_i[1]), .Z(n26760));
    L6MUX21 i18876 (.D0(n21194), .D1(n21195), .SD(index_i[7]), .Z(n21196));
    L6MUX21 i19894 (.D0(n22227), .D1(n22228), .SD(index_i[7]), .Z(n22233));
    L6MUX21 i19895 (.D0(n22229), .D1(n22230), .SD(index_i[7]), .Z(n22234));
    L6MUX21 i20447 (.D0(n22776), .D1(n22777), .SD(index_i[6]), .Z(n22786));
    L6MUX21 i20449 (.D0(n22780), .D1(n22781), .SD(index_i[7]), .Z(n22788));
    L6MUX21 i20450 (.D0(n22782), .D1(n22783), .SD(index_i[7]), .Z(n22789));
    LUT4 mux_193_Mux_0_i363_3_lut_4_lut_3_lut_rep_661 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26621)) /* synthesis lut_function=(A (B+!(C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i363_3_lut_4_lut_3_lut_rep_661.init = 16'hdbdb;
    LUT4 n348_bdd_3_lut_23984_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n25665)) /* synthesis lut_function=(A (B (C)+!B (C+(D)))+!A (B (C)+!B !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n348_bdd_3_lut_23984_4_lut_4_lut_4_lut.init = 16'he3f0;
    LUT4 i19145_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21465)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D))+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19145_3_lut_4_lut.init = 16'hccdb;
    LUT4 i1_4_lut (.A(index_i[6]), .B(n26467), .C(index_i[5]), .D(index_i[4]), 
         .Z(n20076)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i1_4_lut.init = 16'hfffe;
    LUT4 i17413_4_lut (.A(n26638), .B(n892), .C(index_i[6]), .D(index_i[5]), 
         .Z(n19585)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D))))) */ ;
    defparam i17413_4_lut.init = 16'h3a35;
    LUT4 i9603_3_lut_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n12053)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A !(B (C+(D))+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9603_3_lut_3_lut_4_lut_4_lut.init = 16'h44db;
    LUT4 i9374_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n11820)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))+!A !(B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9374_3_lut_4_lut_4_lut.init = 16'hb5b3;
    LUT4 i9377_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n11823)) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B ((D)+!C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9377_3_lut_4_lut_4_lut.init = 16'hcdad;
    LUT4 mux_193_Mux_0_i364_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n364)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A ((C+!(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i364_3_lut_3_lut_4_lut.init = 16'hdb55;
    LUT4 mux_193_Mux_0_i443_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .D(index_i[3]), .Z(n443)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C (D))+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i443_3_lut_4_lut_4_lut_4_lut.init = 16'h0ed5;
    LUT4 i22190_3_lut (.A(n19585), .B(n20076), .C(index_i[7]), .Z(n22188)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22190_3_lut.init = 16'hcaca;
    LUT4 mux_190_i12_3_lut (.A(quarter_wave_sample_register_i[11]), .B(o_val_pipeline_i_0__15__N_2158[11]), 
         .C(phase_negation_i[1]), .Z(n1086[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam mux_190_i12_3_lut.init = 16'hcaca;
    PFUMX i19158 (.BLUT(n21476), .ALUT(n21477), .C0(index_i[4]), .Z(n21478));
    PFUMX i19161 (.BLUT(n21479), .ALUT(n21480), .C0(index_i[4]), .Z(n21481));
    LUT4 mux_190_i11_3_lut (.A(quarter_wave_sample_register_i[10]), .B(o_val_pipeline_i_0__15__N_2158[10]), 
         .C(phase_negation_i[1]), .Z(n1086[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam mux_190_i11_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_5_i397_3_lut (.A(n26661), .B(n332), .C(index_i[3]), 
         .Z(n397)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_5_i397_3_lut.init = 16'hcaca;
    LUT4 mux_190_i10_3_lut (.A(quarter_wave_sample_register_i[9]), .B(o_val_pipeline_i_0__15__N_2158[9]), 
         .C(phase_negation_i[1]), .Z(n1086[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam mux_190_i10_3_lut.init = 16'hcaca;
    LUT4 i9482_3_lut_3_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[0]), .D(index_i[1]), .Z(n762)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C (D)+!C !(D)))+!A !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9482_3_lut_3_lut_4_lut_4_lut.init = 16'h700f;
    LUT4 mux_190_i9_3_lut (.A(quarter_wave_sample_register_i[8]), .B(o_val_pipeline_i_0__15__N_2158[8]), 
         .C(phase_negation_i[1]), .Z(n1086[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam mux_190_i9_3_lut.init = 16'hcaca;
    LUT4 i22108_3_lut (.A(n22168), .B(n25681), .C(index_i[6]), .Z(n22177)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22108_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_0_i428_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[2]), 
         .B(index_i[0]), .C(index_i[1]), .D(index_i[3]), .Z(n428)) /* synthesis lut_function=(A (B (C+!(D))+!B !((D)+!C))+!A (B (D)+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i428_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hd5a9;
    PFUMX i19170 (.BLUT(n21488), .ALUT(n21489), .C0(index_i[4]), .Z(n21490));
    LUT4 index_i_4__bdd_3_lut_22785_4_lut (.A(n26509), .B(index_i[3]), .C(index_i[5]), 
         .D(index_i[4]), .Z(n24371)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam index_i_4__bdd_3_lut_22785_4_lut.init = 16'hf080;
    LUT4 mux_193_Mux_0_i604_3_lut_4_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[1]), .D(index_i[3]), .Z(n604)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A !(B (D)+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i604_3_lut_4_lut_4_lut_4_lut.init = 16'h5439;
    LUT4 mux_190_i8_3_lut (.A(quarter_wave_sample_register_i[7]), .B(o_val_pipeline_i_0__15__N_2158[7]), 
         .C(phase_negation_i[1]), .Z(n1086[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam mux_190_i8_3_lut.init = 16'hcaca;
    LUT4 mux_190_i7_3_lut (.A(quarter_wave_sample_register_i[6]), .B(o_val_pipeline_i_0__15__N_2158[6]), 
         .C(phase_negation_i[1]), .Z(n1086[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam mux_190_i7_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_3_i252_3_lut_4_lut (.A(n26509), .B(index_i[3]), .C(index_i[4]), 
         .D(n14972), .Z(n252)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_3_i252_3_lut_4_lut.init = 16'h08f8;
    LUT4 mux_193_Mux_8_i860_3_lut_4_lut (.A(n26509), .B(index_i[3]), .C(index_i[4]), 
         .D(n26467), .Z(n860)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_8_i860_3_lut_4_lut.init = 16'h08f8;
    LUT4 mux_193_Mux_10_i62_3_lut_3_lut_4_lut (.A(n26509), .B(index_i[3]), 
         .C(n26467), .D(index_i[4]), .Z(n62_adj_2788)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_10_i62_3_lut_3_lut_4_lut.init = 16'hf077;
    LUT4 mux_193_Mux_2_i890_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n890)) /* synthesis lut_function=(A (B (C)+!B !(C+!(D)))+!A !(B (C+(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_2_i890_3_lut_4_lut_4_lut.init = 16'h9394;
    LUT4 mux_193_Mux_6_i955_3_lut_4_lut (.A(n26509), .B(index_i[3]), .C(index_i[4]), 
         .D(n26361), .Z(n955)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_6_i955_3_lut_4_lut.init = 16'h8f80;
    LUT4 i20178_3_lut_4_lut (.A(n26509), .B(index_i[3]), .C(index_i[4]), 
         .D(n364_adj_2789), .Z(n22517)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20178_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_193_Mux_3_i189_3_lut_3_lut_4_lut (.A(n26509), .B(index_i[3]), 
         .C(index_i[4]), .D(n26441), .Z(n189)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_3_i189_3_lut_3_lut_4_lut.init = 16'h08f8;
    LUT4 mux_193_Mux_10_i637_3_lut_4_lut_4_lut (.A(n26510), .B(index_i[4]), 
         .C(index_i[5]), .D(n26416), .Z(n637)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_10_i637_3_lut_4_lut_4_lut.init = 16'h1f1c;
    LUT4 i20551_3_lut (.A(n22887), .B(n22888), .C(index_i[7]), .Z(n22890)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20551_3_lut.init = 16'hcaca;
    LUT4 i9487_3_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[3]), .C(index_i[0]), 
         .D(index_i[1]), .Z(n844)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9487_3_lut_4_lut_4_lut.init = 16'hf00e;
    LUT4 i20176_3_lut_3_lut_4_lut (.A(n26508), .B(index_i[3]), .C(n316), 
         .D(index_i[4]), .Z(n22515)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20176_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 i11210_3_lut_4_lut (.A(n26508), .B(index_i[3]), .C(n9197), .D(index_i[6]), 
         .Z(n765)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11210_3_lut_4_lut.init = 16'hffe0;
    LUT4 mux_193_Mux_10_i317_3_lut_3_lut_4_lut (.A(n26508), .B(index_i[3]), 
         .C(n26441), .D(index_i[4]), .Z(n317)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_10_i317_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 n699_bdd_3_lut_24280_4_lut (.A(n26508), .B(index_i[3]), .C(index_i[4]), 
         .D(n93), .Z(n24426)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n699_bdd_3_lut_24280_4_lut.init = 16'hfe0e;
    LUT4 i18947_3_lut_3_lut_4_lut (.A(n26508), .B(index_i[3]), .C(n93), 
         .D(index_i[4]), .Z(n21267)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18947_3_lut_3_lut_4_lut.init = 16'h11f0;
    LUT4 i19178_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n21498)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B (C+!(D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19178_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h1c18;
    LUT4 i20550_3_lut (.A(n22885), .B(n22886), .C(index_i[7]), .Z(n22889)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20550_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_7_i747_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), 
         .B(index_i[2]), .C(index_i[3]), .D(index_i[0]), .Z(n747)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))+!A (B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_7_i747_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'he1e3;
    LUT4 mux_193_Mux_9_i700_3_lut_4_lut (.A(n26508), .B(index_i[3]), .C(index_i[4]), 
         .D(n26469), .Z(n700)) /* synthesis lut_function=(!(A (C+!(D))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_9_i700_3_lut_4_lut.init = 16'h1f10;
    LUT4 mux_193_Mux_5_i506_3_lut (.A(n26666), .B(n29165), .C(index_i[3]), 
         .Z(n506_adj_2790)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_5_i506_3_lut.init = 16'hcaca;
    LUT4 n172_bdd_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n25219)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n172_bdd_3_lut_4_lut_4_lut_4_lut.init = 16'h1e1c;
    LUT4 mux_193_Mux_7_i762_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), 
         .B(index_i[2]), .C(index_i[3]), .D(index_i[0]), .Z(n762_adj_2791)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B ((D)+!C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_7_i762_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h3878;
    PFUMX i24473 (.BLUT(n26752), .ALUT(n26753), .C0(index_i[1]), .Z(n26754));
    LUT4 mux_193_Mux_7_i891_3_lut_4_lut (.A(n26508), .B(index_i[3]), .C(index_i[4]), 
         .D(n890_adj_2792), .Z(n891)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_7_i891_3_lut_4_lut.init = 16'hfe0e;
    LUT4 mux_193_Mux_9_i316_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), 
         .B(index_i[2]), .C(index_i[3]), .D(index_i[0]), .Z(n316)) /* synthesis lut_function=(!(A (B (C)+!B !(C+(D)))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_9_i316_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h7e7c;
    LUT4 n22_bdd_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n25149)) /* synthesis lut_function=(A (B (C)+!B ((D)+!C))+!A (B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n22_bdd_3_lut_4_lut_4_lut_4_lut.init = 16'he7c7;
    LUT4 i19160_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n21480)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B (C+(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19160_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h7c78;
    LUT4 n301_bdd_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n25146)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A !((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n301_bdd_3_lut_4_lut_4_lut_4_lut.init = 16'h7173;
    PFUMX i19173 (.BLUT(n21491), .ALUT(n21492), .C0(index_i[4]), .Z(n21493));
    LUT4 i18808_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[1]), .Z(n21128)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+!(D)))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18808_3_lut_4_lut_4_lut_4_lut.init = 16'h9399;
    LUT4 mux_193_Mux_5_i475_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[1]), .Z(n475)) /* synthesis lut_function=(A (B ((D)+!C))+!A (B (C)+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_5_i475_3_lut_4_lut_4_lut.init = 16'hd949;
    LUT4 i11182_3_lut_4_lut (.A(n26348), .B(index_i[7]), .C(index_i[8]), 
         .D(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2127[14])) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11182_3_lut_4_lut.init = 16'hffe0;
    LUT4 mux_193_Mux_5_i252_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[4]), .Z(n252_adj_2793)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+(D)))+!A (B (C (D))+!B !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_5_i252_3_lut_4_lut.init = 16'hc993;
    LUT4 i19802_3_lut_4_lut_4_lut (.A(n26467), .B(index_i[4]), .C(index_i[5]), 
         .D(n26402), .Z(n22141)) /* synthesis lut_function=(A ((C+!(D))+!B)+!A (B (C+!(D))+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19802_3_lut_4_lut_4_lut.init = 16'he3ef;
    LUT4 n954_bdd_3_lut_22759 (.A(n19592), .B(n26489), .C(index_i[5]), 
         .Z(n24341)) /* synthesis lut_function=(A (B (C))+!A (B+!(C))) */ ;
    defparam n954_bdd_3_lut_22759.init = 16'hc5c5;
    L6MUX21 i20546 (.D0(n22877), .D1(n22878), .SD(index_i[6]), .Z(n22885));
    L6MUX21 i20549 (.D0(n22883), .D1(n22884), .SD(index_i[6]), .Z(n22888));
    PFUMX i19176 (.BLUT(n21494), .ALUT(n21495), .C0(index_i[4]), .Z(n21496));
    LUT4 i20547_3_lut (.A(n22879), .B(n27969), .C(index_i[6]), .Z(n22886)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20547_3_lut.init = 16'hcaca;
    LUT4 i20548_3_lut (.A(n25254), .B(n22882), .C(index_i[6]), .Z(n22887)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20548_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_0_i379_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n379)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !((D)+!C))+!A !(B ((D)+!C)+!B (D))) */ ;
    defparam mux_193_Mux_0_i379_3_lut_4_lut_4_lut.init = 16'h8079;
    LUT4 mux_193_Mux_8_i443_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n443_adj_2794)) /* synthesis lut_function=(A (B (C+!(D))+!B !((D)+!C))+!A !(B (D)+!B ((D)+!C))) */ ;
    defparam mux_193_Mux_8_i443_3_lut_4_lut_4_lut.init = 16'h80fc;
    LUT4 i19195_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n21515)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B+(C+(D))))) */ ;
    defparam i19195_3_lut_4_lut_4_lut_4_lut.init = 16'h2aab;
    LUT4 i20239_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n22578)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20239_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hf81f;
    LUT4 mux_193_Mux_8_i109_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n109)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C+!(D)))+!A (B (C (D)+!C !(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_8_i109_3_lut_4_lut_4_lut.init = 16'hf83e;
    PFUMX i19179 (.BLUT(n21497), .ALUT(n21498), .C0(index_i[4]), .Z(n21499));
    LUT4 mux_193_Mux_0_i460_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n460)) /* synthesis lut_function=(A (B+(C (D)+!C !(D)))+!A (B (C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i460_3_lut_4_lut_4_lut.init = 16'hf8cb;
    LUT4 i20241_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n22580)) /* synthesis lut_function=(A (B (C+!(D))+!B !((D)+!C))+!A !(B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20241_3_lut_4_lut_4_lut.init = 16'h81f8;
    LUT4 mux_193_Mux_8_i61_3_lut_rep_431_4_lut_4_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[2]), .D(index_i[3]), .Z(n26391)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A (B (C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_8_i61_3_lut_rep_431_4_lut_4_lut_4_lut.init = 16'he0f8;
    LUT4 mux_193_Mux_8_i251_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n251)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_8_i251_3_lut_4_lut_4_lut_4_lut.init = 16'h07e0;
    LUT4 n924_bdd_3_lut_24424 (.A(n924_adj_2795), .B(n24343), .C(index_i[5]), 
         .Z(n24344)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n924_bdd_3_lut_24424.init = 16'hcaca;
    PFUMX i19185 (.BLUT(n21503), .ALUT(n21504), .C0(index_i[4]), .Z(n21505));
    LUT4 i20240_3_lut_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n22579)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C+!(D))+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20240_3_lut_3_lut_4_lut_4_lut.init = 16'h1f81;
    LUT4 i19106_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n21426)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C))+!A (B (C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19106_3_lut_4_lut_4_lut_4_lut.init = 16'he078;
    LUT4 mux_193_Mux_0_i412_3_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[1]), .D(index_i[3]), .Z(n412)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C (D)))+!A (B (C+!(D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i412_3_lut_4_lut_4_lut.init = 16'hf14c;
    LUT4 i18809_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21129)) /* synthesis lut_function=(A (C)+!A !(B (C)+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18809_3_lut_4_lut_4_lut.init = 16'hb4b5;
    LUT4 i19166_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21486)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(D))+!A (B (D)+!B ((D)+!C))) */ ;
    defparam i19166_3_lut_4_lut_4_lut.init = 16'hd52b;
    LUT4 n262_bdd_3_lut_23564 (.A(n26629), .B(n29199), .C(index_i[3]), 
         .Z(n25251)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n262_bdd_3_lut_23564.init = 16'hcaca;
    PFUMX i18807 (.BLUT(n21125), .ALUT(n21126), .C0(index_i[4]), .Z(n21127));
    LUT4 i11433_2_lut_rep_664 (.A(index_i[0]), .B(index_i[1]), .Z(n26624)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11433_2_lut_rep_664.init = 16'heeee;
    LUT4 mux_193_Mux_1_i684_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n684)) /* synthesis lut_function=(A (B ((D)+!C)+!B !((D)+!C))+!A !(B (C+(D))+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_1_i684_3_lut_4_lut_4_lut.init = 16'h992d;
    PFUMX i23293 (.BLUT(n24968), .ALUT(n24964), .C0(index_i[6]), .Z(n24969));
    LUT4 mux_193_Mux_0_i890_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n890_adj_2796)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)+!C !(D)))+!A !(B (C)+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i890_3_lut_4_lut_4_lut.init = 16'h70ca;
    LUT4 mux_193_Mux_1_i716_3_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[1]), .D(index_i[3]), .Z(n716)) /* synthesis lut_function=(!(A (B (D)+!B !(C))+!A !(B (C (D))+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_1_i716_3_lut_4_lut_4_lut.init = 16'h70a9;
    PFUMX i18810 (.BLUT(n21128), .ALUT(n21129), .C0(index_i[4]), .Z(n21130));
    LUT4 mux_193_Mux_11_i445_3_lut_4_lut_4_lut_4_lut (.A(index_i[3]), .B(index_i[4]), 
         .C(index_i[5]), .D(n26498), .Z(n445)) /* synthesis lut_function=(!(A (B (C))+!A !(B+(C+(D))))) */ ;
    defparam mux_193_Mux_11_i445_3_lut_4_lut_4_lut_4_lut.init = 16'h7f7e;
    LUT4 mux_193_Mux_7_i699_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n699)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C+!(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_7_i699_3_lut_4_lut_4_lut.init = 16'hf07e;
    LUT4 mux_193_Mux_8_i101_3_lut_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n101)) /* synthesis lut_function=(!(A (B (C))+!A (B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_8_i101_3_lut_3_lut_3_lut.init = 16'h3e3e;
    LUT4 mux_193_Mux_13_i511_4_lut_4_lut (.A(n26348), .B(index_i[7]), .C(index_i[8]), 
         .D(n254), .Z(n511)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (B (C+!(D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_13_i511_4_lut_4_lut.init = 16'h1c10;
    PFUMX i24520 (.BLUT(n26826), .ALUT(n26827), .C0(index_i[0]), .Z(n26828));
    PFUMX i19191 (.BLUT(n21509), .ALUT(n21510), .C0(index_i[4]), .Z(n21511));
    LUT4 n21224_bdd_4_lut_24039 (.A(n26596), .B(n763), .C(index_i[5]), 
         .D(index_i[4]), .Z(n24191)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam n21224_bdd_4_lut_24039.init = 16'hcfca;
    LUT4 mux_190_i6_3_lut (.A(quarter_wave_sample_register_i[5]), .B(o_val_pipeline_i_0__15__N_2158[5]), 
         .C(phase_negation_i[1]), .Z(n1086[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam mux_190_i6_3_lut.init = 16'hcaca;
    L6MUX21 i20181 (.D0(n22518), .D1(n22519), .SD(index_i[6]), .Z(n382));
    PFUMX i19194 (.BLUT(n21512), .ALUT(n21513), .C0(index_i[4]), .Z(n21514));
    LUT4 index_i_4__bdd_4_lut_22942 (.A(index_i[4]), .B(n26468), .C(index_i[7]), 
         .D(n26469), .Z(n24368)) /* synthesis lut_function=(A (C+!(D))+!A (B+!(C))) */ ;
    defparam index_i_4__bdd_4_lut_22942.init = 16'he5ef;
    LUT4 mux_190_i5_3_lut (.A(quarter_wave_sample_register_i[4]), .B(o_val_pipeline_i_0__15__N_2158[4]), 
         .C(phase_negation_i[1]), .Z(n1086[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam mux_190_i5_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_0_i795_3_lut_3_lut_rep_786 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29165)) /* synthesis lut_function=(A (B+(C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i795_3_lut_3_lut_rep_786.init = 16'hadad;
    LUT4 i11228_2_lut_rep_442_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n26402)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11228_2_lut_rep_442_3_lut_4_lut.init = 16'hfef0;
    LUT4 mux_193_Mux_6_i860_3_lut_3_lut (.A(n26391), .B(index_i[4]), .C(n844_adj_2797), 
         .Z(n860_adj_2798)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam mux_193_Mux_6_i860_3_lut_3_lut.init = 16'h7474;
    LUT4 i18926_3_lut_3_lut (.A(n26391), .B(index_i[4]), .C(n46), .Z(n21246)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam i18926_3_lut_3_lut.init = 16'h7474;
    LUT4 mux_193_Mux_0_i796_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n796)) /* synthesis lut_function=(A (B (C+(D))+!B (C (D)))+!A !(B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i796_3_lut_4_lut_4_lut.init = 16'hadc0;
    LUT4 n773_bdd_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n24789)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n773_bdd_3_lut_4_lut_4_lut.init = 16'ha5ad;
    LUT4 mux_193_Mux_8_i542_3_lut_4_lut (.A(n26641), .B(index_i[3]), .C(index_i[4]), 
         .D(n526_adj_2799), .Z(n542_adj_2800)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_8_i542_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_193_Mux_2_i142_3_lut_4_lut_4_lut_4_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n142)) /* synthesis lut_function=(!(A (B (D)+!B (C (D)+!C !(D)))+!A (B (D)+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_2_i142_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'h03ec;
    LUT4 mux_193_Mux_0_i581_3_lut_3_lut_rep_812 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29191)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i581_3_lut_3_lut_rep_812.init = 16'hc7c7;
    LUT4 i18944_3_lut_4_lut (.A(n26641), .B(index_i[3]), .C(index_i[4]), 
         .D(n635), .Z(n21264)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18944_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_193_Mux_2_i284_rep_787 (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .Z(n29166)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_2_i284_rep_787.init = 16'h4d4d;
    LUT4 i19141_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21461)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+(D)))+!A !(B (D)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19141_3_lut_4_lut_4_lut.init = 16'h99c7;
    LUT4 i21564_3_lut (.A(n21143), .B(n21144), .C(index_i[4]), .Z(n21145)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21564_3_lut.init = 16'hcaca;
    L6MUX21 i20188 (.D0(n22525), .D1(n22526), .SD(index_i[6]), .Z(n509));
    LUT4 i23201_then_4_lut (.A(index_i[6]), .B(index_i[2]), .C(index_i[5]), 
         .D(index_i[0]), .Z(n26785)) /* synthesis lut_function=(A ((C+!(D))+!B)+!A !(B (C (D))+!B !(C+(D)))) */ ;
    defparam i23201_then_4_lut.init = 16'hb7fe;
    PFUMX i19197 (.BLUT(n21515), .ALUT(n21516), .C0(index_i[4]), .Z(n21517));
    LUT4 mux_193_Mux_7_i262_3_lut_rep_814 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29193)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_7_i262_3_lut_rep_814.init = 16'h3838;
    LUT4 n26609_bdd_2_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[4]), .Z(n27967)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C (D)))+!A (B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n26609_bdd_2_lut_4_lut.init = 16'h3800;
    LUT4 mux_190_i4_3_lut (.A(quarter_wave_sample_register_i[3]), .B(o_val_pipeline_i_0__15__N_2158[3]), 
         .C(phase_negation_i[1]), .Z(n1086[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam mux_190_i4_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_3_i653_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n653)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A !(B (D)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_3_i653_3_lut_4_lut_4_lut.init = 16'h4d99;
    LUT4 mux_190_i3_3_lut (.A(quarter_wave_sample_register_i[2]), .B(o_val_pipeline_i_0__15__N_2158[2]), 
         .C(phase_negation_i[1]), .Z(n1086[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam mux_190_i3_3_lut.init = 16'hcaca;
    LUT4 mux_190_i2_3_lut (.A(quarter_wave_sample_register_i[1]), .B(o_val_pipeline_i_0__15__N_2158[1]), 
         .C(phase_negation_i[1]), .Z(n1086[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam mux_190_i2_3_lut.init = 16'hcaca;
    LUT4 mux_190_i1_3_lut (.A(quarter_wave_sample_register_i[0]), .B(o_val_pipeline_i_0__15__N_2158[0]), 
         .C(phase_negation_i[1]), .Z(n1086[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam mux_190_i1_3_lut.init = 16'hcaca;
    LUT4 i18722_3_lut (.A(n26625), .B(n141), .C(index_i[3]), .Z(n21042)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18722_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_0_i397_3_lut (.A(n29191), .B(n26677), .C(index_i[3]), 
         .Z(n397_adj_2801)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i397_3_lut.init = 16'hcaca;
    LUT4 i23201_else_4_lut (.A(index_i[2]), .Z(n26784)) /* synthesis lut_function=(A) */ ;
    defparam i23201_else_4_lut.init = 16'haaaa;
    LUT4 n77_bdd_3_lut_23730 (.A(n26675), .B(n26676), .C(index_i[3]), 
         .Z(n25412)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n77_bdd_3_lut_23730.init = 16'hacac;
    LUT4 i6421_2_lut (.A(phase_i[0]), .B(phase_i[10]), .Z(index_i_9__N_2107[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i6421_2_lut.init = 16'h6666;
    LUT4 i6422_2_lut (.A(phase_i[9]), .B(phase_i[10]), .Z(index_i_9__N_2107[9])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i6422_2_lut.init = 16'h6666;
    LUT4 i6423_2_lut (.A(phase_i[8]), .B(phase_i[10]), .Z(index_i_9__N_2107[8])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i6423_2_lut.init = 16'h6666;
    LUT4 mux_193_Mux_0_i188_3_lut (.A(n26633), .B(n101), .C(index_i[3]), 
         .Z(n188)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i188_3_lut.init = 16'hcaca;
    LUT4 i6424_2_lut (.A(phase_i[7]), .B(phase_i[10]), .Z(index_i_9__N_2107[7])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i6424_2_lut.init = 16'h6666;
    LUT4 i6425_2_lut (.A(phase_i[6]), .B(phase_i[10]), .Z(index_i_9__N_2107[6])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i6425_2_lut.init = 16'h6666;
    PFUMX i15398 (.BLUT(n17546), .ALUT(n17547), .C0(index_i[4]), .Z(n17548));
    LUT4 i6426_2_lut (.A(phase_i[5]), .B(phase_i[10]), .Z(index_i_9__N_2107[5])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i6426_2_lut.init = 16'h6666;
    LUT4 i6427_2_lut (.A(phase_i[4]), .B(phase_i[10]), .Z(index_i_9__N_2107[4])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i6427_2_lut.init = 16'h6666;
    LUT4 i6428_2_lut (.A(phase_i[3]), .B(phase_i[10]), .Z(index_i_9__N_2107[3])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i6428_2_lut.init = 16'h6666;
    LUT4 i19757_3_lut (.A(n25151), .B(n22583), .C(index_i[6]), .Z(n22096)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19757_3_lut.init = 16'hcaca;
    LUT4 i6417_2_lut (.A(phase_i[2]), .B(phase_i[10]), .Z(index_i_9__N_2107[2])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i6417_2_lut.init = 16'h6666;
    LUT4 i6418_2_lut (.A(phase_i[1]), .B(phase_i[10]), .Z(index_i_9__N_2107[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i6418_2_lut.init = 16'h6666;
    LUT4 n21501_bdd_3_lut (.A(n26630), .B(n26664), .C(index_i[3]), .Z(n25436)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n21501_bdd_3_lut.init = 16'hcaca;
    LUT4 i12112_3_lut_rep_820 (.A(index_i[2]), .B(index_i[1]), .C(index_i[0]), 
         .Z(n29199)) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i12112_3_lut_rep_820.init = 16'hc4c4;
    LUT4 i6816_2_lut (.A(index_i[4]), .B(index_i[5]), .Z(n9197)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i6816_2_lut.init = 16'h8888;
    LUT4 mux_193_Mux_2_i189_3_lut_3_lut_4_lut (.A(index_i[1]), .B(n26596), 
         .C(n173), .D(index_i[4]), .Z(n189_adj_2802)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(C+(D)))) */ ;
    defparam mux_193_Mux_2_i189_3_lut_3_lut_4_lut.init = 16'h77f0;
    LUT4 i19118_3_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[1]), .C(index_i[0]), 
         .D(index_i[3]), .Z(n21438)) /* synthesis lut_function=(A (B (C)+!B !(C+!(D)))+!A (B (C+!(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19118_3_lut_4_lut_4_lut.init = 16'hc3c4;
    PFUMX i18816 (.BLUT(n21134), .ALUT(n21135), .C0(index_i[4]), .Z(n21136));
    LUT4 mux_193_Mux_6_i22_rep_789 (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .Z(n29168)) /* synthesis lut_function=(!(A (C)+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_6_i22_rep_789.init = 16'h4a4a;
    LUT4 i11211_4_lut (.A(n14954), .B(index_i[8]), .C(n765), .D(index_i[7]), 
         .Z(n1022)) /* synthesis lut_function=(A (B+(C (D)))+!A (B+(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11211_4_lut.init = 16'hfcdd;
    LUT4 i1_2_lut (.A(index_i[6]), .B(index_i[7]), .Z(n19553)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i1_2_lut.init = 16'heeee;
    LUT4 mux_193_Mux_5_i491_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n491)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A !(B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_5_i491_3_lut_4_lut_4_lut.init = 16'ha54a;
    LUT4 i11217_2_lut_3_lut_4_lut (.A(index_i[1]), .B(n26596), .C(index_i[5]), 
         .D(index_i[4]), .Z(n508)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;
    defparam i11217_2_lut_3_lut_4_lut.init = 16'hf080;
    LUT4 i21678_3_lut (.A(n26086), .B(n124_adj_2803), .C(index_i[4]), 
         .Z(n22864)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21678_3_lut.init = 16'hcaca;
    LUT4 i21710_3_lut (.A(n620), .B(n13842), .C(index_i[4]), .Z(n21282)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21710_3_lut.init = 16'hcaca;
    LUT4 i11316_3_lut_3_lut_rep_790 (.A(index_i[1]), .B(index_i[0]), .C(index_i[2]), 
         .Z(n29169)) /* synthesis lut_function=(!(A+!((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11316_3_lut_3_lut_rep_790.init = 16'h5151;
    PFUMX i18819 (.BLUT(n21137), .ALUT(n21138), .C0(index_i[4]), .Z(n21139));
    LUT4 i19183_3_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[0]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21503)) /* synthesis lut_function=(!(A ((D)+!C)+!A !(B (C (D))+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19183_3_lut_4_lut_4_lut.init = 16'h51a0;
    LUT4 mux_193_Mux_2_i955_then_4_lut (.A(index_i[4]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n26791)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B (C+!(D))+!B !(C (D)))) */ ;
    defparam mux_193_Mux_2_i955_then_4_lut.init = 16'he95d;
    LUT4 mux_193_Mux_0_i475_3_lut_4_lut (.A(n26551), .B(index_i[1]), .C(index_i[3]), 
         .D(n26499), .Z(n475_adj_2804)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i475_3_lut_4_lut.init = 16'h4f40;
    LUT4 mux_193_Mux_3_i491_3_lut_4_lut (.A(n26551), .B(index_i[1]), .C(index_i[3]), 
         .D(n29179), .Z(n491_adj_2805)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_3_i491_3_lut_4_lut.init = 16'h4f40;
    LUT4 mux_193_Mux_2_i955_else_4_lut (.A(index_i[4]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n26790)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+(D)))+!A !(B (C+!(D))+!B !(C+!(D))))) */ ;
    defparam mux_193_Mux_2_i955_else_4_lut.init = 16'h49c6;
    LUT4 i21713_3_lut (.A(n491_adj_2806), .B(n506_adj_2807), .C(index_i[4]), 
         .Z(n21276)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21713_3_lut.init = 16'hcaca;
    LUT4 i18719_3_lut (.A(n26625), .B(n645), .C(index_i[3]), .Z(n21039)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18719_3_lut.init = 16'hcaca;
    LUT4 i18718_3_lut (.A(n26633), .B(n141), .C(index_i[3]), .Z(n21038)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18718_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_7_i173_3_lut (.A(n26659), .B(n645), .C(index_i[3]), 
         .Z(n173_adj_2808)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_7_i173_3_lut.init = 16'hcaca;
    L6MUX21 i20664 (.D0(n22991), .D1(n22992), .SD(index_i[6]), .Z(n23003));
    L6MUX21 i20665 (.D0(n22993), .D1(n22994), .SD(index_i[6]), .Z(n23004));
    L6MUX21 i20666 (.D0(n22995), .D1(n22996), .SD(index_i[6]), .Z(n23005));
    PFUMX i20667 (.BLUT(n22997), .ALUT(n22998), .C0(index_i[6]), .Z(n23006));
    PFUMX i20686 (.BLUT(n732), .ALUT(n763_adj_2809), .C0(index_i[5]), 
          .Z(n23025));
    LUT4 i19850_3_lut (.A(n22185), .B(n22186), .C(index_i[8]), .Z(n22189)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19850_3_lut.init = 16'hcaca;
    LUT4 i19844_3_lut (.A(n22180), .B(n22181), .C(index_i[8]), .Z(n22183)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19844_3_lut.init = 16'hcaca;
    LUT4 i19843_3_lut (.A(n22178), .B(n22179), .C(index_i[8]), .Z(n22182)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19843_3_lut.init = 16'hcaca;
    L6MUX21 i20688 (.D0(n21517), .D1(n891_adj_2810), .SD(index_i[5]), 
            .Z(n23027));
    LUT4 mux_193_Mux_0_i731_3_lut_4_lut (.A(n26627), .B(index_i[2]), .C(index_i[3]), 
         .D(n26625), .Z(n731)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i731_3_lut_4_lut.init = 16'h4f40;
    LUT4 i19193_3_lut_4_lut (.A(n26627), .B(index_i[2]), .C(index_i[3]), 
         .D(n26673), .Z(n21513)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19193_3_lut_4_lut.init = 16'hf404;
    L6MUX21 i20691 (.D0(n23014), .D1(n23015), .SD(index_i[6]), .Z(n23030));
    L6MUX21 i20693 (.D0(n23018), .D1(n23019), .SD(index_i[6]), .Z(n23032));
    L6MUX21 i20694 (.D0(n23020), .D1(n23021), .SD(index_i[6]), .Z(n23033));
    LUT4 n953_bdd_3_lut_23301_4_lut (.A(n26620), .B(index_i[2]), .C(index_i[3]), 
         .D(n26617), .Z(n24796)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n953_bdd_3_lut_23301_4_lut.init = 16'hf606;
    L6MUX21 i20698 (.D0(n23028), .D1(n23029), .SD(index_i[6]), .Z(n23037));
    L6MUX21 i19755 (.D0(n21247), .D1(n21250), .SD(index_i[6]), .Z(n22094));
    LUT4 i19885_3_lut (.A(n190), .B(n25693), .C(index_i[6]), .Z(n22224)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19885_3_lut.init = 16'hcaca;
    LUT4 i19886_3_lut (.A(n22604), .B(n21271), .C(index_i[6]), .Z(n22225)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19886_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_3_i890_3_lut_4_lut (.A(n26620), .B(index_i[2]), .C(index_i[3]), 
         .D(n325), .Z(n890_adj_2811)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_3_i890_3_lut_4_lut.init = 16'h6f60;
    LUT4 i18806_3_lut_4_lut (.A(n26620), .B(index_i[2]), .C(index_i[3]), 
         .D(n26675), .Z(n21126)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18806_3_lut_4_lut.init = 16'hf606;
    L6MUX21 i19758 (.D0(n21259), .D1(n21262), .SD(index_i[6]), .Z(n22097));
    LUT4 mux_193_Mux_0_i348_3_lut_4_lut (.A(n26620), .B(index_i[2]), .C(index_i[3]), 
         .D(n29169), .Z(n348)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i348_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_193_Mux_1_i700_3_lut_4_lut (.A(n26560), .B(index_i[3]), .C(index_i[4]), 
         .D(n684), .Z(n700_adj_2812)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_1_i700_3_lut_4_lut.init = 16'hefe0;
    L6MUX21 i19759 (.D0(n574), .D1(n21265), .SD(index_i[6]), .Z(n22098));
    L6MUX21 i19760 (.D0(n21268), .D1(n764), .SD(index_i[6]), .Z(n22099));
    LUT4 i18844_3_lut (.A(n24373), .B(n21196), .C(index_i[8]), .Z(n21164)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18844_3_lut.init = 16'hcaca;
    LUT4 i12153_3_lut (.A(index_i[2]), .B(index_i[1]), .C(index_i[0]), 
         .Z(n1001)) /* synthesis lut_function=(A (B)+!A (B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i12153_3_lut.init = 16'hdcdc;
    LUT4 i11179_2_lut_rep_388_3_lut_4_lut (.A(n26402), .B(index_i[4]), .C(index_i[6]), 
         .D(index_i[5]), .Z(n26348)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11179_2_lut_rep_388_3_lut_4_lut.init = 16'hf080;
    L6MUX21 i20320 (.D0(n22643), .D1(n22644), .SD(index_i[6]), .Z(n22659));
    L6MUX21 i20321 (.D0(n22645), .D1(n22646), .SD(index_i[6]), .Z(n22660));
    L6MUX21 i20322 (.D0(n22647), .D1(n22648), .SD(index_i[6]), .Z(n22661));
    L6MUX21 i20323 (.D0(n22649), .D1(n22650), .SD(index_i[6]), .Z(n22662));
    L6MUX21 i20324 (.D0(n22651), .D1(n22652), .SD(index_i[6]), .Z(n22663));
    LUT4 i22259_3_lut (.A(n22102), .B(n22103), .C(index_i[8]), .Z(n22106)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22259_3_lut.init = 16'hcaca;
    L6MUX21 i20326 (.D0(n22655), .D1(n22656), .SD(index_i[6]), .Z(n22665));
    LUT4 i21768_3_lut (.A(n109), .B(n124_adj_2813), .C(index_i[4]), .Z(n21249)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21768_3_lut.init = 16'hcaca;
    PFUMX i20307 (.BLUT(n221), .ALUT(n252_adj_2793), .C0(index_i[5]), 
          .Z(n22646));
    PFUMX i23203 (.BLUT(n24877), .ALUT(n26498), .C0(index_i[4]), .Z(n24878));
    PFUMX i19805 (.BLUT(n22140), .ALUT(n22141), .C0(index_i[6]), .Z(n22144));
    PFUMX i19806 (.BLUT(n22142), .ALUT(n22143), .C0(index_i[6]), .Z(n22145));
    LUT4 i20454_3_lut (.A(n22790), .B(n22791), .C(index_i[8]), .Z(n22793)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20454_3_lut.init = 16'hcaca;
    LUT4 i20453_3_lut (.A(n22788), .B(n22789), .C(index_i[8]), .Z(n22792)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20453_3_lut.init = 16'hcaca;
    LUT4 i22284_3_lut (.A(n574_adj_2814), .B(n637), .C(index_i[6]), .Z(n21197)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22284_3_lut.init = 16'hcaca;
    LUT4 i19163_3_lut_4_lut (.A(index_i[0]), .B(n26641), .C(index_i[3]), 
         .D(n26672), .Z(n21483)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19163_3_lut_4_lut.init = 16'hfb0b;
    L6MUX21 i19832 (.D0(n22156), .D1(n22157), .SD(index_i[6]), .Z(n22171));
    L6MUX21 i19833 (.D0(n22158), .D1(n22159), .SD(index_i[6]), .Z(n22172));
    L6MUX21 i19834 (.D0(n22160), .D1(n22161), .SD(index_i[6]), .Z(n22173));
    L6MUX21 i19835 (.D0(n22162), .D1(n22163), .SD(index_i[6]), .Z(n22174));
    L6MUX21 i19836 (.D0(n22164), .D1(n22165), .SD(index_i[6]), .Z(n22175));
    L6MUX21 i20761 (.D0(n23092), .D1(n23093), .SD(index_i[6]), .Z(n23100));
    L6MUX21 i20762 (.D0(n23094), .D1(n23095), .SD(index_i[6]), .Z(n23101));
    L6MUX21 i20763 (.D0(n23096), .D1(n23097), .SD(index_i[6]), .Z(n23102));
    L6MUX21 i20764 (.D0(n23098), .D1(n23099), .SD(index_i[6]), .Z(n23103));
    LUT4 mux_193_Mux_3_i30_3_lut_3_lut_4_lut_3_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n30)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_3_i30_3_lut_3_lut_4_lut_3_lut_4_lut.init = 16'hfe11;
    LUT4 i20704_3_lut (.A(n23040), .B(n23041), .C(index_i[8]), .Z(n23043)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20704_3_lut.init = 16'hcaca;
    LUT4 i20703_3_lut (.A(n23038), .B(n23039), .C(index_i[8]), .Z(n23042)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20703_3_lut.init = 16'hcaca;
    LUT4 n24199_bdd_3_lut_25916 (.A(n24199), .B(n24192), .C(index_i[7]), 
         .Z(n24200)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n24199_bdd_3_lut_25916.init = 16'hcaca;
    PFUMX i18874 (.BLUT(n318), .ALUT(n381), .C0(index_i[6]), .Z(n21194));
    L6MUX21 i20403 (.D0(n22726), .D1(n22727), .SD(index_i[6]), .Z(n22742));
    L6MUX21 i20404 (.D0(n22728), .D1(n22729), .SD(index_i[6]), .Z(n22743));
    LUT4 i19444_3_lut (.A(n26679), .B(n26621), .C(index_i[3]), .Z(n21764)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19444_3_lut.init = 16'hcaca;
    L6MUX21 i20405 (.D0(n22730), .D1(n22731), .SD(index_i[6]), .Z(n22744));
    PFUMX mux_193_Mux_1_i636 (.BLUT(n620_adj_2815), .ALUT(n635_adj_2816), 
          .C0(index_i[4]), .Z(n636)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    PFUMX i20407 (.BLUT(n22734), .ALUT(n22735), .C0(index_i[6]), .Z(n22746));
    L6MUX21 i19884 (.D0(n22590), .D1(n22597), .SD(index_i[6]), .Z(n22223));
    LUT4 index_i_2__bdd_4_lut_25880 (.A(index_i[2]), .B(index_i[0]), .C(index_i[4]), 
         .D(index_i[1]), .Z(n27963)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((C (D))+!B))) */ ;
    defparam index_i_2__bdd_4_lut_25880.init = 16'h0cec;
    L6MUX21 i20408 (.D0(n22736), .D1(n22737), .SD(index_i[6]), .Z(n22747));
    L6MUX21 i20409 (.D0(n22738), .D1(n22739), .SD(index_i[6]), .Z(n22748));
    PFUMX i20410 (.BLUT(n22740), .ALUT(n22741), .C0(index_i[6]), .Z(n22749));
    LUT4 index_i_2__bdd_3_lut_25881 (.A(index_i[2]), .B(index_i[0]), .C(index_i[4]), 
         .Z(n27964)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B (C)+!B !(C)))) */ ;
    defparam index_i_2__bdd_3_lut_25881.init = 16'h6969;
    L6MUX21 i19887 (.D0(n21274), .D1(n21277), .SD(index_i[6]), .Z(n22226));
    L6MUX21 i19888 (.D0(n21280), .D1(n21283), .SD(index_i[6]), .Z(n22227));
    L6MUX21 i19889 (.D0(n21286), .D1(n21289), .SD(index_i[6]), .Z(n22228));
    PFUMX i19890 (.BLUT(n21292), .ALUT(n892_adj_2817), .C0(index_i[6]), 
          .Z(n22229));
    LUT4 i18839_3_lut_4_lut (.A(n26616), .B(index_i[2]), .C(index_i[3]), 
         .D(n26677), .Z(n21159)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18839_3_lut_4_lut.init = 16'h6f60;
    PFUMX i20437 (.BLUT(n797), .ALUT(n828), .C0(index_i[5]), .Z(n22776));
    L6MUX21 i20441 (.D0(n22764), .D1(n22765), .SD(index_i[6]), .Z(n22780));
    L6MUX21 i20442 (.D0(n22766), .D1(n22767), .SD(index_i[6]), .Z(n22781));
    LUT4 mux_193_Mux_6_i285_3_lut_4_lut (.A(n26616), .B(index_i[2]), .C(index_i[3]), 
         .D(n26675), .Z(n285)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_6_i285_3_lut_4_lut.init = 16'hf606;
    LUT4 n26609_bdd_3_lut_25445 (.A(n26499), .B(n29179), .C(index_i[4]), 
         .Z(n27966)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n26609_bdd_3_lut_25445.init = 16'hcaca;
    L6MUX21 i20443 (.D0(n22768), .D1(n22769), .SD(index_i[6]), .Z(n22782));
    L6MUX21 i20444 (.D0(n22770), .D1(n22771), .SD(index_i[6]), .Z(n22783));
    L6MUX21 i20445 (.D0(n22772), .D1(n22773), .SD(index_i[6]), .Z(n22784));
    LUT4 mux_193_Mux_3_i460_3_lut_4_lut (.A(n26616), .B(index_i[2]), .C(index_i[3]), 
         .D(n26681), .Z(n460_adj_2818)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_3_i460_3_lut_4_lut.init = 16'h6f60;
    LUT4 i19154_3_lut_4_lut (.A(n26616), .B(index_i[2]), .C(index_i[3]), 
         .D(n26661), .Z(n21474)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19154_3_lut_4_lut.init = 16'hf606;
    PFUMX mux_193_Mux_2_i891 (.BLUT(n875), .ALUT(n890), .C0(index_i[4]), 
          .Z(n891_adj_2819)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 i15443_4_lut (.A(index_i[0]), .B(index_i[4]), .C(index_i[1]), 
         .D(n26575), .Z(n286)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i15443_4_lut.init = 16'hccc8;
    L6MUX21 i20448 (.D0(n22778), .D1(n22779), .SD(index_i[6]), .Z(n22787));
    PFUMX mux_193_Mux_2_i860 (.BLUT(n844), .ALUT(n859), .C0(index_i[4]), 
          .Z(n860_adj_2820)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 mux_193_Mux_0_i684_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n684_adj_2821)) /* synthesis lut_function=(!(A ((D)+!B)+!A !(B (D)+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i684_3_lut_4_lut_4_lut.init = 16'h5498;
    LUT4 i21324_3_lut (.A(n21446), .B(n26764), .C(index_i[4]), .Z(n21448)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21324_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_3_i924_3_lut (.A(n908), .B(index_i[0]), .C(index_i[4]), 
         .Z(n924_adj_2822)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_3_i924_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_3_i891_3_lut (.A(n541_adj_2823), .B(n890_adj_2811), 
         .C(index_i[4]), .Z(n891_adj_2824)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_3_i891_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_3_i669_3_lut (.A(n653), .B(n668), .C(index_i[4]), 
         .Z(n669)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_3_i669_3_lut.init = 16'hcaca;
    LUT4 i9480_4_lut (.A(n26639), .B(n26499), .C(index_i[3]), .D(index_i[4]), 
         .Z(n11926)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B ((D)+!C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9480_4_lut.init = 16'h3afa;
    LUT4 i21334_3_lut (.A(n21434), .B(n21435), .C(index_i[4]), .Z(n21436)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21334_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_3_i476_3_lut (.A(n460_adj_2818), .B(n285), .C(index_i[4]), 
         .Z(n476_adj_2825)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_3_i476_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_3_i413_3_lut (.A(n397_adj_2826), .B(n26577), .C(index_i[4]), 
         .Z(n413)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_3_i413_3_lut.init = 16'hcaca;
    PFUMX mux_193_Mux_3_i763 (.BLUT(n747_adj_2827), .ALUT(n762), .C0(index_i[4]), 
          .Z(n763_adj_2828)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 mux_193_Mux_3_i286_4_lut (.A(n93_adj_2829), .B(index_i[2]), .C(index_i[4]), 
         .D(n14747), .Z(n286_adj_2830)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_3_i286_4_lut.init = 16'h3aca;
    LUT4 mux_193_Mux_9_i763_3_lut_4_lut (.A(n26627), .B(n26575), .C(index_i[4]), 
         .D(n26467), .Z(n763)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;
    defparam mux_193_Mux_9_i763_3_lut_4_lut.init = 16'hf101;
    LUT4 mux_193_Mux_8_i763_3_lut_4_lut (.A(n26627), .B(n26575), .C(index_i[4]), 
         .D(n26467), .Z(n14970)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam mux_193_Mux_8_i763_3_lut_4_lut.init = 16'hfe0e;
    LUT4 mux_193_Mux_3_i158_3_lut (.A(n142_adj_2831), .B(n26413), .C(index_i[4]), 
         .Z(n158)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_3_i158_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_3_i125_3_lut (.A(n46), .B(n526_adj_2832), .C(index_i[4]), 
         .Z(n125)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_3_i125_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_3_i31_3_lut (.A(n781), .B(n30), .C(index_i[4]), .Z(n31)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_3_i31_3_lut.init = 16'hcaca;
    LUT4 i20524_3_lut_3_lut_4_lut (.A(n26499), .B(index_i[3]), .C(n93_adj_2833), 
         .D(index_i[4]), .Z(n22863)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20524_3_lut_3_lut_4_lut.init = 16'hf077;
    PFUMX i18831 (.BLUT(n21149), .ALUT(n21150), .C0(index_i[4]), .Z(n21151));
    LUT4 n627_bdd_3_lut_23952 (.A(n26617), .B(n26676), .C(index_i[3]), 
         .Z(n25668)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n627_bdd_3_lut_23952.init = 16'hcaca;
    PFUMX i20738 (.BLUT(n557), .ALUT(n572), .C0(index_i[4]), .Z(n23077));
    LUT4 i22700_then_4_lut (.A(index_i[0]), .B(index_i[4]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n26797)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)+!C !(D))+!B (C (D)))) */ ;
    defparam i22700_then_4_lut.init = 16'hda0e;
    LUT4 n262_bdd_3_lut_23958 (.A(n26679), .B(n29199), .C(index_i[3]), 
         .Z(n25677)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n262_bdd_3_lut_23958.init = 16'hcaca;
    LUT4 mux_193_Mux_8_i732_3_lut (.A(index_i[3]), .B(n14970), .C(index_i[5]), 
         .Z(n732_adj_2834)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_8_i732_3_lut.init = 16'h3a3a;
    PFUMX i20739 (.BLUT(n589), .ALUT(n604), .C0(index_i[4]), .Z(n23078));
    LUT4 n62_bdd_3_lut_25655 (.A(n62_adj_2788), .B(n125_adj_2835), .C(index_i[6]), 
         .Z(n28204)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n62_bdd_3_lut_25655.init = 16'hcaca;
    LUT4 n22149_bdd_4_lut_25652 (.A(n252_adj_2836), .B(n26468), .C(index_i[4]), 
         .D(index_i[5]), .Z(n28202)) /* synthesis lut_function=(A (B (D)+!B ((D)+!C))+!A !(B+(C+(D)))) */ ;
    defparam n22149_bdd_4_lut_25652.init = 16'haa03;
    LUT4 n627_bdd_3_lut_23987 (.A(n26617), .B(n588), .C(index_i[3]), .Z(n25679)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n627_bdd_3_lut_23987.init = 16'hacac;
    LUT4 n62_bdd_4_lut_25656 (.A(n26575), .B(n26469), .C(index_i[6]), 
         .D(index_i[4]), .Z(n28205)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C+(D)))+!A (B ((D)+!C)+!B !(C)))) */ ;
    defparam n62_bdd_4_lut_25656.init = 16'h3af0;
    LUT4 i22700_else_4_lut (.A(index_i[0]), .B(index_i[4]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n26796)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C))+!A (B (C)+!B (C+(D)))) */ ;
    defparam i22700_else_4_lut.init = 16'hf178;
    LUT4 i21362_3_lut (.A(n21038), .B(n21039), .C(index_i[4]), .Z(n21040)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i21362_3_lut.init = 16'hcaca;
    LUT4 n21042_bdd_3_lut (.A(n26659), .B(n26611), .C(index_i[3]), .Z(n25689)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n21042_bdd_3_lut.init = 16'hcaca;
    LUT4 i20402_4_lut (.A(n21427), .B(n1002), .C(index_i[5]), .D(index_i[4]), 
         .Z(n22741)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;
    defparam i20402_4_lut.init = 16'hfaca;
    LUT4 mux_193_Mux_4_i860_3_lut (.A(n506_adj_2790), .B(n24792), .C(index_i[4]), 
         .Z(n860_adj_2837)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_4_i860_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_0_i908_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n908_adj_2838)) /* synthesis lut_function=(!(A (B (C (D))+!B !(D))+!A (B+((D)+!C)))) */ ;
    defparam mux_193_Mux_0_i908_3_lut_4_lut_4_lut.init = 16'h2a98;
    LUT4 i18959_3_lut_4_lut_4_lut_4_lut (.A(n26624), .B(index_i[2]), .C(index_i[3]), 
         .D(index_i[4]), .Z(n21279)) /* synthesis lut_function=(A (B)+!A (B (C (D))+!B !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18959_3_lut_4_lut_4_lut_4_lut.init = 16'hc999;
    LUT4 i18824_3_lut_4_lut (.A(n26624), .B(index_i[2]), .C(index_i[3]), 
         .D(n29193), .Z(n21144)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18824_3_lut_4_lut.init = 16'h6f60;
    LUT4 index_i_1__bdd_4_lut_25677 (.A(index_i[1]), .B(index_i[3]), .C(index_i[0]), 
         .D(index_i[2]), .Z(n28346)) /* synthesis lut_function=(A (B (C+(D))+!B (C (D)))+!A !(B (C)+!B !(C+(D)))) */ ;
    defparam index_i_1__bdd_4_lut_25677.init = 16'hbd94;
    LUT4 n28346_bdd_3_lut (.A(n28346), .B(index_i[1]), .C(index_i[4]), 
         .Z(n28347)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n28346_bdd_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_7_i475_3_lut_4_lut (.A(n26624), .B(index_i[2]), .C(index_i[3]), 
         .D(n29191), .Z(n475_adj_2839)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_7_i475_3_lut_4_lut.init = 16'h9f90;
    LUT4 i21383_3_lut (.A(n21416), .B(n21417), .C(index_i[4]), .Z(n21418)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21383_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_7_i653_3_lut_4_lut (.A(n26624), .B(index_i[2]), .C(index_i[3]), 
         .D(n70), .Z(n653_adj_2840)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_7_i653_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_193_Mux_2_i684_3_lut_4_lut (.A(n26624), .B(index_i[2]), .C(index_i[3]), 
         .D(n29169), .Z(n684_adj_2841)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_2_i684_3_lut_4_lut.init = 16'h6f60;
    LUT4 i18961_4_lut_4_lut_4_lut (.A(n26624), .B(index_i[2]), .C(index_i[4]), 
         .D(index_i[3]), .Z(n21281)) /* synthesis lut_function=(A (B)+!A !(B (C+(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18961_4_lut_4_lut_4_lut.init = 16'h999c;
    LUT4 i21385_3_lut (.A(n21413), .B(n21414), .C(index_i[4]), .Z(n21415)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21385_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_4_i700_3_lut (.A(n684_adj_2842), .B(index_i[1]), .C(index_i[4]), 
         .Z(n700_adj_2843)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_4_i700_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_4_i669_3_lut (.A(n781), .B(n668_adj_2844), .C(index_i[4]), 
         .Z(n669_adj_2845)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_4_i669_3_lut.init = 16'hcaca;
    PFUMX i24512 (.BLUT(n26814), .ALUT(n26815), .C0(index_i[8]), .Z(n26816));
    LUT4 mux_193_Mux_3_i221_3_lut_4_lut (.A(n26499), .B(index_i[3]), .C(index_i[4]), 
         .D(n26468), .Z(n221_adj_2846)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_3_i221_3_lut_4_lut.init = 16'h08f8;
    PFUMX i18927 (.BLUT(n21245), .ALUT(n21246), .C0(index_i[5]), .Z(n21247));
    LUT4 mux_193_Mux_4_i542_3_lut (.A(n526_adj_2832), .B(n506), .C(index_i[4]), 
         .Z(n542)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_4_i542_3_lut.init = 16'hcaca;
    LUT4 i20396_4_lut (.A(n26474), .B(n26760), .C(index_i[5]), .D(index_i[4]), 
         .Z(n22735)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam i20396_4_lut.init = 16'hc5ca;
    LUT4 i20523_3_lut_4_lut (.A(n26499), .B(index_i[3]), .C(index_i[4]), 
         .D(n46_adj_2847), .Z(n22862)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20523_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_193_Mux_3_i1018_3_lut_4_lut (.A(index_i[1]), .B(n26575), .C(index_i[4]), 
         .D(n19598), .Z(n1018)) /* synthesis lut_function=(A (C+!(D))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_3_i1018_3_lut_4_lut.init = 16'he0ef;
    PFUMX i20740 (.BLUT(n620_adj_2848), .ALUT(n635_adj_2849), .C0(index_i[4]), 
          .Z(n23079));
    LUT4 mux_193_Mux_2_i700_3_lut_4_lut (.A(index_i[1]), .B(n26575), .C(index_i[4]), 
         .D(n684_adj_2841), .Z(n700_adj_2850)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_2_i700_3_lut_4_lut.init = 16'hefe0;
    LUT4 mux_193_Mux_4_i286_3_lut (.A(n270), .B(n15_adj_2851), .C(index_i[4]), 
         .Z(n286_adj_2852)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_4_i286_3_lut.init = 16'hcaca;
    LUT4 i19804_3_lut_4_lut_4_lut (.A(n26459), .B(index_i[4]), .C(index_i[5]), 
         .D(n26441), .Z(n22143)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C)+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19804_3_lut_4_lut_4_lut.init = 16'h0434;
    LUT4 mux_193_Mux_4_i94_3_lut (.A(n61), .B(n26576), .C(index_i[4]), 
         .Z(n94)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_4_i94_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_8_i460_3_lut_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n460_adj_2853)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_8_i460_3_lut_3_lut_3_lut_4_lut.init = 16'hf10f;
    LUT4 mux_193_Mux_8_i892_3_lut_4_lut (.A(n26459), .B(index_i[4]), .C(index_i[5]), 
         .D(n860), .Z(n892_adj_2854)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_8_i892_3_lut_4_lut.init = 16'h4f40;
    PFUMX i18930 (.BLUT(n21248), .ALUT(n21249), .C0(index_i[5]), .Z(n21250));
    LUT4 mux_190_i16_3_lut (.A(\quarter_wave_sample_register_q[15] ), .B(o_val_pipeline_i_0__15__N_2158[15]), 
         .C(phase_negation_i[1]), .Z(n1086[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam mux_190_i16_3_lut.init = 16'hcaca;
    LUT4 i21413_3_lut (.A(n716_adj_2855), .B(n731_adj_2856), .C(index_i[4]), 
         .Z(n732_adj_2857)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21413_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_2_i669_3_lut (.A(n653_adj_2858), .B(n475_adj_2859), 
         .C(index_i[4]), .Z(n669_adj_2860)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_2_i669_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_10_i125_3_lut_4_lut_4_lut (.A(n26639), .B(index_i[3]), 
         .C(index_i[4]), .D(n26499), .Z(n125_adj_2835)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B (C (D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_10_i125_3_lut_4_lut_4_lut.init = 16'h3efe;
    LUT4 n699_bdd_3_lut_22824_4_lut (.A(n26639), .B(index_i[3]), .C(index_i[4]), 
         .D(n124_adj_2861), .Z(n24425)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n699_bdd_3_lut_22824_4_lut.init = 16'hf101;
    LUT4 mux_193_Mux_2_i605_3_lut (.A(n142_adj_2831), .B(n604_adj_2862), 
         .C(index_i[4]), .Z(n605)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_2_i605_3_lut.init = 16'hcaca;
    PFUMX i20741 (.BLUT(n653_adj_2863), .ALUT(n668_adj_2864), .C0(index_i[4]), 
          .Z(n23080));
    LUT4 i21418_3_lut (.A(n26769), .B(n21465), .C(index_i[4]), .Z(n21466)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21418_3_lut.init = 16'hcaca;
    LUT4 i20175_3_lut_4_lut (.A(n26639), .B(index_i[3]), .C(index_i[4]), 
         .D(n285_adj_2865), .Z(n22514)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20175_3_lut_4_lut.init = 16'hfe0e;
    LUT4 mux_193_Mux_4_i573_3_lut_4_lut_4_lut_4_lut (.A(n26639), .B(index_i[3]), 
         .C(n26498), .D(index_i[4]), .Z(n573)) /* synthesis lut_function=(!(A (B (D)+!B ((D)+!C))+!A (B (D)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_4_i573_3_lut_4_lut_4_lut_4_lut.init = 16'h11fc;
    PFUMX i20742 (.BLUT(n684_adj_2821), .ALUT(n699_adj_2866), .C0(index_i[4]), 
          .Z(n23081));
    LUT4 i21420_3_lut (.A(n21461), .B(n21462), .C(index_i[4]), .Z(n21463)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21420_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_3_i573_3_lut_3_lut_4_lut (.A(n26639), .B(index_i[3]), 
         .C(n460_adj_2853), .D(index_i[4]), .Z(n573_adj_2867)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_3_i573_3_lut_3_lut_4_lut.init = 16'h11f0;
    LUT4 mux_193_Mux_2_i573_3_lut_3_lut_4_lut (.A(n26639), .B(index_i[3]), 
         .C(n557_adj_2868), .D(index_i[4]), .Z(n573_adj_2869)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_2_i573_3_lut_3_lut_4_lut.init = 16'h11f0;
    LUT4 i19810_4_lut_4_lut (.A(n26402), .B(n26510), .C(index_i[5]), .D(index_i[4]), 
         .Z(n22149)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C+(D))+!B !(C (D)+!C !(D)))) */ ;
    defparam i19810_4_lut_4_lut.init = 16'hcf50;
    LUT4 mux_193_Mux_2_i413_3_lut (.A(n397_adj_2870), .B(n954), .C(index_i[4]), 
         .Z(n413_adj_2871)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_2_i413_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_2_i317_3_lut (.A(n668), .B(n316_adj_2872), .C(index_i[4]), 
         .Z(n317_adj_2873)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_2_i317_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_2_i286_3_lut (.A(n270_adj_2874), .B(n653), .C(index_i[4]), 
         .Z(n286_adj_2875)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_2_i286_3_lut.init = 16'hcaca;
    PFUMX i18834 (.BLUT(n21152), .ALUT(n21153), .C0(index_i[4]), .Z(n21154));
    LUT4 i21433_3_lut (.A(n142), .B(n13969), .C(index_i[4]), .Z(n158_adj_2876)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21433_3_lut.init = 16'hcaca;
    LUT4 i19196_3_lut_4_lut (.A(n26624), .B(index_i[2]), .C(index_i[3]), 
         .D(n26660), .Z(n21516)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19196_3_lut_4_lut.init = 16'hdfd0;
    LUT4 mux_193_Mux_4_i62_4_lut (.A(n26640), .B(n61), .C(index_i[4]), 
         .D(index_i[3]), .Z(n62_adj_2877)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_4_i62_4_lut.init = 16'hc5ca;
    PFUMX i18939 (.BLUT(n21257), .ALUT(n21258), .C0(index_i[5]), .Z(n21259));
    PFUMX i20743 (.BLUT(n716_adj_2878), .ALUT(n731), .C0(index_i[4]), 
          .Z(n23082));
    LUT4 i18841_3_lut_4_lut (.A(index_i[0]), .B(n26639), .C(index_i[3]), 
         .D(n26681), .Z(n21161)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A ((D)+!C)) */ ;
    defparam i18841_3_lut_4_lut.init = 16'hfd0d;
    PFUMX mux_193_Mux_5_i732 (.BLUT(n11912), .ALUT(n731_adj_2879), .C0(index_i[4]), 
          .Z(n732_adj_2880)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 mux_193_Mux_4_i31_4_lut (.A(n15_adj_2851), .B(n26454), .C(index_i[4]), 
         .D(index_i[3]), .Z(n31_adj_2881)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_4_i31_4_lut.init = 16'h3aca;
    PFUMX i18942 (.BLUT(n21260), .ALUT(n21261), .C0(index_i[5]), .Z(n21262));
    PFUMX i18945 (.BLUT(n21263), .ALUT(n21264), .C0(index_i[5]), .Z(n21265));
    PFUMX i20744 (.BLUT(n747_adj_2882), .ALUT(n762_adj_2883), .C0(index_i[4]), 
          .Z(n23083));
    PFUMX i18948 (.BLUT(n21266), .ALUT(n21267), .C0(index_i[5]), .Z(n21268));
    PFUMX i18951 (.BLUT(n21269), .ALUT(n21270), .C0(index_i[5]), .Z(n21271));
    PFUMX i18837 (.BLUT(n21155), .ALUT(n21156), .C0(index_i[4]), .Z(n21157));
    LUT4 index_i_6__bdd_4_lut_26001 (.A(index_i[6]), .B(index_i[5]), .C(index_i[1]), 
         .D(index_i[0]), .Z(n28801)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C))+!A (B (C)+!B !(C)))) */ ;
    defparam index_i_6__bdd_4_lut_26001.init = 16'h3cbc;
    PFUMX i20745 (.BLUT(n781_adj_2884), .ALUT(n796), .C0(index_i[4]), 
          .Z(n23084));
    LUT4 n22665_bdd_3_lut_24063 (.A(n22665), .B(n24345), .C(index_i[7]), 
         .Z(n25814)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n22665_bdd_3_lut_24063.init = 16'hcaca;
    LUT4 n22665_bdd_3_lut_25579 (.A(n22663), .B(n22664), .C(index_i[7]), 
         .Z(n25815)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n22665_bdd_3_lut_25579.init = 16'hcaca;
    LUT4 n22668_bdd_3_lut (.A(n22659), .B(n22660), .C(index_i[7]), .Z(n25817)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n22668_bdd_3_lut.init = 16'hcaca;
    LUT4 n25817_bdd_3_lut (.A(n25817), .B(n22668), .C(index_i[8]), .Z(n25818)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n25817_bdd_3_lut.init = 16'hcaca;
    LUT4 n25818_bdd_3_lut (.A(n25818), .B(n25816), .C(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2127[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n25818_bdd_3_lut.init = 16'hcaca;
    LUT4 index_i_6__bdd_1_lut (.A(index_i[5]), .Z(n28800)) /* synthesis lut_function=(!(A)) */ ;
    defparam index_i_6__bdd_1_lut.init = 16'h5555;
    LUT4 index_i_5__bdd_3_lut (.A(index_i[5]), .B(n28802), .C(index_i[3]), 
         .Z(n28803)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam index_i_5__bdd_3_lut.init = 16'hcaca;
    LUT4 n26624_bdd_3_lut (.A(n26508), .B(index_i[6]), .C(index_i[5]), 
         .Z(n28804)) /* synthesis lut_function=(!(A (B)+!A (C))) */ ;
    defparam n26624_bdd_3_lut.init = 16'h2727;
    LUT4 n26624_bdd_4_lut (.A(n26624), .B(index_i[6]), .C(index_i[2]), 
         .D(index_i[5]), .Z(n28805)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A !(B (C+(D))+!B (D)))) */ ;
    defparam n26624_bdd_4_lut.init = 16'h5fe0;
    PFUMX i20746 (.BLUT(n812), .ALUT(n11820), .C0(index_i[4]), .Z(n23085));
    LUT4 n28806_bdd_3_lut (.A(n28806), .B(n28803), .C(index_i[4]), .Z(n28807)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n28806_bdd_3_lut.init = 16'hcaca;
    PFUMX i20748 (.BLUT(n875_adj_2885), .ALUT(n890_adj_2796), .C0(index_i[4]), 
          .Z(n23087));
    PFUMX i20749 (.BLUT(n908_adj_2838), .ALUT(n923), .C0(index_i[4]), 
          .Z(n23088));
    LUT4 n25844_bdd_3_lut (.A(n28207), .B(n22146), .C(index_i[8]), .Z(n25845)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n25844_bdd_3_lut.init = 16'hcaca;
    LUT4 n21197_bdd_3_lut (.A(n26351), .B(n701), .C(index_i[6]), .Z(n25841)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n21197_bdd_3_lut.init = 16'hacac;
    PFUMX i20750 (.BLUT(n939), .ALUT(n954_adj_2886), .C0(index_i[4]), 
          .Z(n23089));
    PFUMX i20751 (.BLUT(n971), .ALUT(n986_adj_2887), .C0(index_i[4]), 
          .Z(n23090));
    LUT4 i9463_2_lut_rep_640 (.A(index_i[3]), .B(index_i[4]), .Z(n26600)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9463_2_lut_rep_640.init = 16'heeee;
    LUT4 i11183_2_lut_rep_538_3_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .Z(n26498)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11183_2_lut_rep_538_3_lut.init = 16'he0e0;
    LUT4 mux_193_Mux_5_i891_3_lut (.A(n875_adj_2888), .B(n379_adj_2889), 
         .C(index_i[4]), .Z(n891_adj_2890)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_5_i891_3_lut.init = 16'hcaca;
    PFUMX i20752 (.BLUT(n1002_adj_2891), .ALUT(n1017), .C0(index_i[4]), 
          .Z(n23091));
    LUT4 mux_193_Mux_5_i860_3_lut (.A(n15), .B(n859_adj_2892), .C(index_i[4]), 
         .Z(n860_adj_2893)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_5_i860_3_lut.init = 16'hcaca;
    PFUMX i18954 (.BLUT(n21272), .ALUT(n21273), .C0(index_i[5]), .Z(n21274));
    LUT4 i21489_3_lut (.A(n21161), .B(n21162), .C(index_i[4]), .Z(n21163)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21489_3_lut.init = 16'hcaca;
    PFUMX i18957 (.BLUT(n21275), .ALUT(n21276), .C0(index_i[5]), .Z(n21277));
    PFUMX i18840 (.BLUT(n21158), .ALUT(n21159), .C0(index_i[4]), .Z(n21160));
    PFUMX i18960 (.BLUT(n21278), .ALUT(n21279), .C0(index_i[5]), .Z(n21280));
    PFUMX i18963 (.BLUT(n21281), .ALUT(n21282), .C0(index_i[5]), .Z(n21283));
    LUT4 i11241_3_lut_4_lut (.A(n26596), .B(index_i[4]), .C(index_i[5]), 
         .D(n26624), .Z(n892)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11241_3_lut_4_lut.init = 16'hf8f0;
    LUT4 mux_193_Mux_5_i636_4_lut (.A(n157), .B(n26480), .C(index_i[4]), 
         .D(index_i[3]), .Z(n636_adj_2894)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_5_i636_4_lut.init = 16'h3aca;
    PFUMX i23141 (.BLUT(n24809), .ALUT(n26586), .C0(index_i[5]), .Z(n24810));
    PFUMX i18966 (.BLUT(n21284), .ALUT(n21285), .C0(index_i[5]), .Z(n21286));
    LUT4 i9460_3_lut_4_lut (.A(n26665), .B(index_i[2]), .C(n26638), .D(n26682), 
         .Z(n444)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9460_3_lut_4_lut.init = 16'h6f60;
    LUT4 i21494_3_lut (.A(n17549), .B(n17550), .C(index_i[4]), .Z(n17551)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21494_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_5_i507_3_lut (.A(n491), .B(n506_adj_2790), .C(index_i[4]), 
         .Z(n507)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_5_i507_3_lut.init = 16'hcaca;
    PFUMX i18969 (.BLUT(n21287), .ALUT(n21288), .C0(index_i[5]), .Z(n21289));
    LUT4 mux_193_Mux_5_i476_3_lut (.A(n460_adj_2895), .B(n475), .C(index_i[4]), 
         .Z(n476_adj_2896)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_5_i476_3_lut.init = 16'hcaca;
    PFUMX i23139 (.BLUT(n26670), .ALUT(n24807), .C0(index_i[2]), .Z(n24808));
    LUT4 mux_193_Mux_4_i747_3_lut_4_lut (.A(n26665), .B(index_i[2]), .C(index_i[3]), 
         .D(n26677), .Z(n747_adj_2897)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_4_i747_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_193_Mux_5_i413_3_lut (.A(n397), .B(n251_adj_2898), .C(index_i[4]), 
         .Z(n413_adj_2899)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_5_i413_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_6_i251_3_lut_4_lut (.A(n26665), .B(index_i[2]), .C(index_i[3]), 
         .D(n26682), .Z(n251_adj_2898)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_6_i251_3_lut_4_lut.init = 16'hf606;
    LUT4 n773_bdd_3_lut_23117_4_lut (.A(n26613), .B(index_i[2]), .C(n26672), 
         .D(index_i[3]), .Z(n24788)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n773_bdd_3_lut_23117_4_lut.init = 16'hf066;
    LUT4 mux_193_Mux_3_i668_3_lut_4_lut (.A(n26613), .B(index_i[2]), .C(index_i[3]), 
         .D(n26669), .Z(n668)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_3_i668_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_193_Mux_4_i763_3_lut_4_lut (.A(n26613), .B(index_i[2]), .C(index_i[4]), 
         .D(n747_adj_2897), .Z(n763_adj_2900)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_4_i763_3_lut_4_lut.init = 16'h6f60;
    L6MUX21 i23137 (.D0(n24805), .D1(n24802), .SD(index_i[5]), .Z(n24806));
    LUT4 i15432_3_lut (.A(n17580), .B(n17581), .C(index_i[4]), .Z(n17582)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15432_3_lut.init = 16'hcaca;
    LUT4 i19117_3_lut_3_lut_4_lut (.A(index_i[2]), .B(n26627), .C(n645), 
         .D(index_i[3]), .Z(n21437)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (B (C (D))+!B (C+!(D)))) */ ;
    defparam i19117_3_lut_3_lut_4_lut.init = 16'hf099;
    LUT4 mux_193_Mux_5_i125_3_lut (.A(n109_adj_2901), .B(n124), .C(index_i[4]), 
         .Z(n125_adj_2902)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_5_i125_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_5_i94_3_lut (.A(n653_adj_2903), .B(n635_adj_2904), 
         .C(index_i[4]), .Z(n94_adj_2905)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_5_i94_3_lut.init = 16'hcaca;
    LUT4 n476_bdd_3_lut_23321_3_lut_4_lut (.A(index_i[2]), .B(n26627), .C(n491_adj_2906), 
         .D(index_i[4]), .Z(n24997)) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))+!A !(B ((D)+!C)+!B !(C+(D)))) */ ;
    defparam n476_bdd_3_lut_23321_3_lut_4_lut.init = 16'h99f0;
    LUT4 mux_193_Mux_5_i31_3_lut (.A(n15), .B(n30_adj_2907), .C(index_i[4]), 
         .Z(n31_adj_2908)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_5_i31_3_lut.init = 16'hcaca;
    LUT4 i18823_3_lut_3_lut_4_lut (.A(index_i[2]), .B(n26627), .C(n26611), 
         .D(index_i[3]), .Z(n21143)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (B (C (D))+!B (C+!(D)))) */ ;
    defparam i18823_3_lut_3_lut_4_lut.init = 16'hf099;
    LUT4 mux_193_Mux_7_i443_3_lut_4_lut (.A(index_i[2]), .B(n26627), .C(index_i[3]), 
         .D(n26611), .Z(n443_adj_2909)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;
    defparam mux_193_Mux_7_i443_3_lut_4_lut.init = 16'h6f60;
    PFUMX i20389 (.BLUT(n158_adj_2910), .ALUT(n189_adj_2911), .C0(index_i[5]), 
          .Z(n22728));
    LUT4 mux_193_Mux_1_i924_3_lut (.A(n316_adj_2912), .B(n412_adj_2913), 
         .C(index_i[4]), .Z(n924_adj_2914)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_1_i924_3_lut.init = 16'hcaca;
    LUT4 n254_bdd_4_lut (.A(index_i[5]), .B(index_i[3]), .C(index_i[6]), 
         .D(index_i[4]), .Z(n25884)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;
    defparam n254_bdd_4_lut.init = 16'hf8f0;
    LUT4 mux_193_Mux_3_i860_3_lut_4_lut (.A(index_i[2]), .B(n26627), .C(index_i[4]), 
         .D(n859_adj_2915), .Z(n860_adj_2916)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam mux_193_Mux_3_i860_3_lut_4_lut.init = 16'hf606;
    LUT4 n25889_bdd_3_lut (.A(n26816), .B(n25885), .C(index_i[7]), .Z(n25890)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n25889_bdd_3_lut.init = 16'hcaca;
    LUT4 i12173_3_lut (.A(index_i[3]), .B(index_i[1]), .C(index_i[0]), 
         .Z(n14741)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i12173_3_lut.init = 16'hecec;
    LUT4 i21518_3_lut (.A(n21506), .B(n21507), .C(index_i[4]), .Z(n21508)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21518_3_lut.init = 16'hcaca;
    LUT4 i19762_3_lut_4_lut (.A(n26406), .B(n26405), .C(index_i[5]), .D(index_i[6]), 
         .Z(n22101)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (B+((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19762_3_lut_4_lut.init = 16'hffc5;
    LUT4 i18830_3_lut_4_lut (.A(n26642), .B(index_i[1]), .C(index_i[3]), 
         .D(n404), .Z(n21150)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18830_3_lut_4_lut.init = 16'hdfd0;
    LUT4 mux_193_Mux_1_i620_3_lut_4_lut (.A(n26642), .B(index_i[1]), .C(index_i[3]), 
         .D(n26662), .Z(n620_adj_2815)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_1_i620_3_lut_4_lut.init = 16'hdfd0;
    PFUMX i23135 (.BLUT(n24804), .ALUT(n475_adj_2859), .C0(index_i[4]), 
          .Z(n24805));
    LUT4 mux_193_Mux_0_i173_3_lut_4_lut (.A(n26642), .B(index_i[1]), .C(index_i[3]), 
         .D(n26669), .Z(n173_adj_2917)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i173_3_lut_4_lut.init = 16'hdfd0;
    L6MUX21 i24278 (.D0(n26105), .D1(n26102), .SD(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2127[4]));
    PFUMX i24276 (.BLUT(n26104), .ALUT(n26103), .C0(index_i[8]), .Z(n26105));
    LUT4 mux_193_Mux_1_i349_3_lut (.A(n506), .B(n348_adj_2918), .C(index_i[4]), 
         .Z(n349)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_1_i349_3_lut.init = 16'hcaca;
    LUT4 i21548_3_lut (.A(n21482), .B(n21483), .C(index_i[4]), .Z(n21484)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21548_3_lut.init = 16'hcaca;
    PFUMX i20538 (.BLUT(n22861), .ALUT(n22862), .C0(index_i[5]), .Z(n22877));
    PFUMX i20539 (.BLUT(n22863), .ALUT(n22864), .C0(index_i[5]), .Z(n22878));
    LUT4 i9493_3_lut (.A(n11938), .B(n26662), .C(index_i[3]), .Z(n11939)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9493_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_1_i94_3_lut (.A(index_i[0]), .B(n93_adj_2919), .C(index_i[4]), 
         .Z(n94_adj_2920)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_1_i94_3_lut.init = 16'hcaca;
    L6MUX21 i20540 (.D0(n22865), .D1(n22866), .SD(index_i[5]), .Z(n22879));
    LUT4 mux_193_Mux_5_i124_3_lut (.A(n645), .B(n26680), .C(index_i[3]), 
         .Z(n124)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_5_i124_3_lut.init = 16'hcaca;
    LUT4 i19082_3_lut (.A(n26669), .B(n26679), .C(index_i[3]), .Z(n21402)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19082_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_6_i636_4_lut_4_lut (.A(index_i[1]), .B(index_i[4]), 
         .C(n635_adj_2904), .D(n14379), .Z(n636_adj_2921)) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_6_i636_4_lut_4_lut.init = 16'hf3d1;
    LUT4 index_i_4__bdd_4_lut (.A(index_i[4]), .B(n26416), .C(n24193), 
         .D(index_i[5]), .Z(n26344)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (B (C (D))+!B (C+!(D)))) */ ;
    defparam index_i_4__bdd_4_lut.init = 16'hf099;
    PFUMX i23132 (.BLUT(n24801), .ALUT(n21141), .C0(index_i[4]), .Z(n24802));
    LUT4 mux_193_Mux_1_i987_3_lut_4_lut (.A(n29193), .B(index_i[3]), .C(index_i[4]), 
         .D(n986), .Z(n987)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_1_i987_3_lut_4_lut.init = 16'hf202;
    L6MUX21 i20543 (.D0(n22871), .D1(n22872), .SD(index_i[5]), .Z(n22882));
    PFUMX i24273 (.BLUT(n26101), .ALUT(n22753), .C0(index_i[8]), .Z(n26102));
    LUT4 mux_193_Mux_6_i891_3_lut (.A(n301), .B(n890_adj_2922), .C(index_i[4]), 
         .Z(n891_adj_2923)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_6_i891_3_lut.init = 16'hcaca;
    L6MUX21 i20544 (.D0(n22873), .D1(n22874), .SD(index_i[5]), .Z(n22883));
    LUT4 mux_193_Mux_6_i828_4_lut (.A(n812_adj_2924), .B(n13872), .C(index_i[4]), 
         .D(index_i[2]), .Z(n828_adj_2925)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_6_i828_4_lut.init = 16'hfaca;
    LUT4 mux_193_Mux_6_i797_3_lut (.A(n781), .B(n26360), .C(index_i[4]), 
         .Z(n797_adj_2926)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_6_i797_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_6_i669_3_lut (.A(n653_adj_2903), .B(n668_adj_2927), 
         .C(index_i[4]), .Z(n669_adj_2928)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_6_i669_3_lut.init = 16'hcaca;
    LUT4 n24800_bdd_3_lut_25422 (.A(n24800), .B(n22988), .C(index_i[6]), 
         .Z(n25942)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n24800_bdd_3_lut_25422.init = 16'hcaca;
    LUT4 index_i_7__bdd_4_lut_24668 (.A(index_i[7]), .B(n14872), .C(n24368), 
         .D(index_i[5]), .Z(n26345)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(B (C+(D))+!B !((D)+!C)))) */ ;
    defparam index_i_7__bdd_4_lut_24668.init = 16'h66f0;
    LUT4 n24800_bdd_3_lut_24149 (.A(n22989), .B(n24806), .C(index_i[6]), 
         .Z(n25941)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n24800_bdd_3_lut_24149.init = 16'hcaca;
    L6MUX21 i20545 (.D0(n22875), .D1(n22876), .SD(index_i[5]), .Z(n22884));
    LUT4 n24794_bdd_3_lut (.A(n24794), .B(n22984), .C(index_i[6]), .Z(n25944)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n24794_bdd_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_6_i542_3_lut (.A(n526_adj_2929), .B(n541_adj_2823), 
         .C(index_i[4]), .Z(n542_adj_2930)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_6_i542_3_lut.init = 16'hcaca;
    PFUMX i24263 (.BLUT(n26085), .ALUT(n29199), .C0(index_i[3]), .Z(n26086));
    LUT4 mux_193_Mux_6_i731_3_lut (.A(n26611), .B(n29193), .C(index_i[3]), 
         .Z(n731_adj_2931)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_6_i731_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_6_i252_4_lut (.A(index_i[2]), .B(n251_adj_2898), .C(index_i[4]), 
         .D(n11082), .Z(n252_adj_2932)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_6_i252_4_lut.init = 16'hc5ca;
    LUT4 i21963_3_lut (.A(n25383), .B(n252_adj_2932), .C(index_i[5]), 
         .Z(n22986)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21963_3_lut.init = 16'hcaca;
    L6MUX21 i23130 (.D0(n24799), .D1(n24797), .SD(index_i[5]), .Z(n24800));
    PFUMX i23128 (.BLUT(n24798), .ALUT(n285), .C0(index_i[4]), .Z(n24799));
    LUT4 mux_193_Mux_6_i844_3_lut_4_lut (.A(n26624), .B(index_i[2]), .C(index_i[3]), 
         .D(n26626), .Z(n844_adj_2797)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_6_i844_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_193_Mux_8_i157_3_lut_4_lut (.A(n26624), .B(index_i[2]), .C(index_i[3]), 
         .D(n26628), .Z(n15_adj_2933)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_8_i157_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_193_Mux_8_i301_3_lut_4_lut (.A(n26624), .B(index_i[2]), .C(index_i[3]), 
         .D(n70), .Z(n301)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_8_i301_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_193_Mux_8_i653_3_lut_rep_401_3_lut_4_lut (.A(n26624), .B(index_i[2]), 
         .C(index_i[3]), .D(n26508), .Z(n26361)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_8_i653_3_lut_rep_401_3_lut_4_lut.init = 16'h08f8;
    LUT4 i12377_2_lut_3_lut_4_lut (.A(n26416), .B(index_i[4]), .C(index_i[6]), 
         .D(index_i[5]), .Z(n14954)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i12377_2_lut_3_lut_4_lut.init = 16'hfef0;
    LUT4 mux_193_Mux_3_i251_3_lut_4_lut (.A(n26624), .B(index_i[2]), .C(index_i[3]), 
         .D(n26509), .Z(n14972)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_3_i251_3_lut_4_lut.init = 16'h8f80;
    PFUMX i23126 (.BLUT(n24796), .ALUT(n24795), .C0(index_i[4]), .Z(n24797));
    LUT4 i22402_2_lut_rep_411_3_lut_4_lut (.A(n26624), .B(index_i[2]), .C(index_i[5]), 
         .D(n26600), .Z(n26371)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i22402_2_lut_rep_411_3_lut_4_lut.init = 16'h0f7f;
    LUT4 n20957_bdd_3_lut_23120 (.A(n29168), .B(n26675), .C(index_i[3]), 
         .Z(n24791)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n20957_bdd_3_lut_23120.init = 16'hcaca;
    LUT4 mux_193_Mux_10_i574_4_lut_4_lut (.A(n26416), .B(index_i[4]), .C(index_i[5]), 
         .D(n26396), .Z(n574_adj_2814)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_10_i574_4_lut_4_lut.init = 16'h1f1c;
    LUT4 i19186_3_lut_3_lut_4_lut (.A(n26624), .B(index_i[2]), .C(n1001), 
         .D(index_i[3]), .Z(n21506)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19186_3_lut_3_lut_4_lut.init = 16'hf077;
    LUT4 mux_193_Mux_9_i364_3_lut_3_lut_4_lut (.A(n26624), .B(index_i[2]), 
         .C(n26509), .D(index_i[3]), .Z(n364_adj_2789)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_9_i364_3_lut_3_lut_4_lut.init = 16'h77f0;
    LUT4 n954_bdd_3_lut_24420_3_lut_4_lut (.A(n26624), .B(index_i[2]), .C(n70), 
         .D(index_i[3]), .Z(n24342)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n954_bdd_3_lut_24420_3_lut_4_lut.init = 16'hf077;
    LUT4 mux_193_Mux_3_i828_3_lut_3_lut_4_lut_4_lut_4_lut (.A(n26624), .B(index_i[2]), 
         .C(index_i[4]), .D(index_i[3]), .Z(n828)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C (D)+!C !(D)))+!A !(B (C+!(D))+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_3_i828_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h70c7;
    LUT4 mux_193_Mux_0_i1002_3_lut_3_lut_4_lut (.A(n26627), .B(index_i[2]), 
         .C(n1001), .D(index_i[3]), .Z(n1002_adj_2891)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i1002_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 mux_193_Mux_7_i890_3_lut_4_lut (.A(n26627), .B(index_i[2]), .C(index_i[3]), 
         .D(n26508), .Z(n890_adj_2792)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_7_i890_3_lut_4_lut.init = 16'hf101;
    L6MUX21 i23123 (.D0(n24793), .D1(n24790), .SD(index_i[5]), .Z(n24794));
    LUT4 n953_bdd_3_lut_23125 (.A(n26614), .B(index_i[3]), .C(n26682), 
         .Z(n24795)) /* synthesis lut_function=(A (B+(C))+!A !(B+!(C))) */ ;
    defparam n953_bdd_3_lut_23125.init = 16'hb8b8;
    LUT4 mux_193_Mux_8_i124_3_lut_3_lut_4_lut (.A(n26627), .B(index_i[2]), 
         .C(n26626), .D(index_i[3]), .Z(n124_adj_2813)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_8_i124_3_lut_3_lut_4_lut.init = 16'h11f0;
    PFUMX i23121 (.BLUT(n24792), .ALUT(n24791), .C0(index_i[4]), .Z(n24793));
    LUT4 mux_193_Mux_9_i124_3_lut_4_lut (.A(n26627), .B(index_i[2]), .C(index_i[3]), 
         .D(n26509), .Z(n124_adj_2861)) /* synthesis lut_function=(!(A (C+!(D))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_9_i124_3_lut_4_lut.init = 16'h1f10;
    LUT4 n285_bdd_3_lut (.A(n26614), .B(n26677), .C(index_i[3]), .Z(n24798)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n285_bdd_3_lut.init = 16'hacac;
    LUT4 mux_193_Mux_6_i890_3_lut_3_lut_4_lut (.A(n26627), .B(index_i[2]), 
         .C(n26629), .D(index_i[3]), .Z(n890_adj_2922)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_6_i890_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 mux_193_Mux_8_i475_3_lut_4_lut (.A(n26627), .B(index_i[2]), .C(index_i[3]), 
         .D(n26509), .Z(n475_adj_2934)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_8_i475_3_lut_4_lut.init = 16'hf101;
    LUT4 mux_193_Mux_7_i333_3_lut (.A(n26630), .B(n645), .C(index_i[3]), 
         .Z(n333)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_7_i333_3_lut.init = 16'hcaca;
    LUT4 n21141_bdd_3_lut_23531 (.A(n26673), .B(n26676), .C(index_i[3]), 
         .Z(n24801)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n21141_bdd_3_lut_23531.init = 16'hcaca;
    LUT4 mux_193_Mux_7_i348_3_lut (.A(n26625), .B(n29191), .C(index_i[3]), 
         .Z(n348_adj_2935)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_7_i348_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_3_i93_3_lut_4_lut (.A(n26627), .B(index_i[2]), .C(index_i[3]), 
         .D(n70), .Z(n93_adj_2829)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_3_i93_3_lut_4_lut.init = 16'hefe0;
    LUT4 n22753_bdd_3_lut (.A(n22746), .B(n22747), .C(index_i[7]), .Z(n26101)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n22753_bdd_3_lut.init = 16'hcaca;
    LUT4 n25002_bdd_3_lut_24275 (.A(n25002), .B(n22744), .C(index_i[7]), 
         .Z(n26103)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n25002_bdd_3_lut_24275.init = 16'hacac;
    PFUMX i23118 (.BLUT(n24789), .ALUT(n24788), .C0(index_i[4]), .Z(n24790));
    LUT4 i20522_3_lut (.A(n15_adj_2936), .B(n30_adj_2937), .C(index_i[4]), 
         .Z(n22861)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20522_3_lut.init = 16'hcaca;
    LUT4 i9492_3_lut_4_lut (.A(index_i[0]), .B(n26641), .C(index_i[4]), 
         .D(n588), .Z(n11938)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9492_3_lut_4_lut.init = 16'h4f40;
    LUT4 n25002_bdd_3_lut_25337 (.A(n22742), .B(n22743), .C(index_i[7]), 
         .Z(n26104)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n25002_bdd_3_lut_25337.init = 16'hcaca;
    LUT4 mux_193_Mux_2_i859_3_lut_4_lut (.A(index_i[0]), .B(n26641), .C(index_i[3]), 
         .D(n26614), .Z(n859)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_2_i859_3_lut_4_lut.init = 16'h4f40;
    LUT4 i19123_3_lut_4_lut (.A(index_i[0]), .B(n26641), .C(index_i[3]), 
         .D(n26678), .Z(n21443)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19123_3_lut_4_lut.init = 16'hf404;
    LUT4 mux_193_Mux_7_i397_3_lut (.A(n26625), .B(n26630), .C(index_i[3]), 
         .Z(n397_adj_2938)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_7_i397_3_lut.init = 16'hcaca;
    LUT4 n308_bdd_3_lut_23534 (.A(n29166), .B(n29179), .C(index_i[3]), 
         .Z(n24804)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n308_bdd_3_lut_23534.init = 16'hacac;
    PFUMX i20179 (.BLUT(n22514), .ALUT(n22515), .C0(index_i[5]), .Z(n22518));
    LUT4 mux_193_Mux_4_i158_3_lut (.A(n142_adj_2939), .B(n157), .C(index_i[4]), 
         .Z(n158_adj_2910)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_4_i158_3_lut.init = 16'hcaca;
    PFUMX i20180 (.BLUT(n22516), .ALUT(n22517), .C0(index_i[5]), .Z(n22519));
    PFUMX i20186 (.BLUT(n22521), .ALUT(n22522), .C0(index_i[5]), .Z(n22525));
    PFUMX i20187 (.BLUT(n22523), .ALUT(n22524), .C0(index_i[5]), .Z(n22526));
    LUT4 mux_193_Mux_7_i892_3_lut (.A(n62), .B(n891), .C(index_i[5]), 
         .Z(n892_adj_2817)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_7_i892_3_lut.init = 16'hcaca;
    LUT4 i18968_3_lut (.A(n747), .B(n762_adj_2791), .C(index_i[4]), .Z(n21288)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18968_3_lut.init = 16'hcaca;
    LUT4 i18967_3_lut (.A(n716_adj_2940), .B(n14714), .C(index_i[4]), 
         .Z(n21287)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18967_3_lut.init = 16'hcaca;
    LUT4 n24808_bdd_3_lut (.A(n24808), .B(n157_adj_2941), .C(index_i[4]), 
         .Z(n24809)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n24808_bdd_3_lut.init = 16'hcaca;
    LUT4 i18965_3_lut (.A(n93_adj_2942), .B(n699), .C(index_i[4]), .Z(n21285)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18965_3_lut.init = 16'hcaca;
    LUT4 i18964_3_lut (.A(n653_adj_2840), .B(n26391), .C(index_i[4]), 
         .Z(n21284)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18964_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_5_i700_3_lut (.A(n460_adj_2895), .B(n26675), .C(index_i[4]), 
         .Z(n700_adj_2943)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_5_i700_3_lut.init = 16'hcaca;
    LUT4 i18838_3_lut (.A(n325), .B(n26621), .C(index_i[3]), .Z(n21158)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18838_3_lut.init = 16'hcaca;
    LUT4 i18958_3_lut (.A(n526_adj_2944), .B(n15_adj_2936), .C(index_i[4]), 
         .Z(n21278)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18958_3_lut.init = 16'hcaca;
    LUT4 i18955_3_lut (.A(n397_adj_2938), .B(n475_adj_2839), .C(index_i[4]), 
         .Z(n21275)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18955_3_lut.init = 16'hcaca;
    LUT4 i18953_3_lut (.A(n348_adj_2935), .B(n443_adj_2909), .C(index_i[4]), 
         .Z(n21273)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18953_3_lut.init = 16'hcaca;
    LUT4 i18952_3_lut (.A(n397_adj_2938), .B(n731_adj_2931), .C(index_i[4]), 
         .Z(n21272)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18952_3_lut.init = 16'hcaca;
    LUT4 index_i_8__bdd_3_lut_then_4_lut (.A(index_i[4]), .B(index_i[6]), 
         .C(index_i[5]), .D(n26402), .Z(n26815)) /* synthesis lut_function=(!(A (B (C+(D)))+!A (B (C)))) */ ;
    defparam index_i_8__bdd_3_lut_then_4_lut.init = 16'h373f;
    LUT4 i19138_3_lut_3_lut_4_lut (.A(index_i[0]), .B(n26639), .C(n26509), 
         .D(index_i[3]), .Z(n21458)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(C+(D)))) */ ;
    defparam i19138_3_lut_3_lut_4_lut.init = 16'h77f0;
    LUT4 mux_193_Mux_0_i30_3_lut (.A(n26626), .B(n26628), .C(index_i[3]), 
         .Z(n30_adj_2937)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i30_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_5_i987_4_lut_4_lut_4_lut (.A(index_i[0]), .B(n26639), 
         .C(index_i[4]), .D(index_i[3]), .Z(n19592)) /* synthesis lut_function=(A (B (C+!(D))+!B (D))+!A (B (C (D)+!C !(D))+!B (D))) */ ;
    defparam mux_193_Mux_5_i987_4_lut_4_lut_4_lut.init = 16'hf38c;
    LUT4 i11214_3_lut_4_lut (.A(index_i[0]), .B(n26639), .C(n26600), .D(index_i[5]), 
         .Z(n318)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (C (D))) */ ;
    defparam i11214_3_lut_4_lut.init = 16'hf800;
    LUT4 i19171_3_lut_3_lut_4_lut (.A(index_i[0]), .B(n26639), .C(index_i[3]), 
         .D(n26509), .Z(n21491)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A !(C+(D))) */ ;
    defparam i19171_3_lut_3_lut_4_lut.init = 16'h808f;
    LUT4 mux_193_Mux_0_i986_3_lut (.A(n26673), .B(n985), .C(index_i[3]), 
         .Z(n986_adj_2887)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i986_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_0_i971_3_lut (.A(n26676), .B(n26629), .C(index_i[3]), 
         .Z(n971)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i971_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_0_i939_4_lut (.A(n588), .B(n26665), .C(index_i[3]), 
         .D(index_i[2]), .Z(n939)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i939_4_lut.init = 16'hfaca;
    LUT4 i22250_3_lut_4_lut (.A(n26507), .B(n19553), .C(index_i[8]), .D(n766), 
         .Z(n21165)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i22250_3_lut_4_lut.init = 16'hefe0;
    LUT4 mux_193_Mux_0_i572_3_lut_4_lut (.A(n26642), .B(index_i[1]), .C(index_i[3]), 
         .D(n26676), .Z(n572)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i572_3_lut_4_lut.init = 16'hefe0;
    LUT4 mux_193_Mux_0_i923_3_lut (.A(n26611), .B(n29191), .C(index_i[3]), 
         .Z(n923)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i923_3_lut.init = 16'hcaca;
    LUT4 i9392_4_lut_4_lut (.A(n26642), .B(index_i[1]), .C(index_i[3]), 
         .D(n20368), .Z(n11838)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A (B (C)+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9392_4_lut_4_lut.init = 16'h0e3e;
    LUT4 index_i_3__bdd_3_lut_22652_3_lut_4_lut (.A(n26642), .B(index_i[1]), 
         .C(index_i[4]), .D(index_i[3]), .Z(n24196)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam index_i_3__bdd_3_lut_22652_3_lut_4_lut.init = 16'hf10f;
    LUT4 i11194_2_lut_rep_417_3_lut_4_lut (.A(n26642), .B(index_i[1]), .C(index_i[4]), 
         .D(index_i[3]), .Z(n26377)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11194_2_lut_rep_417_3_lut_4_lut.init = 16'hfef0;
    LUT4 i20184_3_lut_4_lut (.A(n26498), .B(index_i[3]), .C(index_i[4]), 
         .D(n26459), .Z(n22523)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20184_3_lut_4_lut.init = 16'hfe0e;
    LUT4 i18943_4_lut_4_lut_3_lut_4_lut (.A(n26642), .B(index_i[1]), .C(index_i[4]), 
         .D(index_i[3]), .Z(n21263)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18943_4_lut_4_lut_3_lut_4_lut.init = 16'h11ef;
    LUT4 i12294_1_lut_2_lut_3_lut_4_lut (.A(n26498), .B(index_i[3]), .C(index_i[5]), 
         .D(index_i[4]), .Z(n381)) /* synthesis lut_function=(!(A (C+(D))+!A (B (C+(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i12294_1_lut_2_lut_3_lut_4_lut.init = 16'h010f;
    LUT4 i18836_3_lut (.A(n26661), .B(n26677), .C(index_i[3]), .Z(n21156)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18836_3_lut.init = 16'hcaca;
    LUT4 i9393_3_lut_4_lut_4_lut (.A(n26641), .B(index_i[3]), .C(index_i[5]), 
         .D(n26508), .Z(n11839)) /* synthesis lut_function=(A (B+(C (D)))+!A (B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9393_3_lut_4_lut_4_lut.init = 16'hf8c8;
    LUT4 i18835_3_lut (.A(n26660), .B(n26676), .C(index_i[3]), .Z(n21155)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18835_3_lut.init = 16'hcaca;
    LUT4 i18950_3_lut (.A(n364_adj_2945), .B(n379_adj_2889), .C(index_i[4]), 
         .Z(n21270)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18950_3_lut.init = 16'hcaca;
    LUT4 i18949_3_lut (.A(n333), .B(n348_adj_2935), .C(index_i[4]), .Z(n21269)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18949_3_lut.init = 16'hcaca;
    LUT4 i20177_3_lut_3_lut_4_lut_4_lut (.A(n26641), .B(index_i[3]), .C(index_i[4]), 
         .D(n26498), .Z(n22516)) /* synthesis lut_function=(!(A (B (C)+!B ((D)+!C))+!A (B+((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20177_3_lut_3_lut_4_lut_4_lut.init = 16'h0838;
    LUT4 n62_bdd_3_lut_4_lut (.A(n26641), .B(index_i[3]), .C(index_i[4]), 
         .D(n30_adj_2946), .Z(n24428)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n62_bdd_3_lut_4_lut.init = 16'hf808;
    LUT4 index_i_3__bdd_3_lut_22668_4_lut_4_lut (.A(n26641), .B(index_i[3]), 
         .C(index_i[4]), .D(n26499), .Z(n24197)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C))+!A !(B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam index_i_3__bdd_3_lut_22668_4_lut_4_lut.init = 16'h838f;
    LUT4 mux_193_Mux_10_i413_3_lut_3_lut_4_lut (.A(n26498), .B(index_i[3]), 
         .C(n26441), .D(index_i[4]), .Z(n413_adj_2947)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_10_i413_3_lut_3_lut_4_lut.init = 16'hf011;
    L6MUX21 i20645 (.D0(n21127), .D1(n21130), .SD(index_i[5]), .Z(n22984));
    LUT4 i18941_3_lut (.A(n491_adj_2948), .B(n506), .C(index_i[4]), .Z(n21261)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18941_3_lut.init = 16'hcaca;
    LUT4 i18940_3_lut (.A(n460_adj_2853), .B(n475_adj_2934), .C(index_i[4]), 
         .Z(n21260)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18940_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_5_i731_3_lut (.A(n26621), .B(n26677), .C(index_i[3]), 
         .Z(n731_adj_2879)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_5_i731_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_0_i716_3_lut (.A(n26674), .B(n26656), .C(index_i[3]), 
         .Z(n716_adj_2878)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i716_3_lut.init = 16'hcaca;
    LUT4 i18938_3_lut (.A(n251), .B(n443_adj_2794), .C(index_i[4]), .Z(n21258)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18938_3_lut.init = 16'hcaca;
    LUT4 i18937_3_lut (.A(n460_adj_2853), .B(n14714), .C(index_i[4]), 
         .Z(n21257)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;
    defparam i18937_3_lut.init = 16'h3a3a;
    L6MUX21 i20649 (.D0(n21136), .D1(n17548), .SD(index_i[5]), .Z(n22988));
    LUT4 i20182_3_lut_3_lut_4_lut (.A(n26498), .B(index_i[3]), .C(n412_adj_2913), 
         .D(index_i[4]), .Z(n22521)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20182_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 mux_193_Mux_10_i252_3_lut_4_lut_4_lut (.A(n26498), .B(index_i[3]), 
         .C(index_i[4]), .D(n26499), .Z(n252_adj_2836)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B (C (D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_10_i252_3_lut_4_lut_4_lut.init = 16'h3efe;
    L6MUX21 i20650 (.D0(n21139), .D1(n11888), .SD(index_i[5]), .Z(n22989));
    L6MUX21 i24154 (.D0(n25945), .D1(n25943), .SD(index_i[8]), .Z(n25946));
    LUT4 i18833_3_lut (.A(n29166), .B(n26676), .C(index_i[3]), .Z(n21153)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18833_3_lut.init = 16'hcaca;
    PFUMX i20652 (.BLUT(n542_adj_2930), .ALUT(n573_adj_2949), .C0(index_i[5]), 
          .Z(n22991));
    PFUMX i20653 (.BLUT(n605_adj_2950), .ALUT(n636_adj_2921), .C0(index_i[5]), 
          .Z(n22992));
    LUT4 index_i_8__bdd_3_lut_else_4_lut (.A(n26469), .B(index_i[4]), .C(index_i[6]), 
         .D(index_i[5]), .Z(n26814)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;
    defparam index_i_8__bdd_3_lut_else_4_lut.init = 16'hf080;
    PFUMX i24152 (.BLUT(n25944), .ALUT(n23000), .C0(index_i[7]), .Z(n25945));
    LUT4 mux_193_Mux_0_i653_3_lut (.A(n645), .B(n26666), .C(index_i[3]), 
         .Z(n653_adj_2863)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i653_3_lut.init = 16'hcaca;
    PFUMX i20654 (.BLUT(n669_adj_2928), .ALUT(n700_adj_2951), .C0(index_i[5]), 
          .Z(n22993));
    LUT4 i18928_3_lut (.A(n301), .B(n93_adj_2942), .C(index_i[4]), .Z(n21248)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18928_3_lut.init = 16'hcaca;
    PFUMX i20655 (.BLUT(n732_adj_2952), .ALUT(n21145), .C0(index_i[5]), 
          .Z(n22994));
    LUT4 mux_193_Mux_0_i620_3_lut (.A(n26625), .B(n26662), .C(index_i[3]), 
         .Z(n620_adj_2848)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i620_3_lut.init = 16'hcaca;
    LUT4 i18925_3_lut (.A(n15_adj_2933), .B(n526_adj_2832), .C(index_i[4]), 
         .Z(n21245)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18925_3_lut.init = 16'hcaca;
    PFUMX i20656 (.BLUT(n797_adj_2926), .ALUT(n828_adj_2925), .C0(index_i[5]), 
          .Z(n22995));
    PFUMX i20657 (.BLUT(n860_adj_2798), .ALUT(n891_adj_2923), .C0(index_i[5]), 
          .Z(n22996));
    PFUMX i24150 (.BLUT(n25942), .ALUT(n25941), .C0(index_i[7]), .Z(n25943));
    LUT4 i22231_3_lut_rep_391_4_lut (.A(n26489), .B(index_i[5]), .C(index_i[8]), 
         .D(n1021), .Z(n26351)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i22231_3_lut_rep_391_4_lut.init = 16'hf808;
    L6MUX21 i20244 (.D0(n22581), .D1(n22582), .SD(index_i[5]), .Z(n22583));
    PFUMX i20676 (.BLUT(n94_adj_2920), .ALUT(n21475), .C0(index_i[5]), 
          .Z(n23015));
    LUT4 mux_193_Mux_0_i589_3_lut (.A(n29191), .B(n588), .C(index_i[3]), 
         .Z(n589)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i589_3_lut.init = 16'hcaca;
    L6MUX21 i20251 (.D0(n22588), .D1(n22589), .SD(index_i[5]), .Z(n22590));
    L6MUX21 i20677 (.D0(n21478), .D1(n21481), .SD(index_i[5]), .Z(n23016));
    LUT4 i11652_3_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .Z(n11082)) /* synthesis lut_function=(!((B (C))+!A)) */ ;
    defparam i11652_3_lut.init = 16'h2a2a;
    PFUMX i20675 (.BLUT(n11939), .ALUT(n62_adj_2953), .C0(index_i[5]), 
          .Z(n23014));
    L6MUX21 i20258 (.D0(n22595), .D1(n22596), .SD(index_i[5]), .Z(n22597));
    LUT4 i18829_3_lut (.A(n26679), .B(n26676), .C(index_i[3]), .Z(n21149)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18829_3_lut.init = 16'hcaca;
    PFUMX i20679 (.BLUT(n21484), .ALUT(n317_adj_2954), .C0(index_i[5]), 
          .Z(n23018));
    L6MUX21 i20265 (.D0(n22602), .D1(n22603), .SD(index_i[5]), .Z(n22604));
    PFUMX i20680 (.BLUT(n349), .ALUT(n21487), .C0(index_i[5]), .Z(n23019));
    L6MUX21 i20681 (.D0(n21490), .D1(n21493), .SD(index_i[5]), .Z(n23020));
    LUT4 mux_193_Mux_6_i653_3_lut (.A(n26658), .B(n85), .C(index_i[3]), 
         .Z(n653_adj_2903)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_6_i653_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_6_i668_3_lut (.A(n108), .B(n26633), .C(index_i[3]), 
         .Z(n668_adj_2927)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_6_i668_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_6_i684_3_lut (.A(n645), .B(n29199), .C(index_i[3]), 
         .Z(n684_adj_2955)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_6_i684_3_lut.init = 16'hcaca;
    LUT4 i18827_3_lut (.A(n26680), .B(n29199), .C(index_i[3]), .Z(n21147)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18827_3_lut.init = 16'hcaca;
    L6MUX21 i20682 (.D0(n21496), .D1(n21499), .SD(index_i[5]), .Z(n23021));
    LUT4 i21505_3_lut (.A(n21146), .B(n21147), .C(index_i[4]), .Z(n21148)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21505_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_3_i747_3_lut (.A(n26679), .B(n404), .C(index_i[3]), 
         .Z(n747_adj_2827)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_3_i747_3_lut.init = 16'hcaca;
    LUT4 n187_bdd_4_lut_23266 (.A(n26499), .B(index_i[6]), .C(index_i[5]), 
         .D(n26628), .Z(n24872)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(D))+!A !(B (C+(D))+!B (D)))) */ ;
    defparam n187_bdd_4_lut_23266.init = 16'h7f40;
    LUT4 i21908_3_lut (.A(n286), .B(n317), .C(index_i[5]), .Z(n22140)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21908_3_lut.init = 16'hcaca;
    L6MUX21 i20684 (.D0(n21505), .D1(n636), .SD(index_i[5]), .Z(n23023));
    LUT4 n24875_bdd_3_lut (.A(n26786), .B(n24872), .C(index_i[4]), .Z(n24876)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n24875_bdd_3_lut.init = 16'hcaca;
    PFUMX i20747 (.BLUT(n844_adj_2956), .ALUT(n11823), .C0(index_i[4]), 
          .Z(n23086));
    LUT4 i1_3_lut_rep_529_4_lut (.A(index_i[3]), .B(index_i[4]), .C(index_i[2]), 
         .D(n26627), .Z(n26489)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i1_3_lut_rep_529_4_lut.init = 16'hfffe;
    PFUMX i24111 (.BLUT(n25890), .ALUT(n1022), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2127[12]));
    LUT4 n24878_bdd_3_lut (.A(n24878), .B(n24876), .C(index_i[3]), .Z(n24879)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n24878_bdd_3_lut.init = 16'hcaca;
    PFUMX i20685 (.BLUT(n21508), .ALUT(n700_adj_2812), .C0(index_i[5]), 
          .Z(n23024));
    L6MUX21 i20687 (.D0(n21511), .D1(n21514), .SD(index_i[5]), .Z(n23026));
    PFUMX i20689 (.BLUT(n924_adj_2914), .ALUT(n21520), .C0(index_i[5]), 
          .Z(n23028));
    LUT4 i1_3_lut_4_lut (.A(index_i[3]), .B(index_i[4]), .C(index_i[5]), 
         .D(n26639), .Z(n20077)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i1_3_lut_4_lut.init = 16'hfffe;
    LUT4 mux_193_Mux_5_i859_3_lut (.A(n141), .B(n26659), .C(index_i[3]), 
         .Z(n859_adj_2892)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_5_i859_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_5_i875_3_lut (.A(n645), .B(n26625), .C(index_i[3]), 
         .Z(n875_adj_2888)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_5_i875_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_6_i732_3_lut_4_lut (.A(n26630), .B(index_i[3]), .C(index_i[4]), 
         .D(n731_adj_2931), .Z(n732_adj_2952)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_6_i732_3_lut_4_lut.init = 16'hf909;
    LUT4 i9448_3_lut_4_lut (.A(index_i[3]), .B(index_i[4]), .C(n26654), 
         .D(n29199), .Z(n605_adj_2950)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9448_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i24107 (.BLUT(n254_adj_2787), .ALUT(n25884), .C0(index_i[8]), 
          .Z(n25885));
    LUT4 i20659_3_lut_4_lut_4_lut (.A(n26474), .B(index_i[5]), .C(index_i[4]), 
         .D(n26418), .Z(n22998)) /* synthesis lut_function=(A (B+(C (D)))+!A (B+((D)+!C))) */ ;
    defparam i20659_3_lut_4_lut_4_lut.init = 16'hfdcd;
    PFUMX i20690 (.BLUT(n987), .ALUT(n21523), .C0(index_i[5]), .Z(n23029));
    PFUMX i20304 (.BLUT(n31_adj_2908), .ALUT(n21148), .C0(index_i[5]), 
          .Z(n22643));
    PFUMX i20305 (.BLUT(n94_adj_2905), .ALUT(n125_adj_2902), .C0(index_i[5]), 
          .Z(n22644));
    PFUMX i20306 (.BLUT(n17582), .ALUT(n14378), .C0(index_i[5]), .Z(n22645));
    LUT4 i19081_3_lut (.A(n26614), .B(n325), .C(index_i[3]), .Z(n21401)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19081_3_lut.init = 16'hcaca;
    LUT4 i21395_3_lut (.A(n21401), .B(n21402), .C(index_i[4]), .Z(n21403)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21395_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_6_i700_3_lut_4_lut (.A(n26630), .B(index_i[3]), .C(index_i[4]), 
         .D(n684_adj_2955), .Z(n700_adj_2951)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_6_i700_3_lut_4_lut.init = 16'h9f90;
    L6MUX21 i20308 (.D0(n21151), .D1(n21154), .SD(index_i[5]), .Z(n22647));
    L6MUX21 i20309 (.D0(n21157), .D1(n21160), .SD(index_i[5]), .Z(n22648));
    LUT4 mux_193_Mux_1_i732_3_lut (.A(n716), .B(n491), .C(index_i[4]), 
         .Z(n732)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_1_i732_3_lut.init = 16'hcaca;
    PFUMX i20310 (.BLUT(n413_adj_2899), .ALUT(n444), .C0(index_i[5]), 
          .Z(n22649));
    LUT4 mux_193_Mux_4_i15_3_lut (.A(n29165), .B(n588), .C(index_i[3]), 
         .Z(n15_adj_2851)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_4_i15_3_lut.init = 16'hcaca;
    PFUMX i20311 (.BLUT(n476_adj_2896), .ALUT(n507), .C0(index_i[5]), 
          .Z(n22650));
    LUT4 mux_193_Mux_4_i61_3_lut (.A(n26681), .B(n26656), .C(index_i[3]), 
         .Z(n61)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_4_i61_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_2_i908_3_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n908_adj_2957)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C)+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_2_i908_3_lut_4_lut_4_lut.init = 16'h5a51;
    LUT4 i21957_3_lut (.A(n924_adj_2958), .B(n955), .C(index_i[5]), .Z(n22997)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21957_3_lut.init = 16'hcaca;
    LUT4 i9464_3_lut_3_lut_4_lut (.A(index_i[3]), .B(index_i[4]), .C(n26681), 
         .D(index_i[0]), .Z(n605_adj_2959)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9464_3_lut_3_lut_4_lut.init = 16'h10fe;
    PFUMX i20312 (.BLUT(n17551), .ALUT(n573_adj_2960), .C0(index_i[5]), 
          .Z(n22651));
    LUT4 i22202_3_lut (.A(n24810), .B(n22986), .C(index_i[6]), .Z(n23000)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22202_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_2_i270_3_lut (.A(n26659), .B(n26612), .C(index_i[3]), 
         .Z(n270_adj_2874)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_2_i270_3_lut.init = 16'hcaca;
    LUT4 i18821_3_lut (.A(n404), .B(n26660), .C(index_i[3]), .Z(n21141)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18821_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_2_i316_3_lut (.A(n26663), .B(n26681), .C(index_i[3]), 
         .Z(n316_adj_2872)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_2_i316_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_2_i397_3_lut (.A(n29199), .B(n26611), .C(index_i[3]), 
         .Z(n397_adj_2870)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_2_i397_3_lut.init = 16'hcaca;
    LUT4 i18818_3_lut (.A(n404), .B(n26667), .C(index_i[3]), .Z(n21138)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18818_3_lut.init = 16'hcaca;
    LUT4 i18817_3_lut (.A(n26669), .B(n325), .C(index_i[3]), .Z(n21137)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18817_3_lut.init = 16'hcaca;
    LUT4 i18815_3_lut (.A(n26669), .B(n26667), .C(index_i[3]), .Z(n21135)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18815_3_lut.init = 16'hcaca;
    PFUMX i20313 (.BLUT(n605_adj_2959), .ALUT(n636_adj_2894), .C0(index_i[5]), 
          .Z(n22652));
    LUT4 i18814_3_lut (.A(n325), .B(n332), .C(index_i[3]), .Z(n21134)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18814_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_4_i270_3_lut (.A(n26662), .B(n26666), .C(index_i[3]), 
         .Z(n270)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_4_i270_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_4_i348_3_lut (.A(n26617), .B(n26669), .C(index_i[3]), 
         .Z(n348_adj_2961)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_4_i348_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_4_i684_3_lut (.A(n85), .B(n108), .C(index_i[3]), 
         .Z(n684_adj_2842)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_4_i684_3_lut.init = 16'hcaca;
    LUT4 i15397_3_lut (.A(n26667), .B(n26661), .C(index_i[3]), .Z(n17547)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15397_3_lut.init = 16'hcaca;
    LUT4 i15396_3_lut (.A(n26661), .B(n26669), .C(index_i[3]), .Z(n17546)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15396_3_lut.init = 16'hcaca;
    PFUMX i20314 (.BLUT(n21163), .ALUT(n700_adj_2943), .C0(index_i[5]), 
          .Z(n22653));
    LUT4 i22468_2_lut (.A(index_i[5]), .B(index_i[4]), .Z(n21938)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i22468_2_lut.init = 16'heeee;
    LUT4 i1_3_lut (.A(index_i[0]), .B(index_i[4]), .C(index_i[2]), .Z(n20368)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i1_3_lut.init = 16'hfefe;
    LUT4 i12179_3_lut (.A(index_i[3]), .B(index_i[1]), .C(index_i[0]), 
         .Z(n14747)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i12179_3_lut.init = 16'hc8c8;
    LUT4 mux_193_Mux_3_i348_3_lut (.A(n29179), .B(n26660), .C(index_i[3]), 
         .Z(n348_adj_2962)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_3_i348_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_3_i908_3_lut (.A(n26678), .B(n26656), .C(index_i[3]), 
         .Z(n908)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_3_i908_3_lut.init = 16'hcaca;
    L6MUX21 i20315 (.D0(n732_adj_2880), .D1(n21766), .SD(index_i[5]), 
            .Z(n22654));
    PFUMX i20316 (.BLUT(n797_adj_2963), .ALUT(n828_adj_2964), .C0(index_i[5]), 
          .Z(n22655));
    LUT4 i19201_3_lut (.A(n26666), .B(n26678), .C(index_i[3]), .Z(n21521)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19201_3_lut.init = 16'hcaca;
    PFUMX i20317 (.BLUT(n860_adj_2893), .ALUT(n891_adj_2890), .C0(index_i[5]), 
          .Z(n22656));
    LUT4 i21508_3_lut (.A(n21521), .B(n21522), .C(index_i[4]), .Z(n21523)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21508_3_lut.init = 16'hcaca;
    PFUMX i24078 (.BLUT(n25845), .ALUT(n25843), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2127[10]));
    LUT4 i20699_3_lut (.A(n23030), .B(n23031), .C(index_i[7]), .Z(n23038)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20699_3_lut.init = 16'hcaca;
    LUT4 i20692_3_lut (.A(n23016), .B(n25417), .C(index_i[6]), .Z(n23031)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20692_3_lut.init = 16'hcaca;
    LUT4 i20701_3_lut (.A(n23034), .B(n23035), .C(index_i[7]), .Z(n23040)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20701_3_lut.init = 16'hcaca;
    LUT4 i20695_3_lut (.A(n25438), .B(n23023), .C(index_i[6]), .Z(n23034)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20695_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_6_i924_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[4]), .D(n762_adj_2791), .Z(n924_adj_2958)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_6_i924_3_lut_4_lut.init = 16'h6f60;
    PFUMX i25985 (.BLUT(n28805), .ALUT(n28804), .C0(index_i[3]), .Z(n28806));
    PFUMX i24076 (.BLUT(n21197), .ALUT(n25841), .C0(index_i[7]), .Z(n25842));
    LUT4 i20451_3_lut (.A(n22784), .B(n22785), .C(index_i[7]), .Z(n22790)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20451_3_lut.init = 16'hcaca;
    PFUMX i25983 (.BLUT(n28801), .ALUT(n28800), .C0(index_i[2]), .Z(n28802));
    LUT4 i20446_3_lut (.A(n22774), .B(n22775), .C(index_i[6]), .Z(n22785)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20446_3_lut.init = 16'hcaca;
    PFUMX mux_193_Mux_1_i891 (.BLUT(n882), .ALUT(n890_adj_2965), .C0(n26552), 
          .Z(n891_adj_2810)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 i19198_3_lut (.A(n1001), .B(n588), .C(index_i[3]), .Z(n21518)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19198_3_lut.init = 16'hcaca;
    LUT4 i8618_4_lut_4_lut (.A(index_i[3]), .B(index_i[0]), .C(index_i[1]), 
         .D(index_i[2]), .Z(n11000)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (D)+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i8618_4_lut_4_lut.init = 16'h0bf4;
    LUT4 i21510_3_lut (.A(n21518), .B(n21519), .C(index_i[4]), .Z(n21520)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21510_3_lut.init = 16'hcaca;
    LUT4 i20325_3_lut (.A(n22653), .B(n22654), .C(index_i[6]), .Z(n22664)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20325_3_lut.init = 16'hcaca;
    PFUMX i24064 (.BLUT(n25815), .ALUT(n25814), .C0(index_i[8]), .Z(n25816));
    LUT4 mux_193_Mux_2_i221_4_lut_4_lut (.A(index_i[3]), .B(index_i[4]), 
         .C(n26508), .D(n26396), .Z(n221_adj_2966)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (B+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_2_i221_4_lut_4_lut.init = 16'hf7c4;
    LUT4 i19839_3_lut (.A(n24969), .B(n22171), .C(index_i[7]), .Z(n22178)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19839_3_lut.init = 16'hcaca;
    LUT4 i20183_3_lut_4_lut_3_lut (.A(index_i[3]), .B(index_i[4]), .C(n26499), 
         .Z(n22522)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20183_3_lut_4_lut_3_lut.init = 16'h6464;
    LUT4 i19846_3_lut (.A(n24430), .B(n28807), .C(index_i[7]), .Z(n22185)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19846_3_lut.init = 16'hcaca;
    LUT4 i11132_4_lut_4_lut (.A(index_i[3]), .B(index_i[2]), .C(index_i[0]), 
         .D(index_i[1]), .Z(n875_adj_2885)) /* synthesis lut_function=((B (C)+!B (D))+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11132_4_lut_4_lut.init = 16'hf7d5;
    LUT4 i18971_4_lut_3_lut (.A(index_i[3]), .B(index_i[4]), .C(n26508), 
         .Z(n21291)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18971_4_lut_3_lut.init = 16'h6565;
    LUT4 i9394_3_lut_3_lut (.A(index_i[3]), .B(index_i[4]), .C(n11839), 
         .Z(n11840)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9394_3_lut_3_lut.init = 16'h7474;
    LUT4 i19829_4_lut_4_lut (.A(index_i[4]), .B(index_i[5]), .C(n26792), 
         .D(n908_adj_2957), .Z(n22168)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam i19829_4_lut_4_lut.init = 16'hd1c0;
    LUT4 mux_193_Mux_3_i796_3_lut_3_lut (.A(index_i[4]), .B(n731_adj_2931), 
         .C(index_i[2]), .Z(n796_adj_2967)) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam mux_193_Mux_3_i796_3_lut_3_lut.init = 16'he4e4;
    LUT4 i12113_2_lut_rep_591 (.A(index_i[2]), .B(index_i[0]), .Z(n26551)) /* synthesis lut_function=(A (B)) */ ;
    defparam i12113_2_lut_rep_591.init = 16'h8888;
    LUT4 mux_193_Mux_3_i700_3_lut_4_lut (.A(index_i[4]), .B(index_i[3]), 
         .C(n684_adj_2968), .D(n29168), .Z(n700_adj_2969)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_3_i700_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i22444_2_lut_rep_592 (.A(index_i[4]), .B(index_i[3]), .Z(n26552)) /* synthesis lut_function=((B)+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i22444_2_lut_rep_592.init = 16'hdddd;
    LUT4 mux_193_Mux_3_i797_3_lut_4_lut (.A(index_i[4]), .B(index_i[3]), 
         .C(n796_adj_2967), .D(n70), .Z(n797)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_3_i797_3_lut_4_lut.init = 16'hf2d0;
    LUT4 n25842_bdd_3_lut_3_lut (.A(n1021), .B(index_i[8]), .C(n25842), 
         .Z(n25843)) /* synthesis lut_function=(A (B+(C))+!A !(B+!(C))) */ ;
    defparam n25842_bdd_3_lut_3_lut.init = 16'hb8b8;
    PFUMX i20387 (.BLUT(n31_adj_2881), .ALUT(n62_adj_2877), .C0(index_i[5]), 
          .Z(n22726));
    LUT4 n17754_bdd_4_lut_then_4_lut (.A(index_i[3]), .B(index_i[4]), .C(index_i[1]), 
         .D(index_i[2]), .Z(n26827)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B+(C (D)+!C !(D)))) */ ;
    defparam n17754_bdd_4_lut_then_4_lut.init = 16'hf44f;
    LUT4 n17754_bdd_4_lut_else_4_lut (.A(index_i[3]), .B(index_i[4]), .C(index_i[1]), 
         .D(index_i[2]), .Z(n26826)) /* synthesis lut_function=(!(A (B (D)+!B ((D)+!C))+!A !(B+!((D)+!C)))) */ ;
    defparam n17754_bdd_4_lut_else_4_lut.init = 16'h44fc;
    PFUMX i24501 (.BLUT(n26796), .ALUT(n26797), .C0(index_i[1]), .Z(n26798));
    PFUMX i19817 (.BLUT(n158_adj_2876), .ALUT(n189_adj_2802), .C0(index_i[5]), 
          .Z(n22156));
    PFUMX i19818 (.BLUT(n221_adj_2966), .ALUT(n21454), .C0(index_i[5]), 
          .Z(n22157));
    LUT4 i11429_2_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n635_adj_2816)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A (B (C+!(D))+!B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11429_2_lut_4_lut_4_lut.init = 16'hf1fc;
    LUT4 i19169_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n21489)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B ((D)+!C)+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19169_3_lut_4_lut_4_lut.init = 16'hfc1c;
    PFUMX i19819 (.BLUT(n286_adj_2875), .ALUT(n317_adj_2873), .C0(index_i[5]), 
          .Z(n22158));
    PFUMX i19820 (.BLUT(n349_adj_2970), .ALUT(n21457), .C0(index_i[5]), 
          .Z(n22159));
    PFUMX i19821 (.BLUT(n413_adj_2871), .ALUT(n21460), .C0(index_i[5]), 
          .Z(n22160));
    LUT4 n24963_bdd_3_lut (.A(n24963), .B(n476), .C(index_i[5]), .Z(n24964)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n24963_bdd_3_lut.init = 16'hcaca;
    LUT4 i19190_3_lut (.A(n26681), .B(n26660), .C(index_i[3]), .Z(n21510)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19190_3_lut.init = 16'hcaca;
    PFUMX i19822 (.BLUT(n21463), .ALUT(n507_adj_2971), .C0(index_i[5]), 
          .Z(n22161));
    PFUMX i19823 (.BLUT(n21466), .ALUT(n573_adj_2869), .C0(index_i[5]), 
          .Z(n22162));
    PFUMX i19824 (.BLUT(n605), .ALUT(n21469), .C0(index_i[5]), .Z(n22163));
    PFUMX i19825 (.BLUT(n669_adj_2860), .ALUT(n700_adj_2850), .C0(index_i[5]), 
          .Z(n22164));
    PFUMX i19826 (.BLUT(n732_adj_2857), .ALUT(n763_adj_2972), .C0(index_i[5]), 
          .Z(n22165));
    LUT4 i22323_2_lut_rep_600 (.A(index_i[1]), .B(index_i[2]), .Z(n26560)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i22323_2_lut_rep_600.init = 16'h9999;
    LUT4 n262_bdd_2_lut_23957_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[3]), 
         .Z(n25676)) /* synthesis lut_function=(A (B+(C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n262_bdd_2_lut_23957_3_lut.init = 16'hf9f9;
    LUT4 mux_193_Mux_0_i93_3_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .Z(n93_adj_2833)) /* synthesis lut_function=(A (B)+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i93_3_lut_3_lut.init = 16'h9c9c;
    L6MUX21 i19828 (.D0(n860_adj_2820), .D1(n891_adj_2819), .SD(index_i[5]), 
            .Z(n22167));
    L6MUX21 i20753 (.D0(n23076), .D1(n23077), .SD(index_i[5]), .Z(n23092));
    L6MUX21 i20754 (.D0(n23078), .D1(n23079), .SD(index_i[5]), .Z(n23093));
    L6MUX21 i20755 (.D0(n23080), .D1(n23081), .SD(index_i[5]), .Z(n23094));
    L6MUX21 i20756 (.D0(n23082), .D1(n23083), .SD(index_i[5]), .Z(n23095));
    PFUMX i20388 (.BLUT(n94), .ALUT(n21397), .C0(index_i[5]), .Z(n22727));
    LUT4 i19898_3_lut (.A(n22235), .B(n22236), .C(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2127[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19898_3_lut.init = 16'hcaca;
    LUT4 i20674_3_lut (.A(n25946), .B(n23012), .C(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2127[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20674_3_lut.init = 16'hcaca;
    LUT4 i20673_3_lut (.A(n23009), .B(n23010), .C(index_i[8]), .Z(n23012)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20673_3_lut.init = 16'hcaca;
    L6MUX21 i20757 (.D0(n23084), .D1(n23085), .SD(index_i[5]), .Z(n23096));
    LUT4 i11409_3_lut_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n13969)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11409_3_lut_3_lut_3_lut_4_lut.init = 16'h10ff;
    PFUMX i20390 (.BLUT(n221_adj_2973), .ALUT(n252_adj_2974), .C0(index_i[5]), 
          .Z(n22729));
    LUT4 mux_193_Mux_5_i781_3_lut_4_lut_4_lut_then_4_lut (.A(index_i[3]), 
         .B(index_i[0]), .C(index_i[4]), .D(index_i[2]), .Z(n26753)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_5_i781_3_lut_4_lut_4_lut_then_4_lut.init = 16'hece0;
    LUT4 n24967_bdd_3_lut (.A(n26777), .B(n24965), .C(index_i[5]), .Z(n24968)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n24967_bdd_3_lut.init = 16'hcaca;
    PFUMX i20391 (.BLUT(n286_adj_2852), .ALUT(n21400), .C0(index_i[5]), 
          .Z(n22730));
    LUT4 mux_193_Mux_0_i915_3_lut_rep_651_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26611)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i915_3_lut_rep_651_3_lut.init = 16'he3e3;
    L6MUX21 i20758 (.D0(n23086), .D1(n23087), .SD(index_i[5]), .Z(n23097));
    LUT4 mux_193_Mux_2_i716_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n716_adj_2855)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)+!C !(D)))+!A (B (D)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_2_i716_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h31cf;
    PFUMX i20392 (.BLUT(n349_adj_2975), .ALUT(n21403), .C0(index_i[5]), 
          .Z(n22731));
    LUT4 mux_193_Mux_3_i157_3_lut_3_lut_rep_453_3_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n26413)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_3_i157_3_lut_3_lut_rep_453_3_lut_4_lut.init = 16'h1ff0;
    LUT4 mux_193_Mux_0_i15_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n15_adj_2936)) /* synthesis lut_function=(A (B (D)+!B (C+!(D)))+!A (B (D)+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i15_3_lut_4_lut_4_lut_4_lut.init = 16'hec33;
    LUT4 i19159_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n21479)) /* synthesis lut_function=(A (B (D)+!B ((D)+!C))+!A (B (D)+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19159_3_lut_4_lut_4_lut_4_lut.init = 16'hfe13;
    LUT4 mux_193_Mux_0_i698_3_lut_rep_665 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26625)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i698_3_lut_rep_665.init = 16'h1c1c;
    LUT4 mux_193_Mux_8_i45_3_lut_rep_666 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26626)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_8_i45_3_lut_rep_666.init = 16'hc1c1;
    LUT4 n22_bdd_3_lut_23451_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n25148)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C (D)+!C !(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n22_bdd_3_lut_23451_3_lut_4_lut.init = 16'h0fc1;
    LUT4 i19115_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21435)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19115_3_lut_3_lut_4_lut.init = 16'h0f1c;
    LUT4 i19192_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21512)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C (D)))+!A (B (C+(D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19192_4_lut_4_lut_4_lut.init = 16'h301c;
    L6MUX21 i20759 (.D0(n23088), .D1(n23089), .SD(index_i[5]), .Z(n23098));
    LUT4 mux_193_Mux_0_i699_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n699_adj_2866)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (D))+!A (B (C+!(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i699_3_lut_3_lut_4_lut.init = 16'h1c33;
    LUT4 mux_193_Mux_0_i557_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n557)) /* synthesis lut_function=(A ((D)+!C)+!A !((D)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i557_3_lut_4_lut.init = 16'haa4e;
    LUT4 i11434_2_lut_rep_667 (.A(index_i[0]), .B(index_i[1]), .Z(n26627)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11434_2_lut_rep_667.init = 16'h8888;
    LUT4 i11113_2_lut_rep_653 (.A(index_i[0]), .B(index_i[1]), .Z(n26613)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11113_2_lut_rep_653.init = 16'h4444;
    L6MUX21 i20760 (.D0(n23090), .D1(n23091), .SD(index_i[5]), .Z(n23099));
    LUT4 i11312_2_lut_2_lut_3_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .Z(n13872)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11312_2_lut_2_lut_3_lut.init = 16'h0808;
    LUT4 i19177_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n21497)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A (B (C)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19177_3_lut_4_lut_4_lut.init = 16'h3c8c;
    LUT4 n676_bdd_2_lut_24268_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n25433)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A (B+((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n676_bdd_2_lut_24268_4_lut_4_lut_4_lut.init = 16'h0038;
    LUT4 mux_193_Mux_0_i954_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n954_adj_2886)) /* synthesis lut_function=(A (D)+!A !(B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i954_3_lut_4_lut_4_lut.init = 16'haf40;
    LUT4 n77_bdd_3_lut_24299_3_lut_4_lut_4_lut_3_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n25413)) /* synthesis lut_function=(A (B (C)+!B !(D))+!A !(D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n77_bdd_3_lut_24299_3_lut_4_lut_4_lut_3_lut_4_lut.init = 16'h80f7;
    PFUMX i20397 (.BLUT(n669_adj_2845), .ALUT(n700_adj_2843), .C0(index_i[5]), 
          .Z(n22736));
    LUT4 mux_193_Mux_8_i526_3_lut_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n526_adj_2799)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_8_i526_3_lut_3_lut_3_lut_4_lut.init = 16'h0f70;
    LUT4 i11118_2_lut_rep_436_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n26396)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11118_2_lut_rep_436_3_lut_4_lut.init = 16'hf080;
    LUT4 mux_193_Mux_8_i635_3_lut_4_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n635)) /* synthesis lut_function=(!(A (B (C (D))+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_8_i635_3_lut_4_lut_3_lut_4_lut.init = 16'h0ff8;
    LUT4 i12299_2_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(n26638), 
         .D(index_i[2]), .Z(n14872)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i12299_2_lut_3_lut_4_lut.init = 16'hf080;
    LUT4 i20238_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n22577)) /* synthesis lut_function=(A (B (D)+!B !(C (D)+!C !(D)))+!A !(B (C+!(D))+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20238_3_lut_4_lut_4_lut.init = 16'h8f30;
    LUT4 mux_193_Mux_4_i1002_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n1002)) /* synthesis lut_function=(A (B (C (D))+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_4_i1002_3_lut_3_lut_4_lut.init = 16'hf007;
    LUT4 mux_193_Mux_6_i812_3_lut_4_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n812_adj_2924)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(D))+!A !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_6_i812_3_lut_4_lut_3_lut_4_lut.init = 16'h7780;
    LUT4 i11117_2_lut_rep_539_3_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .Z(n26499)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11117_2_lut_rep_539_3_lut.init = 16'hf8f8;
    PFUMX i20398 (.BLUT(n21415), .ALUT(n763_adj_2900), .C0(index_i[5]), 
          .Z(n22737));
    LUT4 mux_193_Mux_3_i1002_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n19598)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (D))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_3_i1002_3_lut_3_lut_4_lut.init = 16'hf708;
    LUT4 i19172_3_lut_4_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n21492)) /* synthesis lut_function=(!(A (B (D)+!B !((D)+!C))+!A (B (C+(D))+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19172_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'h338f;
    LUT4 mux_193_Mux_1_i348_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n348_adj_2918)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A (B ((D)+!C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_1_i348_3_lut_4_lut_4_lut_4_lut.init = 16'h38f0;
    LUT4 mux_193_Mux_8_i172_rep_34_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n70)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_8_i172_rep_34_3_lut_3_lut.init = 16'h7c7c;
    PFUMX i20399 (.BLUT(n21418), .ALUT(n828_adj_2976), .C0(index_i[5]), 
          .Z(n22738));
    LUT4 mux_193_Mux_7_i491_3_lut_4_lut_4_lut_4_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[2]), .D(index_i[3]), .Z(n491_adj_2806)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A (B ((D)+!C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_7_i491_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'h3870;
    LUT4 i11283_3_lut_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n13842)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (D))+!A (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11283_3_lut_3_lut_3_lut_4_lut.init = 16'h00f7;
    LUT4 i22518_2_lut_rep_499_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n26459)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i22518_2_lut_rep_499_3_lut_4_lut.init = 16'h0007;
    LUT4 mux_193_Mux_7_i141_3_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n141)) /* synthesis lut_function=(A ((C)+!B)+!A (B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_7_i141_3_lut_4_lut_3_lut.init = 16'he7e7;
    CCU2D unary_minus_10_add_3_17 (.A0(\quarter_wave_sample_register_q[15] ), 
          .B0(GND_net), .C0(GND_net), .D0(GND_net), .A1(GND_net), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n17398), .S0(o_val_pipeline_i_0__15__N_2158[15]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam unary_minus_10_add_3_17.INIT0 = 16'hf555;
    defparam unary_minus_10_add_3_17.INIT1 = 16'h0000;
    defparam unary_minus_10_add_3_17.INJECT1_0 = "NO";
    defparam unary_minus_10_add_3_17.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_508_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n26468)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i1_2_lut_rep_508_3_lut_4_lut.init = 16'h8000;
    LUT4 mux_193_Mux_6_i781_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n781)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A (B (C (D)+!C !(D))+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_6_i781_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hc837;
    LUT4 mux_193_Mux_7_i526_3_lut_3_lut_4_lut_4_lut_3_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n526_adj_2944)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(D))+!A !(D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_7_i526_3_lut_3_lut_4_lut_4_lut_3_lut_4_lut.init = 16'h887f;
    LUT4 i19105_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n21425)) /* synthesis lut_function=(!(A (B (D)+!B !(D))+!A (B ((D)+!C)+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19105_3_lut_4_lut_4_lut_4_lut.init = 16'h33c8;
    LUT4 mux_193_Mux_0_i29_3_lut_rep_668 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26628)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i29_3_lut_rep_668.init = 16'h8383;
    LUT4 mux_193_Mux_8_i29_3_lut_rep_669 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26629)) /* synthesis lut_function=(!(A (B (C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_8_i29_3_lut_rep_669.init = 16'h7e7e;
    LUT4 mux_193_Mux_7_i92_3_lut_rep_670 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26630)) /* synthesis lut_function=(A (B+!(C))+!A !((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_7_i92_3_lut_rep_670.init = 16'h8e8e;
    LUT4 mux_193_Mux_5_i781_3_lut_4_lut_4_lut_else_4_lut (.A(index_i[3]), 
         .B(index_i[0]), .C(index_i[4]), .Z(n26752)) /* synthesis lut_function=(!(A (C)+!A (B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_5_i781_3_lut_4_lut_4_lut_else_4_lut.init = 16'h1f1f;
    LUT4 mux_193_Mux_7_i60_3_lut_4_lut_3_lut_rep_673 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26633)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_7_i60_3_lut_4_lut_3_lut_rep_673.init = 16'h1818;
    CCU2D unary_minus_10_add_3_15 (.A0(quarter_wave_sample_register_i[13]), 
          .B0(GND_net), .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[14]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17397), .COUT(n17398), 
          .S0(o_val_pipeline_i_0__15__N_2158[13]), .S1(o_val_pipeline_i_0__15__N_2158[14]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam unary_minus_10_add_3_15.INIT0 = 16'hf555;
    defparam unary_minus_10_add_3_15.INIT1 = 16'hf555;
    defparam unary_minus_10_add_3_15.INJECT1_0 = "NO";
    defparam unary_minus_10_add_3_15.INJECT1_1 = "NO";
    LUT4 i19157_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21477)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A (B (D)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19157_3_lut_4_lut.init = 16'h18cc;
    LUT4 mux_193_Mux_2_i557_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n557_adj_2868)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C+!(D))+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_2_i557_3_lut_3_lut_4_lut.init = 16'h0f18;
    LUT4 mux_193_Mux_7_i716_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n716_adj_2940)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C+!(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_7_i716_3_lut_3_lut_4_lut.init = 16'h0f81;
    LUT4 n262_bdd_3_lut_24192_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n25252)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C))+!A (B (C (D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n262_bdd_3_lut_24192_3_lut_4_lut.init = 16'h0fc7;
    LUT4 i19114_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21434)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)))+!A !(B (C+!(D))+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19114_3_lut_3_lut_4_lut.init = 16'h71cc;
    LUT4 mux_193_Mux_4_i526_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n526_adj_2832)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A !(B ((D)+!C)+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_4_i526_3_lut_3_lut_4_lut.init = 16'h7e0f;
    LUT4 mux_193_Mux_8_i93_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n93_adj_2942)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C))+!A (B (C+!(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_8_i93_3_lut_3_lut_4_lut.init = 16'h0f83;
    LUT4 mux_193_Mux_7_i620_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n620)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B ((D)+!C)+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_7_i620_3_lut_4_lut_4_lut.init = 16'h83c3;
    LUT4 mux_193_Mux_4_i812_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[4]), .D(index_i[3]), .Z(n812_adj_2977)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A !(B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_4_i812_3_lut_4_lut_4_lut.init = 16'ha595;
    PFUMX i20400 (.BLUT(n860_adj_2837), .ALUT(n21421), .C0(index_i[5]), 
          .Z(n22739));
    LUT4 i19175_3_lut (.A(n29165), .B(n26682), .C(index_i[3]), .Z(n21495)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19175_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_4_i142_3_lut_3_lut_3_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[3]), .Z(n142_adj_2939)) /* synthesis lut_function=(A (B (C))+!A !(B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_4_i142_3_lut_3_lut_3_lut.init = 16'h9595;
    L6MUX21 i23963 (.D0(n25692), .D1(n25690), .SD(index_i[5]), .Z(n25693));
    PFUMX i23961 (.BLUT(n25691), .ALUT(n645), .C0(index_i[3]), .Z(n25692));
    CCU2D unary_minus_10_add_3_13 (.A0(quarter_wave_sample_register_i[11]), 
          .B0(GND_net), .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[12]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17396), .COUT(n17397), 
          .S0(o_val_pipeline_i_0__15__N_2158[11]), .S1(o_val_pipeline_i_0__15__N_2158[12]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam unary_minus_10_add_3_13.INIT0 = 16'hf555;
    defparam unary_minus_10_add_3_13.INIT1 = 16'hf555;
    defparam unary_minus_10_add_3_13.INJECT1_0 = "NO";
    defparam unary_minus_10_add_3_13.INJECT1_1 = "NO";
    PFUMX mux_193_Mux_7_i190 (.BLUT(n21040), .ALUT(n173_adj_2808), .C0(index_i[5]), 
          .Z(n190)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    PFUMX i23959 (.BLUT(n25689), .ALUT(n21042), .C0(index_i[4]), .Z(n25690));
    L6MUX21 i23955 (.D0(n25680), .D1(n25678), .SD(index_i[5]), .Z(n25681));
    L6MUX21 i25554 (.D0(n28206), .D1(n28203), .SD(index_i[7]), .Z(n28207));
    PFUMX i25552 (.BLUT(n28205), .ALUT(n28204), .C0(index_i[5]), .Z(n28206));
    PFUMX i23953 (.BLUT(n572_adj_2978), .ALUT(n25679), .C0(index_i[4]), 
          .Z(n25680));
    PFUMX i25550 (.BLUT(n22149), .ALUT(n28202), .C0(index_i[6]), .Z(n28203));
    PFUMX i23950 (.BLUT(n25677), .ALUT(n25676), .C0(index_i[4]), .Z(n25678));
    PFUMX mux_193_Mux_8_i764 (.BLUT(n716_adj_2979), .ALUT(n732_adj_2834), 
          .C0(n21938), .Z(n764)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    L6MUX21 i23943 (.D0(n25669), .D1(n25666), .SD(index_i[5]), .Z(n25670));
    LUT4 i9477_2_lut_rep_678 (.A(index_i[3]), .B(index_i[4]), .Z(n26638)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9477_2_lut_rep_678.init = 16'h8888;
    PFUMX mux_193_Mux_8_i574 (.BLUT(n542_adj_2800), .ALUT(n11838), .C0(index_i[5]), 
          .Z(n574)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    PFUMX i23941 (.BLUT(n25668), .ALUT(n25667), .C0(index_i[4]), .Z(n25669));
    LUT4 i1_2_lut_rep_547_3_lut (.A(index_i[3]), .B(index_i[4]), .C(index_i[5]), 
         .Z(n26507)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i1_2_lut_rep_547_3_lut.init = 16'hf8f8;
    LUT4 i19803_3_lut_3_lut_4_lut (.A(index_i[3]), .B(index_i[4]), .C(n413_adj_2947), 
         .D(index_i[5]), .Z(n22142)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19803_3_lut_3_lut_4_lut.init = 16'h77f0;
    LUT4 i1_2_lut_3_lut (.A(index_i[3]), .B(index_i[4]), .C(index_i[5]), 
         .Z(n20226)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i1_2_lut_3_lut.init = 16'h8080;
    LUT4 i11428_2_lut_rep_679 (.A(index_i[1]), .B(index_i[2]), .Z(n26639)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11428_2_lut_rep_679.init = 16'h8888;
    LUT4 i9484_2_lut_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[3]), 
         .Z(n11930)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9484_2_lut_3_lut.init = 16'h8080;
    LUT4 i19076_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n21396)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C (D)+!C !(D)))+!A !(B (D)+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19076_3_lut_4_lut_4_lut_4_lut.init = 16'h7c03;
    PFUMX i18875 (.BLUT(n445), .ALUT(n508), .C0(index_i[6]), .Z(n21195));
    LUT4 i15399_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n17549)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C (D)+!C !(D)))+!A !(B (D)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i15399_3_lut_4_lut_4_lut_4_lut.init = 16'h83fc;
    LUT4 i19097_3_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[3]), 
         .D(index_i[0]), .Z(n21417)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19097_3_lut_3_lut_4_lut.init = 16'hf80f;
    LUT4 i11815_2_lut_rep_520_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[0]), 
         .Z(n26480)) /* synthesis lut_function=(A (B+!(C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11815_2_lut_rep_520_3_lut.init = 16'h8f8f;
    PFUMX i23938 (.BLUT(n26368), .ALUT(n25665), .C0(index_i[4]), .Z(n25666));
    PFUMX i19891 (.BLUT(n956), .ALUT(n20077), .C0(index_i[6]), .Z(n22230));
    LUT4 i11226_2_lut_rep_514_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[3]), 
         .Z(n26474)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11226_2_lut_rep_514_3_lut.init = 16'hf8f8;
    LUT4 mux_193_Mux_4_i93_3_lut_4_lut_3_lut_rep_616_4_lut (.A(index_i[1]), 
         .B(index_i[2]), .C(index_i[3]), .D(index_i[0]), .Z(n26576)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_4_i93_3_lut_4_lut_3_lut_rep_616_4_lut.init = 16'h07f0;
    PFUMX i20425 (.BLUT(n31), .ALUT(n62_adj_2980), .C0(index_i[5]), .Z(n22764));
    LUT4 i11752_2_lut_rep_548_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[0]), 
         .Z(n26508)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11752_2_lut_rep_548_3_lut.init = 16'h8080;
    LUT4 i19139_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .D(index_i[3]), .Z(n21459)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(D))+!A (B+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19139_3_lut_4_lut_4_lut_4_lut.init = 16'h3380;
    PFUMX i20426 (.BLUT(n94_adj_2981), .ALUT(n125), .C0(index_i[5]), .Z(n22765));
    LUT4 mux_193_Mux_3_i142_3_lut_3_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .Z(n142_adj_2831)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_3_i142_3_lut_3_lut_3_lut.init = 16'h3838;
    LUT4 i11209_2_lut_rep_458_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n26418)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11209_2_lut_rep_458_3_lut_4_lut.init = 16'hf8f0;
    LUT4 i19168_3_lut (.A(n26681), .B(n26621), .C(index_i[3]), .Z(n21488)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19168_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_8_i491_3_lut_3_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n491_adj_2948)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_8_i491_3_lut_3_lut_3_lut_4_lut.init = 16'h7870;
    LUT4 mux_193_Mux_9_i30_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .D(index_i[3]), .Z(n30_adj_2946)) /* synthesis lut_function=(A (B (C (D))+!B !(D))+!A !(B+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_9_i30_3_lut_4_lut_4_lut_4_lut.init = 16'h8033;
    PFUMX i20427 (.BLUT(n158), .ALUT(n189), .C0(index_i[5]), .Z(n22766));
    LUT4 i11749_2_lut_rep_680 (.A(index_i[1]), .B(index_i[2]), .C(index_i[0]), 
         .Z(n26640)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11749_2_lut_rep_680.init = 16'h7070;
    LUT4 i21545_3_lut (.A(n21485), .B(n21486), .C(index_i[4]), .Z(n21487)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21545_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_0_i1017_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .D(index_i[3]), .Z(n1017)) /* synthesis lut_function=(A (B (D)+!B !((D)+!C))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i1017_4_lut_4_lut_4_lut.init = 16'hdd70;
    LUT4 i11437_2_lut_rep_681 (.A(index_i[1]), .B(index_i[2]), .Z(n26641)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11437_2_lut_rep_681.init = 16'heeee;
    LUT4 mux_193_Mux_8_i412_3_lut_4_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .Z(n14714)) /* synthesis lut_function=(A (B+!(C))+!A !((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_8_i412_3_lut_4_lut_3_lut.init = 16'h8e8e;
    LUT4 i11751_2_lut_rep_494_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[0]), 
         .Z(n26454)) /* synthesis lut_function=(A (C)+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11751_2_lut_rep_494_3_lut.init = 16'hf1f1;
    LUT4 mux_193_Mux_9_i93_3_lut_3_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .Z(n93)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_9_i93_3_lut_3_lut_3_lut.init = 16'hc1c1;
    PFUMX i20428 (.BLUT(n221_adj_2846), .ALUT(n252), .C0(index_i[5]), 
          .Z(n22767));
    LUT4 mux_193_Mux_4_i236_3_lut_4_lut_3_lut_rep_617_4_lut (.A(index_i[1]), 
         .B(index_i[2]), .C(index_i[3]), .D(index_i[0]), .Z(n26577)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_4_i236_3_lut_4_lut_3_lut_rep_617_4_lut.init = 16'hf01f;
    LUT4 mux_193_Mux_9_i412_3_lut_3_lut_4_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .Z(n412_adj_2913)) /* synthesis lut_function=(!(A (B (C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_9_i412_3_lut_3_lut_4_lut_3_lut.init = 16'h7e7e;
    PFUMX i20429 (.BLUT(n286_adj_2830), .ALUT(n21430), .C0(index_i[5]), 
          .Z(n22768));
    LUT4 i11218_2_lut_rep_550_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[3]), 
         .Z(n26510)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11218_2_lut_rep_550_3_lut.init = 16'he0e0;
    LUT4 i19075_3_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[3]), 
         .D(index_i[0]), .Z(n21395)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19075_3_lut_3_lut_4_lut.init = 16'h0fe0;
    LUT4 n476_bdd_3_lut_24678 (.A(n476), .B(n24997), .C(index_i[5]), .Z(n24998)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n476_bdd_3_lut_24678.init = 16'hcaca;
    LUT4 i19202_3_lut_3_lut_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[3]), 
         .Z(n21522)) /* synthesis lut_function=(A (C)+!A (B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19202_3_lut_3_lut_3_lut.init = 16'he5e5;
    LUT4 i11219_2_lut_rep_457_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[4]), .D(index_i[3]), .Z(n26417)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11219_2_lut_rep_457_3_lut_4_lut.init = 16'hfef0;
    LUT4 mux_193_Mux_1_i317_3_lut (.A(n301_adj_2982), .B(n908_adj_2957), 
         .C(index_i[4]), .Z(n317_adj_2954)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_1_i317_3_lut.init = 16'hcaca;
    LUT4 n9680_bdd_3_lut_24042_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[4]), .D(index_i[3]), .Z(n24193)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C+(D)))+!A (B (C (D)+!C !(D))+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n9680_bdd_3_lut_24042_4_lut_4_lut_4_lut.init = 16'hc10f;
    PFUMX i20430 (.BLUT(n349_adj_2983), .ALUT(n21433), .C0(index_i[5]), 
          .Z(n22769));
    LUT4 i12174_2_lut_rep_682 (.A(index_i[2]), .B(index_i[0]), .Z(n26642)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i12174_2_lut_rep_682.init = 16'heeee;
    LUT4 i19079_3_lut (.A(n26672), .B(n26666), .C(index_i[3]), .Z(n21399)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19079_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_2_i173_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[2]), 
         .B(index_i[0]), .C(index_i[3]), .D(index_i[1]), .Z(n173)) /* synthesis lut_function=(!(A (C)+!A (B (C+!(D))+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_2_i173_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h0f1a;
    PFUMX i20431 (.BLUT(n413), .ALUT(n444_adj_2984), .C0(index_i[5]), 
          .Z(n22770));
    LUT4 i1_2_lut_rep_549_3_lut (.A(index_i[2]), .B(index_i[0]), .C(index_i[1]), 
         .Z(n26509)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i1_2_lut_rep_549_3_lut.init = 16'hfefe;
    LUT4 mux_193_Mux_0_i46_3_lut_4_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[1]), .D(index_i[3]), .Z(n46_adj_2847)) /* synthesis lut_function=(A (D)+!A (B+(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i46_3_lut_4_lut_4_lut_4_lut.init = 16'hfe55;
    LUT4 mux_193_Mux_8_i716_3_lut_4_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[1]), .D(index_i[3]), .Z(n716_adj_2979)) /* synthesis lut_function=(!(A (D)+!A !(B+(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_8_i716_3_lut_4_lut_4_lut_4_lut.init = 16'h55fe;
    PFUMX i20432 (.BLUT(n476_adj_2825), .ALUT(n507_adj_2985), .C0(index_i[5]), 
          .Z(n22771));
    LUT4 i11193_2_lut_rep_456_3_lut_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[1]), .Z(n26416)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11193_2_lut_rep_456_3_lut_4_lut.init = 16'hf0e0;
    LUT4 mux_193_Mux_9_i285_3_lut_3_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[1]), .Z(n285_adj_2865)) /* synthesis lut_function=(A (C)+!A !(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_9_i285_3_lut_3_lut_4_lut_4_lut.init = 16'ha0a1;
    PFUMX i20433 (.BLUT(n21436), .ALUT(n573_adj_2867), .C0(index_i[5]), 
          .Z(n22772));
    LUT4 mux_193_Mux_5_i954_3_lut_3_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[1]), .Z(n954)) /* synthesis lut_function=(!(A (C)+!A (B+((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_5_i954_3_lut_3_lut_4_lut_4_lut.init = 16'h0a1a;
    PFUMX i20434 (.BLUT(n11926), .ALUT(n21439), .C0(index_i[5]), .Z(n22773));
    LUT4 n172_bdd_2_lut_3_lut_3_lut_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[1]), .D(index_i[3]), .Z(n25218)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n172_bdd_2_lut_3_lut_3_lut_4_lut.init = 16'h00fe;
    LUT4 i19156_3_lut (.A(n900), .B(n26660), .C(index_i[3]), .Z(n21476)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19156_3_lut.init = 16'hcaca;
    PFUMX i20435 (.BLUT(n669), .ALUT(n700_adj_2969), .C0(index_i[5]), 
          .Z(n22774));
    L6MUX21 i20436 (.D0(n21442), .D1(n763_adj_2828), .SD(index_i[5]), 
            .Z(n22775));
    PFUMX i20438 (.BLUT(n860_adj_2916), .ALUT(n891_adj_2824), .C0(index_i[5]), 
          .Z(n22777));
    PFUMX i20439 (.BLUT(n924_adj_2822), .ALUT(n21445), .C0(index_i[5]), 
          .Z(n22778));
    PFUMX i20440 (.BLUT(n21448), .ALUT(n1018), .C0(index_i[5]), .Z(n22779));
    LUT4 i21399_3_lut (.A(n21398), .B(n21399), .C(index_i[4]), .Z(n21400)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21399_3_lut.init = 16'hcaca;
    LUT4 i18946_3_lut_4_lut_4_lut (.A(n26508), .B(index_i[4]), .C(index_i[3]), 
         .D(n26498), .Z(n21266)) /* synthesis lut_function=(A (B (C)+!B !(C+!(D)))+!A (B (C)+!B (C+(D)))) */ ;
    defparam i18946_3_lut_4_lut_4_lut.init = 16'hd3d0;
    LUT4 i7339_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n157)) /* synthesis lut_function=(!(A (C (D))+!A !(B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i7339_3_lut_4_lut_4_lut.init = 16'h4aaa;
    LUT4 i11224_2_lut_rep_615 (.A(index_i[2]), .B(index_i[3]), .Z(n26575)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11224_2_lut_rep_615.init = 16'heeee;
    L6MUX21 i25350 (.D0(n27968), .D1(n27965), .SD(index_i[5]), .Z(n27969));
    PFUMX i25348 (.BLUT(n27967), .ALUT(n27966), .C0(index_i[3]), .Z(n27968));
    PFUMX i25346 (.BLUT(n27964), .ALUT(n27963), .C0(index_i[3]), .Z(n27965));
    LUT4 i20246_3_lut_3_lut (.A(n26630), .B(index_i[3]), .C(n29199), .Z(n22585)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam i20246_3_lut_3_lut.init = 16'h7474;
    CCU2D unary_minus_10_add_3_11 (.A0(quarter_wave_sample_register_i[9]), 
          .B0(GND_net), .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[10]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17395), .COUT(n17396), 
          .S0(o_val_pipeline_i_0__15__N_2158[9]), .S1(o_val_pipeline_i_0__15__N_2158[10]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam unary_minus_10_add_3_11.INIT0 = 16'hf555;
    defparam unary_minus_10_add_3_11.INIT1 = 16'hf555;
    defparam unary_minus_10_add_3_11.INJECT1_0 = "NO";
    defparam unary_minus_10_add_3_11.INJECT1_1 = "NO";
    LUT4 i21556_3_lut (.A(n26773), .B(n21474), .C(index_i[4]), .Z(n21475)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21556_3_lut.init = 16'hcaca;
    LUT4 i19092_then_4_lut (.A(index_i[0]), .B(index_i[4]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n26759)) /* synthesis lut_function=(A (B (C)+!B (C (D)+!C !(D)))+!A !(B (C+!(D))+!B !(C+!(D)))) */ ;
    defparam i19092_then_4_lut.init = 16'hb493;
    LUT4 mux_193_Mux_7_i364_3_lut_3_lut (.A(n26630), .B(index_i[3]), .C(n26625), 
         .Z(n364_adj_2945)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;
    defparam mux_193_Mux_7_i364_3_lut_3_lut.init = 16'hd1d1;
    LUT4 i11760_2_lut_rep_509_3_lut (.A(index_i[2]), .B(index_i[3]), .C(index_i[1]), 
         .Z(n26469)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11760_2_lut_rep_509_3_lut.init = 16'hfefe;
    LUT4 i19147_3_lut (.A(n404), .B(n26614), .C(index_i[3]), .Z(n21467)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19147_3_lut.init = 16'hcaca;
    LUT4 i20766_3_lut (.A(n23102), .B(n23103), .C(index_i[7]), .Z(n23105)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20766_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_4_i668_3_lut_3_lut (.A(n26630), .B(index_i[3]), .C(n29199), 
         .Z(n668_adj_2844)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;
    defparam mux_193_Mux_4_i668_3_lut_3_lut.init = 16'hd1d1;
    PFUMX i19446 (.BLUT(n21764), .ALUT(n21765), .C0(index_i[4]), .Z(n21766));
    LUT4 mux_193_Mux_7_i379_3_lut_3_lut (.A(n26630), .B(index_i[3]), .C(n29191), 
         .Z(n379_adj_2889)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam mux_193_Mux_7_i379_3_lut_3_lut.init = 16'h7474;
    LUT4 i19088_3_lut_3_lut (.A(n26630), .B(index_i[3]), .C(n1001), .Z(n21408)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam i19088_3_lut_3_lut.init = 16'h7474;
    LUT4 i21416_3_lut (.A(n21467), .B(n21468), .C(index_i[4]), .Z(n21469)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21416_3_lut.init = 16'hcaca;
    PFUMX i20705 (.BLUT(n23042), .ALUT(n23043), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2127[1]));
    LUT4 i19092_else_4_lut (.A(index_i[0]), .B(index_i[4]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n26758)) /* synthesis lut_function=(!(A (B (C)+!B !(C+!(D)))+!A (B (C)+!B (D)))) */ ;
    defparam i19092_else_4_lut.init = 16'h2c3f;
    LUT4 i20765_3_lut (.A(n23100), .B(n23101), .C(index_i[7]), .Z(n23104)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20765_3_lut.init = 16'hcaca;
    LUT4 i19142_3_lut (.A(n404), .B(n29166), .C(index_i[3]), .Z(n21462)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19142_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_2_i763_4_lut_4_lut (.A(index_i[0]), .B(n11930), .C(index_i[4]), 
         .D(n157_adj_2941), .Z(n763_adj_2972)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_2_i763_4_lut_4_lut.init = 16'hdfd0;
    LUT4 mux_193_Mux_5_i573_3_lut_3_lut (.A(index_i[0]), .B(index_i[4]), 
         .C(n572_adj_2978), .Z(n573_adj_2960)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_5_i573_3_lut_3_lut.init = 16'hd1d1;
    LUT4 mux_193_Mux_2_i507_3_lut_3_lut (.A(index_i[0]), .B(index_i[4]), 
         .C(n491_adj_2986), .Z(n507_adj_2971)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_2_i507_3_lut_3_lut.init = 16'h7474;
    LUT4 i21422_3_lut (.A(n21458), .B(n21459), .C(index_i[4]), .Z(n21460)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21422_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_0_i953_rep_654 (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .Z(n26614)) /* synthesis lut_function=(A (C)+!A !((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i953_rep_654.init = 16'ha4a4;
    PFUMX i9442 (.BLUT(n12052), .ALUT(n12053), .C0(n22053), .Z(n11888));
    LUT4 i19187_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21507)) /* synthesis lut_function=(!(A ((D)+!C)+!A !(B ((D)+!C)+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19187_3_lut_3_lut_4_lut.init = 16'h55a4;
    LUT4 mux_193_Mux_4_i221_3_lut_3_lut (.A(index_i[0]), .B(index_i[4]), 
         .C(n205), .Z(n221_adj_2973)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_4_i221_3_lut_3_lut.init = 16'h7474;
    L6MUX21 i22655 (.D0(n24198), .D1(n26344), .SD(index_i[6]), .Z(n24199));
    LUT4 mux_193_Mux_0_i781_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n781_adj_2884)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A (B (C)+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i781_4_lut_4_lut_4_lut.init = 16'h0cb4;
    LUT4 mux_193_Mux_1_i890_4_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[3]), 
         .C(n645), .D(index_i[4]), .Z(n890_adj_2965)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (D))+!A !((C+(D))+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_1_i890_4_lut_4_lut_4_lut_4_lut.init = 16'h55f3;
    PFUMX i20455 (.BLUT(n22792), .ALUT(n22793), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2127[3]));
    LUT4 mux_193_Mux_2_i349_3_lut_3_lut (.A(index_i[0]), .B(index_i[4]), 
         .C(n348_adj_2987), .Z(n349_adj_2970)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_2_i349_3_lut_3_lut.init = 16'hd1d1;
    LUT4 mux_193_Mux_4_i252_4_lut_4_lut (.A(index_i[0]), .B(index_i[3]), 
         .C(n26641), .D(index_i[4]), .Z(n252_adj_2974)) /* synthesis lut_function=(!(A (B (D)+!B !(D))+!A !(B ((D)+!C)+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_4_i252_4_lut_4_lut.init = 16'h669d;
    LUT4 mux_193_Mux_3_i444_3_lut_4_lut (.A(index_i[0]), .B(index_i[3]), 
         .C(n26639), .D(index_i[4]), .Z(n444_adj_2984)) /* synthesis lut_function=(!(A (B (D)+!B (C (D)))+!A !(B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_3_i444_3_lut_4_lut.init = 16'h46aa;
    LUT4 i19136_3_lut (.A(n29166), .B(n26680), .C(index_i[3]), .Z(n21456)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19136_3_lut.init = 16'hcaca;
    LUT4 i22327_2_lut_rep_694 (.A(index_i[0]), .B(index_i[1]), .Z(n26654)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i22327_2_lut_rep_694.init = 16'h9999;
    LUT4 mux_193_Mux_6_i498_3_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n404)) /* synthesis lut_function=(A (B+!(C))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_6_i498_3_lut_4_lut_3_lut.init = 16'h9b9b;
    LUT4 n25000_bdd_3_lut (.A(n26767), .B(n444_adj_2988), .C(index_i[5]), 
         .Z(n25001)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n25000_bdd_3_lut.init = 16'hcaca;
    LUT4 i11131_2_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n844_adj_2956)) /* synthesis lut_function=(A (B+!(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11131_2_lut_3_lut_4_lut.init = 16'h9ff9;
    LUT4 mux_193_Mux_2_i604_3_lut_4_lut_4_lut_4_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n604_adj_2862)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)+!C !(D)))+!A (B (C)+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_2_i604_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'h3c9f;
    LUT4 i19174_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n21494)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !(B (C+!(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19174_3_lut_4_lut_4_lut.init = 16'ha5a9;
    LUT4 i9476_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(n26596), .D(index_i[4]), .Z(n189_adj_2911)) /* synthesis lut_function=(A (B (C (D)))+!A !(B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9476_3_lut_4_lut_4_lut_4_lut.init = 16'h9555;
    LUT4 i19837_3_lut (.A(n25670), .B(n22167), .C(index_i[6]), .Z(n22176)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19837_3_lut.init = 16'hcaca;
    LUT4 i9446_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n541_adj_2823)) /* synthesis lut_function=(A (B (C (D))+!B !(C (D)))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9446_3_lut_4_lut_4_lut_4_lut.init = 16'h9333;
    LUT4 i21424_3_lut (.A(n21455), .B(n21456), .C(index_i[4]), .Z(n21457)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21424_3_lut.init = 16'hcaca;
    LUT4 i21403_3_lut (.A(n21395), .B(n21396), .C(index_i[4]), .Z(n21397)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21403_3_lut.init = 16'hcaca;
    PFUMX i19769 (.BLUT(n22106), .ALUT(n22107), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2127[8]));
    LUT4 i11125_2_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n668_adj_2864)) /* synthesis lut_function=(!(A ((D)+!B)+!A (B ((D)+!C)+!B (C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11125_2_lut_4_lut_4_lut_4_lut.init = 16'h00c9;
    LUT4 i15430_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n17580)) /* synthesis lut_function=(A (B)+!A !(B (C (D))+!B !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i15430_3_lut_4_lut_4_lut.init = 16'h9ccc;
    LUT4 i11114_2_lut_rep_656 (.A(index_i[0]), .B(index_i[1]), .Z(n26616)) /* synthesis lut_function=((B)+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11114_2_lut_rep_656.init = 16'hdddd;
    LUT4 i21431_3_lut (.A(n21452), .B(n21453), .C(index_i[4]), .Z(n21454)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21431_3_lut.init = 16'hcaca;
    LUT4 i15431_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n17581)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i15431_3_lut_4_lut_4_lut_4_lut.init = 16'h3999;
    LUT4 i20262_3_lut (.A(n141), .B(n29193), .C(index_i[3]), .Z(n22601)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20262_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_6_i573_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[4]), .D(n572_adj_2989), .Z(n573_adj_2949)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_6_i573_3_lut_4_lut.init = 16'hf909;
    LUT4 i20261_3_lut (.A(n85), .B(n26625), .C(index_i[3]), .Z(n22600)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20261_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_7_i45_3_lut_3_lut_rep_652_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26612)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_7_i45_3_lut_3_lut_rep_652_3_lut.init = 16'h3939;
    LUT4 i20260_3_lut (.A(n29169), .B(n26630), .C(index_i[3]), .Z(n22599)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20260_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_8_i46_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n46)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (B (C)+!B !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_8_i46_3_lut_4_lut_4_lut_4_lut.init = 16'hc1f0;
    LUT4 mux_193_Mux_5_i109_3_lut_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .Z(n109_adj_2901)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_5_i109_3_lut_3_lut_3_lut.init = 16'h3939;
    LUT4 mux_193_Mux_5_i572_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n572_adj_2978)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A !(B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_5_i572_3_lut_4_lut_4_lut.init = 16'ha9a5;
    PFUMX i24497 (.BLUT(n26790), .ALUT(n26791), .C0(index_i[0]), .Z(n26792));
    LUT4 mux_193_Mux_0_i635_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n635_adj_2849)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i635_3_lut_4_lut_4_lut.init = 16'hfd0a;
    LUT4 i20259_3_lut (.A(n29193), .B(n29191), .C(index_i[3]), .Z(n22598)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20259_3_lut.init = 16'hcaca;
    PFUMX i22653 (.BLUT(n24197), .ALUT(n24196), .C0(index_i[5]), .Z(n24198));
    LUT4 n133_bdd_3_lut_23801_4_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .Z(n24807)) /* synthesis lut_function=(A (B)+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n133_bdd_3_lut_23801_4_lut_3_lut.init = 16'hd9d9;
    LUT4 n627_bdd_3_lut_23940_4_lut_4_lut (.A(index_i[2]), .B(n85), .C(index_i[3]), 
         .D(n26624), .Z(n25667)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B ((D)+!C)+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n627_bdd_3_lut_23940_4_lut_4_lut.init = 16'h5c0c;
    LUT4 mux_193_Mux_9_i62_3_lut_4_lut_then_4_lut (.A(index_i[4]), .B(index_i[2]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n26859)) /* synthesis lut_function=(!(A (B (C+(D)))+!A (B+(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_9_i62_3_lut_4_lut_then_4_lut.init = 16'h222b;
    LUT4 mux_193_Mux_0_i316_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n316_adj_2912)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+(D)))+!A (B (C+(D))+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i316_3_lut_4_lut_4_lut_4_lut.init = 16'h332d;
    LUT4 mux_193_Mux_0_i715_3_lut_3_lut_rep_696 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26656)) /* synthesis lut_function=(A (B (C))+!A !(B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i715_3_lut_3_lut_rep_696.init = 16'h9595;
    L6MUX21 i12933359_i1 (.D0(n22891), .D1(n23106), .SD(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2127[0]));
    LUT4 mux_193_Mux_9_i62_3_lut_4_lut_else_4_lut (.A(index_i[4]), .B(index_i[2]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n26858)) /* synthesis lut_function=((B+(C (D)))+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_9_i62_3_lut_4_lut_else_4_lut.init = 16'hfddd;
    LUT4 mux_193_Mux_6_i645_3_lut_4_lut_3_lut_rep_698 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26658)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_6_i645_3_lut_4_lut_3_lut_rep_698.init = 16'h1919;
    LUT4 mux_193_Mux_7_i77_3_lut_3_lut_rep_699 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26659)) /* synthesis lut_function=(A (B)+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_7_i77_3_lut_3_lut_rep_699.init = 16'h9c9c;
    LUT4 mux_193_Mux_0_i660_3_lut_rep_700 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26660)) /* synthesis lut_function=(A (B)+!A (B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i660_3_lut_rep_700.init = 16'hc9c9;
    LUT4 mux_193_Mux_4_i491_3_lut_4_lut_4_lut (.A(index_i[2]), .B(n26625), 
         .C(index_i[3]), .D(n26627), .Z(n491_adj_2906)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_4_i491_3_lut_4_lut_4_lut.init = 16'hfc5c;
    LUT4 mux_193_Mux_6_i356_3_lut_4_lut_3_lut_rep_701 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26661)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_6_i356_3_lut_4_lut_3_lut_rep_701.init = 16'h4949;
    LUT4 mux_193_Mux_4_i262_3_lut_3_lut_rep_702 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26662)) /* synthesis lut_function=(A (B+(C))+!A !(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_4_i262_3_lut_3_lut_rep_702.init = 16'ha9a9;
    LUT4 mux_193_Mux_3_i676_3_lut_4_lut_3_lut_rep_703 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26663)) /* synthesis lut_function=(A (B (C))+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_3_i676_3_lut_4_lut_3_lut_rep_703.init = 16'h9494;
    LUT4 mux_193_Mux_6_i564_3_lut_4_lut_3_lut_rep_704 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26664)) /* synthesis lut_function=(A (B)+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_6_i564_3_lut_4_lut_3_lut_rep_704.init = 16'hd9d9;
    LUT4 i22122_3_lut (.A(n11840), .B(n892_adj_2854), .C(index_i[6]), 
         .Z(n22100)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22122_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_6_i572_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n572_adj_2989)) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_6_i572_3_lut_4_lut.init = 16'hccd9;
    LUT4 index_i_6__bdd_4_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[6]), 
         .C(index_i[5]), .D(n26498), .Z(n24877)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (D))+!A (B (C (D))+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam index_i_6__bdd_4_lut_4_lut_4_lut.init = 16'h04f7;
    LUT4 n676_bdd_3_lut_24001_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n25434)) /* synthesis lut_function=(A (B (C+(D)))+!A (B ((D)+!C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n676_bdd_3_lut_24001_4_lut.init = 16'hcc94;
    LUT4 mux_193_Mux_3_i684_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[4]), .Z(n684_adj_2968)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A !(B ((D)+!C)+!B (C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_3_i684_3_lut_3_lut_4_lut.init = 16'h5594;
    LUT4 mux_193_Mux_2_i653_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n653_adj_2858)) /* synthesis lut_function=(A (B (C+!(D))+!B !(D))+!A !(B (C+!(D))+!B !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_2_i653_3_lut_4_lut.init = 16'h94aa;
    PFUMX i18846 (.BLUT(n21164), .ALUT(n21165), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2127[11]));
    LUT4 mux_193_Mux_3_i397_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n397_adj_2826)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !(B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_3_i397_3_lut_4_lut_4_lut.init = 16'ha95a;
    LUT4 i19120_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21440)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A !(B (D)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19120_3_lut_3_lut_4_lut.init = 16'ha955;
    LUT4 i19165_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21485)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (D))+!A !(B (C (D))+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19165_3_lut_3_lut_4_lut.init = 16'h4933;
    LUT4 i19199_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21519)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C+(D)))+!A (B (C)+!B !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19199_3_lut_4_lut_4_lut.init = 16'hc95a;
    LUT4 n12049_bdd_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[4]), 
         .D(index_i[2]), .Z(n25691)) /* synthesis lut_function=(A (B)+!A !(B (D)+!B !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n12049_bdd_3_lut_4_lut.init = 16'h98cc;
    LUT4 i19133_3_lut_4_lut_4_lut (.A(index_i[2]), .B(n141), .C(index_i[3]), 
         .D(n26624), .Z(n21453)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19133_3_lut_4_lut_4_lut.init = 16'hc5c0;
    LUT4 mux_193_Mux_3_i859_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n859_adj_2915)) /* synthesis lut_function=(!(A (B (D)+!B !(D))+!A (B (C+(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_3_i859_3_lut_3_lut_4_lut.init = 16'h339c;
    LUT4 i18826_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21146)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(D))+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18826_3_lut_3_lut_4_lut.init = 16'h3319;
    LUT4 mux_193_Mux_0_i762_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n762_adj_2883)) /* synthesis lut_function=(A (B+!((D)+!C))+!A !(B (D)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i762_3_lut_4_lut_4_lut.init = 16'h98fc;
    LUT4 mux_193_Mux_1_i93_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n93_adj_2919)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C+(D)))+!A !(B (C (D)+!C !(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_1_i93_3_lut_4_lut_4_lut.init = 16'h955a;
    LUT4 i19189_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21509)) /* synthesis lut_function=(A (B (C)+!B (C (D)+!C !(D)))+!A !(B (C+!(D))+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19189_3_lut_4_lut_4_lut.init = 16'ha593;
    LUT4 i11435_2_lut_rep_705 (.A(index_i[0]), .B(index_i[1]), .Z(n26665)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11435_2_lut_rep_705.init = 16'h2222;
    LUT4 mux_193_Mux_6_i157_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n157_adj_2941)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (D))+!A !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_6_i157_3_lut_4_lut_4_lut_4_lut.init = 16'h5d22;
    PFUMX i19845 (.BLUT(n22182), .ALUT(n22183), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2127[2]));
    LUT4 mux_193_Mux_4_i205_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n205)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_4_i205_3_lut_4_lut_4_lut.init = 16'h5a2a;
    LUT4 mux_193_Mux_4_i900_3_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n900)) /* synthesis lut_function=(A ((C)+!B)+!A !(B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_4_i900_3_lut_4_lut_3_lut.init = 16'hb2b2;
    LUT4 mux_193_Mux_7_i506_3_lut_4_lut_4_lut (.A(index_i[2]), .B(n26625), 
         .C(index_i[3]), .D(n26624), .Z(n506_adj_2807)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B ((D)+!C)+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_7_i506_3_lut_4_lut_4_lut.init = 16'h5c0c;
    LUT4 i19124_3_lut (.A(n325), .B(n26660), .C(index_i[3]), .Z(n21444)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19124_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_0_i985_3_lut_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n985)) /* synthesis lut_function=(!(A (B+!(C))+!A (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i985_3_lut_3_lut_3_lut.init = 16'h2525;
    LUT4 i21327_3_lut (.A(n21443), .B(n21444), .C(index_i[4]), .Z(n21445)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21327_3_lut.init = 16'hcaca;
    LUT4 i19121_3_lut (.A(n26663), .B(n26677), .C(index_i[3]), .Z(n21441)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19121_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_5_i924_4_lut_3_lut (.A(index_i[2]), .B(n14741), .C(index_i[4]), 
         .Z(n924_adj_2795)) /* synthesis lut_function=(!(A (B+(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_5_i924_4_lut_3_lut.init = 16'h5656;
    LUT4 mux_193_Mux_6_i70_3_lut_rep_706 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26666)) /* synthesis lut_function=(!(A (B+(C))+!A !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_6_i70_3_lut_rep_706.init = 16'h5252;
    PFUMX i19852 (.BLUT(n22189), .ALUT(n22190), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2127[9]));
    LUT4 mux_193_Mux_0_i490_3_lut_4_lut_3_lut_rep_707 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26667)) /* synthesis lut_function=(!(A (B+!(C))+!A ((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i490_3_lut_4_lut_3_lut_rep_707.init = 16'h2424;
    LUT4 mux_193_Mux_0_i627_3_lut_rep_657 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26617)) /* synthesis lut_function=(A (B+!(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i627_3_lut_rep_657.init = 16'hdada;
    LUT4 mux_193_Mux_0_i165_3_lut_4_lut_3_lut_rep_709 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26669)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i165_3_lut_4_lut_3_lut_rep_709.init = 16'h9292;
    LUT4 i19135_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21455)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C))+!A !(B ((D)+!C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19135_3_lut_4_lut_4_lut.init = 16'h925a;
    LUT4 mux_193_Mux_0_i812_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n812)) /* synthesis lut_function=(A (B (C+(D))+!B !(C))+!A (B (D)+!B !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i812_3_lut_4_lut_4_lut_4_lut.init = 16'hcf92;
    LUT4 i19078_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21398)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A !(B (C+!(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19078_3_lut_4_lut_4_lut.init = 16'ha52b;
    LUT4 mux_193_Mux_0_i491_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n491_adj_2990)) /* synthesis lut_function=(!(A (B (D)+!B !(C+!(D)))+!A ((C+!(D))+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i491_3_lut_4_lut.init = 16'h24aa;
    LUT4 i19162_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21482)) /* synthesis lut_function=(!(A (B (C (D))+!B (C (D)+!C !(D)))+!A !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19162_3_lut_4_lut_4_lut.init = 16'h5aad;
    LUT4 i19184_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21504)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C))+!A !(B (C)+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19184_3_lut_4_lut_4_lut.init = 16'h5ad3;
    LUT4 i22247_3_lut (.A(n24200), .B(n22188), .C(index_i[8]), .Z(n22190)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22247_3_lut.init = 16'hcaca;
    LUT4 i21332_3_lut (.A(n21437), .B(n21438), .C(index_i[4]), .Z(n21439)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21332_3_lut.init = 16'hcaca;
    LUT4 n316_bdd_3_lut_24411_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n25249)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A !(B ((D)+!C)+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n316_bdd_3_lut_24411_3_lut_4_lut.init = 16'h552c;
    CCU2D unary_minus_10_add_3_9 (.A0(quarter_wave_sample_register_i[7]), 
          .B0(GND_net), .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[8]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17394), .COUT(n17395), 
          .S0(o_val_pipeline_i_0__15__N_2158[7]), .S1(o_val_pipeline_i_0__15__N_2158[8]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam unary_minus_10_add_3_9.INIT0 = 16'hf555;
    defparam unary_minus_10_add_3_9.INIT1 = 16'hf555;
    defparam unary_minus_10_add_3_9.INJECT1_0 = "NO";
    defparam unary_minus_10_add_3_9.INJECT1_1 = "NO";
    LUT4 mux_193_Mux_3_i62_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[4]), .D(n812_adj_2924), .Z(n62_adj_2980)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_3_i62_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_193_Mux_3_i94_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[4]), .D(n93_adj_2829), .Z(n94_adj_2981)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_3_i94_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_193_Mux_2_i348_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n348_adj_2987)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_2_i348_3_lut_4_lut_4_lut.init = 16'h52a5;
    LUT4 i18805_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21125)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C))+!A !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18805_3_lut_4_lut_4_lut.init = 16'h5a52;
    LUT4 index_i_1__bdd_4_lut_25416 (.A(index_i[1]), .B(index_i[0]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n26773)) /* synthesis lut_function=(!(A (B (D)+!B (C+!(D)))+!A !(B (C (D)+!C !(D))+!B !((D)+!C)))) */ ;
    defparam index_i_1__bdd_4_lut_25416.init = 16'h429c;
    LUT4 mux_193_Mux_11_i766_3_lut (.A(n638), .B(n765), .C(index_i[7]), 
         .Z(n766)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_11_i766_3_lut.init = 16'h3a3a;
    LUT4 i4410_2_lut_rep_710 (.A(index_i[0]), .B(index_i[1]), .Z(n26670)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i4410_2_lut_rep_710.init = 16'h6666;
    LUT4 index_i_0__bdd_4_lut_25039 (.A(index_i[0]), .B(index_i[3]), .C(index_i[1]), 
         .D(index_i[2]), .Z(n26769)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C (D)))+!A !(B (C+!(D))+!B !(C+(D))))) */ ;
    defparam index_i_0__bdd_4_lut_25039.init = 16'h4ae7;
    LUT4 i12116_2_lut (.A(index_i[1]), .B(index_i[3]), .Z(n541)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i12116_2_lut.init = 16'h1111;
    LUT4 mux_193_Mux_0_i157_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n157_adj_2991)) /* synthesis lut_function=(A (B (C+!(D))+!B !(D))+!A (B (D)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i157_3_lut_4_lut.init = 16'hd4aa;
    LUT4 i9458_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(n26596), .D(index_i[4]), .Z(n221)) /* synthesis lut_function=(!(A (B)+!A (B (C+(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9458_3_lut_4_lut_4_lut_4_lut.init = 16'h3336;
    LUT4 i9478_3_lut_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[4]), .D(index_i[3]), .Z(n444_adj_2988)) /* synthesis lut_function=(!(A (B)+!A !(B (C (D))+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9478_3_lut_3_lut_4_lut_4_lut.init = 16'h6333;
    LUT4 mux_190_i15_3_lut (.A(quarter_wave_sample_register_i[14]), .B(o_val_pipeline_i_0__15__N_2158[14]), 
         .C(phase_negation_i[1]), .Z(n1086[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam mux_190_i15_3_lut.init = 16'hcaca;
    LUT4 i19099_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21419)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19099_3_lut_4_lut_4_lut.init = 16'hda5a;
    LUT4 i9444_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n526_adj_2929)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+(D)))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9444_3_lut_4_lut_4_lut.init = 16'h666c;
    LUT4 mux_193_Mux_7_i108_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n108)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_7_i108_3_lut_3_lut.init = 16'hc6c6;
    LUT4 mux_193_Mux_5_i828_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[4]), .D(n26575), .Z(n828_adj_2964)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_5_i828_4_lut_4_lut.init = 16'hc66c;
    LUT4 n61_bdd_3_lut_24080_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n25415)) /* synthesis lut_function=(!(A (B)+!A !(B (C+(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n61_bdd_3_lut_24080_4_lut_4_lut_4_lut.init = 16'h6663;
    LUT4 i11436_2_lut_rep_660 (.A(index_i[0]), .B(index_i[1]), .Z(n26620)) /* synthesis lut_function=(A+!(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11436_2_lut_rep_660.init = 16'hbbbb;
    LUT4 mux_193_Mux_0_i645_3_lut_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n645)) /* synthesis lut_function=(!(A (B)+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i645_3_lut_3_lut_3_lut.init = 16'h6363;
    LUT4 mux_193_Mux_1_i882_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n882)) /* synthesis lut_function=(A ((C)+!B)+!A !((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_1_i882_3_lut_3_lut.init = 16'ha6a6;
    LUT4 i4399_2_lut_rep_626 (.A(index_i[0]), .B(index_i[2]), .Z(n26586)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i4399_2_lut_rep_626.init = 16'h6666;
    LUT4 mux_193_Mux_2_i731_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n731_adj_2856)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_2_i731_3_lut_4_lut_4_lut.init = 16'h6cc6;
    LUT4 i19112_3_lut (.A(n26621), .B(n26666), .C(index_i[3]), .Z(n21432)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19112_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_1_i62_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[4]), .D(index_i[3]), .Z(n62_adj_2953)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))+!A !(B (C)+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_1_i62_3_lut_4_lut_4_lut.init = 16'ha5a6;
    LUT4 i19111_3_lut (.A(n26676), .B(n26661), .C(index_i[3]), .Z(n21431)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19111_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_4_i349_3_lut_4_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[4]), .D(n348_adj_2961), .Z(n349_adj_2975)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_4_i349_3_lut_4_lut.init = 16'hf606;
    LUT4 i9602_3_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[4]), 
         .Z(n12052)) /* synthesis lut_function=(!(A (B)+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9602_3_lut_4_lut_3_lut.init = 16'h6262;
    LUT4 mux_193_Mux_3_i507_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[4]), .D(n491_adj_2805), .Z(n507_adj_2985)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_3_i507_3_lut_4_lut.init = 16'h6f60;
    LUT4 i21338_3_lut (.A(n21431), .B(n21432), .C(index_i[4]), .Z(n21433)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21338_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_0_i588_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n588)) /* synthesis lut_function=(!(A (B+(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i588_3_lut_3_lut.init = 16'h5656;
    LUT4 mux_193_Mux_6_i325_3_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n325)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_6_i325_3_lut_4_lut_3_lut.init = 16'h6d6d;
    LUT4 i15400_3_lut_3_lut (.A(index_i[0]), .B(index_i[2]), .C(index_i[3]), 
         .Z(n17550)) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i15400_3_lut_3_lut.init = 16'h6a6a;
    LUT4 n273_bdd_3_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .Z(n26085)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n273_bdd_3_lut_4_lut_3_lut.init = 16'h6161;
    LUT4 i19109_3_lut (.A(n29199), .B(n26658), .C(index_i[3]), .Z(n21429)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19109_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_0_i747_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n747_adj_2882)) /* synthesis lut_function=(!(A (B+!(C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i747_3_lut_4_lut_4_lut_4_lut.init = 16'h6556;
    LUT4 mux_193_Mux_4_i828_3_lut_4_lut (.A(index_i[4]), .B(index_i[3]), 
         .C(n812_adj_2977), .D(n29168), .Z(n828_adj_2976)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_4_i828_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i19108_3_lut (.A(n26630), .B(n85), .C(index_i[3]), .Z(n21428)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19108_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_5_i797_3_lut_4_lut (.A(index_i[4]), .B(index_i[3]), 
         .C(n26754), .D(n26679), .Z(n797_adj_2963)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_5_i797_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_193_Mux_1_i763_3_lut_4_lut (.A(index_i[4]), .B(index_i[3]), 
         .C(n26828), .D(n26679), .Z(n763_adj_2809)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_1_i763_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i21340_3_lut (.A(n21428), .B(n21429), .C(index_i[4]), .Z(n21430)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21340_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_6_i7_3_lut_4_lut_3_lut_rep_712 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26672)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_6_i7_3_lut_4_lut_3_lut_rep_712.init = 16'hd6d6;
    LUT4 mux_193_Mux_0_i123_3_lut_3_lut_rep_713 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26673)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i123_3_lut_3_lut_rep_713.init = 16'h6c6c;
    LUT4 mux_193_Mux_5_i754_3_lut_4_lut_3_lut_rep_714 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26674)) /* synthesis lut_function=(!(A (B)+!A ((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_5_i754_3_lut_4_lut_3_lut_rep_714.init = 16'h2626;
    LUT4 mux_193_Mux_0_i134_3_lut_4_lut_3_lut_rep_715 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26675)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i134_3_lut_4_lut_3_lut_rep_715.init = 16'h6969;
    LUT4 mux_193_Mux_0_i963_3_lut_3_lut_3_lut_rep_716 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26676)) /* synthesis lut_function=(!(A (B)+!A (B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i963_3_lut_3_lut_3_lut_rep_716.init = 16'h3636;
    LUT4 mux_193_Mux_0_i396_3_lut_4_lut_3_lut_rep_717 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26677)) /* synthesis lut_function=(A ((C)+!B)+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i396_3_lut_4_lut_3_lut_rep_717.init = 16'hb6b6;
    LUT4 mux_193_Mux_5_i459_3_lut_4_lut_3_lut_rep_718 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26678)) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_5_i459_3_lut_4_lut_3_lut_rep_718.init = 16'h6b6b;
    LUT4 mux_193_Mux_6_i442_rep_719 (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .Z(n26679)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_6_i442_rep_719.init = 16'h6464;
    PFUMX i20526 (.BLUT(n142_adj_2992), .ALUT(n157_adj_2991), .C0(index_i[4]), 
          .Z(n22865));
    LUT4 mux_193_Mux_5_i53_3_lut_4_lut_3_lut_rep_720 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26680)) /* synthesis lut_function=(A ((C)+!B)+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_5_i53_3_lut_4_lut_3_lut_rep_720.init = 16'he6e6;
    L6MUX21 i23754 (.D0(n25437), .D1(n25435), .SD(index_i[5]), .Z(n25438));
    LUT4 mux_193_Mux_0_i525_3_lut_3_lut_rep_721 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26681)) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i525_3_lut_3_lut_rep_721.init = 16'h6a6a;
    PFUMX i23752 (.BLUT(n25436), .ALUT(n21501), .C0(index_i[4]), .Z(n25437));
    PFUMX i24493 (.BLUT(n26784), .ALUT(n26785), .C0(index_i[1]), .Z(n26786));
    LUT4 mux_193_Mux_6_i134_3_lut_4_lut_3_lut_rep_722 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26682)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_6_i134_3_lut_4_lut_3_lut_rep_722.init = 16'h9696;
    LUT4 i19181_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21501)) /* synthesis lut_function=(A (B (C+(D))+!B ((D)+!C))+!A !(B (C+(D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19181_3_lut_4_lut.init = 16'haa96;
    LUT4 mux_193_Mux_2_i491_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n491_adj_2986)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A !(B (C)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_2_i491_3_lut_4_lut_4_lut.init = 16'h6a5a;
    LUT4 mux_193_Mux_6_i635_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n635_adj_2904)) /* synthesis lut_function=(A (B (C+(D))+!B !(D))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_6_i635_3_lut_4_lut.init = 16'hcce6;
    PFUMX i23750 (.BLUT(n25434), .ALUT(n25433), .C0(index_i[4]), .Z(n25435));
    L6MUX21 i22829 (.D0(n24429), .D1(n24427), .SD(index_i[6]), .Z(n24430));
    LUT4 i19093_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21413)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19093_3_lut_4_lut.init = 16'h64cc;
    PFUMX i20527 (.BLUT(n173_adj_2917), .ALUT(n188), .C0(index_i[4]), 
          .Z(n22866));
    LUT4 mux_193_Mux_5_i460_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n460_adj_2895)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A !(B (C)+!B !(C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_5_i460_3_lut_4_lut_4_lut.init = 16'h6b5a;
    LUT4 mux_193_Mux_1_i301_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n301_adj_2982)) /* synthesis lut_function=(A (B (C+(D))+!B !(D))+!A !(B (C+(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_1_i301_3_lut_4_lut_4_lut.init = 16'h99b6;
    PFUMX i22827 (.BLUT(n24428), .ALUT(n62), .C0(index_i[5]), .Z(n24429));
    LUT4 mux_193_Mux_6_i475_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n475_adj_2859)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A !(B (C+(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_6_i475_3_lut_4_lut_4_lut.init = 16'h9936;
    LUT4 mux_193_Mux_0_i142_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n142_adj_2992)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C))+!A !(B (C (D)+!C !(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i142_3_lut_4_lut_4_lut.init = 16'ha569;
    LUT4 i20255_3_lut (.A(n26612), .B(n29191), .C(index_i[3]), .Z(n22594)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20255_3_lut.init = 16'hcaca;
    LUT4 i19126_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21446)) /* synthesis lut_function=(!(A (B)+!A (B (C+(D))+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19126_3_lut_3_lut_4_lut.init = 16'h3326;
    LUT4 mux_193_Mux_0_i124_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n124_adj_2803)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A !(B (D)+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i124_3_lut_4_lut_4_lut.init = 16'h6c99;
    LUT4 i1_3_lut_4_lut_adj_86 (.A(n26377), .B(index_i[5]), .C(index_i[8]), 
         .D(n19553), .Z(n19900)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i1_3_lut_4_lut_adj_86.init = 16'hfff8;
    LUT4 n20957_bdd_3_lut_23638_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n24792)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C))+!A !(B (C+!(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n20957_bdd_3_lut_23638_4_lut_4_lut.init = 16'h5ad6;
    LUT4 i20254_3_lut (.A(n29169), .B(n108), .C(index_i[3]), .Z(n22593)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20254_3_lut.init = 16'hcaca;
    PFUMX i20532 (.BLUT(n333_adj_2993), .ALUT(n348), .C0(index_i[4]), 
          .Z(n22871));
    LUT4 i18842_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21162)) /* synthesis lut_function=(A (B (C)+!B !(C (D)+!C !(D)))+!A (B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18842_3_lut_4_lut_4_lut.init = 16'hd6a5;
    L6MUX21 i23735 (.D0(n25416), .D1(n25414), .SD(index_i[4]), .Z(n25417));
    PFUMX i23733 (.BLUT(n26396), .ALUT(n25415), .C0(index_i[5]), .Z(n25416));
    LUT4 i9466_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n11912)) /* synthesis lut_function=(!(A (B (D)+!B (C+!(D)))+!A !(B (D)+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9466_3_lut_4_lut_4_lut.init = 16'h4699;
    PFUMX i20533 (.BLUT(n364), .ALUT(n379), .C0(index_i[4]), .Z(n22872));
    PFUMX i23731 (.BLUT(n25413), .ALUT(n25412), .C0(index_i[5]), .Z(n25414));
    LUT4 mux_193_Mux_5_i30_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n30_adj_2907)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A (B+!(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_5_i30_3_lut_4_lut.init = 16'hcc67;
    PFUMX i20534 (.BLUT(n397_adj_2801), .ALUT(n412), .C0(index_i[4]), 
          .Z(n22873));
    PFUMX i20535 (.BLUT(n428), .ALUT(n443), .C0(index_i[4]), .Z(n22874));
    LUT4 i20253_3_lut (.A(n85), .B(n26630), .C(index_i[3]), .Z(n22592)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20253_3_lut.init = 16'hcaca;
    PFUMX i20536 (.BLUT(n460), .ALUT(n475_adj_2804), .C0(index_i[4]), 
          .Z(n22875));
    PFUMX i20537 (.BLUT(n491_adj_2990), .ALUT(n11000), .C0(index_i[4]), 
          .Z(n22876));
    LUT4 i20252_3_lut (.A(n645), .B(n26659), .C(index_i[3]), .Z(n22591)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20252_3_lut.init = 16'hcaca;
    LUT4 i19764_3_lut (.A(n22096), .B(n22097), .C(index_i[7]), .Z(n22103)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19764_3_lut.init = 16'hcaca;
    PFUMX i22648 (.BLUT(n21224), .ALUT(n24191), .C0(index_i[6]), .Z(n24192));
    LUT4 i19763_3_lut (.A(n22094), .B(n24879), .C(index_i[7]), .Z(n22102)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19763_3_lut.init = 16'hcaca;
    LUT4 index_i_0__bdd_4_lut_24483 (.A(index_i[0]), .B(index_i[3]), .C(index_i[1]), 
         .D(index_i[2]), .Z(n26764)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C))+!A (B (C (D)+!C !(D))+!B !(C+!(D))))) */ ;
    defparam index_i_0__bdd_4_lut_24483.init = 16'h16d3;
    PFUMX mux_193_Mux_13_i1023 (.BLUT(n511), .ALUT(n19900), .C0(index_i[9]), 
          .Z(quarter_wave_sample_register_i_15__N_2127[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 i19100_3_lut (.A(n26677), .B(n325), .C(index_i[3]), .Z(n21420)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19100_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_0_i219_3_lut_3_lut_3_lut_rep_800 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29179)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i219_3_lut_3_lut_3_lut_rep_800.init = 16'h9393;
    PFUMX i22825 (.BLUT(n24426), .ALUT(n24425), .C0(index_i[5]), .Z(n24427));
    PFUMX i23700 (.BLUT(n25382), .ALUT(n26586), .C0(index_i[4]), .Z(n25383));
    LUT4 i21371_3_lut (.A(n21419), .B(n21420), .C(index_i[4]), .Z(n21421)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21371_3_lut.init = 16'hcaca;
    LUT4 i19096_3_lut (.A(n588), .B(n26681), .C(index_i[3]), .Z(n21416)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19096_3_lut.init = 16'hcaca;
    LUT4 i19768_3_lut (.A(n22104), .B(n22105), .C(index_i[8]), .Z(n22107)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19768_3_lut.init = 16'hcaca;
    LUT4 i11284_2_lut_rep_636 (.A(index_i[2]), .B(index_i[3]), .Z(n26596)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11284_2_lut_rep_636.init = 16'h8888;
    LUT4 i23322_then_4_lut (.A(index_i[0]), .B(index_i[4]), .C(index_i[1]), 
         .D(index_i[3]), .Z(n26766)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam i23322_then_4_lut.init = 16'h3c69;
    LUT4 i11816_2_lut_rep_481_3_lut (.A(index_i[2]), .B(index_i[3]), .C(index_i[1]), 
         .Z(n26441)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11816_2_lut_rep_481_3_lut.init = 16'h8080;
    LUT4 i20185_3_lut_3_lut_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[4]), .D(index_i[1]), .Z(n22524)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20185_3_lut_3_lut_3_lut_4_lut.init = 16'h878f;
    LUT4 mux_190_i13_3_lut (.A(quarter_wave_sample_register_i[12]), .B(o_val_pipeline_i_0__15__N_2158[12]), 
         .C(phase_negation_i[1]), .Z(n1086[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam mux_190_i13_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_7_i924_3_lut_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[4]), .D(n26624), .Z(n924)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_7_i924_3_lut_3_lut_4_lut.init = 16'h878f;
    LUT4 i11231_2_lut_rep_446_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[4]), .D(n26624), .Z(n26406)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11231_2_lut_rep_446_3_lut_4_lut.init = 16'hf8f0;
    LUT4 i19714_1_lut_2_lut (.A(index_i[2]), .B(index_i[3]), .Z(n22053)) /* synthesis lut_function=(!(A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19714_1_lut_2_lut.init = 16'h7777;
    LUT4 i11213_2_lut_rep_445_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[4]), .D(n26627), .Z(n26405)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11213_2_lut_rep_445_3_lut_4_lut.init = 16'hf8f0;
    LUT4 i11819_2_lut_2_lut_3_lut (.A(index_i[2]), .B(index_i[3]), .C(index_i[0]), 
         .Z(n14379)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11819_2_lut_2_lut_3_lut.init = 16'h0808;
    L6MUX21 i22783 (.D0(n24372), .D1(n26345), .SD(index_i[6]), .Z(n24373));
    LUT4 i11310_3_lut_3_lut (.A(index_i[1]), .B(index_i[0]), .C(index_i[2]), 
         .Z(n85)) /* synthesis lut_function=(!(A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11310_3_lut_3_lut.init = 16'h7575;
    PFUMX i22781 (.BLUT(n24371), .ALUT(n26371), .C0(index_i[7]), .Z(n24372));
    LUT4 i12291_2_lut_rep_507_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n26467)) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i12291_2_lut_rep_507_3_lut_4_lut.init = 16'he000;
    LUT4 mux_193_Mux_0_i333_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n333_adj_2993)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_0_i333_3_lut_3_lut_4_lut.init = 16'hf10e;
    LUT4 mux_193_Mux_3_i349_3_lut_3_lut (.A(index_i[1]), .B(index_i[4]), 
         .C(n348_adj_2962), .Z(n349_adj_2983)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_3_i349_3_lut_3_lut.init = 16'hd1d1;
    LUT4 n21450_bdd_3_lut_3_lut (.A(index_i[1]), .B(n526_adj_2929), .C(index_i[4]), 
         .Z(n24965)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n21450_bdd_3_lut_3_lut.init = 16'h5c5c;
    LUT4 i11242_4_lut (.A(n26507), .B(index_i[7]), .C(n892), .D(index_i[6]), 
         .Z(n1021)) /* synthesis lut_function=(A (B+(C (D)))+!A (B+(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11242_4_lut.init = 16'hfcdd;
    LUT4 i18832_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21152)) /* synthesis lut_function=(A (B (C (D))+!B !(C (D)))+!A !(B (D)+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18832_3_lut_4_lut_4_lut.init = 16'h9366;
    LUT4 i19094_3_lut (.A(n900), .B(n325), .C(index_i[3]), .Z(n21414)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19094_3_lut.init = 16'hcaca;
    LUT4 i11818_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(n26596), .C(index_i[4]), 
         .D(index_i[0]), .Z(n14378)) /* synthesis lut_function=(!(A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11818_3_lut_4_lut_4_lut_4_lut.init = 16'h55d5;
    LUT4 i20671_3_lut (.A(n23005), .B(n23006), .C(index_i[7]), .Z(n23010)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20671_3_lut.init = 16'hcaca;
    LUT4 i19087_3_lut (.A(n29199), .B(n29169), .C(index_i[3]), .Z(n21407)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19087_3_lut.init = 16'hcaca;
    LUT4 i20248_3_lut (.A(n29191), .B(n26633), .C(index_i[3]), .Z(n22587)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20248_3_lut.init = 16'hcaca;
    LUT4 i20247_3_lut (.A(n1001), .B(n26612), .C(index_i[3]), .Z(n22586)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20247_3_lut.init = 16'hcaca;
    LUT4 i20245_3_lut (.A(n26633), .B(n645), .C(index_i[3]), .Z(n22584)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20245_3_lut.init = 16'hcaca;
    L6MUX21 i23567 (.D0(n25253), .D1(n25250), .SD(index_i[5]), .Z(n25254));
    PFUMX i23565 (.BLUT(n25252), .ALUT(n25251), .C0(index_i[4]), .Z(n25253));
    LUT4 i19893_3_lut (.A(n22225), .B(n22226), .C(index_i[7]), .Z(n22232)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19893_3_lut.init = 16'hcaca;
    PFUMX i23562 (.BLUT(n25249), .ALUT(n316_adj_2912), .C0(index_i[4]), 
          .Z(n25250));
    PFUMX i22762 (.BLUT(n24344), .ALUT(n24341), .C0(index_i[6]), .Z(n24345));
    PFUMX i22760 (.BLUT(n24342), .ALUT(n954), .C0(index_i[4]), .Z(n24343));
    LUT4 i12126_1_lut_rep_408_2_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n26368)) /* synthesis lut_function=(!(A (C+(D))+!A (B (C+(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i12126_1_lut_rep_408_2_lut_3_lut_4_lut.init = 16'h010f;
    LUT4 mux_193_Mux_11_i638_4_lut_4_lut (.A(n26377), .B(index_i[5]), .C(index_i[6]), 
         .D(n26417), .Z(n638)) /* synthesis lut_function=(A (B (C (D))+!B !(C))+!A (B ((D)+!C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_11_i638_4_lut_4_lut.init = 16'hc707;
    CCU2D unary_minus_10_add_3_7 (.A0(quarter_wave_sample_register_i[5]), 
          .B0(GND_net), .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[6]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17393), .COUT(n17394), 
          .S0(o_val_pipeline_i_0__15__N_2158[5]), .S1(o_val_pipeline_i_0__15__N_2158[6]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam unary_minus_10_add_3_7.INIT0 = 16'hf555;
    defparam unary_minus_10_add_3_7.INIT1 = 16'hf555;
    defparam unary_minus_10_add_3_7.INJECT1_0 = "NO";
    defparam unary_minus_10_add_3_7.INJECT1_1 = "NO";
    PFUMX i23529 (.BLUT(n25219), .ALUT(n25218), .C0(index_i[4]), .Z(n25220));
    CCU2D unary_minus_10_add_3_5 (.A0(quarter_wave_sample_register_i[3]), 
          .B0(GND_net), .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[4]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17392), .COUT(n17393), 
          .S0(o_val_pipeline_i_0__15__N_2158[3]), .S1(o_val_pipeline_i_0__15__N_2158[4]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam unary_minus_10_add_3_5.INIT0 = 16'hf555;
    defparam unary_minus_10_add_3_5.INIT1 = 16'hf555;
    defparam unary_minus_10_add_3_5.INJECT1_0 = "NO";
    defparam unary_minus_10_add_3_5.INJECT1_1 = "NO";
    CCU2D unary_minus_10_add_3_3 (.A0(quarter_wave_sample_register_i[1]), 
          .B0(GND_net), .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[2]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17391), .COUT(n17392), 
          .S0(o_val_pipeline_i_0__15__N_2158[1]), .S1(o_val_pipeline_i_0__15__N_2158[2]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam unary_minus_10_add_3_3.INIT0 = 16'hf555;
    defparam unary_minus_10_add_3_3.INIT1 = 16'hf555;
    defparam unary_minus_10_add_3_3.INJECT1_0 = "NO";
    defparam unary_minus_10_add_3_3.INJECT1_1 = "NO";
    LUT4 mux_193_Mux_7_i572_3_lut_rep_400_3_lut_3_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n26360)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_193_Mux_7_i572_3_lut_rep_400_3_lut_3_lut_4_lut.init = 16'hfe01;
    CCU2D unary_minus_10_add_3_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(quarter_wave_sample_register_i[0]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .COUT(n17391), .S1(o_val_pipeline_i_0__15__N_2158[0]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam unary_minus_10_add_3_1.INIT0 = 16'hF000;
    defparam unary_minus_10_add_3_1.INIT1 = 16'h0aaa;
    defparam unary_minus_10_add_3_1.INJECT1_0 = "NO";
    defparam unary_minus_10_add_3_1.INJECT1_1 = "NO";
    FD1S3BX quarter_wave_sample_register_i_i14 (.D(quarter_wave_sample_register_i_15__N_2127[14]), 
            .CK(dac_clk_p_c), .PD(n26683), .Q(quarter_wave_sample_register_i[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i14.GSR = "DISABLED";
    L6MUX21 i23454 (.D0(n25150), .D1(n25147), .SD(index_i[5]), .Z(n25151));
    PFUMX i23452 (.BLUT(n25149), .ALUT(n25148), .C0(index_i[4]), .Z(n25150));
    FD1S3BX quarter_wave_sample_register_i_i13 (.D(quarter_wave_sample_register_i_15__N_2127[13]), 
            .CK(dac_clk_p_c), .PD(n26683), .Q(quarter_wave_sample_register_i[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i13.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i12 (.D(quarter_wave_sample_register_i_15__N_2127[12]), 
            .CK(dac_clk_p_c), .PD(n26683), .Q(quarter_wave_sample_register_i[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i12.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i11 (.D(quarter_wave_sample_register_i_15__N_2127[11]), 
            .CK(dac_clk_p_c), .PD(n26683), .Q(quarter_wave_sample_register_i[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i11.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i10 (.D(quarter_wave_sample_register_i_15__N_2127[10]), 
            .CK(dac_clk_p_c), .PD(n26683), .Q(quarter_wave_sample_register_i[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i10.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i9 (.D(quarter_wave_sample_register_i_15__N_2127[9]), 
            .CK(dac_clk_p_c), .PD(n26683), .Q(quarter_wave_sample_register_i[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i9.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i8 (.D(quarter_wave_sample_register_i_15__N_2127[8]), 
            .CK(dac_clk_p_c), .PD(n26683), .Q(quarter_wave_sample_register_i[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i8.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i7 (.D(quarter_wave_sample_register_i_15__N_2127[7]), 
            .CK(dac_clk_p_c), .PD(n26683), .Q(quarter_wave_sample_register_i[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i7.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i6 (.D(quarter_wave_sample_register_i_15__N_2127[6]), 
            .CK(dac_clk_p_c), .PD(n26683), .Q(quarter_wave_sample_register_i[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i6.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i5 (.D(quarter_wave_sample_register_i_15__N_2127[5]), 
            .CK(dac_clk_p_c), .PD(n26683), .Q(quarter_wave_sample_register_i[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i5.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i4 (.D(quarter_wave_sample_register_i_15__N_2127[4]), 
            .CK(dac_clk_p_c), .PD(n26683), .Q(quarter_wave_sample_register_i[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i4.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i3 (.D(quarter_wave_sample_register_i_15__N_2127[3]), 
            .CK(dac_clk_p_c), .PD(n26683), .Q(quarter_wave_sample_register_i[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i3.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i2 (.D(quarter_wave_sample_register_i_15__N_2127[2]), 
            .CK(dac_clk_p_c), .PD(n26683), .Q(quarter_wave_sample_register_i[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i2.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i1 (.D(quarter_wave_sample_register_i_15__N_2127[1]), 
            .CK(dac_clk_p_c), .PD(n26683), .Q(quarter_wave_sample_register_i[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i1.GSR = "DISABLED";
    PFUMX i23449 (.BLUT(n301), .ALUT(n25146), .C0(index_i[4]), .Z(n25147));
    
endmodule
//
// Verilog Description of module \nco(OW=12) 
//

module \nco(OW=12)  (dac_clk_p_c, n26683, increment, o_phase, GND_net) /* synthesis syn_module_defined=1 */ ;
    input dac_clk_p_c;
    input n26683;
    input [30:0]increment;
    output [11:0]o_phase;
    input GND_net;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(29[49:58])
    wire [31:0]n233;
    wire [31:0]n133;
    
    wire n17445, n17444, n17443, n17442, n17441, n17440, n17439, 
        n17438, n17437, n17436, n17435, n17434, n17433, n17432, 
        n17431;
    
    FD1S3DX phase_register_547__i0 (.D(n133[0]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(n233[0])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i0.GSR = "DISABLED";
    CCU2D phase_register_547_add_4_32 (.A0(increment[30]), .B0(o_phase[10]), 
          .C0(GND_net), .D0(GND_net), .A1(o_phase[11]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n17445), .S0(n133[30]), .S1(n133[31]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547_add_4_32.INIT0 = 16'h5666;
    defparam phase_register_547_add_4_32.INIT1 = 16'hfaaa;
    defparam phase_register_547_add_4_32.INJECT1_0 = "NO";
    defparam phase_register_547_add_4_32.INJECT1_1 = "NO";
    CCU2D phase_register_547_add_4_30 (.A0(increment[28]), .B0(o_phase[8]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[29]), .B1(o_phase[9]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17444), .COUT(n17445), .S0(n133[28]), 
          .S1(n133[29]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547_add_4_30.INIT0 = 16'h5666;
    defparam phase_register_547_add_4_30.INIT1 = 16'h5666;
    defparam phase_register_547_add_4_30.INJECT1_0 = "NO";
    defparam phase_register_547_add_4_30.INJECT1_1 = "NO";
    CCU2D phase_register_547_add_4_28 (.A0(increment[26]), .B0(o_phase[6]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[27]), .B1(o_phase[7]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17443), .COUT(n17444), .S0(n133[26]), 
          .S1(n133[27]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547_add_4_28.INIT0 = 16'h5666;
    defparam phase_register_547_add_4_28.INIT1 = 16'h5666;
    defparam phase_register_547_add_4_28.INJECT1_0 = "NO";
    defparam phase_register_547_add_4_28.INJECT1_1 = "NO";
    CCU2D phase_register_547_add_4_26 (.A0(increment[24]), .B0(o_phase[4]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[25]), .B1(o_phase[5]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17442), .COUT(n17443), .S0(n133[24]), 
          .S1(n133[25]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547_add_4_26.INIT0 = 16'h5666;
    defparam phase_register_547_add_4_26.INIT1 = 16'h5666;
    defparam phase_register_547_add_4_26.INJECT1_0 = "NO";
    defparam phase_register_547_add_4_26.INJECT1_1 = "NO";
    CCU2D phase_register_547_add_4_24 (.A0(increment[22]), .B0(o_phase[2]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[23]), .B1(o_phase[3]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17441), .COUT(n17442), .S0(n133[22]), 
          .S1(n133[23]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547_add_4_24.INIT0 = 16'h5666;
    defparam phase_register_547_add_4_24.INIT1 = 16'h5666;
    defparam phase_register_547_add_4_24.INJECT1_0 = "NO";
    defparam phase_register_547_add_4_24.INJECT1_1 = "NO";
    CCU2D phase_register_547_add_4_22 (.A0(increment[20]), .B0(o_phase[0]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[21]), .B1(o_phase[1]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17440), .COUT(n17441), .S0(n133[20]), 
          .S1(n133[21]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547_add_4_22.INIT0 = 16'h5666;
    defparam phase_register_547_add_4_22.INIT1 = 16'h5666;
    defparam phase_register_547_add_4_22.INJECT1_0 = "NO";
    defparam phase_register_547_add_4_22.INJECT1_1 = "NO";
    CCU2D phase_register_547_add_4_20 (.A0(increment[18]), .B0(n233[18]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[19]), .B1(n233[19]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17439), .COUT(n17440), .S0(n133[18]), 
          .S1(n133[19]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547_add_4_20.INIT0 = 16'h5666;
    defparam phase_register_547_add_4_20.INIT1 = 16'h5666;
    defparam phase_register_547_add_4_20.INJECT1_0 = "NO";
    defparam phase_register_547_add_4_20.INJECT1_1 = "NO";
    CCU2D phase_register_547_add_4_18 (.A0(increment[16]), .B0(n233[16]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[17]), .B1(n233[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17438), .COUT(n17439), .S0(n133[16]), 
          .S1(n133[17]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547_add_4_18.INIT0 = 16'h5666;
    defparam phase_register_547_add_4_18.INIT1 = 16'h5666;
    defparam phase_register_547_add_4_18.INJECT1_0 = "NO";
    defparam phase_register_547_add_4_18.INJECT1_1 = "NO";
    CCU2D phase_register_547_add_4_16 (.A0(increment[14]), .B0(n233[14]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[15]), .B1(n233[15]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17437), .COUT(n17438), .S0(n133[14]), 
          .S1(n133[15]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547_add_4_16.INIT0 = 16'h5666;
    defparam phase_register_547_add_4_16.INIT1 = 16'h5666;
    defparam phase_register_547_add_4_16.INJECT1_0 = "NO";
    defparam phase_register_547_add_4_16.INJECT1_1 = "NO";
    CCU2D phase_register_547_add_4_14 (.A0(increment[12]), .B0(n233[12]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[13]), .B1(n233[13]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17436), .COUT(n17437), .S0(n133[12]), 
          .S1(n133[13]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547_add_4_14.INIT0 = 16'h5666;
    defparam phase_register_547_add_4_14.INIT1 = 16'h5666;
    defparam phase_register_547_add_4_14.INJECT1_0 = "NO";
    defparam phase_register_547_add_4_14.INJECT1_1 = "NO";
    CCU2D phase_register_547_add_4_12 (.A0(increment[10]), .B0(n233[10]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[11]), .B1(n233[11]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17435), .COUT(n17436), .S0(n133[10]), 
          .S1(n133[11]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547_add_4_12.INIT0 = 16'h5666;
    defparam phase_register_547_add_4_12.INIT1 = 16'h5666;
    defparam phase_register_547_add_4_12.INJECT1_0 = "NO";
    defparam phase_register_547_add_4_12.INJECT1_1 = "NO";
    CCU2D phase_register_547_add_4_10 (.A0(increment[8]), .B0(n233[8]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[9]), .B1(n233[9]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17434), .COUT(n17435), .S0(n133[8]), 
          .S1(n133[9]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547_add_4_10.INIT0 = 16'h5666;
    defparam phase_register_547_add_4_10.INIT1 = 16'h5666;
    defparam phase_register_547_add_4_10.INJECT1_0 = "NO";
    defparam phase_register_547_add_4_10.INJECT1_1 = "NO";
    CCU2D phase_register_547_add_4_8 (.A0(increment[6]), .B0(n233[6]), .C0(GND_net), 
          .D0(GND_net), .A1(increment[7]), .B1(n233[7]), .C1(GND_net), 
          .D1(GND_net), .CIN(n17433), .COUT(n17434), .S0(n133[6]), .S1(n133[7]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547_add_4_8.INIT0 = 16'h5666;
    defparam phase_register_547_add_4_8.INIT1 = 16'h5666;
    defparam phase_register_547_add_4_8.INJECT1_0 = "NO";
    defparam phase_register_547_add_4_8.INJECT1_1 = "NO";
    CCU2D phase_register_547_add_4_6 (.A0(increment[4]), .B0(n233[4]), .C0(GND_net), 
          .D0(GND_net), .A1(increment[5]), .B1(n233[5]), .C1(GND_net), 
          .D1(GND_net), .CIN(n17432), .COUT(n17433), .S0(n133[4]), .S1(n133[5]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547_add_4_6.INIT0 = 16'h5666;
    defparam phase_register_547_add_4_6.INIT1 = 16'h5666;
    defparam phase_register_547_add_4_6.INJECT1_0 = "NO";
    defparam phase_register_547_add_4_6.INJECT1_1 = "NO";
    CCU2D phase_register_547_add_4_4 (.A0(increment[2]), .B0(n233[2]), .C0(GND_net), 
          .D0(GND_net), .A1(increment[3]), .B1(n233[3]), .C1(GND_net), 
          .D1(GND_net), .CIN(n17431), .COUT(n17432), .S0(n133[2]), .S1(n133[3]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547_add_4_4.INIT0 = 16'h5666;
    defparam phase_register_547_add_4_4.INIT1 = 16'h5666;
    defparam phase_register_547_add_4_4.INJECT1_0 = "NO";
    defparam phase_register_547_add_4_4.INJECT1_1 = "NO";
    CCU2D phase_register_547_add_4_2 (.A0(increment[0]), .B0(n233[0]), .C0(GND_net), 
          .D0(GND_net), .A1(increment[1]), .B1(n233[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n17431), .S1(n133[1]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547_add_4_2.INIT0 = 16'h7000;
    defparam phase_register_547_add_4_2.INIT1 = 16'h5666;
    defparam phase_register_547_add_4_2.INJECT1_0 = "NO";
    defparam phase_register_547_add_4_2.INJECT1_1 = "NO";
    LUT4 i15348_2_lut (.A(increment[0]), .B(n233[0]), .Z(n133[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i15348_2_lut.init = 16'h6666;
    FD1S3DX phase_register_547__i31 (.D(n133[31]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(o_phase[11])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i31.GSR = "DISABLED";
    FD1S3DX phase_register_547__i30 (.D(n133[30]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(o_phase[10])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i30.GSR = "DISABLED";
    FD1S3DX phase_register_547__i29 (.D(n133[29]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(o_phase[9])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i29.GSR = "DISABLED";
    FD1S3DX phase_register_547__i28 (.D(n133[28]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(o_phase[8])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i28.GSR = "DISABLED";
    FD1S3DX phase_register_547__i27 (.D(n133[27]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(o_phase[7])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i27.GSR = "DISABLED";
    FD1S3DX phase_register_547__i26 (.D(n133[26]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(o_phase[6])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i26.GSR = "DISABLED";
    FD1S3DX phase_register_547__i25 (.D(n133[25]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(o_phase[5])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i25.GSR = "DISABLED";
    FD1S3DX phase_register_547__i24 (.D(n133[24]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(o_phase[4])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i24.GSR = "DISABLED";
    FD1S3DX phase_register_547__i23 (.D(n133[23]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(o_phase[3])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i23.GSR = "DISABLED";
    FD1S3DX phase_register_547__i22 (.D(n133[22]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(o_phase[2])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i22.GSR = "DISABLED";
    FD1S3DX phase_register_547__i21 (.D(n133[21]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(o_phase[1])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i21.GSR = "DISABLED";
    FD1S3DX phase_register_547__i20 (.D(n133[20]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(o_phase[0])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i20.GSR = "DISABLED";
    FD1S3DX phase_register_547__i19 (.D(n133[19]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(n233[19])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i19.GSR = "DISABLED";
    FD1S3DX phase_register_547__i18 (.D(n133[18]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(n233[18])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i18.GSR = "DISABLED";
    FD1S3DX phase_register_547__i17 (.D(n133[17]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(n233[17])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i17.GSR = "DISABLED";
    FD1S3DX phase_register_547__i16 (.D(n133[16]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(n233[16])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i16.GSR = "DISABLED";
    FD1S3DX phase_register_547__i15 (.D(n133[15]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(n233[15])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i15.GSR = "DISABLED";
    FD1S3DX phase_register_547__i14 (.D(n133[14]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(n233[14])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i14.GSR = "DISABLED";
    FD1S3DX phase_register_547__i13 (.D(n133[13]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(n233[13])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i13.GSR = "DISABLED";
    FD1S3DX phase_register_547__i12 (.D(n133[12]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(n233[12])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i12.GSR = "DISABLED";
    FD1S3DX phase_register_547__i11 (.D(n133[11]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(n233[11])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i11.GSR = "DISABLED";
    FD1S3DX phase_register_547__i10 (.D(n133[10]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(n233[10])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i10.GSR = "DISABLED";
    FD1S3DX phase_register_547__i9 (.D(n133[9]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(n233[9])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i9.GSR = "DISABLED";
    FD1S3DX phase_register_547__i8 (.D(n133[8]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(n233[8])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i8.GSR = "DISABLED";
    FD1S3DX phase_register_547__i7 (.D(n133[7]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(n233[7])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i7.GSR = "DISABLED";
    FD1S3DX phase_register_547__i6 (.D(n133[6]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(n233[6])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i6.GSR = "DISABLED";
    FD1S3DX phase_register_547__i5 (.D(n133[5]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(n233[5])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i5.GSR = "DISABLED";
    FD1S3DX phase_register_547__i4 (.D(n133[4]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(n233[4])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i4.GSR = "DISABLED";
    FD1S3DX phase_register_547__i3 (.D(n133[3]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(n233[3])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i3.GSR = "DISABLED";
    FD1S3DX phase_register_547__i2 (.D(n133[2]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(n233[2])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i2.GSR = "DISABLED";
    FD1S3DX phase_register_547__i1 (.D(n133[1]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(n233[1])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i1.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module dds_U2
//

module dds_U2 (dac_clk_p_c, n26683, carrier_increment, o_dac_cw_b_c_c, 
            o_dac_b_c_7, \o_sample_i[7] , \o_sample_i[15] , \o_sample_i[14] , 
            \o_sample_i[13] , \o_sample_i[12] , \o_sample_i[11] , \o_sample_i[10] , 
            \o_sample_i[9] , \o_sample_i[8] , \quarter_wave_sample_register_q[15] , 
            n29209, o_dac_b_c_15, o_dac_b_c_14, o_dac_b_c_13, o_dac_b_c_12, 
            o_dac_b_c_11, o_dac_b_c_10, n3537, o_dac_b_c_8, GND_net) /* synthesis syn_module_defined=1 */ ;
    input dac_clk_p_c;
    input n26683;
    input [30:0]carrier_increment;
    input o_dac_cw_b_c_c;
    output o_dac_b_c_7;
    output \o_sample_i[7] ;
    output \o_sample_i[15] ;
    output \o_sample_i[14] ;
    output \o_sample_i[13] ;
    output \o_sample_i[12] ;
    output \o_sample_i[11] ;
    output \o_sample_i[10] ;
    output \o_sample_i[9] ;
    output \o_sample_i[8] ;
    output \quarter_wave_sample_register_q[15] ;
    input n29209;
    output o_dac_b_c_15;
    output o_dac_b_c_14;
    output o_dac_b_c_13;
    output o_dac_b_c_12;
    output o_dac_b_c_11;
    output o_dac_b_c_10;
    output n3537;
    output o_dac_b_c_8;
    input GND_net;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(29[49:58])
    wire o_dac_b_c_7 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire \o_sample_i[7]  /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[39:49])
    wire \o_sample_i[15]  /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[39:49])
    wire \o_sample_i[14]  /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[39:49])
    wire \o_sample_i[13]  /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[39:49])
    wire \o_sample_i[12]  /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[39:49])
    wire \o_sample_i[11]  /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[39:49])
    wire \o_sample_i[10]  /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[39:49])
    wire \o_sample_i[9]  /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[39:49])
    wire \o_sample_i[8]  /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[39:49])
    wire o_dac_b_c_15 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire o_dac_b_c_14 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire o_dac_b_c_13 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire o_dac_b_c_12 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire o_dac_b_c_11 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire o_dac_b_c_10 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire n3537 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire o_dac_b_c_8 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire [30:0]increment;   // d:/documents/git_local/fm_modulator/rtl/dds.v(14[31:40])
    wire [11:0]o_phase;   // d:/documents/git_local/fm_modulator/rtl/dds.v(18[26:33])
    
    FD1S3DX increment_i0 (.D(carrier_increment[0]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(increment[0])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i0.GSR = "DISABLED";
    FD1S3DX increment_i30 (.D(carrier_increment[30]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(increment[30])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i30.GSR = "DISABLED";
    FD1S3DX increment_i29 (.D(carrier_increment[29]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(increment[29])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i29.GSR = "DISABLED";
    FD1S3DX increment_i28 (.D(carrier_increment[28]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(increment[28])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i28.GSR = "DISABLED";
    FD1S3DX increment_i27 (.D(carrier_increment[27]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(increment[27])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i27.GSR = "DISABLED";
    FD1S3DX increment_i26 (.D(carrier_increment[26]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(increment[26])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i26.GSR = "DISABLED";
    FD1S3DX increment_i25 (.D(carrier_increment[25]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(increment[25])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i25.GSR = "DISABLED";
    FD1S3DX increment_i24 (.D(carrier_increment[24]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(increment[24])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i24.GSR = "DISABLED";
    FD1S3DX increment_i23 (.D(carrier_increment[23]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(increment[23])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i23.GSR = "DISABLED";
    FD1S3DX increment_i22 (.D(carrier_increment[22]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(increment[22])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i22.GSR = "DISABLED";
    FD1S3DX increment_i21 (.D(carrier_increment[21]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(increment[21])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i21.GSR = "DISABLED";
    FD1S3DX increment_i20 (.D(carrier_increment[20]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(increment[20])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i20.GSR = "DISABLED";
    FD1S3DX increment_i19 (.D(carrier_increment[19]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(increment[19])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i19.GSR = "DISABLED";
    FD1S3DX increment_i18 (.D(carrier_increment[18]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(increment[18])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i18.GSR = "DISABLED";
    FD1S3DX increment_i17 (.D(carrier_increment[17]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(increment[17])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i17.GSR = "DISABLED";
    FD1S3DX increment_i16 (.D(carrier_increment[16]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(increment[16])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i16.GSR = "DISABLED";
    FD1S3DX increment_i15 (.D(carrier_increment[15]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(increment[15])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i15.GSR = "DISABLED";
    FD1S3DX increment_i14 (.D(carrier_increment[14]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(increment[14])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i14.GSR = "DISABLED";
    FD1S3DX increment_i13 (.D(carrier_increment[13]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(increment[13])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i13.GSR = "DISABLED";
    FD1S3DX increment_i12 (.D(carrier_increment[12]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(increment[12])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i12.GSR = "DISABLED";
    FD1S3DX increment_i11 (.D(carrier_increment[11]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(increment[11])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i11.GSR = "DISABLED";
    FD1S3DX increment_i10 (.D(carrier_increment[10]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(increment[10])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i10.GSR = "DISABLED";
    FD1S3DX increment_i9 (.D(carrier_increment[9]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(increment[9])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i9.GSR = "DISABLED";
    FD1S3DX increment_i8 (.D(carrier_increment[8]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(increment[8])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i8.GSR = "DISABLED";
    FD1S3DX increment_i7 (.D(carrier_increment[7]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(increment[7])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i7.GSR = "DISABLED";
    FD1S3DX increment_i6 (.D(carrier_increment[6]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(increment[6])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i6.GSR = "DISABLED";
    FD1S3DX increment_i5 (.D(carrier_increment[5]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(increment[5])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i5.GSR = "DISABLED";
    FD1S3DX increment_i4 (.D(carrier_increment[4]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(increment[4])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i4.GSR = "DISABLED";
    FD1S3DX increment_i3 (.D(carrier_increment[3]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(increment[3])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i3.GSR = "DISABLED";
    FD1S3DX increment_i2 (.D(carrier_increment[2]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(increment[2])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i2.GSR = "DISABLED";
    FD1S3DX increment_i1 (.D(carrier_increment[1]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(increment[1])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=78, LSE_RLINE=78 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i1.GSR = "DISABLED";
    quarter_wave_sine_lookup_U0 qtr_inst (.dac_clk_p_c(dac_clk_p_c), .n26683(n26683), 
            .o_dac_cw_b_c_c(o_dac_cw_b_c_c), .o_phase({o_phase}), .o_dac_b_c_7(o_dac_b_c_7), 
            .\o_sample_i[7] (\o_sample_i[7] ), .\o_sample_i[15] (\o_sample_i[15] ), 
            .\o_sample_i[14] (\o_sample_i[14] ), .\o_sample_i[13] (\o_sample_i[13] ), 
            .\o_sample_i[12] (\o_sample_i[12] ), .\o_sample_i[11] (\o_sample_i[11] ), 
            .\o_sample_i[10] (\o_sample_i[10] ), .\o_sample_i[9] (\o_sample_i[9] ), 
            .\o_sample_i[8] (\o_sample_i[8] ), .\quarter_wave_sample_register_q[15] (\quarter_wave_sample_register_q[15] ), 
            .n29209(n29209), .o_dac_b_c_15(o_dac_b_c_15), .o_dac_b_c_14(o_dac_b_c_14), 
            .o_dac_b_c_13(o_dac_b_c_13), .o_dac_b_c_12(o_dac_b_c_12), .o_dac_b_c_11(o_dac_b_c_11), 
            .o_dac_b_c_10(o_dac_b_c_10), .n3537(n3537), .o_dac_b_c_8(o_dac_b_c_8), 
            .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(21[70:134])
    \nco(OW=12)_U1  nco_inst (.increment({increment}), .GND_net(GND_net), 
            .o_phase({o_phase}), .dac_clk_p_c(dac_clk_p_c), .n26683(n26683)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(20[49:100])
    
endmodule
//
// Verilog Description of module quarter_wave_sine_lookup_U0
//

module quarter_wave_sine_lookup_U0 (dac_clk_p_c, n26683, o_dac_cw_b_c_c, 
            o_phase, o_dac_b_c_7, \o_sample_i[7] , \o_sample_i[15] , 
            \o_sample_i[14] , \o_sample_i[13] , \o_sample_i[12] , \o_sample_i[11] , 
            \o_sample_i[10] , \o_sample_i[9] , \o_sample_i[8] , \quarter_wave_sample_register_q[15] , 
            n29209, o_dac_b_c_15, o_dac_b_c_14, o_dac_b_c_13, o_dac_b_c_12, 
            o_dac_b_c_11, o_dac_b_c_10, n3537, o_dac_b_c_8, GND_net) /* synthesis syn_module_defined=1 */ ;
    input dac_clk_p_c;
    input n26683;
    input o_dac_cw_b_c_c;
    input [11:0]o_phase;
    output o_dac_b_c_7;
    output \o_sample_i[7] ;
    output \o_sample_i[15] ;
    output \o_sample_i[14] ;
    output \o_sample_i[13] ;
    output \o_sample_i[12] ;
    output \o_sample_i[11] ;
    output \o_sample_i[10] ;
    output \o_sample_i[9] ;
    output \o_sample_i[8] ;
    output \quarter_wave_sample_register_q[15] ;
    input n29209;
    output o_dac_b_c_15;
    output o_dac_b_c_14;
    output o_dac_b_c_13;
    output o_dac_b_c_12;
    output o_dac_b_c_11;
    output o_dac_b_c_10;
    output n3537;
    output o_dac_b_c_8;
    input GND_net;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(29[49:58])
    wire o_dac_b_c_7 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire [15:0]\o_val_pipeline_q[0]  /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(16[24:40])
    wire \o_sample_i[7]  /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[39:49])
    wire [15:0]\o_val_pipeline_i[0]  /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(15[24:40])
    wire \o_sample_i[15]  /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[39:49])
    wire \o_sample_i[14]  /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[39:49])
    wire \o_sample_i[13]  /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[39:49])
    wire \o_sample_i[12]  /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[39:49])
    wire \o_sample_i[11]  /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[39:49])
    wire \o_sample_i[10]  /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[39:49])
    wire \o_sample_i[9]  /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[39:49])
    wire \o_sample_i[8]  /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[39:49])
    wire o_dac_b_c_15 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire o_dac_b_c_14 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire o_dac_b_c_13 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire o_dac_b_c_12 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire o_dac_b_c_11 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire o_dac_b_c_10 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire n3537 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire o_dac_b_c_8 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(24[51:61])
    wire [9:0]index_i;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(31[17:24])
    
    wire n29180, n24310, n24308, n24311, n22330, n22331, n22334, 
        n541, n890;
    wire [9:0]index_q;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(31[26:33])
    
    wire n891, n22332, n22333, n22335, n26496, n26482, n62, n22421, 
        n22422, n22426, n22858, n22859, n22860, n900, n22483, 
        n22484, n22488, n26430, n9970, n765, n93, n24456, n924, 
        n24309, n22920, n22921, n22922, n25085, n25082, n25086, 
        n22507, n22508, n22511, n14728, n252, n25553, n541_adj_2251, 
        n26697, n26709, n526, n26607, n29194, n22684, n26604, 
        n108, n22683, n22509, n22510, n22512, n653, n668, n669, 
        n70, n26541, n23107, n26538, n29190, n11873;
    wire [15:0]quarter_wave_sample_register_i;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(22[24:54])
    wire [14:0]quarter_wave_sample_register_i_15__N_2127;
    
    wire n21371, n21372, n21373, n26734, n26770, n26771, n26772, 
        n26438, n26519, n21314, n21083, n21084, n21085, n301, 
        n21047, n660, n26735, n460, n285, n476, n25072, n25069, 
        n25073, n25071, n25070, n26547, n221, n526_adj_2252, n541_adj_2253, 
        n23045, n21569, n397, n26582, n413, n26521, n316, n325;
    wire [11:0]phase_q;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(12[17:24])
    
    wire n23135, n23136, n23137, n619, n26650, n22682, n882, n860;
    wire [1:0]phase_negation_i;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(23[12:28])
    wire [11:0]phase_i;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(11[17:24])
    wire [1:0]phase_negation_q;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(23[30:46])
    wire [9:0]index_i_9__N_2107;
    wire [9:0]index_q_9__N_2117;
    wire [15:0]quarter_wave_sample_register_q;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(22[56:86])
    wire [14:0]quarter_wave_sample_register_q_15__N_2142;
    
    wire n93_adj_2254, n13857, n286, n21383, n21384, n21385, n26691, 
        n22681, n21086, n21087, n21088, n28444, n26851, n22252, 
        o_val_pipeline_i_0__15__N_2157, n24920, o_val_pipeline_i_0__15__N_2159, 
        o_val_pipeline_i_0__15__N_2161, o_val_pipeline_i_0__15__N_2163, 
        n635, n21363, n24307, n26478, o_val_pipeline_i_0__15__N_2165, 
        o_val_pipeline_i_0__15__N_2167, o_val_pipeline_i_0__15__N_2169, 
        n173, n70_adj_2255, n21386, n21387, n21388, n26736, n491, 
        n507, o_val_pipeline_i_0__15__N_2171, n542, n573, n22246, 
        n26647, n301_adj_2256, o_val_pipeline_i_0__15__N_2173, n26719, 
        n26728, n270, n23073, n23074, n23075, n747, n891_adj_2257, 
        n22717, n22718, n22722, n12058, n26737, n26740, n26720, 
        n29197, n316_adj_2258, n26485, n26820, n29200, n29182, n397_adj_2259, 
        n22501, n22502, n26649, n844, n26477, n700, n620, n635_adj_2260, 
        n636, n21033, n26750, n26605, n157, n412, n526_adj_2261, 
        n29176, n21081, n796, n931, n25068, n26648, n22677, n21114, 
        n364, n882_adj_2262, n38, n22676, n12047, n475, n396, 
        n954, n22674, n22322, n22323, n157_adj_2263;
    wire [14:0]n1703;
    
    wire n954_adj_2264, n12065, n26695, n26687, n17568, n572, n17567, 
        n26585, n828, n22281, n22282, n22291, n22285, n22286, 
        n22293, n22287, n22288, n22294, n875, n890_adj_2265, n891_adj_2266, 
        n22304, n22305, n22310, n844_adj_2267, n859, n860_adj_2268, 
        n22499, n22500, n285_adj_2269, n26598;
    wire [11:0]phase_q_11__N_2233;
    
    wire n25067, n29198, n26724, n21080, n444, n22306, n22307, 
        n22311, n21554, n21555, n21556, n26741, n26571, n781, 
        n732, n21065, n21082, n684, n700_adj_2270, n21710, n382, 
        n509, n22316, n21203, n21204, n21205, n22326, n22327, 
        n21036, n22328, n22329, n21212, n21213, n21214, n26861, 
        n26862, n62_adj_2271, n25583, n22820, n22821, n22822, n22353, 
        n22354, n22361, n22355, n22356, n22362, n26373, n20230, 
        n26486, n254, n22411, n22412, n22415, n22416, n22423, 
        n22417, n22418, n22424, n22448, n22449, n22455, n22450, 
        n22451, n22456, n22452, n22453, n22457, n22471, n22472, 
        n22482, n22473, n22474, n22479, n22480, n22486, n382_adj_2272, 
        n509_adj_2273, n22493, n22503, n22504, n22505, n22506, n21089, 
        n21090, n21091, n26761, n26762, n26763, n22943, n22944, 
        n22949, n22958, n22959, n22964, n22960, n22961, n22965, 
        n26372, n20234, n254_adj_2274, n22973, n22974, n22975, n22623, 
        n22624, n22630, n22625, n22626, n22631, n22627, n22628, 
        n22632, n26599, n22918, n22919, n22129, n22130, n22135, 
        n26748, n444_adj_2275, n22705, n22706, n22716, n22707, n22708, 
        n26855, n26856, n26857, n22713, n22714, n22720, n26718, 
        n21078, n676, n21077, n21079, n26411, n22208, n22209, 
        n22216, n22210, n22211, n22217, n747_adj_2276, n762, n763, 
        n23129, n23130, n23134, n26721, n797, n828_adj_2277, n22269, 
        n22270, n22271, n22272, n22273, n22274, n29196, n985, 
        n986, n22275, n22276, n812, n22277, n22278, n22289, n22283, 
        n22284, n22292, n12014, n21349, n22301, n29185, n971, 
        n26711, n939, n22916, n22917, n21355, n21358, n22303, 
        n574, n21361, n21364, n764, n22680, n22687, n21322, n21325, 
        n22325, n21328, n21331, n21334, n21337, n21340, n892, 
        n26584, n20006, n17544, n26849, n26850, n22816, n22817, 
        n22818, n22819, n29189, n923, n62_adj_2278, n491_adj_2279, 
        n22337, n22338, n11815, n11812, n109, n124, n21345, n21642, 
        n890_adj_2280, n364_adj_2281, n22559, n26842, n26843, n26844, 
        n844_adj_2282, n22339, n22340, n12009, n22341, n22342, n21696, 
        n26457, n189, n491_adj_2283, n22343, n22344, n11856, n26497, 
        n637, n29181, n443, n620_adj_2284, n14085, n21330, n142, 
        n716, n21063, n30, n26755, n26756, n26757, n781_adj_2285, 
        n25592, n22345, n22346, n22357, n526_adj_2286, n908, n46, 
        n428, n716_adj_2287, n541_adj_2288, n1017, n22636, n604, 
        n26622, n348, n21798, n21108, n635_adj_2289, n22349, n22350, 
        n22359, n26505, n26472, n860_adj_2290, n25274, n364_adj_2291, 
        n22538, n26593, n21621, n62_adj_2292, n21690, n12012, n404, 
        n21549, n812_adj_2293, n26835, n26836, n26837, n26359, n955, 
        n15026, n252_adj_2294, n17573, n26354, n26470, n189_adj_2295, 
        n24169, n22495, n22497, n26506, n26414, n637_adj_2296, n491_adj_2297, 
        n507_adj_2298, n26583, n21548, n26495, n22368, n22369, n22384, 
        n747_adj_2299, n22370, n22371, n22385, n22372, n22373, n22386, 
        n21663, n25272, n635_adj_2300, n30_adj_2301, n526_adj_2302, 
        n26832, n26833, n26834, n22376, n22377, n22388, n781_adj_2303, 
        n26542, n25594, n26539, n221_adj_2304, n21056, n25447, n908_adj_2305, 
        n26653, n25206, n443_adj_2306, n21807, n173_adj_2307, n22378, 
        n22379, n22389, n763_adj_2308, n24125, n25584, n22380, n22381, 
        n22390, n22382, n22383, n22391, n348_adj_2309, n349, n747_adj_2310, 
        n797_adj_2311, n828_adj_2312, n26685, n25216, n413_adj_2313, 
        n773, n25328, n173_adj_2314, n747_adj_2315, n25227, n26455, 
        n22544, n26587, n26710, n25229, n252_adj_2316, n157_adj_2317, 
        n15, n21600, n251, n413_adj_2318, n412_adj_2319, n22542, 
        n26700, n25233, n844_adj_2320, n22758, n26387, n26652, n364_adj_2321, 
        n22399, n22400, n21630, n22856, n22857, n21045, n22401, 
        n22402, n22403, n22404, n22637, n22405, n22406, n26595, 
        n22407, n22408, n22419, n22846, n22847, n22854, n22413, 
        n22414, n22852, n22853, n26388, n22638, n22432, n22433, 
        n22447, n22434, n22435, n22436, n22437, n251_adj_2322, n890_adj_2323, 
        n22438, n22439, n22440, n22441, n890_adj_2324, n22848, n27931, 
        n22855, n25209, n22851, n26725, n699, n732_adj_2325, n763_adj_2326, 
        n381, n26523, n252_adj_2327, n21721, n891_adj_2328, n22461, 
        n22462, n22477, n22465, n22466, n22467, n22468, n22475, 
        n22476, n22908, n22909, n22395, n24133, n24126, n24134, 
        n22914, n22915, n25235, n22801, n22808, n26623, n763_adj_2329, 
        n24160, n684_adj_2330, n22566, n460_adj_2331, n109_adj_2332, 
        n22639, n716_adj_2333, n491_adj_2334, n732_adj_2335, n1001, 
        n21057, n668_adj_2336, n21370, n21376, n604_adj_2337, n890_adj_2338, 
        n21379, n21382, n460_adj_2339, n11979, n731, n732_adj_2340, 
        n22796, n29187, n364_adj_2341, n22302, n22309, n26526, n445, 
        n26384, n22124, n157_adj_2342, n21544, n21559, n21562, n892_adj_2343, 
        n397_adj_2344, n252_adj_2345, n26749, n428_adj_2346, n716_adj_2347, 
        n445_adj_2348, n21537, n684_adj_2349, n22300, n22308, n21570, 
        n22313, n443_adj_2350, n29202, n21711, n379, n412_adj_2351, 
        n21719, n699_adj_2352, n26699, n25271, n24290, n26334, n24291, 
        n890_adj_2353, n443_adj_2354, n379_adj_2355, n21789, n684_adj_2356, 
        n29183, n26727, n21032, n29192, n939_adj_2357, n24360, n24168, 
        n24161, n557, n29201, n716_adj_2358, n25309, n26528, n27995, 
        n29161, n24289, n24358, n318, n731_adj_2359, n22910, n27998, 
        n25312, n22913, n21797, n22759, n21107, n26357, n506, 
        n21324, n190, n253, n22815, n21367, n526_adj_2360, n26349, 
        n26646, n700_adj_2361, n25354, n24949, n24946, n24950, n24948, 
        n24947, n25336, n21546, n699_adj_2362, n21069, n26548, n26702, 
        n21717, n731_adj_2363, n620_adj_2364, n25338, n25335, n25339, 
        n379_adj_2365, n26637, n526_adj_2366, n542_adj_2367, n21312, 
        n26823, n26824, n26825, n24945, n24944, n93_adj_2368, n24922, 
        n24923, n24921, n26545, n700_adj_2369, n25310, n204, n21545, 
        n26644, n21360, n21110, n526_adj_2370, n542_adj_2371, n931_adj_2372, 
        n188, n27993, n668_adj_2373, n24918, n24915, n24919, n21612, 
        n22675, n24917, n24916, n22931, n22932, n26701, n21687, 
        n125, n24286, n26546, n908_adj_2374, n29171, n26543, n21051, 
        n29195, n21050, n21052, n24914, n21012, n25207, n21665, 
        n22933, n22934, n22935, n22936, n22945, n22214, n24362, 
        n22219, n25265, n22642, n22956, n26167, n124_adj_2375, n22895, 
        n22937, n22938, n22946, n24912, n24910, n24913, n26732, 
        n29164, n24909, n21567, n348_adj_2376, n21819, n21662, n62_adj_2377, 
        n22212, n22213, n22218, n29162, n21048, n22221, n24911, 
        n15006, n1022, n21049, n24908, n21044, n21046, n890_adj_2378, 
        n21695, n781_adj_2379, n318_adj_2380, n14982, n765_adj_2381, 
        n1022_adj_2382, n25935, n22952, n22950, n254_adj_2383, n511;
    wire [15:0]o_val_pipeline_i_0__15__N_2158;
    
    wire n491_adj_2384, n29167, n21307, n21310, n22957, n316_adj_2385, 
        n22536, n26712, n29175, n716_adj_2386, n124_adj_2387, n21297, 
        n22539, n22540, n574_adj_2388, n21313, n491_adj_2389, n21316, 
        n764_adj_2390, n747_adj_2391, n763_adj_2392, n28282, n28283, 
        n26550, n475_adj_2393, n22546, n22547, n954_adj_2394, n22969, 
        n22970, n460_adj_2395, n22971, n22972, n25450, n9807, n26601, 
        n828_adj_2396, n444_adj_2397, n251_adj_2398, n475_adj_2399, 
        n25465, n17352, n21768, n21030, n22560, n22561, n25467, 
        n26597, n668_adj_2400, n317, n747_adj_2401, n763_adj_2402, 
        n22567, n22568, n21176, n19545, n29170, n25983, n22138, 
        n22136, n24250, n21170, n26606, n25483, n21295, n21298, 
        n22954, n22605, n22606, n22621, n22607, n22608, n22622, 
        n17351, n22609, n22610;
    wire [15:0]o_val_pipeline_q_0__15__N_2190;
    
    wire n22611, n22612, n22613, n22614, n22615, n22616, n21533, 
        n21534, n21535, n17350, n15_adj_2403, n20039, n26706, n397_adj_2404, 
        n21104, n93_adj_2405, n24441, n26561, n475_adj_2406, n29178, 
        n21035, n26794, n21327, n684_adj_2407, n29174, n476_adj_2408, 
        n24490, n24491, n931_adj_2409, n188_adj_2410, n21315, n29172, 
        n475_adj_2411, n22640, n22634, n22629, n22633, n653_adj_2412, 
        n891_adj_2413, n21329, n26845, n124_adj_2414, n22833, n22641, 
        n22962, n22963, n22966, n22117, n22118, n22119, n22120, 
        n700_adj_2415, n557_adj_2416, n572_adj_2417, n23046, n142_adj_2418, 
        n157_adj_2419, n158, n22121, n22122, n22131, n17349, n22123, 
        n22132, n24494, n557_adj_2420, n573_adj_2421, n22492, n22496, 
        n700_adj_2422, n285_adj_2423, n22535, n22459, n23061, n23062, 
        n23069, n22454, n22458, n589, n23047, n21536, n21538, 
        n125_adj_2424, n23063, n23064, n23070, n23065, n23066, n23071, 
        n23067, n23068, n23072, n21008, n21009, n21010, n124_adj_2425, 
        n24440, n157_adj_2426, n620_adj_2427, n23048, n1017_adj_2428, 
        n22364, n954_adj_2429, n22358, n22363, n22366, n22315, n22319, 
        n26821, n26822, n573_adj_2430, n17348, n29163, n21801, n22312, 
        n653_adj_2431, n397_adj_2432, n573_adj_2433, n22220, n574_adj_2434, 
        n21215, n574_adj_2435, n21206, n668_adj_2436, n23049, n23050, 
        n731_adj_2437, n23051, n21791, n763_adj_2438, n22721, n22724, 
        n21547, n762_adj_2439, n23052, n23053, n22719, n22723, n891_adj_2440, 
        n22695, n22696, n22711, n22699, n22700, n22701, n22702, 
        n22709, n22710, n21788, n21790, n812_adj_2441, n23054, n26793, 
        n21550, n498, n29173, n875_adj_2442, n23056, n26437, n924_adj_2443, 
        n956, n27885, n17347, n27886, n25591, n908_adj_2444, n23057, 
        n317_adj_2445, n15024, n23058, n21029, n381_adj_2446, n21027, 
        n21026, n22487, n22490, n22485, n22489, n21024, n23059, 
        n22425, n22428, n26569, n21015, n22427, n1002, n23060, 
        n21020, n21378, n27925, n604_adj_2447, n21773, n27926, n22365, 
        n142_adj_2448, n22295, n22296, n22298, n22297, n26841, n21769, 
        n21343, n21346, n26714, n17541, n17569, n17540, n27928, 
        n475_adj_2449, n250, n22812, n21597, n22811, n26350, n22678, 
        n22810, n22809, n684_adj_2450, n142_adj_2451, n157_adj_2452, 
        n158_adj_2453, n22679, n109_adj_2454, n125_adj_2455, n25632, 
        n22192, n22193, n22194, n22195, n22196, n22197, n22198, 
        n22199, n653_adj_2456, n22200, n22201, n22204, n22205, n21380, 
        n26745, n1002_adj_2457, n22253, n21233, n26429, n21242, 
        n506_adj_2458, n860_adj_2459, n93_adj_2460, n26746, n26747, 
        n26393, n701, n22238, n22239, n22254, n21066, n21067, 
        n27992, n22240, n22241, n22255, n22242, n22243, n22256, 
        n21062, n21064, n22247, n22258, n684_adj_2461, n700_adj_2462, 
        n669_adj_2463, n21566, n21568, n189_adj_2464, n22248, n22249, 
        n22259, n22250, n22251, n22260, n22261, n25633, n22685, 
        n23123, n23124, n23131, n23125, n23126, n23132, n508, 
        n23127, n23128, n23133, n254_adj_2465, n511_adj_2466, n349_adj_2467, 
        n270_adj_2468, n15_adj_2469, n286_adj_2470, n61, n94, n26451, 
        n444_adj_2471, n21571, n573_adj_2472, n22686, n700_adj_2473, 
        n22279, n763_adj_2474, n22280, n860_adj_2475, n620_adj_2476, 
        n924_adj_2477, n21094, n29205, n21097, n1018, n173_adj_2478, 
        n22813, n22814, n21021, n508_adj_2479, n22688, n22689, n22692, 
        n26817, n26818, n26819, n20003, n24537, n24538, n125_adj_2480, 
        n28120, n22690, n22691, n22693, n21575, n21576, n21577, 
        n94_adj_2481, n125_adj_2482, n17585, n14366, n21782, n26567, 
        n21583, n21586, n252_adj_2483, n28118, n21581, n21582, n21589, 
        n21592, n15038, n28121, n21584, n21585, n796_adj_2484, n21068, 
        n413_adj_2485, n444_adj_2486, n476_adj_2487, n507_adj_2488, 
        n24539, n24542, n28177, n28179, n17575, n573_adj_2489, n28180, 
        n875_adj_2490, n891_adj_2491, n15_adj_2492, n859_adj_2493, n860_adj_2494, 
        n605, n636_adj_2495, n62_adj_2496, n21595, n700_adj_2497, 
        n22347, n26513, n31, n29207, n21034, n21598, n22348, n797_adj_2498, 
        n26426, n636_adj_2499, n17543, n17545, n12030, n21733, n124_adj_2500, 
        n507_adj_2501, n860_adj_2502, n891_adj_2503, n476_adj_2504, 
        n22042, n397_adj_2505, n413_adj_2506, n17577, n17578, n17579, 
        n475_adj_2507, n28280, n21730, n173_adj_2508, n30_adj_2509, 
        n31_adj_2510, n109_adj_2511, n124_adj_2512, n125_adj_2513, n653_adj_2514, 
        n635_adj_2515, n94_adj_2516, n30_adj_2517, n31_adj_2518, n28281, 
        n26419, n22978, n15_adj_2519, n30_adj_2520, n31_adj_2521, 
        n26435, n61_adj_2522, n62_adj_2523, n15_adj_2524, n26433, 
        n31_adj_2525, n22760, n781_adj_2526, n30_adj_2527, n31_adj_2528, 
        n12003, n26686, n12004, n21587, n21588, n94_adj_2529, n21601, 
        n14783, n21590, n21591, n221_adj_2530, n252_adj_2531, n28443, 
        n286_adj_2532, n21604, n26688, n21720, n25215, n26703, n24594, 
        n308, n21657, n349_adj_2533, n21607, n635_adj_2534, n636_adj_2535, 
        n26602, n24595, n189_adj_2536, n890_adj_2537, n21596, n26634, 
        n19979, n24597, n731_adj_2538, n796_adj_2539, n22061, n26707, 
        n124_adj_2540, n17346, n24245, n348_adj_2541, n892_adj_2542, 
        n700_adj_2543, n29206, n29208, n19590, n923_adj_2544, n924_adj_2545, 
        n892_adj_2546, n93_adj_2547, n22832, n25806, n24637, n26694, 
        n251_adj_2548, n26635, n669_adj_2549, n700_adj_2550, n24636, 
        n28701, n46_adj_2551, n22831, n21619, n221_adj_2552, n21818, 
        n21820, n28702, n28703, n28700, n21622, n828_adj_2553, n29177, 
        n24640, n860_adj_2554, n21625, n28704, n28705, n28706, n28707, 
        n348_adj_2555, n349_adj_2556, n732_adj_2557, n22040, n21783, 
        n21784, n892_adj_2558, n28762, n28761, n28763, n28764, n28765, 
        n94_adj_2559, n125_adj_2560, n28766, n94_adj_2561, n14450, 
        n21381, n25807, n25812, n28767, n28768, n158_adj_2562, n11915, 
        n11916, n908_adj_2563, n21558, n14848, n21557, n286_adj_2564, 
        n21634, n25822, n349_adj_2565, n21637, n21611, n413_adj_2566, 
        n444_adj_2567, n700_adj_2568, n701_adj_2569, n476_adj_2570, 
        n875_adj_2571, n891_adj_2572, n25823, n25828, n19612, n1018_adj_2573, 
        n22830, n812_adj_2574, n13827, n828_adj_2575, n21640, n26356, 
        n797_adj_2576, n11991, n21643, n669_adj_2577, n700_adj_2578, 
        n22409, n668_adj_2579, n669_adj_2580, n21646, n22410, n22834, 
        n22835, n860_adj_2581, n891_adj_2582, n812_adj_2583, n542_adj_2584, 
        n26352, n25853, n26800, n11010, n252_adj_2585, n25554, n22112, 
        n12017, n28182, n25857, n26183, n26180, n26799, n21543, 
        n21542, n26182, n26181, n17344, n924_adj_2586, n21649, n21390, 
        n21652, n93_adj_2587, n22840, n22841, n22842, n22843, n17343, 
        n22844, n22845, n475_adj_2588, n1002_adj_2589, n26353, n25863, 
        n890_adj_2590, n732_adj_2591, n17342, n158_adj_2592, n28123, 
        n25867, n21629, n21631, n26811, n26812, n26813, n26179, 
        n22265, n221_adj_2593, n21658, n21524, n21525, n21526, n286_adj_2594, 
        n317_adj_2595, n349_adj_2596, n21661, n26410, n22825, n875_adj_2597, 
        n891_adj_2598, n413_adj_2599, n21664, n26570, n21293, n21294, 
        n15074, n26340, n26594, n26802, n286_adj_2600, n21296, n460_adj_2601, 
        n859_adj_2602, n860_adj_2603, n731_adj_2604, n732_adj_2605, 
        n653_adj_2606, n669_adj_2607, n605_adj_2608, n26407, n26394, 
        n26774, n21115, n26408, n26386, n21667, n507_adj_2609, n21111, 
        n21112, n26166, n413_adj_2610, n21678, n24495, n25914, n24760, 
        n26803, n21670, n317_adj_2611, n286_adj_2612, n22805, n22804, 
        n22803, n605_adj_2613, n21673, n22802, n21018, n13863, n158_adj_2614, 
        n21017, n21019, n22798, n22797, n25912, n669_adj_2615, n22795, 
        n732_adj_2616, n763_adj_2617, n25915, n94_adj_2618, n476_adj_2619, 
        n24764, n22443, n21732, n24599, n22928, n25930, n25932, 
        n21731, n26804, n21644, n21645, n21729, n24165, n20372, 
        n21728, n22924, n25933, n285_adj_2620, n26744, n924_adj_2621, 
        n956_adj_2622, n26743, n24766, n24767, n142_adj_2623, n158_adj_2624, 
        n26592, n26708, n21725, n21726, n21727, n21722, n21723, 
        n21724, n21305, n21306, n747_adj_2625, n762_adj_2626, n21308, 
        n21309, n94_adj_2627, n21679, n13839, n26544, n21682, n21685, 
        n22463, n985_adj_2628, n986_adj_2629, n971_adj_2630, n26375, 
        n21359, n24458, n21377, n21688, n317_adj_2631, n939_adj_2632, 
        n22110, n25981, n349_adj_2633, n21691, n24166, n22558, n12018, 
        n923_adj_2634, n26401, n24162, n26346, n21311, n397_adj_2635, 
        n21374, n348_adj_2636, n443_adj_2637, n21369, n21368, n348_adj_2638, 
        n21694, n21697, n21317, n21318, n21319, n21366, n333, 
        n21365, n21700, n21703, n21320, n21321, n557_adj_2639, n572_adj_2640, 
        n23108, n21714, n21706, n573_adj_2641, n22469, n93_adj_2642, 
        n22894, n908_adj_2643, n22114, n25979, n24127, n26347, n26397, 
        n21709, n22470, n22115, n25978, n21712, n26689, n653_adj_2644, 
        n26591, n21699, n21715, n21718, n924_adj_2645, n221_adj_2646, 
        n17341, n397_adj_2647, n27929, n987, n26705, n26588, n716_adj_2648, 
        n891_adj_2649, n812_adj_2650, n14092, n828_adj_2651, n26358, 
        n797_adj_2652, n506_adj_2653, n21323, n26608, n21692, n668_adj_2654, 
        n669_adj_2655, n26808, n26809, n26810, n21689, n301_adj_2656, 
        n908_adj_2657, n22892, n22893, n541_adj_2658, n542_adj_2659, 
        n21357, n557_adj_2660, n21356, n859_adj_2661, n875_adj_2662, 
        n22896, n22897, n589_adj_2663, n23109, n828_adj_2664, n26806, 
        n21354, n653_adj_2665, n21353, n22902, n22903, n723, n21680, 
        n26805, n22904, n22905, n29204, n26807, n22906, n22907, 
        n21344, n21326, n21341, n620_adj_2666, n635_adj_2667, n23110, 
        n762_adj_2668, n21336, n716_adj_2669, n14770, n21335, n17340, 
        n270_adj_2670, n93_adj_2671, n21333, n731_adj_2672, n21332, 
        n732_adj_2673, n17339, n348_adj_2674, n541_adj_2675, n21362, 
        n684_adj_2676, n21671, n21681, n21672, n397_adj_2677, n21342, 
        n21666, n17338, n955_adj_2678, n21705, n348_adj_2679, n443_adj_2680, 
        n11955, n22929, n668_adj_2681, n23111, n333_adj_2682, n21660, 
        n21683, n21684, n21659, n14791, n21656, n506_adj_2683, n348_adj_2684, 
        n22318, n22320, n21686, n573_adj_2685, n93_adj_2686, n491_adj_2687, 
        n605_adj_2688, n636_adj_2689, n30_adj_2690, n26636, n700_adj_2691, 
        n21648, n173_adj_2692, n21647, n21693, n26692, n21641, n732_adj_2693, 
        n908_adj_2694, n21014, n21016, n716_adj_2695, n653_adj_2696, 
        n475_adj_2697, n142_adj_2698, n604_adj_2699, n25982, n25980, 
        n684_adj_2700, n699_adj_2701, n23112, n860_adj_2702, n21669, 
        n23113, n20376, n11946, n24130, n26376, n270_adj_2703, n762_adj_2704, 
        n23114, n22126, n24443, n22537, n316_adj_2705, n397_adj_2706, 
        n21636, n21635, n30_adj_2707, n24131, n653_adj_2708, n21698, 
        n11947, n21633, n21632, n21701, n21702, n797_adj_2709, n21070, 
        n142_adj_2710, n14127, n21707, n21708, n22543, n21624, n22545, 
        n21623, n21650, n21713, n860_adj_2711, n22757, n22761, n22762, 
        n766, n21177, n21620, n21638, n21639, n21618, n796_adj_2712, 
        n23115, n397_adj_2713, n26590, n986_adj_2714, n21716, n22556, 
        n22557, n46_adj_2715, n812_adj_2716, n23116, n190_adj_2717, 
        n25487, n21375, n491_adj_2718, n875_adj_2719, n23118, n22694, 
        n22324, n1002_adj_2720, n23119, n22563, n22564, n22565, 
        n23120, n21606, n21605, n21603, n21617, n21602, n859_adj_2721, 
        n21599, n23121, n542_adj_2722, n26795, n26460, n23122, n892_adj_2723, 
        n684_adj_2724, n890_adj_2725, n26562, n460_adj_2726, n26412, 
        n638, n25934, n25931, n189_adj_2727, n1021, n24765, n21593, 
        n21594, n19899, n26436, n17574, n26476, n1021_adj_2728, 
        n22942, n25916, n25913, n22799, n21579, n316_adj_2729, n17583, 
        n17584, n21578, n21580, n109_adj_2730, n635_adj_2731, n204_adj_2732, 
        n22800, n317_adj_2733, n221_adj_2734, n21103, n22806, n286_adj_2735, 
        n22807, n21095, n26768, n349_adj_2736, n21106, n844_adj_2737, 
        n23055, n25232, n21109, n22013, n507_adj_2738, n573_adj_2739, 
        n21118, n844_adj_2740, n23117, n763_adj_2741, n924_adj_2742, 
        n11995, n22618, n21023, n24455, n22619, n25469, n25630, 
        n26801, n62_adj_2743, n21528, n173_adj_2744, n25865, n491_adj_2745, 
        n22047, n986_adj_2746, n25263, n25260, n716_adj_2747, n24249, 
        n25864, n22290, n25855, n22420, n22478, n25276, n17542, 
        n11827, n924_adj_2748, n573_adj_2749, n22481, n25854, n605_adj_2750, 
        n636_adj_2751, n22712, n22697, n25596, n22715, n25635, n22704, 
        n22054, n24445, n24543, n24460, n684_adj_2752, n21775, n21781, 
        n22202, n22203, n890_adj_2753, n26565, n157_adj_2754, n25357, 
        n22763, n557_adj_2755, n24641, n24638, n24642, n21793, n21799, 
        n21802, n21808, n11225, n21817, n21339, n21391, n987_adj_2756, 
        n21394, n11948, n26415, n638_adj_2757, n859_adj_2758, n24598, 
        n24596, n21816, n22444, n684_adj_2759, n25585, n21561, n11249, 
        n12019, n142_adj_2760, n25449, n491_adj_2761, n26385, n25355, 
        n19975, n62_adj_2762, n25081, n19624, n62_adj_2763, n21102, 
        n21806, n20065, n14756, n25237, n62_adj_2764, n14391, n21022, 
        n21025, n21028, n21031, n491_adj_2765, n25327, n25352, n573_adj_2766, 
        n605_adj_2767, n25217, n21037, n333_adj_2768, n28181, n28178, 
        n21101, n26370, n21116, n21779, n21117, n21780, n28122, 
        n28119, n21792, n506_adj_2769, n21774, n221_adj_2770, n252_adj_2771, 
        n25634, n25631, n27994, n21105, n14395, n21393, n94_adj_2772, 
        n924_adj_2773, n21815, n27930, n27927, n29203, n25595, n25593, 
        n25464, n25329, n19605, n205, n333_adj_2774, n26367, n25226, 
        n12046, n12064, n12059, n21800, n491_adj_2775, n25307, n348_adj_2776, 
        n25262, n572_adj_2777, n189_adj_2778, n22967, n11877, n21092, 
        n21093, n21392, n766_adj_2779, n21171, n364_adj_2780, n25452, 
        n25486, n25484, n26717, n491_adj_2781, n25485, n24459, n24457, 
        n25468, n25466, n24444, n24442, n25231, n25451, n25448, 
        n205_adj_2782, n21389, n14367, n348_adj_2783, n572_adj_2784, 
        n157_adj_2785, n26684, n572_adj_2786, n25337, n25356, n25353, 
        n24361, n24359, n25311, n25308, n24167, n25275, n25273, 
        n25264, n25261, n25236, n25234, n24132, n25230, n25228, 
        n25208, n25205, n25204;
    
    LUT4 i12204_3_lut_3_lut_rep_801 (.A(index_i[2]), .B(index_i[0]), .C(index_i[1]), 
         .Z(n29180)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i12204_3_lut_3_lut_rep_801.init = 16'hd0d0;
    L6MUX21 i22735 (.D0(n24310), .D1(n24308), .SD(index_i[6]), .Z(n24311));
    PFUMX i19995 (.BLUT(n22330), .ALUT(n22331), .C0(index_i[8]), .Z(n22334));
    LUT4 mux_192_Mux_3_i891_3_lut (.A(n541), .B(n890), .C(index_q[4]), 
         .Z(n891)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_3_i891_3_lut.init = 16'hcaca;
    L6MUX21 i19996 (.D0(n22332), .D1(n22333), .SD(index_i[8]), .Z(n22335));
    LUT4 mux_192_Mux_10_i62_3_lut_3_lut_4_lut (.A(n26496), .B(index_q[3]), 
         .C(n26482), .D(index_q[4]), .Z(n62)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_10_i62_3_lut_3_lut_4_lut.init = 16'hf077;
    L6MUX21 i20087 (.D0(n22421), .D1(n22422), .SD(index_i[7]), .Z(n22426));
    PFUMX i20521 (.BLUT(n22858), .ALUT(n22859), .C0(index_i[8]), .Z(n22860));
    LUT4 mux_192_Mux_4_i900_3_lut_4_lut_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n900)) /* synthesis lut_function=(A ((C)+!B)+!A !(B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_4_i900_3_lut_4_lut_3_lut.init = 16'hb2b2;
    L6MUX21 i20149 (.D0(n22483), .D1(n22484), .SD(index_i[7]), .Z(n22488));
    LUT4 i11497_3_lut_4_lut (.A(n26430), .B(index_q[3]), .C(n9970), .D(index_q[6]), 
         .Z(n765)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11497_3_lut_4_lut.init = 16'hffe0;
    LUT4 n124_bdd_3_lut_24220_4_lut (.A(n26430), .B(index_q[3]), .C(index_q[4]), 
         .D(n93), .Z(n24456)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n124_bdd_3_lut_24220_4_lut.init = 16'hfe0e;
    PFUMX i22733 (.BLUT(n924), .ALUT(n24309), .C0(index_i[5]), .Z(n24310));
    PFUMX i20583 (.BLUT(n22920), .ALUT(n22921), .C0(index_q[8]), .Z(n22922));
    PFUMX i23396 (.BLUT(n25085), .ALUT(n25082), .C0(index_q[6]), .Z(n25086));
    PFUMX i20172 (.BLUT(n22507), .ALUT(n22508), .C0(index_q[8]), .Z(n22511));
    LUT4 mux_192_Mux_3_i252_3_lut_4_lut (.A(n26496), .B(index_q[3]), .C(index_q[4]), 
         .D(n14728), .Z(n252)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_3_i252_3_lut_4_lut.init = 16'h08f8;
    LUT4 n624_bdd_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n25553)) /* synthesis lut_function=(!(A (D)+!A !(B (D)+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n624_bdd_4_lut_4_lut_4_lut.init = 16'h54bb;
    LUT4 i12225_2_lut (.A(index_i[1]), .B(index_i[3]), .Z(n541_adj_2251)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i12225_2_lut.init = 16'h1111;
    LUT4 mux_191_Mux_0_i526_3_lut (.A(n26697), .B(n26709), .C(index_i[3]), 
         .Z(n526)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_0_i526_3_lut.init = 16'hcaca;
    LUT4 i20345_3_lut (.A(n26607), .B(n29194), .C(index_i[3]), .Z(n22684)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20345_3_lut.init = 16'hcaca;
    LUT4 i20344_3_lut (.A(n26604), .B(n108), .C(index_i[3]), .Z(n22683)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20344_3_lut.init = 16'hcaca;
    L6MUX21 i20173 (.D0(n22509), .D1(n22510), .SD(index_q[8]), .Z(n22512));
    LUT4 mux_192_Mux_3_i669_3_lut (.A(n653), .B(n668), .C(index_q[4]), 
         .Z(n669)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_3_i669_3_lut.init = 16'hcaca;
    LUT4 mux_191_Mux_7_i156_3_lut_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n70)) /* synthesis lut_function=(!(A (B)+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_7_i156_3_lut_3_lut_3_lut.init = 16'h6363;
    LUT4 i3502_2_lut_rep_581 (.A(index_q[0]), .B(index_q[1]), .Z(n26541)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i3502_2_lut_rep_581.init = 16'h6666;
    PFUMX i20768 (.BLUT(n526), .ALUT(n541_adj_2251), .C0(index_i[4]), 
          .Z(n23107));
    LUT4 i9427_4_lut (.A(n26538), .B(n29190), .C(index_q[3]), .D(index_q[4]), 
         .Z(n11873)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B ((D)+!C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9427_4_lut.init = 16'h3afa;
    FD1S3BX quarter_wave_sample_register_i_i14 (.D(quarter_wave_sample_register_i_15__N_2127[14]), 
            .CK(dac_clk_p_c), .PD(n26683), .Q(quarter_wave_sample_register_i[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i14.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i13 (.D(quarter_wave_sample_register_i_15__N_2127[13]), 
            .CK(dac_clk_p_c), .PD(n26683), .Q(quarter_wave_sample_register_i[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i13.GSR = "DISABLED";
    PFUMX i19053 (.BLUT(n21371), .ALUT(n21372), .C0(index_q[4]), .Z(n21373));
    LUT4 mux_192_Mux_0_i396_3_lut_4_lut_3_lut_rep_774 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n26734)) /* synthesis lut_function=(A ((C)+!B)+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_0_i396_3_lut_4_lut_3_lut_rep_774.init = 16'hb6b6;
    PFUMX i24484 (.BLUT(n26770), .ALUT(n26771), .C0(index_q[1]), .Z(n26772));
    LUT4 i18994_3_lut_4_lut_4_lut (.A(n26438), .B(index_i[4]), .C(index_i[3]), 
         .D(n26519), .Z(n21314)) /* synthesis lut_function=(A (B (C)+!B !(C+!(D)))+!A (B (C)+!B (C+(D)))) */ ;
    defparam i18994_3_lut_4_lut_4_lut.init = 16'hd3d0;
    FD1S3BX quarter_wave_sample_register_i_i12 (.D(quarter_wave_sample_register_i_15__N_2127[12]), 
            .CK(dac_clk_p_c), .PD(n26683), .Q(quarter_wave_sample_register_i[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i12.GSR = "DISABLED";
    LUT4 i21817_3_lut (.A(n21083), .B(n21084), .C(index_q[4]), .Z(n21085)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21817_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_1_i301_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n301)) /* synthesis lut_function=(A (B (C+(D))+!B !(D))+!A !(B (C+(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_1_i301_3_lut_4_lut_4_lut.init = 16'h99b6;
    LUT4 i18727_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21047)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A !(B (C+!(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18727_3_lut_4_lut_4_lut.init = 16'ha52b;
    LUT4 mux_192_Mux_6_i660_3_lut_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n660)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_6_i660_3_lut_3_lut.init = 16'hc6c6;
    LUT4 i11069_2_lut_rep_775 (.A(index_q[0]), .B(index_q[1]), .Z(n26735)) /* synthesis lut_function=((B)+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11069_2_lut_rep_775.init = 16'hdddd;
    LUT4 mux_192_Mux_3_i476_3_lut (.A(n460), .B(n285), .C(index_q[4]), 
         .Z(n476)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_3_i476_3_lut.init = 16'hcaca;
    L6MUX21 i23383 (.D0(n25072), .D1(n25069), .SD(index_q[5]), .Z(n25073));
    PFUMX i23381 (.BLUT(n25071), .ALUT(n25070), .C0(index_q[4]), .Z(n25072));
    LUT4 i9525_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(n26547), .D(index_i[4]), .Z(n221)) /* synthesis lut_function=(!(A (B)+!A (B (C+(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9525_3_lut_4_lut_4_lut_4_lut.init = 16'h3336;
    FD1S3BX quarter_wave_sample_register_i_i11 (.D(quarter_wave_sample_register_i_15__N_2127[11]), 
            .CK(dac_clk_p_c), .PD(n26683), .Q(quarter_wave_sample_register_i[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i11.GSR = "DISABLED";
    PFUMX i20706 (.BLUT(n526_adj_2252), .ALUT(n541_adj_2253), .C0(index_q[4]), 
          .Z(n23045));
    LUT4 i19249_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n21569)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (D))+!A !(D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19249_3_lut_4_lut_4_lut_4_lut.init = 16'ha25d;
    LUT4 mux_192_Mux_3_i413_3_lut (.A(n397), .B(n26582), .C(index_q[4]), 
         .Z(n413)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_3_i413_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_3_i619_3_lut_rep_561_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n26521)) /* synthesis lut_function=(!(A (B)+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_3_i619_3_lut_rep_561_3_lut.init = 16'h6363;
    FD1S3BX quarter_wave_sample_register_i_i10 (.D(quarter_wave_sample_register_i_15__N_2127[10]), 
            .CK(dac_clk_p_c), .PD(n26683), .Q(quarter_wave_sample_register_i[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i10.GSR = "DISABLED";
    LUT4 mux_192_Mux_0_i316_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n316)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+(D)))+!A (B (C+(D))+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_0_i316_3_lut_4_lut_4_lut_4_lut.init = 16'h332d;
    LUT4 mux_192_Mux_5_i356_3_lut_4_lut_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n325)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_5_i356_3_lut_4_lut_3_lut.init = 16'h6d6d;
    FD1S3BX quarter_wave_sample_register_i_i9 (.D(quarter_wave_sample_register_i_15__N_2127[9]), 
            .CK(dac_clk_p_c), .PD(n26683), .Q(quarter_wave_sample_register_i[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i9.GSR = "DISABLED";
    FD1P3AX phase_q__i1 (.D(o_phase[0]), .SP(o_dac_cw_b_c_c), .CK(dac_clk_p_c), 
            .Q(phase_q[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_q__i1.GSR = "DISABLED";
    PFUMX i20798 (.BLUT(n23135), .ALUT(n23136), .C0(index_i[8]), .Z(n23137));
    LUT4 i20343_3_lut (.A(n619), .B(n26650), .C(index_i[3]), .Z(n22682)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20343_3_lut.init = 16'hcaca;
    FD1S3BX quarter_wave_sample_register_i_i8 (.D(quarter_wave_sample_register_i_15__N_2127[8]), 
            .CK(dac_clk_p_c), .PD(n26683), .Q(quarter_wave_sample_register_i[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i8.GSR = "DISABLED";
    LUT4 mux_191_Mux_1_i882_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n882)) /* synthesis lut_function=(A ((C)+!B)+!A !((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_1_i882_3_lut_3_lut.init = 16'ha6a6;
    LUT4 mux_192_Mux_8_i860_3_lut_4_lut (.A(n26496), .B(index_q[3]), .C(index_q[4]), 
         .D(n26482), .Z(n860)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_8_i860_3_lut_4_lut.init = 16'h08f8;
    FD1S3DX o_val_pipeline_q_1__i1 (.D(\o_val_pipeline_q[0] [7]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(o_dac_b_c_7)) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_q_1__i1.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i7 (.D(quarter_wave_sample_register_i_15__N_2127[7]), 
            .CK(dac_clk_p_c), .PD(n26683), .Q(quarter_wave_sample_register_i[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i7.GSR = "DISABLED";
    FD1S3DX phase_negation_i_i0 (.D(phase_i[11]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(phase_negation_i[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_negation_i_i0.GSR = "DISABLED";
    FD1S3DX phase_negation_q_i0 (.D(phase_q[11]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(phase_negation_q[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_negation_q_i0.GSR = "DISABLED";
    FD1S3DX index_i_i0 (.D(index_i_9__N_2107[0]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(index_i[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_i_i0.GSR = "DISABLED";
    FD1S3DX index_q_i0 (.D(index_q_9__N_2117[0]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(index_q[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_q_i0.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i0 (.D(quarter_wave_sample_register_q_15__N_2142[0]), 
            .CK(dac_clk_p_c), .PD(n26683), .Q(quarter_wave_sample_register_q[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_q_i0.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i1 (.D(\o_val_pipeline_i[0] [7]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(\o_sample_i[7] )) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i1.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i0 (.D(quarter_wave_sample_register_i_15__N_2127[0]), 
            .CK(dac_clk_p_c), .PD(n26683), .Q(quarter_wave_sample_register_i[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i0.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i6 (.D(quarter_wave_sample_register_i_15__N_2127[6]), 
            .CK(dac_clk_p_c), .PD(n26683), .Q(quarter_wave_sample_register_i[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i6.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i5 (.D(quarter_wave_sample_register_i_15__N_2127[5]), 
            .CK(dac_clk_p_c), .PD(n26683), .Q(quarter_wave_sample_register_i[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i5.GSR = "DISABLED";
    LUT4 mux_192_Mux_3_i286_4_lut (.A(n93_adj_2254), .B(index_q[2]), .C(index_q[4]), 
         .D(n13857), .Z(n286)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_3_i286_4_lut.init = 16'h3aca;
    FD1S3BX quarter_wave_sample_register_i_i4 (.D(quarter_wave_sample_register_i_15__N_2127[4]), 
            .CK(dac_clk_p_c), .PD(n26683), .Q(quarter_wave_sample_register_i[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i4.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i3 (.D(quarter_wave_sample_register_i_15__N_2127[3]), 
            .CK(dac_clk_p_c), .PD(n26683), .Q(quarter_wave_sample_register_i[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i3.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i2 (.D(quarter_wave_sample_register_i_15__N_2127[2]), 
            .CK(dac_clk_p_c), .PD(n26683), .Q(quarter_wave_sample_register_i[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i2.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i1 (.D(quarter_wave_sample_register_i_15__N_2127[1]), 
            .CK(dac_clk_p_c), .PD(n26683), .Q(quarter_wave_sample_register_i[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i1.GSR = "DISABLED";
    PFUMX i19065 (.BLUT(n21383), .ALUT(n21384), .C0(index_q[4]), .Z(n21385));
    LUT4 i20342_3_lut (.A(n70), .B(n26691), .C(index_i[3]), .Z(n22681)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20342_3_lut.init = 16'hcaca;
    LUT4 i21815_3_lut (.A(n21086), .B(n21087), .C(index_q[4]), .Z(n21088)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21815_3_lut.init = 16'hcaca;
    LUT4 i21828_3_lut (.A(n28444), .B(n26851), .C(index_q[5]), .Z(n22252)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21828_3_lut.init = 16'hcaca;
    FD1S3DX o_val_pipeline_i_1__i18 (.D(o_val_pipeline_i_0__15__N_2157), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(\o_val_pipeline_i[0] [15])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i18.GSR = "DISABLED";
    LUT4 n28_bdd_3_lut_23761_4_lut_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .Z(n24920)) /* synthesis lut_function=(A (B)+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n28_bdd_3_lut_23761_4_lut_3_lut.init = 16'hd9d9;
    FD1S3DX o_val_pipeline_i_1__i17 (.D(o_val_pipeline_i_0__15__N_2159), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(\o_val_pipeline_i[0] [14])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i17.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i16 (.D(o_val_pipeline_i_0__15__N_2161), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(\o_val_pipeline_i[0] [13])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i16.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i15 (.D(o_val_pipeline_i_0__15__N_2163), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(\o_val_pipeline_i[0] [12])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i15.GSR = "DISABLED";
    LUT4 mux_192_Mux_0_i635_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n635)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_0_i635_3_lut_4_lut_4_lut.init = 16'hfd0a;
    LUT4 i19043_3_lut_3_lut_4_lut (.A(n26430), .B(index_q[3]), .C(n93), 
         .D(index_q[4]), .Z(n21363)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19043_3_lut_3_lut_4_lut.init = 16'h11f0;
    PFUMX i22731 (.BLUT(n24307), .ALUT(n26478), .C0(index_i[5]), .Z(n24308));
    LUT4 mux_191_Mux_6_i660_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n108)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_6_i660_3_lut_3_lut.init = 16'hc6c6;
    FD1S3DX o_val_pipeline_i_1__i14 (.D(o_val_pipeline_i_0__15__N_2165), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(\o_val_pipeline_i[0] [11])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i14.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i13 (.D(o_val_pipeline_i_0__15__N_2167), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(\o_val_pipeline_i[0] [10])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i13.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i12 (.D(o_val_pipeline_i_0__15__N_2169), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(\o_val_pipeline_i[0] [9])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i12.GSR = "DISABLED";
    LUT4 n173_bdd_4_lut (.A(n173), .B(n70_adj_2255), .C(index_i[4]), .D(index_i[3]), 
         .Z(n24309)) /* synthesis lut_function=(A (B+(C+!(D)))+!A !((C+!(D))+!B)) */ ;
    defparam n173_bdd_4_lut.init = 16'hacaa;
    PFUMX i19068 (.BLUT(n21386), .ALUT(n21387), .C0(index_q[4]), .Z(n21388));
    LUT4 mux_192_Mux_6_i564_3_lut_4_lut_3_lut_rep_776 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n26736)) /* synthesis lut_function=(A (B)+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_6_i564_3_lut_4_lut_3_lut_rep_776.init = 16'hd9d9;
    LUT4 mux_192_Mux_3_i507_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[4]), .D(n491), .Z(n507)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_3_i507_3_lut_4_lut.init = 16'h6f60;
    FD1S3DX o_val_pipeline_i_1__i11 (.D(o_val_pipeline_i_0__15__N_2171), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(\o_val_pipeline_i[0] [8])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i11.GSR = "DISABLED";
    LUT4 i21832_3_lut (.A(n542), .B(n573), .C(index_q[5]), .Z(n22246)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21832_3_lut.init = 16'hcaca;
    LUT4 mux_191_Mux_8_i301_3_lut_4_lut (.A(n26647), .B(index_i[2]), .C(index_i[3]), 
         .D(n70_adj_2255), .Z(n301_adj_2256)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_8_i301_3_lut_4_lut.init = 16'h8f80;
    FD1S3DX o_val_pipeline_i_1__i10 (.D(o_val_pipeline_i_0__15__N_2173), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(\o_val_pipeline_i[0] [7])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i10.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i9 (.D(\o_val_pipeline_i[0] [15]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(\o_sample_i[15] )) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i9.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i8 (.D(\o_val_pipeline_i[0] [14]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(\o_sample_i[14] )) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i8.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i7 (.D(\o_val_pipeline_i[0] [13]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(\o_sample_i[13] )) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i7.GSR = "DISABLED";
    LUT4 mux_192_Mux_2_i270_3_lut (.A(n26719), .B(n26728), .C(index_q[3]), 
         .Z(n270)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_2_i270_3_lut.init = 16'hcaca;
    PFUMX i20736 (.BLUT(n23073), .ALUT(n23074), .C0(index_q[8]), .Z(n23075));
    LUT4 mux_191_Mux_0_i747_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n747)) /* synthesis lut_function=(!(A (B+!(C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_0_i747_3_lut_4_lut_4_lut_4_lut.init = 16'h6556;
    FD1S3DX o_val_pipeline_i_1__i6 (.D(\o_val_pipeline_i[0] [12]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(\o_sample_i[12] )) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i6.GSR = "DISABLED";
    LUT4 mux_192_Mux_7_i891_3_lut_4_lut_4_lut (.A(n29190), .B(index_q[3]), 
         .C(n26430), .D(index_q[4]), .Z(n891_adj_2257)) /* synthesis lut_function=(A (B (C+!(D))+!B !((D)+!C))+!A (B (C+!(D))+!B (C+(D)))) */ ;
    defparam mux_192_Mux_7_i891_3_lut_4_lut_4_lut.init = 16'hd1fc;
    L6MUX21 i20383 (.D0(n22717), .D1(n22718), .SD(index_q[7]), .Z(n22722));
    LUT4 i9608_3_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[4]), 
         .Z(n12058)) /* synthesis lut_function=(!(A (B)+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9608_3_lut_4_lut_3_lut.init = 16'h6262;
    FD1S3DX o_val_pipeline_i_1__i5 (.D(\o_val_pipeline_i[0] [11]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(\o_sample_i[11] )) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i5.GSR = "DISABLED";
    LUT4 mux_192_Mux_0_i363_3_lut_4_lut_3_lut_rep_777 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n26737)) /* synthesis lut_function=(A (B+!(C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_0_i363_3_lut_4_lut_3_lut_rep_777.init = 16'hdbdb;
    LUT4 mux_192_Mux_6_i459_rep_780 (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .Z(n26740)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_6_i459_rep_780.init = 16'h4d4d;
    LUT4 mux_192_Mux_2_i316_3_lut (.A(n26720), .B(n29197), .C(index_q[3]), 
         .Z(n316_adj_2258)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_2_i316_3_lut.init = 16'hcaca;
    LUT4 index_i_8__bdd_3_lut_24177_else_4_lut (.A(n26485), .B(index_i[4]), 
         .C(index_i[6]), .D(index_i[5]), .Z(n26820)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;
    defparam index_i_8__bdd_3_lut_24177_else_4_lut.init = 16'hf080;
    LUT4 mux_192_Mux_2_i397_3_lut (.A(n29200), .B(n29182), .C(index_q[3]), 
         .Z(n397_adj_2259)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_2_i397_3_lut.init = 16'hcaca;
    LUT4 i20169_3_lut (.A(n22501), .B(n22502), .C(index_q[7]), .Z(n22508)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20169_3_lut.init = 16'hcaca;
    LUT4 mux_191_Mux_6_i844_3_lut_4_lut (.A(n26647), .B(index_i[2]), .C(index_i[3]), 
         .D(n26649), .Z(n844)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_6_i844_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_192_Mux_9_i700_3_lut_4_lut (.A(n26430), .B(index_q[3]), .C(index_q[4]), 
         .D(n26477), .Z(n700)) /* synthesis lut_function=(!(A (C+!(D))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_9_i700_3_lut_4_lut.init = 16'h1f10;
    PFUMX mux_191_Mux_1_i636 (.BLUT(n620), .ALUT(n635_adj_2260), .C0(index_i[4]), 
          .Z(n636)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    FD1S3DX o_val_pipeline_i_1__i4 (.D(\o_val_pipeline_i[0] [10]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(\o_sample_i[10] )) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i4.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i3 (.D(\o_val_pipeline_i[0] [9]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(\o_sample_i[9] )) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i3.GSR = "DISABLED";
    LUT4 mux_192_Mux_3_i653_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n653)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A !(B (D)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_3_i653_3_lut_4_lut_4_lut.init = 16'h4d99;
    FD1S3DX o_val_pipeline_i_1__i2 (.D(\o_val_pipeline_i[0] [8]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(\o_sample_i[8] )) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i2.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i11 (.D(o_phase[11]), .SP(o_dac_cw_b_c_c), .CK(dac_clk_p_c), 
            .Q(phase_i[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i11.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i10 (.D(o_phase[10]), .SP(o_dac_cw_b_c_c), .CK(dac_clk_p_c), 
            .Q(phase_i[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i10.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i9 (.D(o_phase[9]), .SP(o_dac_cw_b_c_c), .CK(dac_clk_p_c), 
            .Q(phase_i[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i9.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i8 (.D(o_phase[8]), .SP(o_dac_cw_b_c_c), .CK(dac_clk_p_c), 
            .Q(phase_i[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i8.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i7 (.D(o_phase[7]), .SP(o_dac_cw_b_c_c), .CK(dac_clk_p_c), 
            .Q(phase_i[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i7.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i6 (.D(o_phase[6]), .SP(o_dac_cw_b_c_c), .CK(dac_clk_p_c), 
            .Q(phase_i[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i6.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i5 (.D(o_phase[5]), .SP(o_dac_cw_b_c_c), .CK(dac_clk_p_c), 
            .Q(phase_i[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i5.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i4 (.D(o_phase[4]), .SP(o_dac_cw_b_c_c), .CK(dac_clk_p_c), 
            .Q(phase_i[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i4.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i3 (.D(o_phase[3]), .SP(o_dac_cw_b_c_c), .CK(dac_clk_p_c), 
            .Q(phase_i[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i3.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i2 (.D(o_phase[2]), .SP(o_dac_cw_b_c_c), .CK(dac_clk_p_c), 
            .Q(phase_i[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i2.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i1 (.D(o_phase[1]), .SP(o_dac_cw_b_c_c), .CK(dac_clk_p_c), 
            .Q(phase_i[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i1.GSR = "DISABLED";
    LUT4 i18713_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21033)) /* synthesis lut_function=(A (B (C)+!B !(C (D)+!C !(D)))+!A (B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18713_3_lut_4_lut_4_lut.init = 16'hd6a5;
    LUT4 mux_192_Mux_9_i62_3_lut_4_lut_then_4_lut (.A(index_q[4]), .B(index_q[2]), 
         .C(index_q[1]), .D(index_q[0]), .Z(n26750)) /* synthesis lut_function=(!(A (B (C+(D)))+!A (B+(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_9_i62_3_lut_4_lut_then_4_lut.init = 16'h222b;
    LUT4 mux_191_Mux_8_i157_3_lut_4_lut (.A(n26647), .B(index_i[2]), .C(index_i[3]), 
         .D(n26605), .Z(n157)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_8_i157_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_192_Mux_0_i412_3_lut_4_lut_4_lut (.A(index_q[2]), .B(index_q[0]), 
         .C(index_q[1]), .D(index_q[3]), .Z(n412)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C (D)))+!A (B (C+!(D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_0_i412_3_lut_4_lut_4_lut.init = 16'hf14c;
    LUT4 i9511_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n526_adj_2261)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+(D)))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9511_3_lut_4_lut_4_lut.init = 16'h666c;
    LUT4 i18761_3_lut (.A(n26737), .B(n29176), .C(index_q[3]), .Z(n21081)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18761_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_0_i796_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n796)) /* synthesis lut_function=(A (B (C+(D))+!B (C (D)))+!A !(B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_0_i796_3_lut_4_lut_4_lut.init = 16'hadc0;
    LUT4 mux_192_Mux_0_i931_3_lut_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n931)) /* synthesis lut_function=(!(A (B+(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_0_i931_3_lut_3_lut.init = 16'h5656;
    LUT4 n53_bdd_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n25068)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n53_bdd_3_lut_4_lut_4_lut.init = 16'ha5ad;
    LUT4 i20338_3_lut (.A(n29194), .B(n26648), .C(index_i[3]), .Z(n22677)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20338_3_lut.init = 16'hcaca;
    FD1S3BX quarter_wave_sample_register_q_i15 (.D(n29209), .CK(dac_clk_p_c), 
            .PD(n26683), .Q(\quarter_wave_sample_register_q[15] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_q_i15.GSR = "DISABLED";
    LUT4 i18794_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21114)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D))+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18794_3_lut_4_lut.init = 16'hccdb;
    LUT4 mux_192_Mux_0_i364_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n364)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A ((C+!(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_0_i364_3_lut_3_lut_4_lut.init = 16'hdb55;
    LUT4 mux_192_Mux_1_i882_3_lut_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n882_adj_2262)) /* synthesis lut_function=(A ((C)+!B)+!A !((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_1_i882_3_lut_3_lut.init = 16'ha6a6;
    LUT4 i20337_3_lut (.A(n38), .B(n26607), .C(index_i[3]), .Z(n22676)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20337_3_lut.init = 16'hcaca;
    LUT4 i9597_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n12047)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A !(B (C+(D))+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9597_3_lut_4_lut_4_lut_4_lut.init = 16'h44db;
    LUT4 mux_192_Mux_5_i475_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n475)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_5_i475_3_lut_4_lut_4_lut.init = 16'hd4a5;
    FD1S3BX quarter_wave_sample_register_q_i14 (.D(quarter_wave_sample_register_q_15__N_2142[14]), 
            .CK(dac_clk_p_c), .PD(n26683), .Q(quarter_wave_sample_register_q[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_q_i14.GSR = "DISABLED";
    LUT4 mux_191_Mux_5_i356_3_lut_4_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n396)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_5_i356_3_lut_4_lut_4_lut_3_lut.init = 16'h6d6d;
    FD1S3BX quarter_wave_sample_register_q_i13 (.D(quarter_wave_sample_register_q_15__N_2142[13]), 
            .CK(dac_clk_p_c), .PD(n26683), .Q(quarter_wave_sample_register_q[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_q_i13.GSR = "DISABLED";
    LUT4 mux_192_Mux_3_i676_3_lut_4_lut_3_lut_rep_760 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n26720)) /* synthesis lut_function=(A (B (C))+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_3_i676_3_lut_4_lut_3_lut_rep_760.init = 16'h9494;
    LUT4 mux_191_Mux_0_i954_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n954)) /* synthesis lut_function=(A (D)+!A !(B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_0_i954_3_lut_4_lut_4_lut.init = 16'haf40;
    FD1S3BX quarter_wave_sample_register_q_i12 (.D(quarter_wave_sample_register_q_15__N_2142[12]), 
            .CK(dac_clk_p_c), .PD(n26683), .Q(quarter_wave_sample_register_q[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_q_i12.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i11 (.D(quarter_wave_sample_register_q_15__N_2142[11]), 
            .CK(dac_clk_p_c), .PD(n26683), .Q(quarter_wave_sample_register_q[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_q_i11.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i10 (.D(quarter_wave_sample_register_q_15__N_2142[10]), 
            .CK(dac_clk_p_c), .PD(n26683), .Q(quarter_wave_sample_register_q[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_q_i10.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i9 (.D(quarter_wave_sample_register_q_15__N_2142[9]), 
            .CK(dac_clk_p_c), .PD(n26683), .Q(quarter_wave_sample_register_q[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_q_i9.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i8 (.D(quarter_wave_sample_register_q_15__N_2142[8]), 
            .CK(dac_clk_p_c), .PD(n26683), .Q(quarter_wave_sample_register_q[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_q_i8.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i7 (.D(quarter_wave_sample_register_q_15__N_2142[7]), 
            .CK(dac_clk_p_c), .PD(n26683), .Q(quarter_wave_sample_register_q[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_q_i7.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i6 (.D(quarter_wave_sample_register_q_15__N_2142[6]), 
            .CK(dac_clk_p_c), .PD(n26683), .Q(quarter_wave_sample_register_q[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_q_i6.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i5 (.D(quarter_wave_sample_register_q_15__N_2142[5]), 
            .CK(dac_clk_p_c), .PD(n26683), .Q(quarter_wave_sample_register_q[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_q_i5.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i4 (.D(quarter_wave_sample_register_q_15__N_2142[4]), 
            .CK(dac_clk_p_c), .PD(n26683), .Q(quarter_wave_sample_register_q[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_q_i4.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i3 (.D(quarter_wave_sample_register_q_15__N_2142[3]), 
            .CK(dac_clk_p_c), .PD(n26683), .Q(quarter_wave_sample_register_q[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_q_i3.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i2 (.D(quarter_wave_sample_register_q_15__N_2142[2]), 
            .CK(dac_clk_p_c), .PD(n26683), .Q(quarter_wave_sample_register_q[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_q_i2.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i1 (.D(quarter_wave_sample_register_q_15__N_2142[1]), 
            .CK(dac_clk_p_c), .PD(n26683), .Q(quarter_wave_sample_register_q[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_q_i1.GSR = "DISABLED";
    LUT4 i20335_3_lut (.A(n26648), .B(n70), .C(index_i[3]), .Z(n22674)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20335_3_lut.init = 16'hcaca;
    FD1S3DX index_q_i9 (.D(index_q_9__N_2117[9]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(index_q[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_q_i9.GSR = "DISABLED";
    FD1S3DX index_q_i8 (.D(index_q_9__N_2117[8]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(index_q[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_q_i8.GSR = "DISABLED";
    FD1S3DX index_q_i7 (.D(index_q_9__N_2117[7]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(index_q[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_q_i7.GSR = "DISABLED";
    FD1S3DX index_q_i6 (.D(index_q_9__N_2117[6]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(index_q[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_q_i6.GSR = "DISABLED";
    FD1S3DX index_q_i5 (.D(index_q_9__N_2117[5]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(index_q[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_q_i5.GSR = "DISABLED";
    FD1S3DX index_q_i4 (.D(index_q_9__N_2117[4]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(index_q[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_q_i4.GSR = "DISABLED";
    FD1S3DX index_q_i3 (.D(index_q_9__N_2117[3]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(index_q[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_q_i3.GSR = "DISABLED";
    FD1S3DX index_q_i2 (.D(index_q_9__N_2117[2]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(index_q[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_q_i2.GSR = "DISABLED";
    FD1S3DX index_q_i1 (.D(index_q_9__N_2117[1]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(index_q[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_q_i1.GSR = "DISABLED";
    FD1S3DX index_i_i9 (.D(index_i_9__N_2107[9]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(index_i[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_i_i9.GSR = "DISABLED";
    FD1S3DX index_i_i8 (.D(index_i_9__N_2107[8]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(index_i[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_i_i8.GSR = "DISABLED";
    LUT4 i19991_3_lut (.A(n22322), .B(n22323), .C(index_i[7]), .Z(n22330)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19991_3_lut.init = 16'hcaca;
    FD1S3DX index_i_i7 (.D(index_i_9__N_2107[7]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(index_i[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_i_i7.GSR = "DISABLED";
    FD1S3DX index_i_i6 (.D(index_i_9__N_2107[6]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(index_i[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_i_i6.GSR = "DISABLED";
    FD1S3DX index_i_i5 (.D(index_i_9__N_2107[5]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(index_i[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_i_i5.GSR = "DISABLED";
    FD1S3DX index_i_i4 (.D(index_i_9__N_2107[4]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(index_i[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_i_i4.GSR = "DISABLED";
    FD1S3DX index_i_i3 (.D(index_i_9__N_2107[3]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(index_i[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_i_i3.GSR = "DISABLED";
    FD1S3DX index_i_i2 (.D(index_i_9__N_2107[2]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(index_i[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_i_i2.GSR = "DISABLED";
    LUT4 mux_192_Mux_0_i157_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n157_adj_2263)) /* synthesis lut_function=(A (B (C+!(D))+!B !(D))+!A (B (D)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_0_i157_3_lut_4_lut.init = 16'hd4aa;
    FD1S3DX index_i_i1 (.D(index_i_9__N_2107[1]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(index_i[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_i_i1.GSR = "DISABLED";
    FD1S3DX phase_negation_q_i1 (.D(phase_negation_q[0]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(phase_negation_q[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_negation_q_i1.GSR = "DISABLED";
    FD1S3DX phase_negation_i_i1 (.D(phase_negation_i[0]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(phase_negation_i[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_negation_i_i1.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i18 (.D(n1703[14]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(\o_val_pipeline_q[0] [15])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_q_1__i18.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i17 (.D(n1703[13]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(\o_val_pipeline_q[0] [14])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_q_1__i17.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i16 (.D(n1703[12]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(\o_val_pipeline_q[0] [13])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_q_1__i16.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i15 (.D(n1703[11]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(\o_val_pipeline_q[0] [12])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_q_1__i15.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i14 (.D(n1703[10]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(\o_val_pipeline_q[0] [11])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_q_1__i14.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i13 (.D(n1703[9]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(\o_val_pipeline_q[0] [10])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_q_1__i13.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i12 (.D(n1703[8]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(\o_val_pipeline_q[0] [9])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_q_1__i12.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i11 (.D(n1703[7]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(\o_val_pipeline_q[0] [8])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_q_1__i11.GSR = "DISABLED";
    LUT4 mux_191_Mux_8_i173_3_lut_3_lut_4_lut (.A(n26647), .B(index_i[2]), 
         .C(n954_adj_2264), .D(index_i[4]), .Z(n173)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_8_i173_3_lut_3_lut_4_lut.init = 16'hf077;
    FD1S3DX o_val_pipeline_q_1__i10 (.D(n1703[6]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(\o_val_pipeline_q[0] [7])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_q_1__i10.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i9 (.D(\o_val_pipeline_q[0] [15]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(o_dac_b_c_15)) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_q_1__i9.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i8 (.D(\o_val_pipeline_q[0] [14]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(o_dac_b_c_14)) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_q_1__i8.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i7 (.D(\o_val_pipeline_q[0] [13]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(o_dac_b_c_13)) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_q_1__i7.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i6 (.D(\o_val_pipeline_q[0] [12]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(o_dac_b_c_12)) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_q_1__i6.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i5 (.D(\o_val_pipeline_q[0] [11]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(o_dac_b_c_11)) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_q_1__i5.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i4 (.D(\o_val_pipeline_q[0] [10]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(o_dac_b_c_10)) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_q_1__i4.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i3 (.D(\o_val_pipeline_q[0] [9]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(n3537)) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_q_1__i3.GSR = "DISABLED";
    LUT4 i9615_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n12065)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B ((D)+!C)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9615_3_lut_4_lut_4_lut.init = 16'h6c3c;
    FD1S3DX o_val_pipeline_q_1__i2 (.D(\o_val_pipeline_q[0] [8]), .CK(dac_clk_p_c), 
            .CD(n26683), .Q(o_dac_b_c_8)) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_q_1__i2.GSR = "DISABLED";
    LUT4 i15418_3_lut (.A(n26695), .B(n26687), .C(index_i[3]), .Z(n17568)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15418_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_6_i572_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n572)) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_6_i572_3_lut_4_lut.init = 16'hccd9;
    LUT4 i15417_3_lut (.A(n26687), .B(n26697), .C(index_i[3]), .Z(n17567)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15417_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_5_i828_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[4]), .D(n26585), .Z(n828)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_5_i828_4_lut_4_lut.init = 16'hc66c;
    L6MUX21 i19952 (.D0(n22281), .D1(n22282), .SD(index_q[6]), .Z(n22291));
    L6MUX21 i19954 (.D0(n22285), .D1(n22286), .SD(index_q[7]), .Z(n22293));
    L6MUX21 i19955 (.D0(n22287), .D1(n22288), .SD(index_q[7]), .Z(n22294));
    PFUMX mux_191_Mux_2_i891 (.BLUT(n875), .ALUT(n890_adj_2265), .C0(index_i[4]), 
          .Z(n891_adj_2266)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    L6MUX21 i19971 (.D0(n22304), .D1(n22305), .SD(index_q[7]), .Z(n22310));
    PFUMX mux_191_Mux_2_i860 (.BLUT(n844_adj_2267), .ALUT(n859), .C0(index_i[4]), 
          .Z(n860_adj_2268)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 i20168_3_lut (.A(n22499), .B(n22500), .C(index_q[7]), .Z(n22507)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20168_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_9_i285_3_lut_4_lut_4_lut (.A(index_q[2]), .B(index_q[0]), 
         .C(index_q[3]), .D(index_q[1]), .Z(n285_adj_2269)) /* synthesis lut_function=(A (C)+!A !(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_9_i285_3_lut_4_lut_4_lut.init = 16'ha0a1;
    LUT4 mux_191_Mux_6_i22_rep_638 (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .Z(n26598)) /* synthesis lut_function=(!(A (C)+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_6_i22_rep_638.init = 16'h4a4a;
    FD1P3AX phase_q__i11 (.D(phase_q_11__N_2233[11]), .SP(o_dac_cw_b_c_c), 
            .CK(dac_clk_p_c), .Q(phase_q[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_q__i11.GSR = "DISABLED";
    PFUMX i23378 (.BLUT(n25068), .ALUT(n25067), .C0(index_q[4]), .Z(n25069));
    LUT4 i18760_3_lut (.A(n29198), .B(n26724), .C(index_q[3]), .Z(n21080)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18760_3_lut.init = 16'hcaca;
    LUT4 i9543_3_lut_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[4]), .D(index_i[3]), .Z(n444)) /* synthesis lut_function=(!(A (B)+!A !(B (C (D))+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9543_3_lut_3_lut_4_lut_4_lut.init = 16'h6333;
    PFUMX i19972 (.BLUT(n22306), .ALUT(n22307), .C0(index_q[7]), .Z(n22311));
    LUT4 i21603_3_lut (.A(n21554), .B(n21555), .C(index_i[4]), .Z(n21556)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21603_3_lut.init = 16'hcaca;
    LUT4 i3591_2_lut_rep_781 (.A(index_q[0]), .B(index_q[2]), .Z(n26741)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i3591_2_lut_rep_781.init = 16'h6666;
    LUT4 mux_192_Mux_6_i732_3_lut_4_lut (.A(n26571), .B(index_q[3]), .C(index_q[4]), 
         .D(n781), .Z(n732)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_6_i732_3_lut_4_lut.init = 16'hf909;
    LUT4 i18745_3_lut (.A(n931), .B(n29197), .C(index_q[3]), .Z(n21065)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18745_3_lut.init = 16'hcaca;
    LUT4 i21821_3_lut (.A(n21080), .B(n21081), .C(index_q[4]), .Z(n21082)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21821_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_6_i700_3_lut_4_lut (.A(n26571), .B(index_q[3]), .C(index_q[4]), 
         .D(n684), .Z(n700_adj_2270)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_6_i700_3_lut_4_lut.init = 16'h9f90;
    LUT4 i19390_3_lut_3_lut_4_lut (.A(n26647), .B(index_i[2]), .C(n38), 
         .D(index_i[3]), .Z(n21710)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19390_3_lut_3_lut_4_lut.init = 16'hf077;
    L6MUX21 i19977 (.D0(n382), .D1(n509), .SD(index_i[7]), .Z(n22316));
    L6MUX21 i18885 (.D0(n21203), .D1(n21204), .SD(index_i[7]), .Z(n21205));
    L6MUX21 i19993 (.D0(n22326), .D1(n22327), .SD(index_i[7]), .Z(n22332));
    LUT4 i18716_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21036)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A (B (C (D)+!C !(D))+!B (D))) */ ;
    defparam i18716_3_lut_4_lut.init = 16'hd926;
    L6MUX21 i19994 (.D0(n22328), .D1(n22329), .SD(index_i[7]), .Z(n22333));
    L6MUX21 i18894 (.D0(n21212), .D1(n21213), .SD(index_q[7]), .Z(n21214));
    PFUMX i24543 (.BLUT(n26861), .ALUT(n26862), .C0(index_i[3]), .Z(n62_adj_2271));
    LUT4 n708_bdd_2_lut_3_lut_3_lut_4_lut (.A(index_q[2]), .B(index_q[0]), 
         .C(index_q[1]), .D(index_q[3]), .Z(n25583)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n708_bdd_2_lut_3_lut_3_lut_4_lut.init = 16'h00fe;
    L6MUX21 i20483 (.D0(n22820), .D1(n22821), .SD(index_q[7]), .Z(n22822));
    L6MUX21 i20022 (.D0(n22353), .D1(n22354), .SD(index_i[7]), .Z(n22361));
    L6MUX21 i20023 (.D0(n22355), .D1(n22356), .SD(index_i[7]), .Z(n22362));
    LUT4 mux_191_Mux_12_i254_4_lut (.A(n26373), .B(n20230), .C(index_i[6]), 
         .D(n26486), .Z(n254)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_12_i254_4_lut.init = 16'hca0a;
    L6MUX21 i20082 (.D0(n22411), .D1(n22412), .SD(index_i[6]), .Z(n22421));
    L6MUX21 i20084 (.D0(n22415), .D1(n22416), .SD(index_i[7]), .Z(n22423));
    L6MUX21 i20085 (.D0(n22417), .D1(n22418), .SD(index_i[7]), .Z(n22424));
    L6MUX21 i20116 (.D0(n22448), .D1(n22449), .SD(index_i[7]), .Z(n22455));
    L6MUX21 i20117 (.D0(n22450), .D1(n22451), .SD(index_i[7]), .Z(n22456));
    PFUMX i20118 (.BLUT(n22452), .ALUT(n22453), .C0(index_i[7]), .Z(n22457));
    L6MUX21 i20143 (.D0(n22471), .D1(n22472), .SD(index_i[6]), .Z(n22482));
    L6MUX21 i20144 (.D0(n22473), .D1(n22474), .SD(index_i[6]), .Z(n22483));
    L6MUX21 i20147 (.D0(n22479), .D1(n22480), .SD(index_i[7]), .Z(n22486));
    L6MUX21 i20154 (.D0(n382_adj_2272), .D1(n509_adj_2273), .SD(index_q[7]), 
            .Z(n22493));
    LUT4 i11662_2_lut_rep_470_3_lut (.A(index_q[1]), .B(index_q[2]), .C(index_q[0]), 
         .Z(n26430)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11662_2_lut_rep_470_3_lut.init = 16'h8080;
    L6MUX21 i20170 (.D0(n22503), .D1(n22504), .SD(index_q[7]), .Z(n22509));
    L6MUX21 i20171 (.D0(n22505), .D1(n22506), .SD(index_q[7]), .Z(n22510));
    PFUMX i18771 (.BLUT(n21089), .ALUT(n21090), .C0(index_q[4]), .Z(n21091));
    PFUMX i24479 (.BLUT(n26761), .ALUT(n26762), .C0(index_i[0]), .Z(n26763));
    L6MUX21 i20610 (.D0(n22943), .D1(n22944), .SD(index_i[7]), .Z(n22949));
    L6MUX21 i20625 (.D0(n22958), .D1(n22959), .SD(index_i[7]), .Z(n22964));
    PFUMX i20626 (.BLUT(n22960), .ALUT(n22961), .C0(index_i[7]), .Z(n22965));
    LUT4 mux_192_Mux_12_i254_4_lut (.A(n26372), .B(n20234), .C(index_q[6]), 
         .D(n29190), .Z(n254_adj_2274)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_12_i254_4_lut.init = 16'hca0a;
    L6MUX21 i20636 (.D0(n22973), .D1(n22974), .SD(index_i[7]), .Z(n22975));
    L6MUX21 i20291 (.D0(n22623), .D1(n22624), .SD(index_q[7]), .Z(n22630));
    L6MUX21 i20292 (.D0(n22625), .D1(n22626), .SD(index_q[7]), .Z(n22631));
    PFUMX i20293 (.BLUT(n22627), .ALUT(n22628), .C0(index_q[7]), .Z(n22632));
    LUT4 mux_191_Mux_6_i269_rep_639 (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .Z(n26599)) /* synthesis lut_function=(A (C)+!A !((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_6_i269_rep_639.init = 16'ha4a4;
    LUT4 i20582_3_lut (.A(n22918), .B(n22919), .C(index_q[7]), .Z(n22921)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20582_3_lut.init = 16'hcaca;
    L6MUX21 i19796 (.D0(n22129), .D1(n22130), .SD(index_q[7]), .Z(n22135));
    LUT4 n25084_bdd_3_lut (.A(n26748), .B(n444_adj_2275), .C(index_q[5]), 
         .Z(n25085)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n25084_bdd_3_lut.init = 16'hcaca;
    L6MUX21 i20377 (.D0(n22705), .D1(n22706), .SD(index_q[6]), .Z(n22716));
    L6MUX21 i20378 (.D0(n22707), .D1(n22708), .SD(index_q[6]), .Z(n22717));
    PFUMX i24539 (.BLUT(n26855), .ALUT(n26856), .C0(index_q[0]), .Z(n26857));
    L6MUX21 i20381 (.D0(n22713), .D1(n22714), .SD(index_q[7]), .Z(n22720));
    LUT4 i18758_3_lut (.A(n29200), .B(n26718), .C(index_q[3]), .Z(n21078)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18758_3_lut.init = 16'hcaca;
    LUT4 i18757_3_lut (.A(n26571), .B(n676), .C(index_q[3]), .Z(n21077)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18757_3_lut.init = 16'hcaca;
    LUT4 i21823_3_lut (.A(n21077), .B(n21078), .C(index_q[4]), .Z(n21079)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21823_3_lut.init = 16'hcaca;
    LUT4 i11271_2_lut_rep_451_3_lut_4_lut (.A(index_q[2]), .B(index_q[0]), 
         .C(index_q[3]), .D(index_q[1]), .Z(n26411)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11271_2_lut_rep_451_3_lut_4_lut.init = 16'hf0e0;
    L6MUX21 i19877 (.D0(n22208), .D1(n22209), .SD(index_q[7]), .Z(n22216));
    L6MUX21 i19878 (.D0(n22210), .D1(n22211), .SD(index_q[7]), .Z(n22217));
    PFUMX mux_191_Mux_3_i763 (.BLUT(n747_adj_2276), .ALUT(n762), .C0(index_i[4]), 
          .Z(n763)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    L6MUX21 i20795 (.D0(n23129), .D1(n23130), .SD(index_i[6]), .Z(n23134));
    LUT4 mux_192_Mux_6_i540_3_lut_3_lut_rep_761 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n26721)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_6_i540_3_lut_3_lut_rep_761.init = 16'h9393;
    PFUMX i19942 (.BLUT(n797), .ALUT(n828_adj_2277), .C0(index_q[5]), 
          .Z(n22281));
    L6MUX21 i19946 (.D0(n22269), .D1(n22270), .SD(index_q[6]), .Z(n22285));
    L6MUX21 i19947 (.D0(n22271), .D1(n22272), .SD(index_q[6]), .Z(n22286));
    L6MUX21 i19948 (.D0(n22273), .D1(n22274), .SD(index_q[6]), .Z(n22287));
    LUT4 mux_192_Mux_0_i986_3_lut (.A(n29196), .B(n985), .C(index_q[3]), 
         .Z(n986)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_0_i986_3_lut.init = 16'hcaca;
    L6MUX21 i19949 (.D0(n22275), .D1(n22276), .SD(index_q[6]), .Z(n22288));
    LUT4 mux_192_Mux_4_i812_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[2]), 
         .C(index_q[4]), .D(index_q[3]), .Z(n812)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A !(B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_4_i812_3_lut_4_lut_4_lut.init = 16'ha595;
    L6MUX21 i19950 (.D0(n22277), .D1(n22278), .SD(index_q[6]), .Z(n22289));
    L6MUX21 i19953 (.D0(n22283), .D1(n22284), .SD(index_q[6]), .Z(n22292));
    PFUMX i19962 (.BLUT(n12014), .ALUT(n21349), .C0(index_q[6]), .Z(n22301));
    LUT4 mux_192_Mux_0_i971_3_lut (.A(n29198), .B(n29185), .C(index_q[3]), 
         .Z(n971)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_0_i971_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_0_i939_4_lut (.A(n931), .B(n26711), .C(index_q[3]), 
         .D(index_q[2]), .Z(n939)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_0_i939_4_lut.init = 16'hfaca;
    LUT4 i20581_3_lut (.A(n22916), .B(n22917), .C(index_q[7]), .Z(n22920)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20581_3_lut.init = 16'hcaca;
    L6MUX21 i19964 (.D0(n21355), .D1(n21358), .SD(index_q[6]), .Z(n22303));
    L6MUX21 i19965 (.D0(n574), .D1(n21361), .SD(index_q[6]), .Z(n22304));
    L6MUX21 i19966 (.D0(n21364), .D1(n764), .SD(index_q[6]), .Z(n22305));
    L6MUX21 i19983 (.D0(n22680), .D1(n22687), .SD(index_i[6]), .Z(n22322));
    L6MUX21 i19986 (.D0(n21322), .D1(n21325), .SD(index_i[6]), .Z(n22325));
    L6MUX21 i19987 (.D0(n21328), .D1(n21331), .SD(index_i[6]), .Z(n22326));
    L6MUX21 i19988 (.D0(n21334), .D1(n21337), .SD(index_i[6]), .Z(n22327));
    PFUMX i19989 (.BLUT(n21340), .ALUT(n892), .C0(index_i[6]), .Z(n22328));
    LUT4 i1_3_lut_4_lut (.A(index_q[1]), .B(index_q[2]), .C(index_q[5]), 
         .D(n26584), .Z(n20006)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_3_lut_4_lut.init = 16'hfff8;
    LUT4 i15394_3_lut_3_lut (.A(index_q[0]), .B(index_q[2]), .C(index_q[3]), 
         .Z(n17544)) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i15394_3_lut_3_lut.init = 16'h6a6a;
    PFUMX i24535 (.BLUT(n26849), .ALUT(n26850), .C0(index_q[1]), .Z(n26851));
    PFUMX i20481 (.BLUT(n22816), .ALUT(n22817), .C0(index_q[6]), .Z(n22820));
    PFUMX i20482 (.BLUT(n22818), .ALUT(n22819), .C0(index_q[6]), .Z(n22821));
    LUT4 mux_192_Mux_0_i923_3_lut (.A(n29182), .B(n29189), .C(index_q[3]), 
         .Z(n923)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_0_i923_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_1_i62_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[2]), 
         .C(index_q[4]), .D(index_q[3]), .Z(n62_adj_2278)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))+!A !(B (C)+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_1_i62_3_lut_4_lut_4_lut.init = 16'ha5a6;
    LUT4 mux_192_Mux_8_i491_3_lut_4_lut_3_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[0]), .D(index_q[3]), .Z(n491_adj_2279)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(D))+!A !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_8_i491_3_lut_4_lut_3_lut_4_lut.init = 16'h7780;
    L6MUX21 i20014 (.D0(n22337), .D1(n22338), .SD(index_i[6]), .Z(n22353));
    LUT4 i9369_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n11815)) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B ((D)+!C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9369_3_lut_4_lut_4_lut.init = 16'hcdad;
    LUT4 i9366_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n11812)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))+!A !(B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9366_3_lut_4_lut_4_lut.init = 16'hb5b3;
    LUT4 i21619_3_lut (.A(n109), .B(n124), .C(index_q[4]), .Z(n21345)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21619_3_lut.init = 16'hcaca;
    LUT4 i19322_3_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[0]), .C(index_i[1]), 
         .D(index_i[3]), .Z(n21642)) /* synthesis lut_function=(A (B (C)+!B !(C+!(D)))+!A (B (C)+!B !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19322_3_lut_4_lut_4_lut.init = 16'hc3d0;
    LUT4 mux_192_Mux_2_i890_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n890_adj_2280)) /* synthesis lut_function=(A (B (C)+!B !(C+!(D)))+!A !(B (C+(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_2_i890_3_lut_4_lut_4_lut.init = 16'h9394;
    LUT4 i20220_3_lut_4_lut (.A(n26496), .B(index_q[3]), .C(index_q[4]), 
         .D(n364_adj_2281), .Z(n22559)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20220_3_lut_4_lut.init = 16'h8f80;
    PFUMX i24530 (.BLUT(n26842), .ALUT(n26843), .C0(index_i[2]), .Z(n26844));
    LUT4 i9434_3_lut_4_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n844_adj_2282)) /* synthesis lut_function=(A (B)+!A !(B+!(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9434_3_lut_4_lut_3_lut_4_lut.init = 16'h9998;
    L6MUX21 i20015 (.D0(n22339), .D1(n22340), .SD(index_i[6]), .Z(n22354));
    LUT4 i9563_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n12009)) /* synthesis lut_function=(A (B (D)+!B !((D)+!C))+!A (((D)+!C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9563_3_lut_4_lut_4_lut_4_lut.init = 16'hdd35;
    L6MUX21 i20016 (.D0(n22341), .D1(n22342), .SD(index_i[6]), .Z(n22355));
    LUT4 i19376_3_lut_4_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n21696)) /* synthesis lut_function=(!(A (B (C)+!B (C+(D)))+!A !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19376_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'h585f;
    LUT4 mux_192_Mux_3_i189_3_lut_3_lut_4_lut (.A(n26496), .B(index_q[3]), 
         .C(index_q[4]), .D(n26457), .Z(n189)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_3_i189_3_lut_3_lut_4_lut.init = 16'h08f8;
    LUT4 mux_191_Mux_7_i491_3_lut_4_lut_4_lut_4_lut_4_lut (.A(index_i[1]), 
         .B(index_i[3]), .C(index_i[2]), .D(index_i[0]), .Z(n491_adj_2283)) /* synthesis lut_function=(!(A (B (C+!(D))+!B ((D)+!C))+!A !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_7_i491_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'h5870;
    L6MUX21 i20017 (.D0(n22343), .D1(n22344), .SD(index_i[6]), .Z(n22356));
    LUT4 i9410_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n11856)) /* synthesis lut_function=(!(A (B (C)+!B ((D)+!C))+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9410_3_lut_4_lut_4_lut.init = 16'h4969;
    LUT4 mux_192_Mux_10_i637_3_lut_4_lut_4_lut (.A(n26497), .B(index_q[4]), 
         .C(index_q[5]), .D(n26411), .Z(n637)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_10_i637_3_lut_4_lut_4_lut.init = 16'h1f1c;
    LUT4 i9554_3_lut_4_lut_3_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n875)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(D))+!A (B (C+!(D))+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9554_3_lut_4_lut_3_lut_3_lut_4_lut.init = 16'hc07f;
    LUT4 i11289_3_lut_3_lut_3_lut_rep_802 (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[0]), .Z(n29181)) /* synthesis lut_function=(!(A+!(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11289_3_lut_3_lut_3_lut_rep_802.init = 16'h4545;
    LUT4 mux_191_Mux_0_i443_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .D(index_i[3]), .Z(n443)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C (D))+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_0_i443_3_lut_4_lut_4_lut_4_lut.init = 16'h0ed5;
    LUT4 i21626_3_lut (.A(n620_adj_2284), .B(n14085), .C(index_i[4]), 
         .Z(n21330)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21626_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_2_i142_3_lut_4_lut_4_lut_4_lut_4_lut (.A(index_q[1]), 
         .B(index_q[2]), .C(index_q[0]), .D(index_q[3]), .Z(n142)) /* synthesis lut_function=(!(A (B)+!A (B (D)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_2_i142_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'h3266;
    LUT4 mux_192_Mux_2_i716_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), 
         .B(index_q[2]), .C(index_q[3]), .D(index_q[0]), .Z(n716)) /* synthesis lut_function=(!(A (B)+!A !(B (C+!(D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_2_i716_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h6367;
    LUT4 i18743_3_lut (.A(n900), .B(n325), .C(index_q[3]), .Z(n21063)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18743_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_9_i30_3_lut_4_lut_4_lut_4_lut (.A(index_q[2]), .B(index_q[3]), 
         .C(index_q[1]), .D(index_q[0]), .Z(n30)) /* synthesis lut_function=(A (B (C (D)))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_9_i30_3_lut_4_lut_4_lut_4_lut.init = 16'h9111;
    PFUMX i24475 (.BLUT(n26755), .ALUT(n26756), .C0(index_i[1]), .Z(n26757));
    LUT4 mux_192_Mux_0_i781_4_lut_4_lut_4_lut (.A(index_q[2]), .B(index_q[3]), 
         .C(index_q[1]), .D(index_q[0]), .Z(n781_adj_2285)) /* synthesis lut_function=(!(A (B+!((D)+!C))+!A !(B (C)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_0_i781_4_lut_4_lut_4_lut.init = 16'h6252;
    LUT4 n77_bdd_3_lut_24032_3_lut_4_lut_4_lut_3_lut_4_lut (.A(index_q[2]), 
         .B(index_q[3]), .C(index_q[0]), .D(index_q[1]), .Z(n25592)) /* synthesis lut_function=(A (B (C (D)))+!A (B+!(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n77_bdd_3_lut_24032_3_lut_4_lut_4_lut_3_lut_4_lut.init = 16'hc555;
    L6MUX21 i20018 (.D0(n22345), .D1(n22346), .SD(index_i[6]), .Z(n22357));
    LUT4 mux_192_Mux_7_i526_3_lut_3_lut_4_lut_4_lut_3_lut_4_lut (.A(index_q[2]), 
         .B(index_q[3]), .C(index_q[0]), .D(index_q[1]), .Z(n526_adj_2286)) /* synthesis lut_function=(A (C (D))+!A !(B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_7_i526_3_lut_3_lut_4_lut_4_lut_3_lut_4_lut.init = 16'hb555;
    LUT4 mux_191_Mux_1_i908_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[3]), 
         .C(index_i[2]), .D(index_i[0]), .Z(n908)) /* synthesis lut_function=(!(A (B+(C))+!A !(B+(C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_1_i908_3_lut_4_lut_4_lut_4_lut.init = 16'h5647;
    LUT4 mux_192_Mux_0_i46_3_lut_4_lut_4_lut_4_lut (.A(index_q[2]), .B(index_q[3]), 
         .C(index_q[1]), .D(index_q[0]), .Z(n46)) /* synthesis lut_function=(A (B)+!A ((C+(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_0_i46_3_lut_4_lut_4_lut_4_lut.init = 16'hddd9;
    LUT4 mux_192_Mux_0_i428_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_q[2]), 
         .B(index_q[0]), .C(index_q[1]), .D(index_q[3]), .Z(n428)) /* synthesis lut_function=(A (B (C+!(D))+!B !((D)+!C))+!A (B (D)+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_0_i428_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hd5a9;
    LUT4 mux_192_Mux_8_i716_3_lut_4_lut_4_lut_4_lut (.A(index_q[2]), .B(index_q[3]), 
         .C(index_q[1]), .D(index_q[0]), .Z(n716_adj_2287)) /* synthesis lut_function=(!(A (B)+!A !(B+(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_8_i716_3_lut_4_lut_4_lut_4_lut.init = 16'h7776;
    LUT4 mux_192_Mux_4_i541_3_lut_4_lut_3_lut_4_lut (.A(index_q[2]), .B(index_q[3]), 
         .C(index_q[0]), .D(index_q[1]), .Z(n541_adj_2288)) /* synthesis lut_function=(!(A (B+!(C+(D)))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_4_i541_3_lut_4_lut_3_lut_4_lut.init = 16'h6664;
    LUT4 mux_191_Mux_0_i1017_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n1017)) /* synthesis lut_function=(A (B (C)+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_0_i1017_4_lut_4_lut_4_lut.init = 16'hd7d0;
    LUT4 i20297_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[3]), 
         .C(index_i[2]), .D(index_i[0]), .Z(n22636)) /* synthesis lut_function=(A (B (C (D))+!B (C))+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20297_3_lut_4_lut_4_lut_4_lut.init = 16'hb434;
    LUT4 mux_192_Mux_0_i604_3_lut_4_lut_4_lut_4_lut (.A(index_q[2]), .B(index_q[0]), 
         .C(index_q[1]), .D(index_q[3]), .Z(n604)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A !(B (D)+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_0_i604_3_lut_4_lut_4_lut_4_lut.init = 16'h5439;
    LUT4 i7656_2_lut_rep_662 (.A(index_q[3]), .B(index_q[4]), .Z(n26622)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i7656_2_lut_rep_662.init = 16'h8888;
    LUT4 mux_191_Mux_1_i348_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[3]), 
         .C(index_i[2]), .D(index_i[0]), .Z(n348)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_1_i348_3_lut_4_lut_4_lut_4_lut.init = 16'h7870;
    LUT4 i19478_3_lut_4_lut_4_lut_4_lut_4_lut (.A(index_q[2]), .B(index_q[0]), 
         .C(index_q[1]), .D(index_q[3]), .Z(n21798)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19478_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'h0fd5;
    LUT4 i18788_3_lut_4_lut_4_lut_4_lut (.A(index_q[2]), .B(index_q[3]), 
         .C(index_q[1]), .D(index_q[0]), .Z(n21108)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18788_3_lut_4_lut_4_lut_4_lut.init = 16'h6444;
    LUT4 mux_192_Mux_8_i635_3_lut_4_lut_3_lut_4_lut (.A(index_q[2]), .B(index_q[3]), 
         .C(index_q[0]), .D(index_q[1]), .Z(n635_adj_2289)) /* synthesis lut_function=(!(A (B)+!A !(B+(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_8_i635_3_lut_4_lut_3_lut_4_lut.init = 16'h7666;
    LUT4 mux_191_Mux_2_i890_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n890_adj_2265)) /* synthesis lut_function=(A (B (C)+!B !(C+!(D)))+!A !(B (C+(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_2_i890_3_lut_4_lut_4_lut.init = 16'h9394;
    L6MUX21 i20020 (.D0(n22349), .D1(n22350), .SD(index_i[6]), .Z(n22359));
    LUT4 mux_191_Mux_8_i860_3_lut_4_lut (.A(n26505), .B(index_i[3]), .C(index_i[4]), 
         .D(n26472), .Z(n860_adj_2290)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_8_i860_3_lut_4_lut.init = 16'h08f8;
    LUT4 n526_bdd_3_lut_24088_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n25274)) /* synthesis lut_function=(!(A (B)+!A !(B (C+(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n526_bdd_3_lut_24088_4_lut_4_lut_4_lut.init = 16'h6663;
    LUT4 i20199_3_lut_4_lut (.A(n26505), .B(index_i[3]), .C(index_i[4]), 
         .D(n364_adj_2291), .Z(n22538)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20199_3_lut_4_lut.init = 16'h8f80;
    LUT4 i9552_3_lut_4_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n844_adj_2267)) /* synthesis lut_function=(A (B)+!A !(B+!(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9552_3_lut_4_lut_3_lut_4_lut.init = 16'h9998;
    LUT4 mux_191_Mux_4_i93_3_lut_4_lut_3_lut_rep_633_4_lut (.A(index_i[0]), 
         .B(index_i[3]), .C(index_i[1]), .D(index_i[2]), .Z(n26593)) /* synthesis lut_function=(!(A (B+(C (D)))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_4_i93_3_lut_4_lut_3_lut_rep_633_4_lut.init = 16'h4666;
    LUT4 i19301_3_lut_4_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[3]), 
         .C(index_i[1]), .D(index_i[2]), .Z(n21621)) /* synthesis lut_function=(A (B+(C (D)))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19301_3_lut_4_lut_3_lut_4_lut.init = 16'hb999;
    LUT4 mux_191_Mux_10_i62_3_lut_3_lut_4_lut (.A(n26505), .B(index_i[3]), 
         .C(n26472), .D(index_i[4]), .Z(n62_adj_2292)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_10_i62_3_lut_3_lut_4_lut.init = 16'hf077;
    LUT4 i19370_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n21690)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(D))+!A (B (D)+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19370_3_lut_4_lut_4_lut_4_lut.init = 16'hd52b;
    LUT4 i9566_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n12012)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D))+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9566_3_lut_4_lut_4_lut_4_lut.init = 16'hcadd;
    LUT4 i19229_3_lut (.A(n404), .B(n26695), .C(index_i[3]), .Z(n21549)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19229_3_lut.init = 16'hcaca;
    LUT4 mux_191_Mux_4_i812_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[4]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n812_adj_2293)) /* synthesis lut_function=(A (B (C+(D)))+!A !(B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_4_i812_3_lut_3_lut_4_lut.init = 16'h9995;
    PFUMX i24526 (.BLUT(n26835), .ALUT(n26836), .C0(index_i[1]), .Z(n26837));
    LUT4 mux_191_Mux_6_i955_3_lut_4_lut (.A(n26505), .B(index_i[3]), .C(index_i[4]), 
         .D(n26359), .Z(n955)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_6_i955_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_191_Mux_3_i252_3_lut_4_lut (.A(n26505), .B(index_i[3]), .C(index_i[4]), 
         .D(n15026), .Z(n252_adj_2294)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_3_i252_3_lut_4_lut.init = 16'h08f8;
    LUT4 i15423_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[1]), .Z(n17573)) /* synthesis lut_function=(A (B (C (D))+!B !(C))+!A (B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i15423_3_lut_4_lut_4_lut_4_lut.init = 16'hd656;
    LUT4 i11369_2_lut_rep_394_3_lut_4_lut (.A(n26505), .B(index_i[3]), .C(index_i[5]), 
         .D(index_i[4]), .Z(n26354)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11369_2_lut_rep_394_3_lut_4_lut.init = 16'hf080;
    LUT4 mux_191_Mux_3_i189_3_lut_3_lut_4_lut (.A(n26505), .B(index_i[3]), 
         .C(index_i[4]), .D(n26470), .Z(n189_adj_2295)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_3_i189_3_lut_3_lut_4_lut.init = 16'h08f8;
    LUT4 i22266_3_lut (.A(n24169), .B(n22495), .C(index_q[8]), .Z(n22497)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22266_3_lut.init = 16'hcaca;
    LUT4 mux_191_Mux_10_i637_3_lut_4_lut_4_lut (.A(n26506), .B(index_i[4]), 
         .C(index_i[5]), .D(n26414), .Z(n637_adj_2296)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_10_i637_3_lut_4_lut_4_lut.init = 16'h1f1c;
    LUT4 mux_191_Mux_3_i507_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[4]), .D(n491_adj_2297), .Z(n507_adj_2298)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_3_i507_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_192_Mux_4_i93_3_lut_4_lut_3_lut_rep_623_4_lut (.A(index_q[0]), 
         .B(index_q[3]), .C(index_q[1]), .D(index_q[2]), .Z(n26583)) /* synthesis lut_function=(!(A (B+(C (D)))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_4_i93_3_lut_4_lut_3_lut_rep_623_4_lut.init = 16'h4666;
    LUT4 i19228_3_lut (.A(n26697), .B(n396), .C(index_i[3]), .Z(n21548)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19228_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_535_3_lut (.A(index_q[3]), .B(index_q[4]), .C(index_q[5]), 
         .Z(n26495)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_2_lut_rep_535_3_lut.init = 16'hf8f8;
    L6MUX21 i20045 (.D0(n22368), .D1(n22369), .SD(index_i[6]), .Z(n22384));
    LUT4 mux_192_Mux_0_i747_3_lut_4_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[2]), 
         .C(index_q[3]), .D(index_q[1]), .Z(n747_adj_2299)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C+(D)))+!A !(B ((D)+!C)+!B (C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_0_i747_3_lut_4_lut_3_lut_4_lut.init = 16'h5596;
    L6MUX21 i20046 (.D0(n22370), .D1(n22371), .SD(index_i[6]), .Z(n22385));
    L6MUX21 i20047 (.D0(n22372), .D1(n22373), .SD(index_i[6]), .Z(n22386));
    LUT4 i19343_3_lut_4_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n21663)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19343_3_lut_4_lut_4_lut_4_lut.init = 16'h6444;
    LUT4 n518_bdd_3_lut_4_lut_4_lut_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[0]), .D(index_i[1]), .Z(n25272)) /* synthesis lut_function=(A (B (C (D)))+!A (B+!(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n518_bdd_3_lut_4_lut_4_lut_3_lut_4_lut.init = 16'hc555;
    LUT4 mux_191_Mux_8_i635_3_lut_4_lut_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[0]), .D(index_i[1]), .Z(n635_adj_2300)) /* synthesis lut_function=(!(A (B)+!A !(B+(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_8_i635_3_lut_4_lut_3_lut_4_lut.init = 16'h7666;
    LUT4 mux_191_Mux_9_i30_3_lut_4_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n30_adj_2301)) /* synthesis lut_function=(A (B (C (D)))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_9_i30_3_lut_4_lut_4_lut_4_lut.init = 16'h9111;
    LUT4 mux_191_Mux_7_i526_3_lut_3_lut_4_lut_4_lut_3_lut_4_lut (.A(index_i[2]), 
         .B(index_i[3]), .C(index_i[0]), .D(index_i[1]), .Z(n526_adj_2302)) /* synthesis lut_function=(A (C (D))+!A !(B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_7_i526_3_lut_3_lut_4_lut_4_lut_3_lut_4_lut.init = 16'hb555;
    PFUMX i24524 (.BLUT(n26832), .ALUT(n26833), .C0(index_i[0]), .Z(n26834));
    PFUMX i20049 (.BLUT(n22376), .ALUT(n22377), .C0(index_i[6]), .Z(n22388));
    LUT4 mux_192_Mux_6_i781_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), 
         .B(index_q[2]), .C(index_q[3]), .D(index_q[0]), .Z(n781_adj_2303)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+(D)))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_6_i781_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h9993;
    LUT4 i11058_2_lut_rep_582 (.A(index_q[0]), .B(index_q[1]), .Z(n26542)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11058_2_lut_rep_582.init = 16'h4444;
    LUT4 n205_bdd_3_lut_24036_4_lut_3_lut_4_lut (.A(index_q[1]), .B(index_q[3]), 
         .C(index_q[2]), .D(index_q[0]), .Z(n25594)) /* synthesis lut_function=(!(A (B (D)+!B ((D)+!C))+!A !(B (D)+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n205_bdd_3_lut_24036_4_lut_3_lut_4_lut.init = 16'h55a9;
    LUT4 i9402_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[0]), 
         .C(index_q[4]), .D(n26539), .Z(n221_adj_2304)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A !(B+(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9402_3_lut_4_lut_4_lut_4_lut.init = 16'h5556;
    LUT4 i9425_3_lut_4_lut_3_lut_4_lut (.A(index_q[1]), .B(index_q[3]), 
         .C(index_q[4]), .D(index_q[0]), .Z(n444_adj_2275)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A !(((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9425_3_lut_4_lut_3_lut_4_lut.init = 16'h5595;
    LUT4 i18736_3_lut (.A(n29200), .B(n29181), .C(index_q[3]), .Z(n21056)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18736_3_lut.init = 16'hcaca;
    LUT4 n812_bdd_3_lut_24256_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[3]), 
         .C(index_q[2]), .D(index_q[0]), .Z(n25447)) /* synthesis lut_function=(A (C)+!A (B ((D)+!C)+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n812_bdd_3_lut_24256_4_lut_4_lut_4_lut.init = 16'hf4b4;
    LUT4 mux_192_Mux_2_i908_3_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[0]), .D(index_q[3]), .Z(n908_adj_2305)) /* synthesis lut_function=(!(A (B+!(D))+!A !(B+!(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_2_i908_3_lut_4_lut_4_lut.init = 16'h6645;
    LUT4 n53_bdd_3_lut_23515 (.A(n26653), .B(n29180), .C(index_i[3]), 
         .Z(n25206)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n53_bdd_3_lut_23515.init = 16'hcaca;
    LUT4 mux_192_Mux_0_i443_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[0]), .D(index_q[3]), .Z(n443_adj_2306)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C (D))+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_0_i443_3_lut_4_lut_4_lut_4_lut.init = 16'h0ed5;
    LUT4 i19487_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .D(index_q[0]), .Z(n21807)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B (C+!(D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19487_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h1c18;
    LUT4 mux_192_Mux_2_i173_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .D(index_q[0]), .Z(n173_adj_2307)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_2_i173_3_lut_4_lut_4_lut_4_lut.init = 16'h0e1e;
    L6MUX21 i20050 (.D0(n22378), .D1(n22379), .SD(index_i[6]), .Z(n22389));
    LUT4 n21233_bdd_4_lut_24430 (.A(n26547), .B(n763_adj_2308), .C(index_i[5]), 
         .D(index_i[4]), .Z(n24125)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam n21233_bdd_4_lut_24430.init = 16'hcfca;
    LUT4 n708_bdd_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .D(index_q[0]), .Z(n25584)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n708_bdd_3_lut_4_lut_4_lut_4_lut.init = 16'h1e1c;
    L6MUX21 i20051 (.D0(n22380), .D1(n22381), .SD(index_i[6]), .Z(n22390));
    PFUMX i20052 (.BLUT(n22382), .ALUT(n22383), .C0(index_i[6]), .Z(n22391));
    LUT4 mux_192_Mux_4_i349_3_lut_4_lut (.A(index_q[0]), .B(index_q[2]), 
         .C(index_q[4]), .D(n348_adj_2309), .Z(n349)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_4_i349_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_192_Mux_7_i747_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), 
         .B(index_q[2]), .C(index_q[3]), .D(index_q[0]), .Z(n747_adj_2310)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))+!A (B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_7_i747_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'he1e3;
    LUT4 mux_192_Mux_0_i14_3_lut_rep_803 (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[0]), .Z(n29182)) /* synthesis lut_function=(A (B)+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_0_i14_3_lut_rep_803.init = 16'hd9d9;
    PFUMX i20072 (.BLUT(n797_adj_2311), .ALUT(n828_adj_2312), .C0(index_i[5]), 
          .Z(n22411));
    LUT4 n953_bdd_3_lut (.A(n26685), .B(n619), .C(index_i[3]), .Z(n25216)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n953_bdd_3_lut.init = 16'hcaca;
    LUT4 i20479_3_lut_3_lut_4_lut (.A(index_q[3]), .B(index_q[4]), .C(n413_adj_2313), 
         .D(index_q[5]), .Z(n22818)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20479_3_lut_3_lut_4_lut.init = 16'h77f0;
    LUT4 mux_191_Mux_4_i773_3_lut_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n773)) /* synthesis lut_function=(!(A (B+(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_4_i773_3_lut_3_lut_3_lut.init = 16'h5656;
    LUT4 n45_bdd_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n25328)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n45_bdd_3_lut_4_lut_4_lut_4_lut.init = 16'h1e1c;
    LUT4 mux_191_Mux_2_i173_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n173_adj_2314)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_2_i173_3_lut_4_lut_4_lut_4_lut.init = 16'h0e1e;
    LUT4 i1_2_lut_3_lut (.A(index_q[3]), .B(index_q[4]), .C(index_q[5]), 
         .Z(n20234)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_2_lut_3_lut.init = 16'h8080;
    LUT4 mux_191_Mux_7_i747_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n747_adj_2315)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))+!A (B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_7_i747_3_lut_4_lut_4_lut_4_lut.init = 16'he1e3;
    LUT4 index_i_5__bdd_4_lut_23648 (.A(n619), .B(index_i[2]), .C(index_i[3]), 
         .D(n26647), .Z(n25227)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (B+!(C (D))))) */ ;
    defparam index_i_5__bdd_4_lut_23648.init = 16'h3a0a;
    LUT4 i20205_3_lut_4_lut (.A(n26519), .B(index_i[3]), .C(index_i[4]), 
         .D(n26455), .Z(n22544)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20205_3_lut_4_lut.init = 16'hfe0e;
    LUT4 n300_bdd_3_lut_23546 (.A(n26587), .B(n26710), .C(index_i[3]), 
         .Z(n25229)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n300_bdd_3_lut_23546.init = 16'hcaca;
    LUT4 mux_191_Mux_10_i252_3_lut_4_lut_4_lut (.A(n26519), .B(index_i[3]), 
         .C(index_i[4]), .D(n26486), .Z(n252_adj_2316)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B (C (D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_10_i252_3_lut_4_lut_4_lut.init = 16'h3efe;
    LUT4 mux_191_Mux_3_i828_3_lut_3_lut_4_lut (.A(n26519), .B(index_i[3]), 
         .C(n157_adj_2317), .D(index_i[4]), .Z(n828_adj_2312)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_3_i828_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 mux_192_Mux_0_i15_3_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[0]), .D(index_q[3]), .Z(n15)) /* synthesis lut_function=(A (B)+!A ((C (D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_0_i15_3_lut_4_lut_4_lut.init = 16'hd999;
    LUT4 i19280_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[1]), .Z(n21600)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C))+!A (B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19280_3_lut_4_lut_4_lut_4_lut.init = 16'h29a9;
    LUT4 mux_192_Mux_8_i251_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), 
         .B(index_q[1]), .C(index_q[2]), .D(index_q[3]), .Z(n251)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_8_i251_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h07e0;
    LUT4 mux_191_Mux_10_i413_3_lut_3_lut_4_lut (.A(n26519), .B(index_i[3]), 
         .C(n26470), .D(index_i[4]), .Z(n413_adj_2318)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_10_i413_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 i20203_3_lut_3_lut_4_lut (.A(n26519), .B(index_i[3]), .C(n412_adj_2319), 
         .D(index_i[4]), .Z(n22542)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20203_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 n442_bdd_3_lut_23552 (.A(n26700), .B(n29180), .C(index_i[3]), 
         .Z(n25233)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n442_bdd_3_lut_23552.init = 16'hcaca;
    LUT4 mux_192_Mux_6_i844_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n844_adj_2320)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (B (C)+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_6_i844_3_lut_4_lut_4_lut.init = 16'hc1e0;
    LUT4 i20419_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n22758)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20419_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hf81f;
    LUT4 mux_192_Mux_6_i859_3_lut_rep_427_4_lut_4_lut_4_lut (.A(index_q[0]), 
         .B(index_q[1]), .C(index_q[2]), .D(index_q[3]), .Z(n26387)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A (B (C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_6_i859_3_lut_rep_427_4_lut_4_lut_4_lut.init = 16'he0f8;
    LUT4 mux_191_Mux_7_i364_3_lut_3_lut (.A(n26650), .B(index_i[3]), .C(n26652), 
         .Z(n364_adj_2321)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;
    defparam mux_191_Mux_7_i364_3_lut_3_lut.init = 16'hd1d1;
    LUT4 i9547_3_lut_3_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[0]), .D(index_i[1]), .Z(n762)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C (D)+!C !(D)))+!A !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9547_3_lut_3_lut_4_lut_4_lut.init = 16'h700f;
    L6MUX21 i20076 (.D0(n22399), .D1(n22400), .SD(index_i[6]), .Z(n22415));
    LUT4 i19310_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n21630)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C))+!A (B (C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19310_3_lut_4_lut_4_lut_4_lut.init = 16'he078;
    LUT4 i20520_3_lut (.A(n22856), .B(n22857), .C(index_i[7]), .Z(n22859)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20520_3_lut.init = 16'hcaca;
    LUT4 i18725_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[2]), 
         .C(index_q[3]), .D(index_q[1]), .Z(n21045)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C))+!A (B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18725_3_lut_4_lut_4_lut_4_lut.init = 16'h29a9;
    L6MUX21 i20077 (.D0(n22401), .D1(n22402), .SD(index_i[6]), .Z(n22416));
    L6MUX21 i20078 (.D0(n22403), .D1(n22404), .SD(index_i[6]), .Z(n22417));
    LUT4 i20298_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n22637)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20298_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hf81f;
    L6MUX21 i20079 (.D0(n22405), .D1(n22406), .SD(index_i[6]), .Z(n22418));
    LUT4 i22411_2_lut_rep_413_3_lut_4_lut (.A(n26647), .B(index_i[2]), .C(index_i[5]), 
         .D(n26595), .Z(n26373)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i22411_2_lut_rep_413_3_lut_4_lut.init = 16'h0f7f;
    L6MUX21 i20080 (.D0(n22407), .D1(n22408), .SD(index_i[6]), .Z(n22419));
    L6MUX21 i20515 (.D0(n22846), .D1(n22847), .SD(index_i[6]), .Z(n22854));
    L6MUX21 i20083 (.D0(n22413), .D1(n22414), .SD(index_i[6]), .Z(n22422));
    L6MUX21 i20518 (.D0(n22852), .D1(n22853), .SD(index_i[6]), .Z(n22857));
    LUT4 mux_191_Mux_8_i61_3_lut_rep_428_4_lut_4_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[2]), .D(index_i[3]), .Z(n26388)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A (B (C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_8_i61_3_lut_rep_428_4_lut_4_lut_4_lut.init = 16'he0f8;
    LUT4 i11266_3_lut (.A(index_q[2]), .B(index_q[1]), .C(index_q[0]), 
         .Z(n676)) /* synthesis lut_function=(!(A (B (C))+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11266_3_lut.init = 16'h3b3b;
    LUT4 i20299_3_lut_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n22638)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C+!(D))+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20299_3_lut_3_lut_4_lut_4_lut.init = 16'h1f81;
    L6MUX21 i20108 (.D0(n22432), .D1(n22433), .SD(index_i[6]), .Z(n22447));
    L6MUX21 i20109 (.D0(n22434), .D1(n22435), .SD(index_i[6]), .Z(n22448));
    L6MUX21 i20110 (.D0(n22436), .D1(n22437), .SD(index_i[6]), .Z(n22449));
    LUT4 mux_191_Mux_8_i251_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n251_adj_2322)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_8_i251_3_lut_4_lut_4_lut_4_lut.init = 16'h07e0;
    LUT4 mux_192_Mux_0_i890_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n890_adj_2323)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)+!C !(D)))+!A !(B (C)+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_0_i890_3_lut_4_lut_4_lut.init = 16'h70ca;
    L6MUX21 i20111 (.D0(n22438), .D1(n22439), .SD(index_i[6]), .Z(n22450));
    L6MUX21 i20112 (.D0(n22440), .D1(n22441), .SD(index_i[6]), .Z(n22451));
    LUT4 mux_192_Mux_6_i890_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), 
         .B(index_q[1]), .C(index_q[2]), .D(index_q[3]), .Z(n890_adj_2324)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !((D)+!C))+!A !(B ((D)+!C)+!B (C (D)+!C !(D))))) */ ;
    defparam mux_192_Mux_6_i890_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h7e07;
    LUT4 mux_192_Mux_6_i378_3_lut_4_lut_3_lut_rep_764 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n26724)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_6_i378_3_lut_4_lut_3_lut_rep_764.init = 16'h4949;
    LUT4 i20516_3_lut (.A(n22848), .B(n27931), .C(index_i[6]), .Z(n22855)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20516_3_lut.init = 16'hcaca;
    LUT4 i20517_3_lut (.A(n25209), .B(n22851), .C(index_i[6]), .Z(n22856)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20517_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_6_i308_3_lut_4_lut_3_lut_rep_765 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n26725)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_6_i308_3_lut_4_lut_3_lut_rep_765.init = 16'h9696;
    LUT4 i20519_3_lut (.A(n22854), .B(n22855), .C(index_i[7]), .Z(n22858)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20519_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_7_i699_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n699)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (D))) */ ;
    defparam mux_192_Mux_7_i699_3_lut_4_lut_4_lut_4_lut.init = 16'hf70e;
    PFUMX i20133 (.BLUT(n732_adj_2325), .ALUT(n763_adj_2326), .C0(index_i[5]), 
          .Z(n22472));
    LUT4 i12488_1_lut_2_lut_3_lut_4_lut (.A(n26519), .B(index_i[3]), .C(index_i[5]), 
         .D(index_i[4]), .Z(n381)) /* synthesis lut_function=(!(A (C+(D))+!A (B (C+(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i12488_1_lut_2_lut_3_lut_4_lut.init = 16'h010f;
    LUT4 i19066_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n21386)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B+(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19066_3_lut_4_lut_4_lut_4_lut.init = 16'h2aab;
    LUT4 i11291_2_lut_rep_563_3_lut (.A(index_q[1]), .B(index_q[2]), .C(index_q[3]), 
         .Z(n26523)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11291_2_lut_rep_563_3_lut.init = 16'hf8f8;
    LUT4 mux_192_Mux_5_i252_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[4]), .Z(n252_adj_2327)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+(D)))+!A (B (C (D))+!B !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_5_i252_3_lut_4_lut.init = 16'hc993;
    L6MUX21 i20135 (.D0(n21721), .D1(n891_adj_2328), .SD(index_i[5]), 
            .Z(n22474));
    L6MUX21 i20138 (.D0(n22461), .D1(n22462), .SD(index_i[6]), .Z(n22477));
    L6MUX21 i20140 (.D0(n22465), .D1(n22466), .SD(index_i[6]), .Z(n22479));
    L6MUX21 i20141 (.D0(n22467), .D1(n22468), .SD(index_i[6]), .Z(n22480));
    L6MUX21 i20145 (.D0(n22475), .D1(n22476), .SD(index_i[6]), .Z(n22484));
    L6MUX21 i20577 (.D0(n22908), .D1(n22909), .SD(index_q[6]), .Z(n22916));
    LUT4 i9382_2_lut_rep_579 (.A(index_q[2]), .B(index_q[3]), .Z(n26539)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9382_2_lut_rep_579.init = 16'h8888;
    LUT4 i20056_3_lut (.A(n22390), .B(n22391), .C(index_i[7]), .Z(n22395)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20056_3_lut.init = 16'hcaca;
    LUT4 n24133_bdd_3_lut_25793 (.A(n24133), .B(n24126), .C(index_i[7]), 
         .Z(n24134)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n24133_bdd_3_lut_25793.init = 16'hcaca;
    L6MUX21 i20580 (.D0(n22914), .D1(n22915), .SD(index_q[6]), .Z(n22919));
    LUT4 n300_bdd_3_lut_24427 (.A(n26587), .B(n773), .C(index_i[3]), .Z(n25235)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n300_bdd_3_lut_24427.init = 16'hacac;
    L6MUX21 i20160 (.D0(n22801), .D1(n22808), .SD(index_q[6]), .Z(n22499));
    LUT4 i12093_2_lut_rep_663 (.A(index_q[2]), .B(index_q[0]), .Z(n26623)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12093_2_lut_rep_663.init = 16'heeee;
    LUT4 n21242_bdd_4_lut_24387 (.A(n26539), .B(n763_adj_2329), .C(index_q[5]), 
         .D(index_q[4]), .Z(n24160)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam n21242_bdd_4_lut_24387.init = 16'hcfca;
    LUT4 mux_191_Mux_1_i684_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n684_adj_2330)) /* synthesis lut_function=(A (B ((D)+!C)+!B !((D)+!C))+!A !(B (C+(D))+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_1_i684_3_lut_4_lut_4_lut.init = 16'h992d;
    LUT4 i20227_3_lut_3_lut_3_lut_4_lut (.A(index_q[2]), .B(index_q[3]), 
         .C(index_q[4]), .D(index_q[1]), .Z(n22566)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20227_3_lut_3_lut_3_lut_4_lut.init = 16'h878f;
    LUT4 mux_191_Mux_0_i460_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n460_adj_2331)) /* synthesis lut_function=(A (B+(C (D)+!C !(D)))+!A (B (C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_0_i460_3_lut_4_lut_4_lut.init = 16'hf8cb;
    LUT4 mux_191_Mux_8_i109_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n109_adj_2332)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C+!(D)))+!A (B (C (D)+!C !(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_8_i109_3_lut_4_lut_4_lut.init = 16'hf83e;
    LUT4 i20300_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n22639)) /* synthesis lut_function=(A (B (C+!(D))+!B !((D)+!C))+!A !(B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20300_3_lut_4_lut_4_lut.init = 16'h81f8;
    LUT4 mux_192_Mux_1_i732_3_lut (.A(n716_adj_2333), .B(n491_adj_2334), 
         .C(index_q[4]), .Z(n732_adj_2335)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_1_i732_3_lut.init = 16'hcaca;
    LUT4 i18737_3_lut_3_lut (.A(n26571), .B(index_q[3]), .C(n1001), .Z(n21057)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam i18737_3_lut_3_lut.init = 16'h7474;
    LUT4 mux_192_Mux_4_i668_3_lut_3_lut (.A(n26571), .B(index_q[3]), .C(n29200), 
         .Z(n668_adj_2336)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;
    defparam mux_192_Mux_4_i668_3_lut_3_lut.init = 16'hd1d1;
    L6MUX21 i20163 (.D0(n21370), .D1(n21376), .SD(index_q[6]), .Z(n22502));
    LUT4 mux_191_Mux_0_i604_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n604_adj_2337)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)+!C !(D)))+!A (B (C (D))+!B (C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_0_i604_3_lut_4_lut_4_lut.init = 16'h0e65;
    LUT4 mux_192_Mux_5_i890_3_lut_3_lut (.A(n26571), .B(index_q[3]), .C(n29189), 
         .Z(n890_adj_2338)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam mux_192_Mux_5_i890_3_lut_3_lut.init = 16'h7474;
    L6MUX21 i20164 (.D0(n21379), .D1(n21382), .SD(index_q[6]), .Z(n22503));
    LUT4 mux_192_Mux_0_i460_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n460_adj_2339)) /* synthesis lut_function=(A (B+(C (D)+!C !(D)))+!A (B (C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_0_i460_3_lut_4_lut_4_lut.init = 16'hf8cb;
    PFUMX mux_191_Mux_5_i732 (.BLUT(n11979), .ALUT(n731), .C0(index_i[4]), 
          .Z(n732_adj_2340)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 i20457_3_lut_3_lut (.A(n26571), .B(index_q[3]), .C(n29200), .Z(n22796)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam i20457_3_lut_3_lut.init = 16'h7474;
    LUT4 mux_192_Mux_7_i364_3_lut_3_lut (.A(n26571), .B(index_q[3]), .C(n29187), 
         .Z(n364_adj_2341)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;
    defparam mux_192_Mux_7_i364_3_lut_3_lut.init = 16'hd1d1;
    LUT4 mux_192_Mux_8_i109_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n109)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C+!(D)))+!A (B (C (D)+!C !(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_8_i109_3_lut_4_lut_4_lut.init = 16'hf83e;
    LUT4 i19970_3_lut (.A(n22302), .B(n22303), .C(index_q[7]), .Z(n22309)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19970_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_11_i445_3_lut_4_lut_4_lut_4_lut (.A(index_q[3]), .B(index_q[4]), 
         .C(index_q[5]), .D(n26526), .Z(n445)) /* synthesis lut_function=(!(A (B (C))+!A !(B+(C+(D))))) */ ;
    defparam mux_192_Mux_11_i445_3_lut_4_lut_4_lut_4_lut.init = 16'h7f7e;
    LUT4 i19785_3_lut_4_lut_4_lut (.A(n26523), .B(index_q[5]), .C(index_q[4]), 
         .D(n26384), .Z(n22124)) /* synthesis lut_function=(A (B+(C (D)))+!A (B+((D)+!C))) */ ;
    defparam i19785_3_lut_4_lut_4_lut.init = 16'hfdcd;
    LUT4 i7141_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n157_adj_2342)) /* synthesis lut_function=(!(A (C (D))+!A !(B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i7141_3_lut_4_lut_4_lut.init = 16'h4aaa;
    L6MUX21 i20165 (.D0(n21544), .D1(n21559), .SD(index_q[6]), .Z(n22504));
    PFUMX i20166 (.BLUT(n21562), .ALUT(n892_adj_2343), .C0(index_q[6]), 
          .Z(n22505));
    LUT4 mux_192_Mux_0_i397_3_lut (.A(n29189), .B(n26734), .C(index_q[3]), 
         .Z(n397_adj_2344)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_0_i397_3_lut.init = 16'hcaca;
    LUT4 mux_191_Mux_5_i252_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[4]), .Z(n252_adj_2345)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+(D)))+!A (B (C (D))+!B !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_5_i252_3_lut_4_lut.init = 16'hc993;
    LUT4 mux_192_Mux_9_i62_3_lut_4_lut_else_4_lut (.A(index_q[4]), .B(index_q[2]), 
         .C(index_q[1]), .D(index_q[0]), .Z(n26749)) /* synthesis lut_function=((B+(C (D)))+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_9_i62_3_lut_4_lut_else_4_lut.init = 16'hfddd;
    LUT4 mux_191_Mux_0_i428_3_lut_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n428_adj_2346)) /* synthesis lut_function=(A (B (C+(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B (C))) */ ;
    defparam mux_191_Mux_0_i428_3_lut_3_lut_4_lut_4_lut.init = 16'h8fe1;
    LUT4 mux_191_Mux_1_i716_3_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[1]), .D(index_i[3]), .Z(n716_adj_2347)) /* synthesis lut_function=(!(A (B (D)+!B !(C))+!A !(B (C (D))+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_1_i716_3_lut_4_lut_4_lut.init = 16'h70a9;
    LUT4 mux_191_Mux_11_i445_3_lut_4_lut_4_lut_4_lut (.A(index_i[3]), .B(index_i[4]), 
         .C(index_i[5]), .D(n26519), .Z(n445_adj_2348)) /* synthesis lut_function=(!(A (B (C))+!A !(B+(C+(D))))) */ ;
    defparam mux_191_Mux_11_i445_3_lut_4_lut_4_lut_4_lut.init = 16'h7f7e;
    LUT4 i19217_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21537)) /* synthesis lut_function=(A (C)+!A !(B (C)+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19217_3_lut_4_lut_4_lut.init = 16'hb4b5;
    LUT4 mux_192_Mux_1_i684_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n684_adj_2349)) /* synthesis lut_function=(A (B ((D)+!C)+!B !((D)+!C))+!A !(B (C+(D))+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_1_i684_3_lut_4_lut_4_lut.init = 16'h992d;
    LUT4 i19969_3_lut (.A(n22300), .B(n22301), .C(index_q[7]), .Z(n22308)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19969_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_1_i716_3_lut_4_lut_4_lut (.A(index_q[2]), .B(index_q[0]), 
         .C(index_q[1]), .D(index_q[3]), .Z(n716_adj_2333)) /* synthesis lut_function=(!(A (B (D)+!B !(C))+!A !(B (C (D))+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_1_i716_3_lut_4_lut_4_lut.init = 16'h70a9;
    LUT4 i19250_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21570)) /* synthesis lut_function=(A (C)+!A !(B (C)+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19250_3_lut_4_lut_4_lut.init = 16'hb4b5;
    LUT4 i19974_3_lut (.A(n22310), .B(n22311), .C(index_q[8]), .Z(n22313)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19974_3_lut.init = 16'hcaca;
    LUT4 mux_191_Mux_8_i443_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n443_adj_2350)) /* synthesis lut_function=(A (B (C+!(D))+!B !((D)+!C))+!A !(B (D)+!B ((D)+!C))) */ ;
    defparam mux_191_Mux_8_i443_3_lut_4_lut_4_lut.init = 16'h80fc;
    LUT4 i19027_3_lut_else_4_lut (.A(index_q[4]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n29202)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C+!(D)))+!A !(B ((D)+!C)+!B (C (D)+!C !(D))))) */ ;
    defparam i19027_3_lut_else_4_lut.init = 16'h5685;
    LUT4 i19391_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21711)) /* synthesis lut_function=(!(A ((D)+!C)+!A !(B ((D)+!C)+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19391_3_lut_3_lut_4_lut.init = 16'h55a4;
    LUT4 mux_191_Mux_0_i379_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n379)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !((D)+!C))+!A !(B ((D)+!C)+!B (D))) */ ;
    defparam mux_191_Mux_0_i379_3_lut_4_lut_4_lut.init = 16'h8079;
    LUT4 mux_191_Mux_0_i412_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n412_adj_2351)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(D))+!A (B (D)+!B !(C+!(D)))) */ ;
    defparam mux_191_Mux_0_i412_3_lut_4_lut_4_lut.init = 16'hcd2a;
    LUT4 i19399_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n21719)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B+(C+(D))))) */ ;
    defparam i19399_3_lut_4_lut_4_lut_4_lut.init = 16'h2aab;
    LUT4 mux_191_Mux_7_i699_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n699_adj_2352)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C+!(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_7_i699_3_lut_4_lut_4_lut.init = 16'hf07e;
    LUT4 n518_bdd_3_lut_23586 (.A(n26710), .B(n26699), .C(index_i[3]), 
         .Z(n25271)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n518_bdd_3_lut_23586.init = 16'hcaca;
    L6MUX21 i22716 (.D0(n24290), .D1(n26334), .SD(index_q[6]), .Z(n24291));
    LUT4 mux_191_Mux_0_i890_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n890_adj_2353)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)+!C !(D)))+!A !(B (C)+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_0_i890_3_lut_4_lut_4_lut.init = 16'h70ca;
    LUT4 mux_192_Mux_8_i443_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n443_adj_2354)) /* synthesis lut_function=(A (B (C+!(D))+!B !((D)+!C))+!A !(B (D)+!B ((D)+!C))) */ ;
    defparam mux_192_Mux_8_i443_3_lut_4_lut_4_lut.init = 16'h80fc;
    LUT4 mux_192_Mux_0_i379_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n379_adj_2355)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !((D)+!C))+!A !(B ((D)+!C)+!B (D))) */ ;
    defparam mux_192_Mux_0_i379_3_lut_4_lut_4_lut.init = 16'h8079;
    LUT4 i19469_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21789)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(D))+!A (B (D)+!B ((D)+!C))) */ ;
    defparam i19469_3_lut_4_lut_4_lut.init = 16'hd52b;
    LUT4 mux_192_Mux_0_i684_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n684_adj_2356)) /* synthesis lut_function=(!(A ((D)+!B)+!A !(B (D)+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_0_i684_3_lut_4_lut_4_lut_4_lut.init = 16'h5498;
    LUT4 mux_192_Mux_2_i549_3_lut_4_lut_3_lut_rep_804 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29183)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_2_i549_3_lut_4_lut_3_lut_rep_804.init = 16'h1818;
    LUT4 mux_192_Mux_0_i134_3_lut_4_lut_3_lut_rep_767 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n26727)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_0_i134_3_lut_4_lut_3_lut_rep_767.init = 16'h6969;
    LUT4 i18712_3_lut_4_lut (.A(index_q[0]), .B(n26538), .C(index_q[3]), 
         .D(n29197), .Z(n21032)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A ((D)+!C)) */ ;
    defparam i18712_3_lut_4_lut.init = 16'hfd0d;
    LUT4 n867_bdd_4_lut (.A(n29192), .B(n939_adj_2357), .C(index_q[4]), 
         .D(index_q[3]), .Z(n24360)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D)))) */ ;
    defparam n867_bdd_4_lut.init = 16'hcacc;
    LUT4 n24168_bdd_3_lut_25810 (.A(n24168), .B(n24161), .C(index_q[7]), 
         .Z(n24169)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n24168_bdd_3_lut_25810.init = 16'hcaca;
    LUT4 mux_192_Mux_2_i557_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n557)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C+!(D))+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_2_i557_3_lut_3_lut_4_lut.init = 16'h0f18;
    LUT4 index_q_1__bdd_4_lut (.A(index_q[1]), .B(index_q[0]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n29201)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A !(B ((D)+!C)+!B (D))) */ ;
    defparam index_q_1__bdd_4_lut.init = 16'h8a51;
    LUT4 mux_192_Mux_7_i716_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n716_adj_2358)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C+!(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_7_i716_3_lut_3_lut_4_lut.init = 16'h0f81;
    LUT4 n970_bdd_3_lut_23625 (.A(n29185), .B(n29200), .C(index_q[3]), 
         .Z(n25309)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n970_bdd_3_lut_23625.init = 16'hcaca;
    LUT4 n26528_bdd_4_lut (.A(n26528), .B(index_q[4]), .C(n27995), .D(index_q[5]), 
         .Z(n29161)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C (D))) */ ;
    defparam n26528_bdd_4_lut.init = 16'hf088;
    PFUMX i22714 (.BLUT(n24289), .ALUT(n26372), .C0(index_q[7]), .Z(n24290));
    LUT4 n986_bdd_4_lut_4_lut_4_lut (.A(index_q[0]), .B(n26538), .C(index_q[4]), 
         .D(index_q[3]), .Z(n24358)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (D))+!A (B (C (D)+!C !(D))+!B (D)))) */ ;
    defparam n986_bdd_4_lut_4_lut_4_lut.init = 16'h0c73;
    LUT4 i11509_3_lut_4_lut (.A(index_q[0]), .B(n26538), .C(n26584), .D(index_q[5]), 
         .Z(n318)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (C (D))) */ ;
    defparam i11509_3_lut_4_lut.init = 16'hf800;
    LUT4 mux_191_Mux_2_i731_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n731_adj_2359)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_2_i731_3_lut_4_lut_4_lut.init = 16'h6cc6;
    LUT4 i20578_3_lut (.A(n22910), .B(n27998), .C(index_q[6]), .Z(n22917)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20578_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_2_i269_3_lut_3_lut_3_lut_rep_768 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n26728)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_2_i269_3_lut_3_lut_3_lut_rep_768.init = 16'h3939;
    LUT4 i20579_3_lut (.A(n25312), .B(n22913), .C(index_q[6]), .Z(n22918)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20579_3_lut.init = 16'hcaca;
    LUT4 i19477_3_lut_3_lut_4_lut (.A(index_q[0]), .B(n26538), .C(index_q[3]), 
         .D(n26496), .Z(n21797)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A !(C+(D))) */ ;
    defparam i19477_3_lut_3_lut_4_lut.init = 16'h808f;
    LUT4 i20420_3_lut_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n22759)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C+!(D))+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20420_3_lut_3_lut_4_lut_4_lut.init = 16'h1f81;
    LUT4 i18787_3_lut_3_lut_4_lut (.A(index_q[0]), .B(n26538), .C(n26496), 
         .D(index_q[3]), .Z(n21107)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(C+(D)))) */ ;
    defparam i18787_3_lut_3_lut_4_lut.init = 16'h77f0;
    LUT4 mux_192_Mux_6_i939_3_lut_rep_397_3_lut_4_lut (.A(index_q[0]), .B(n26538), 
         .C(n26526), .D(index_q[3]), .Z(n26357)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(C+(D)))) */ ;
    defparam mux_192_Mux_6_i939_3_lut_rep_397_3_lut_4_lut.init = 16'h77f0;
    LUT4 i21639_3_lut (.A(n491_adj_2283), .B(n506), .C(index_i[4]), .Z(n21324)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21639_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_0_i970_3_lut_rep_806 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29185)) /* synthesis lut_function=(!(A (B (C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_0_i970_3_lut_rep_806.init = 16'h7e7e;
    LUT4 i20161_3_lut (.A(n190), .B(n253), .C(index_q[6]), .Z(n22500)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20161_3_lut.init = 16'hcaca;
    LUT4 i20162_3_lut (.A(n22815), .B(n21367), .C(index_q[6]), .Z(n22501)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20162_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_4_i526_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n526_adj_2360)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A !(B ((D)+!C)+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_4_i526_3_lut_3_lut_4_lut.init = 16'h7e0f;
    LUT4 i11485_3_lut_4_lut (.A(n26349), .B(index_q[7]), .C(index_q[8]), 
         .D(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_2142[14])) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11485_3_lut_4_lut.init = 16'hffe0;
    LUT4 mux_192_Mux_1_i700_3_lut_4_lut (.A(n26646), .B(index_q[3]), .C(index_q[4]), 
         .D(n684_adj_2349), .Z(n700_adj_2361)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_1_i700_3_lut_4_lut.init = 16'hefe0;
    LUT4 n10961_bdd_3_lut_23670_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n25354)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C (D)+!C !(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n10961_bdd_3_lut_23670_3_lut_4_lut.init = 16'h0fc1;
    LUT4 mux_192_Mux_0_i723_3_lut_rep_808 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29187)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_0_i723_3_lut_rep_808.init = 16'h1c1c;
    L6MUX21 i23279 (.D0(n24949), .D1(n24946), .SD(index_i[5]), .Z(n24950));
    LUT4 i18764_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21084)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18764_3_lut_3_lut_4_lut.init = 16'h0f1c;
    PFUMX i23277 (.BLUT(n24948), .ALUT(n24947), .C0(index_i[4]), .Z(n24949));
    LUT4 i19063_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21383)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C (D)))+!A (B (C+(D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19063_4_lut_4_lut_4_lut.init = 16'h301c;
    LUT4 index_i_5__bdd_4_lut_23653 (.A(index_i[2]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[0]), .Z(n25336)) /* synthesis lut_function=(A (B (C+!(D))+!B !(D))+!A !(B (C+!(D))+!B !(D))) */ ;
    defparam index_i_5__bdd_4_lut_23653.init = 16'h95aa;
    LUT4 i19226_3_lut (.A(n26697), .B(n26695), .C(index_i[3]), .Z(n21546)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19226_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_0_i699_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n699_adj_2362)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (D))+!A (B (C+!(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_0_i699_3_lut_3_lut_4_lut.init = 16'h1c33;
    LUT4 mux_192_Mux_8_i124_3_lut_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n124)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C+!(D)))+!A (B (C (D)+!C !(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_8_i124_3_lut_3_lut_4_lut_4_lut.init = 16'h07c1;
    LUT4 i18749_3_lut (.A(n26734), .B(n325), .C(index_q[3]), .Z(n21069)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18749_3_lut.init = 16'hcaca;
    LUT4 i19397_3_lut_4_lut (.A(n26548), .B(index_i[2]), .C(index_i[3]), 
         .D(n26702), .Z(n21717)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19397_3_lut_4_lut.init = 16'hf404;
    LUT4 mux_191_Mux_0_i731_3_lut_4_lut (.A(n26548), .B(index_i[2]), .C(index_i[3]), 
         .D(n26652), .Z(n731_adj_2363)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_0_i731_3_lut_4_lut.init = 16'h4f40;
    LUT4 mux_192_Mux_7_i620_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n620_adj_2364)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B ((D)+!C)+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_7_i620_3_lut_4_lut_4_lut.init = 16'h83c3;
    LUT4 n25338_bdd_3_lut (.A(n25338), .B(n25335), .C(index_i[4]), .Z(n25339)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n25338_bdd_3_lut.init = 16'hcaca;
    LUT4 mux_191_Mux_7_i379_3_lut_3_lut (.A(n26650), .B(index_i[3]), .C(n29194), 
         .Z(n379_adj_2365)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam mux_191_Mux_7_i379_3_lut_3_lut.init = 16'h7474;
    LUT4 mux_191_Mux_8_i542_3_lut_4_lut (.A(n26637), .B(index_i[3]), .C(index_i[4]), 
         .D(n526_adj_2366), .Z(n542_adj_2367)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_8_i542_3_lut_4_lut.init = 16'h6f60;
    LUT4 i18992_3_lut_4_lut (.A(n26637), .B(index_i[3]), .C(index_i[4]), 
         .D(n635_adj_2300), .Z(n21312)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18992_3_lut_4_lut.init = 16'hf606;
    PFUMX i24518 (.BLUT(n26823), .ALUT(n26824), .C0(index_q[8]), .Z(n26825));
    PFUMX i23274 (.BLUT(n24945), .ALUT(n24944), .C0(index_i[4]), .Z(n24946));
    LUT4 mux_192_Mux_8_i93_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n93_adj_2368)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C))+!A (B (C+!(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_8_i93_3_lut_3_lut_4_lut.init = 16'h0f83;
    PFUMX i23251 (.BLUT(n24922), .ALUT(n26741), .C0(index_q[5]), .Z(n24923));
    LUT4 mux_192_Mux_5_i882_3_lut_3_lut_3_lut_rep_810 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29189)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_5_i882_3_lut_3_lut_3_lut_rep_810.init = 16'hc7c7;
    PFUMX i23249 (.BLUT(n26541), .ALUT(n24920), .C0(index_q[2]), .Z(n24921));
    LUT4 mux_191_Mux_1_i700_3_lut_4_lut (.A(n26545), .B(index_i[3]), .C(index_i[4]), 
         .D(n684_adj_2330), .Z(n700_adj_2369)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_1_i700_3_lut_4_lut.init = 16'hefe0;
    LUT4 n970_bdd_3_lut_24383_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n25310)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C))+!A (B (C (D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n970_bdd_3_lut_24383_3_lut_4_lut.init = 16'h0fc7;
    LUT4 i19225_3_lut (.A(n396), .B(n204), .C(index_i[3]), .Z(n21545)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19225_3_lut.init = 16'hcaca;
    LUT4 i19040_3_lut_4_lut (.A(n26644), .B(index_q[3]), .C(index_q[4]), 
         .D(n635_adj_2289), .Z(n21360)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19040_3_lut_4_lut.init = 16'hf606;
    LUT4 i18790_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21110)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+(D)))+!A !(B (D)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18790_3_lut_4_lut_4_lut.init = 16'h99c7;
    LUT4 mux_192_Mux_8_i542_3_lut_4_lut (.A(n26644), .B(index_q[3]), .C(index_q[4]), 
         .D(n526_adj_2370), .Z(n542_adj_2371)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_8_i542_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_192_Mux_0_i188_3_lut (.A(n29183), .B(n931_adj_2372), .C(index_q[3]), 
         .Z(n188)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_0_i188_3_lut.init = 16'hcaca;
    LUT4 i11061_2_lut_rep_811 (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .Z(n29190)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11061_2_lut_rep_811.init = 16'hf8f8;
    LUT4 n26462_bdd_3_lut_25712_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[5]), .Z(n27993)) /* synthesis lut_function=(A (B+(C+(D)))+!A !((D)+!C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n26462_bdd_3_lut_25712_4_lut.init = 16'haaf8;
    LUT4 mux_191_Mux_4_i668_3_lut_3_lut (.A(n26650), .B(index_i[3]), .C(n29180), 
         .Z(n668_adj_2373)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;
    defparam mux_191_Mux_4_i668_3_lut_3_lut.init = 16'hd1d1;
    L6MUX21 i23247 (.D0(n24918), .D1(n24915), .SD(index_q[5]), .Z(n24919));
    LUT4 i19292_3_lut_3_lut (.A(n26650), .B(index_i[3]), .C(n38), .Z(n21612)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam i19292_3_lut_3_lut.init = 16'h7474;
    LUT4 mux_192_Mux_3_i788_rep_813 (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .Z(n29192)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_3_i788_rep_813.init = 16'h7c7c;
    LUT4 i20336_3_lut_3_lut (.A(n26650), .B(index_i[3]), .C(n29180), .Z(n22675)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam i20336_3_lut_3_lut.init = 16'h7474;
    PFUMX i23245 (.BLUT(n24917), .ALUT(n24916), .C0(index_q[4]), .Z(n24918));
    L6MUX21 i20604 (.D0(n22931), .D1(n22932), .SD(index_i[6]), .Z(n22943));
    LUT4 i19367_3_lut_4_lut (.A(index_i[0]), .B(n26637), .C(index_i[3]), 
         .D(n26701), .Z(n21687)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19367_3_lut_4_lut.init = 16'hfb0b;
    LUT4 index_q_7__bdd_4_lut_24624 (.A(index_q[7]), .B(n125), .C(n24286), 
         .D(index_q[5]), .Z(n26334)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(B (C+(D))+!B !((D)+!C)))) */ ;
    defparam index_q_7__bdd_4_lut_24624.init = 16'h66f0;
    LUT4 mux_191_Mux_0_i908_3_lut_4_lut (.A(index_i[0]), .B(n26546), .C(index_i[3]), 
         .D(n26685), .Z(n908_adj_2374)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (C+!(D)))) */ ;
    defparam mux_191_Mux_0_i908_3_lut_4_lut.init = 16'h2f20;
    LUT4 i18731_3_lut (.A(n29171), .B(n26543), .C(index_q[3]), .Z(n21051)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18731_3_lut.init = 16'hcaca;
    LUT4 i18730_3_lut (.A(n29195), .B(n325), .C(index_q[3]), .Z(n21050)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18730_3_lut.init = 16'hcaca;
    LUT4 i21316_3_lut (.A(n21050), .B(n21051), .C(index_q[4]), .Z(n21052)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21316_3_lut.init = 16'hcaca;
    PFUMX i23242 (.BLUT(n24914), .ALUT(n21012), .C0(index_q[4]), .Z(n24915));
    LUT4 mux_191_Mux_7_i123_3_lut_3_lut_rep_815 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29194)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_7_i123_3_lut_3_lut_rep_815.init = 16'hc7c7;
    LUT4 n53_bdd_3_lut_24454_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n25207)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C))+!A (B (C (D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n53_bdd_3_lut_24454_3_lut_4_lut.init = 16'h0fc7;
    LUT4 i19345_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21665)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+(D)))+!A !(B (D)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19345_3_lut_4_lut_4_lut.init = 16'h99c7;
    L6MUX21 i20605 (.D0(n22933), .D1(n22934), .SD(index_i[6]), .Z(n22944));
    L6MUX21 i20606 (.D0(n22935), .D1(n22936), .SD(index_i[6]), .Z(n22945));
    LUT4 i19880_3_lut (.A(n22214), .B(n24362), .C(index_q[7]), .Z(n22219)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19880_3_lut.init = 16'hcaca;
    LUT4 i20617_3_lut (.A(n25265), .B(n22642), .C(index_i[6]), .Z(n22956)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20617_3_lut.init = 16'hcaca;
    LUT4 i21636_3_lut (.A(n26167), .B(n124_adj_2375), .C(index_q[4]), 
         .Z(n22895)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21636_3_lut.init = 16'hcaca;
    PFUMX i20607 (.BLUT(n22937), .ALUT(n22938), .C0(index_i[6]), .Z(n22946));
    L6MUX21 i23240 (.D0(n24912), .D1(n24910), .SD(index_q[5]), .Z(n24913));
    LUT4 n315_bdd_3_lut_23777_4_lut (.A(n26732), .B(index_q[2]), .C(index_q[3]), 
         .D(n29164), .Z(n24909)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n315_bdd_3_lut_23777_4_lut.init = 16'hf606;
    LUT4 mux_192_Mux_3_i890_3_lut_4_lut (.A(n26732), .B(index_q[2]), .C(index_q[3]), 
         .D(n325), .Z(n890)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_3_i890_3_lut_4_lut.init = 16'h6f60;
    LUT4 i19247_3_lut_4_lut (.A(n26732), .B(index_q[2]), .C(index_q[3]), 
         .D(n26727), .Z(n21567)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19247_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_192_Mux_0_i348_3_lut_4_lut (.A(n26732), .B(index_q[2]), .C(index_q[3]), 
         .D(n29181), .Z(n348_adj_2376)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_0_i348_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_192_Mux_6_i269_rep_816 (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .Z(n29195)) /* synthesis lut_function=(A (C)+!A !((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_6_i269_rep_816.init = 16'ha4a4;
    LUT4 i19499_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21819)) /* synthesis lut_function=(!(A ((D)+!C)+!A !(B ((D)+!C)+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19499_3_lut_3_lut_4_lut.init = 16'h55a4;
    LUT4 i19342_3_lut_3_lut_4_lut (.A(index_i[0]), .B(n26546), .C(n26505), 
         .D(index_i[3]), .Z(n21662)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(C+(D)))) */ ;
    defparam i19342_3_lut_3_lut_4_lut.init = 16'h77f0;
    LUT4 mux_192_Mux_0_i123_3_lut_3_lut_rep_817 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29196)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_0_i123_3_lut_3_lut_rep_817.init = 16'h6c6c;
    LUT4 mux_192_Mux_0_i124_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n124_adj_2375)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A !(B (D)+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_0_i124_3_lut_4_lut_4_lut.init = 16'h6c99;
    PFUMX i24471 (.BLUT(n26749), .ALUT(n26750), .C0(index_q[3]), .Z(n62_adj_2377));
    LUT4 i19879_3_lut (.A(n22212), .B(n22213), .C(index_q[7]), .Z(n22218)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19879_3_lut.init = 16'hcaca;
    LUT4 i18728_3_lut (.A(n29162), .B(n29176), .C(index_q[3]), .Z(n21048)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18728_3_lut.init = 16'hcaca;
    LUT4 i22278_3_lut (.A(n22218), .B(n22219), .C(index_q[8]), .Z(n22221)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22278_3_lut.init = 16'hcaca;
    PFUMX i23238 (.BLUT(n24911), .ALUT(n285), .C0(index_q[4]), .Z(n24912));
    LUT4 i11498_4_lut (.A(n15006), .B(index_q[8]), .C(n765), .D(index_q[7]), 
         .Z(n1022)) /* synthesis lut_function=(A (B+(C (D)))+!A (B+(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11498_4_lut.init = 16'hfcdd;
    LUT4 i21318_3_lut (.A(n21047), .B(n21048), .C(index_q[4]), .Z(n21049)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21318_3_lut.init = 16'hcaca;
    PFUMX i23236 (.BLUT(n24909), .ALUT(n24908), .C0(index_q[4]), .Z(n24910));
    LUT4 i21322_3_lut (.A(n21044), .B(n21045), .C(index_q[4]), .Z(n21046)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21322_3_lut.init = 16'hcaca;
    LUT4 mux_191_Mux_7_i890_3_lut_4_lut (.A(index_i[0]), .B(n26546), .C(index_i[3]), 
         .D(n26486), .Z(n890_adj_2378)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A !(C+(D))) */ ;
    defparam mux_191_Mux_7_i890_3_lut_4_lut.init = 16'h808f;
    LUT4 i19375_3_lut_3_lut_4_lut (.A(index_i[0]), .B(n26546), .C(index_i[3]), 
         .D(n26505), .Z(n21695)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A !(C+(D))) */ ;
    defparam i19375_3_lut_3_lut_4_lut.init = 16'h808f;
    LUT4 mux_191_Mux_0_i781_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n781_adj_2379)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A (B (C)+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_0_i781_4_lut_4_lut_4_lut.init = 16'h0cb4;
    LUT4 mux_191_Mux_8_i653_3_lut_rep_399_3_lut_4_lut (.A(index_i[0]), .B(n26546), 
         .C(n26519), .D(index_i[3]), .Z(n26359)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(C+(D)))) */ ;
    defparam mux_191_Mux_8_i653_3_lut_rep_399_3_lut_4_lut.init = 16'h77f0;
    LUT4 i11440_3_lut_4_lut (.A(index_i[0]), .B(n26546), .C(n26595), .D(index_i[5]), 
         .Z(n318_adj_2380)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (C (D))) */ ;
    defparam i11440_3_lut_4_lut.init = 16'hf800;
    LUT4 i11425_4_lut (.A(n14982), .B(index_i[8]), .C(n765_adj_2381), 
         .D(index_i[7]), .Z(n1022_adj_2382)) /* synthesis lut_function=(A (B+(C (D)))+!A (B+(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11425_4_lut.init = 16'hfcdd;
    LUT4 i19997_3_lut (.A(n22334), .B(n22335), .C(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2127[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19997_3_lut.init = 16'hcaca;
    LUT4 i6419_2_lut (.A(phase_q[0]), .B(phase_i[10]), .Z(index_i_9__N_2107[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i6419_2_lut.init = 16'h6666;
    LUT4 i22297_2_lut (.A(phase_q[0]), .B(phase_i[10]), .Z(index_q_9__N_2117[0])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i22297_2_lut.init = 16'h9999;
    LUT4 i20614_3_lut (.A(n25935), .B(n22952), .C(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2127[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20614_3_lut.init = 16'hcaca;
    LUT4 n699_bdd_4_lut_4_lut_4_lut (.A(index_i[0]), .B(n26546), .C(index_i[4]), 
         .D(index_i[3]), .Z(n24307)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (D))+!A (B (C (D)+!C !(D))+!B (D)))) */ ;
    defparam n699_bdd_4_lut_4_lut_4_lut.init = 16'h0c73;
    LUT4 i20613_3_lut (.A(n22949), .B(n22950), .C(index_i[8]), .Z(n22952)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20613_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_0_i525_3_lut_3_lut_rep_818 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29197)) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_0_i525_3_lut_3_lut_rep_818.init = 16'h6a6a;
    LUT4 mux_192_Mux_14_i511_4_lut_4_lut (.A(n26349), .B(index_q[7]), .C(index_q[8]), 
         .D(n254_adj_2383), .Z(n511)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (B (C+!(D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_14_i511_4_lut_4_lut.init = 16'h1c10;
    LUT4 i1_2_lut_rep_536_3_lut (.A(index_q[2]), .B(index_q[0]), .C(index_q[1]), 
         .Z(n26496)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_2_lut_rep_536_3_lut.init = 16'hfefe;
    LUT4 quarter_wave_sample_register_i_15__I_0_3_lut (.A(\quarter_wave_sample_register_q[15] ), 
         .B(o_val_pipeline_i_0__15__N_2158[15]), .C(phase_negation_i[1]), 
         .Z(o_val_pipeline_i_0__15__N_2157)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[14] 77[8])
    defparam quarter_wave_sample_register_i_15__I_0_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_2_i491_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n491_adj_2384)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A !(B (C)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_2_i491_3_lut_4_lut_4_lut.init = 16'h6a5a;
    LUT4 mux_192_Mux_5_i459_3_lut_4_lut_3_lut_rep_788 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29167)) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_5_i459_3_lut_4_lut_3_lut_rep_788.init = 16'h6b6b;
    LUT4 quarter_wave_sample_register_i_14__I_0_3_lut (.A(quarter_wave_sample_register_i[14]), 
         .B(o_val_pipeline_i_0__15__N_2158[14]), .C(phase_negation_i[1]), 
         .Z(o_val_pipeline_i_0__15__N_2159)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[14] 77[8])
    defparam quarter_wave_sample_register_i_14__I_0_3_lut.init = 16'hcaca;
    L6MUX21 i20618 (.D0(n21307), .D1(n21310), .SD(index_i[6]), .Z(n22957));
    LUT4 quarter_wave_sample_register_i_13__I_0_3_lut (.A(quarter_wave_sample_register_i[13]), 
         .B(o_val_pipeline_i_0__15__N_2158[13]), .C(phase_negation_i[1]), 
         .Z(o_val_pipeline_i_0__15__N_2161)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[14] 77[8])
    defparam quarter_wave_sample_register_i_13__I_0_3_lut.init = 16'hcaca;
    LUT4 quarter_wave_sample_register_i_12__I_0_3_lut (.A(quarter_wave_sample_register_i[12]), 
         .B(o_val_pipeline_i_0__15__N_2158[12]), .C(phase_negation_i[1]), 
         .Z(o_val_pipeline_i_0__15__N_2163)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[14] 77[8])
    defparam quarter_wave_sample_register_i_12__I_0_3_lut.init = 16'hcaca;
    LUT4 i20197_3_lut_3_lut_4_lut (.A(n26438), .B(index_i[3]), .C(n316_adj_2385), 
         .D(index_i[4]), .Z(n22536)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20197_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 mux_192_Mux_0_i716_3_lut (.A(n26712), .B(n29175), .C(index_q[3]), 
         .Z(n716_adj_2386)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_0_i716_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_0_i963_3_lut_3_lut_rep_819 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29198)) /* synthesis lut_function=(!(A (B)+!A (B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_0_i963_3_lut_3_lut_rep_819.init = 16'h3636;
    LUT4 i21694_3_lut (.A(n109_adj_2332), .B(n124_adj_2387), .C(index_i[4]), 
         .Z(n21297)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21694_3_lut.init = 16'hcaca;
    L6MUX21 i20202 (.D0(n22539), .D1(n22540), .SD(index_i[6]), .Z(n382));
    L6MUX21 i20619 (.D0(n574_adj_2388), .D1(n21313), .SD(index_i[6]), 
            .Z(n22958));
    LUT4 quarter_wave_sample_register_i_11__I_0_3_lut (.A(quarter_wave_sample_register_i[11]), 
         .B(o_val_pipeline_i_0__15__N_2158[11]), .C(phase_negation_i[1]), 
         .Z(o_val_pipeline_i_0__15__N_2165)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[14] 77[8])
    defparam quarter_wave_sample_register_i_11__I_0_3_lut.init = 16'hcaca;
    LUT4 quarter_wave_sample_register_i_10__I_0_3_lut (.A(quarter_wave_sample_register_i[10]), 
         .B(o_val_pipeline_i_0__15__N_2158[10]), .C(phase_negation_i[1]), 
         .Z(o_val_pipeline_i_0__15__N_2167)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[14] 77[8])
    defparam quarter_wave_sample_register_i_10__I_0_3_lut.init = 16'hcaca;
    LUT4 quarter_wave_sample_register_i_9__I_0_3_lut (.A(quarter_wave_sample_register_i[9]), 
         .B(o_val_pipeline_i_0__15__N_2158[9]), .C(phase_negation_i[1]), 
         .Z(o_val_pipeline_i_0__15__N_2169)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[14] 77[8])
    defparam quarter_wave_sample_register_i_9__I_0_3_lut.init = 16'hcaca;
    LUT4 n53_bdd_3_lut_23377_4_lut (.A(n26542), .B(index_q[2]), .C(n29162), 
         .D(index_q[3]), .Z(n25067)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n53_bdd_3_lut_23377_4_lut.init = 16'hf066;
    LUT4 n308_bdd_3_lut_23244_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n24916)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A !(B (C+(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n308_bdd_3_lut_23244_4_lut_4_lut.init = 16'h9936;
    LUT4 mux_191_Mux_5_i491_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n491_adj_2389)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A !(B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_5_i491_3_lut_4_lut_4_lut.init = 16'ha54a;
    LUT4 quarter_wave_sample_register_i_8__I_0_3_lut (.A(quarter_wave_sample_register_i[8]), 
         .B(o_val_pipeline_i_0__15__N_2158[8]), .C(phase_negation_i[1]), 
         .Z(o_val_pipeline_i_0__15__N_2171)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[14] 77[8])
    defparam quarter_wave_sample_register_i_8__I_0_3_lut.init = 16'hcaca;
    LUT4 quarter_wave_sample_register_i_7__I_0_3_lut (.A(quarter_wave_sample_register_i[7]), 
         .B(o_val_pipeline_i_0__15__N_2158[7]), .C(phase_negation_i[1]), 
         .Z(o_val_pipeline_i_0__15__N_2173)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[14] 77[8])
    defparam quarter_wave_sample_register_i_7__I_0_3_lut.init = 16'hcaca;
    L6MUX21 i20620 (.D0(n21316), .D1(n764_adj_2390), .SD(index_i[6]), 
            .Z(n22959));
    LUT4 mux_192_Mux_3_i668_3_lut_4_lut (.A(n26542), .B(index_q[2]), .C(index_q[3]), 
         .D(n29171), .Z(n668)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_3_i668_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_192_Mux_4_i763_3_lut_4_lut (.A(n26542), .B(index_q[2]), .C(index_q[4]), 
         .D(n747_adj_2391), .Z(n763_adj_2392)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_4_i763_3_lut_4_lut.init = 16'h6f60;
    LUT4 n28282_bdd_3_lut_4_lut (.A(index_i[0]), .B(index_i[2]), .C(index_i[5]), 
         .D(n28282), .Z(n28283)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;
    defparam n28282_bdd_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_192_Mux_0_i475_3_lut_4_lut (.A(n26550), .B(index_q[1]), .C(index_q[3]), 
         .D(n29190), .Z(n475_adj_2393)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_0_i475_3_lut_4_lut.init = 16'h4f40;
    LUT4 mux_192_Mux_3_i491_3_lut_4_lut (.A(n26550), .B(index_q[1]), .C(index_q[3]), 
         .D(n26721), .Z(n491)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_3_i491_3_lut_4_lut.init = 16'h4f40;
    L6MUX21 i20209 (.D0(n22546), .D1(n22547), .SD(index_i[6]), .Z(n509));
    LUT4 mux_192_Mux_0_i954_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n954_adj_2394)) /* synthesis lut_function=(A (D)+!A !(B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_0_i954_3_lut_4_lut_4_lut.init = 16'haf40;
    PFUMX i20634 (.BLUT(n22969), .ALUT(n22970), .C0(index_i[6]), .Z(n22973));
    LUT4 mux_192_Mux_5_i460_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n460_adj_2395)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A !(B (C)+!B !(C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_5_i460_3_lut_4_lut_4_lut.init = 16'h6b5a;
    LUT4 i12092_3_lut_rep_821 (.A(index_q[2]), .B(index_q[1]), .C(index_q[0]), 
         .Z(n29200)) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12092_3_lut_rep_821.init = 16'hc4c4;
    PFUMX i20635 (.BLUT(n22971), .ALUT(n22972), .C0(index_i[6]), .Z(n22974));
    LUT4 i18767_3_lut_4_lut_4_lut (.A(index_q[2]), .B(index_q[1]), .C(index_q[0]), 
         .D(index_q[3]), .Z(n21087)) /* synthesis lut_function=(A (B (C)+!B !(C+!(D)))+!A (B (C+!(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18767_3_lut_4_lut_4_lut.init = 16'hc3c4;
    LUT4 n627_bdd_3_lut_23785 (.A(n29164), .B(n29198), .C(index_q[3]), 
         .Z(n25450)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n627_bdd_3_lut_23785.init = 16'hcaca;
    LUT4 i7426_2_lut (.A(index_i[4]), .B(index_i[5]), .Z(n9807)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i7426_2_lut.init = 16'h8888;
    LUT4 mux_191_Mux_5_i828_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[4]), .D(n26601), .Z(n828_adj_2396)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_5_i828_4_lut_4_lut.init = 16'hc66c;
    LUT4 i9404_3_lut_4_lut (.A(n26711), .B(index_q[2]), .C(n26622), .D(n26725), 
         .Z(n444_adj_2397)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9404_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_192_Mux_6_i251_3_lut_4_lut (.A(n26711), .B(index_q[2]), .C(index_q[3]), 
         .D(n26725), .Z(n251_adj_2398)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_6_i251_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_192_Mux_4_i747_3_lut_4_lut (.A(n26711), .B(index_q[2]), .C(index_q[3]), 
         .D(n26734), .Z(n747_adj_2391)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_4_i747_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_191_Mux_5_i475_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n475_adj_2399)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_5_i475_3_lut_4_lut_4_lut.init = 16'hd4a5;
    LUT4 n378_bdd_3_lut_23791 (.A(n26543), .B(n29200), .C(index_q[3]), 
         .Z(n25465)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n378_bdd_3_lut_23791.init = 16'hcaca;
    LUT4 mux_192_Mux_6_i285_3_lut_4_lut (.A(n26735), .B(index_q[2]), .C(index_q[3]), 
         .D(n26727), .Z(n285)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_6_i285_3_lut_4_lut.init = 16'hf606;
    CCU2D add_371_15 (.A0(quarter_wave_sample_register_i[14]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(\quarter_wave_sample_register_q[15] ), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17352), .S0(o_val_pipeline_i_0__15__N_2158[14]), 
          .S1(o_val_pipeline_i_0__15__N_2158[15]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam add_371_15.INIT0 = 16'hf555;
    defparam add_371_15.INIT1 = 16'hf555;
    defparam add_371_15.INJECT1_0 = "NO";
    defparam add_371_15.INJECT1_1 = "NO";
    LUT4 i19448_3_lut_4_lut (.A(n26735), .B(index_q[2]), .C(index_q[3]), 
         .D(n26724), .Z(n21768)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19448_3_lut_4_lut.init = 16'hf606;
    LUT4 i18710_3_lut_4_lut (.A(n26735), .B(index_q[2]), .C(index_q[3]), 
         .D(n26734), .Z(n21030)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18710_3_lut_4_lut.init = 16'h6f60;
    L6MUX21 i20223 (.D0(n22560), .D1(n22561), .SD(index_q[6]), .Z(n382_adj_2272));
    LUT4 mux_192_Mux_3_i460_3_lut_4_lut (.A(n26735), .B(index_q[2]), .C(index_q[3]), 
         .D(n29197), .Z(n460)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_3_i460_3_lut_4_lut.init = 16'h6f60;
    LUT4 n627_bdd_3_lut_24259 (.A(n29164), .B(n931), .C(index_q[3]), .Z(n25467)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n627_bdd_3_lut_24259.init = 16'hacac;
    LUT4 i7589_2_lut (.A(index_q[4]), .B(index_q[5]), .Z(n9970)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i7589_2_lut.init = 16'h8888;
    LUT4 mux_191_Mux_3_i668_3_lut_4_lut (.A(n26597), .B(index_i[2]), .C(index_i[3]), 
         .D(n26697), .Z(n668_adj_2400)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_3_i668_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_191_Mux_10_i317_3_lut_3_lut_4_lut (.A(n26438), .B(index_i[3]), 
         .C(n26470), .D(index_i[4]), .Z(n317)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_10_i317_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 n53_bdd_3_lut_23273_4_lut (.A(n26597), .B(index_i[2]), .C(n26701), 
         .D(index_i[3]), .Z(n24944)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n53_bdd_3_lut_23273_4_lut.init = 16'hf066;
    LUT4 mux_191_Mux_4_i763_3_lut_4_lut (.A(n26597), .B(index_i[2]), .C(index_i[4]), 
         .D(n747_adj_2401), .Z(n763_adj_2402)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_4_i763_3_lut_4_lut.init = 16'h6f60;
    L6MUX21 i20230 (.D0(n22567), .D1(n22568), .SD(index_q[6]), .Z(n509_adj_2273));
    LUT4 i18856_3_lut (.A(n24291), .B(n21214), .C(index_q[8]), .Z(n21176)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18856_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut (.A(index_q[6]), .B(index_q[7]), .Z(n19545)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_2_lut.init = 16'heeee;
    LUT4 mux_192_Mux_4_i262_3_lut_3_lut_rep_791 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29170)) /* synthesis lut_function=(A (B+(C))+!A !(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_4_i262_3_lut_3_lut_rep_791.init = 16'ha9a9;
    LUT4 mux_192_Mux_3_i397_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n397)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !(B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_3_i397_3_lut_4_lut_4_lut.init = 16'ha95a;
    LUT4 i20174_3_lut (.A(n22511), .B(n22512), .C(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_2142[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20174_3_lut.init = 16'hcaca;
    LUT4 i19800_3_lut (.A(n25983), .B(n22138), .C(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_2142[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19800_3_lut.init = 16'hcaca;
    LUT4 i19799_3_lut (.A(n22135), .B(n22136), .C(index_q[8]), .Z(n22138)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19799_3_lut.init = 16'hcaca;
    LUT4 i18850_3_lut (.A(n24250), .B(n21205), .C(index_i[8]), .Z(n21170)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18850_3_lut.init = 16'hcaca;
    LUT4 i22299_2_lut (.A(phase_i[9]), .B(phase_i[10]), .Z(index_q_9__N_2117[9])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i22299_2_lut.init = 16'h9999;
    LUT4 i22301_2_lut (.A(phase_i[8]), .B(phase_i[10]), .Z(index_q_9__N_2117[8])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i22301_2_lut.init = 16'h9999;
    LUT4 n21528_bdd_3_lut (.A(n26691), .B(n26606), .C(index_i[3]), .Z(n25483)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n21528_bdd_3_lut.init = 16'hcaca;
    L6MUX21 i20615 (.D0(n21295), .D1(n21298), .SD(index_i[6]), .Z(n22954));
    LUT4 i22303_2_lut (.A(phase_i[7]), .B(phase_i[10]), .Z(index_q_9__N_2117[7])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i22303_2_lut.init = 16'h9999;
    LUT4 i22305_2_lut (.A(phase_i[6]), .B(phase_i[10]), .Z(index_q_9__N_2117[6])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i22305_2_lut.init = 16'h9999;
    LUT4 i22307_2_lut (.A(phase_i[5]), .B(phase_i[10]), .Z(index_q_9__N_2117[5])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i22307_2_lut.init = 16'h9999;
    LUT4 i22309_2_lut (.A(phase_i[4]), .B(phase_i[10]), .Z(index_q_9__N_2117[4])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i22309_2_lut.init = 16'h9999;
    LUT4 i22311_2_lut (.A(phase_i[3]), .B(phase_i[10]), .Z(index_q_9__N_2117[3])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i22311_2_lut.init = 16'h9999;
    LUT4 i22313_2_lut (.A(phase_i[2]), .B(phase_i[10]), .Z(index_q_9__N_2117[2])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i22313_2_lut.init = 16'h9999;
    LUT4 i22315_2_lut (.A(phase_i[1]), .B(phase_i[10]), .Z(index_q_9__N_2117[1])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i22315_2_lut.init = 16'h9999;
    LUT4 i6438_2_lut (.A(phase_i[9]), .B(phase_i[10]), .Z(index_i_9__N_2107[9])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i6438_2_lut.init = 16'h6666;
    LUT4 i6439_2_lut (.A(phase_i[8]), .B(phase_i[10]), .Z(index_i_9__N_2107[8])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i6439_2_lut.init = 16'h6666;
    LUT4 i6440_2_lut (.A(phase_i[7]), .B(phase_i[10]), .Z(index_i_9__N_2107[7])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i6440_2_lut.init = 16'h6666;
    LUT4 i6441_2_lut (.A(phase_i[6]), .B(phase_i[10]), .Z(index_i_9__N_2107[6])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i6441_2_lut.init = 16'h6666;
    PFUMX i20282 (.BLUT(n22605), .ALUT(n22606), .C0(index_q[6]), .Z(n22621));
    LUT4 i6442_2_lut (.A(phase_i[5]), .B(phase_i[10]), .Z(index_i_9__N_2107[5])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i6442_2_lut.init = 16'h6666;
    LUT4 i6443_2_lut (.A(phase_i[4]), .B(phase_i[10]), .Z(index_i_9__N_2107[4])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i6443_2_lut.init = 16'h6666;
    LUT4 i6444_2_lut (.A(phase_i[3]), .B(phase_i[10]), .Z(index_i_9__N_2107[3])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i6444_2_lut.init = 16'h6666;
    L6MUX21 i20283 (.D0(n22607), .D1(n22608), .SD(index_q[6]), .Z(n22622));
    CCU2D add_371_13 (.A0(quarter_wave_sample_register_i[12]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[13]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17351), .COUT(n17352), 
          .S0(o_val_pipeline_i_0__15__N_2158[12]), .S1(o_val_pipeline_i_0__15__N_2158[13]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam add_371_13.INIT0 = 16'hf555;
    defparam add_371_13.INIT1 = 16'hf555;
    defparam add_371_13.INJECT1_0 = "NO";
    defparam add_371_13.INJECT1_1 = "NO";
    LUT4 i6445_2_lut (.A(phase_i[2]), .B(phase_i[10]), .Z(index_i_9__N_2107[2])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i6445_2_lut.init = 16'h6666;
    L6MUX21 i20284 (.D0(n22609), .D1(n22610), .SD(index_q[6]), .Z(n22623));
    LUT4 i6446_2_lut (.A(phase_i[1]), .B(phase_i[10]), .Z(index_i_9__N_2107[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i6446_2_lut.init = 16'h6666;
    LUT4 mux_412_i9_3_lut (.A(\quarter_wave_sample_register_q[15] ), .B(o_val_pipeline_q_0__15__N_2190[15]), 
         .C(phase_negation_q[1]), .Z(n1703[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(80[29:60])
    defparam mux_412_i9_3_lut.init = 16'hcaca;
    L6MUX21 i20285 (.D0(n22611), .D1(n22612), .SD(index_q[6]), .Z(n22624));
    L6MUX21 i20286 (.D0(n22613), .D1(n22614), .SD(index_q[6]), .Z(n22625));
    LUT4 mux_412_i8_3_lut (.A(quarter_wave_sample_register_q[14]), .B(o_val_pipeline_q_0__15__N_2190[14]), 
         .C(phase_negation_q[1]), .Z(n1703[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(80[29:60])
    defparam mux_412_i8_3_lut.init = 16'hcaca;
    LUT4 mux_412_i7_3_lut (.A(quarter_wave_sample_register_q[13]), .B(o_val_pipeline_q_0__15__N_2190[13]), 
         .C(phase_negation_q[1]), .Z(n1703[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(80[29:60])
    defparam mux_412_i7_3_lut.init = 16'hcaca;
    LUT4 mux_412_i6_3_lut (.A(quarter_wave_sample_register_q[12]), .B(o_val_pipeline_q_0__15__N_2190[12]), 
         .C(phase_negation_q[1]), .Z(n1703[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(80[29:60])
    defparam mux_412_i6_3_lut.init = 16'hcaca;
    L6MUX21 i20287 (.D0(n22615), .D1(n22616), .SD(index_q[6]), .Z(n22626));
    LUT4 mux_412_i5_3_lut (.A(quarter_wave_sample_register_q[11]), .B(o_val_pipeline_q_0__15__N_2190[11]), 
         .C(phase_negation_q[1]), .Z(n1703[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(80[29:60])
    defparam mux_412_i5_3_lut.init = 16'hcaca;
    LUT4 mux_412_i4_3_lut (.A(quarter_wave_sample_register_q[10]), .B(o_val_pipeline_q_0__15__N_2190[10]), 
         .C(phase_negation_q[1]), .Z(n1703[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(80[29:60])
    defparam mux_412_i4_3_lut.init = 16'hcaca;
    PFUMX i19215 (.BLUT(n21533), .ALUT(n21534), .C0(index_i[4]), .Z(n21535));
    LUT4 mux_412_i3_3_lut (.A(quarter_wave_sample_register_q[9]), .B(o_val_pipeline_q_0__15__N_2190[9]), 
         .C(phase_negation_q[1]), .Z(n1703[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(80[29:60])
    defparam mux_412_i3_3_lut.init = 16'hcaca;
    LUT4 mux_412_i2_3_lut (.A(quarter_wave_sample_register_q[8]), .B(o_val_pipeline_q_0__15__N_2190[8]), 
         .C(phase_negation_q[1]), .Z(n1703[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(80[29:60])
    defparam mux_412_i2_3_lut.init = 16'hcaca;
    LUT4 mux_412_i1_3_lut (.A(quarter_wave_sample_register_q[7]), .B(o_val_pipeline_q_0__15__N_2190[7]), 
         .C(phase_negation_q[1]), .Z(n1703[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(80[29:60])
    defparam mux_412_i1_3_lut.init = 16'hcaca;
    CCU2D add_371_11 (.A0(quarter_wave_sample_register_i[10]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[11]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17350), .COUT(n17351), 
          .S0(o_val_pipeline_i_0__15__N_2158[10]), .S1(o_val_pipeline_i_0__15__N_2158[11]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam add_371_11.INIT0 = 16'hf555;
    defparam add_371_11.INIT1 = 16'hf555;
    defparam add_371_11.INJECT1_0 = "NO";
    defparam add_371_11.INJECT1_1 = "NO";
    LUT4 mux_192_Mux_8_i15_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n15_adj_2403)) /* synthesis lut_function=(A (B (C)+!B !(C (D)+!C !(D)))+!A !(B ((D)+!C)+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_8_i15_3_lut_4_lut_4_lut.init = 16'h83e0;
    LUT4 i1_4_lut (.A(index_i[7]), .B(n26354), .C(index_i[6]), .D(index_i[8]), 
         .Z(n20039)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i1_4_lut.init = 16'hfffe;
    LUT4 mux_192_Mux_6_i340_3_lut_4_lut_3_lut_rep_792 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29171)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_6_i340_3_lut_4_lut_3_lut_rep_792.init = 16'h9292;
    LUT4 mux_191_Mux_0_i397_3_lut (.A(n29194), .B(n26706), .C(index_i[3]), 
         .Z(n397_adj_2404)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_0_i397_3_lut.init = 16'hcaca;
    LUT4 i18784_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21104)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C))+!A !(B ((D)+!C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18784_3_lut_4_lut_4_lut.init = 16'h925a;
    LUT4 i11424_3_lut_4_lut (.A(n26438), .B(index_i[3]), .C(n9807), .D(index_i[6]), 
         .Z(n765_adj_2381)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11424_3_lut_4_lut.init = 16'hffe0;
    LUT4 n699_bdd_3_lut_24250_4_lut (.A(n26438), .B(index_i[3]), .C(index_i[4]), 
         .D(n93_adj_2405), .Z(n24441)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n699_bdd_3_lut_24250_4_lut.init = 16'hfe0e;
    LUT4 mux_191_Mux_0_i475_3_lut_4_lut (.A(n26561), .B(index_i[1]), .C(index_i[3]), 
         .D(n26486), .Z(n475_adj_2406)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_0_i475_3_lut_4_lut.init = 16'h4f40;
    LUT4 mux_191_Mux_3_i491_3_lut_4_lut (.A(n26561), .B(index_i[1]), .C(index_i[3]), 
         .D(n29178), .Z(n491_adj_2297)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_3_i491_3_lut_4_lut.init = 16'h4f40;
    LUT4 i18715_3_lut (.A(n26543), .B(n26737), .C(index_q[3]), .Z(n21035)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18715_3_lut.init = 16'hcaca;
    LUT4 i19296_then_4_lut (.A(index_i[2]), .B(index_i[1]), .C(index_i[4]), 
         .D(index_i[3]), .Z(n26794)) /* synthesis lut_function=(A (B (C+(D))+!B !(C))+!A !(B (C+(D))+!B !(C+!(D)))) */ ;
    defparam i19296_then_4_lut.init = 16'h9a97;
    LUT4 i19007_3_lut_4_lut_4_lut_4_lut (.A(n26647), .B(index_i[2]), .C(index_i[3]), 
         .D(index_i[4]), .Z(n21327)) /* synthesis lut_function=(A (B)+!A (B (C (D))+!B !(C (D)))) */ ;
    defparam i19007_3_lut_4_lut_4_lut_4_lut.init = 16'hc999;
    LUT4 mux_191_Mux_2_i684_3_lut_4_lut (.A(n26647), .B(index_i[2]), .C(index_i[3]), 
         .D(n26604), .Z(n684_adj_2407)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;
    defparam mux_191_Mux_2_i684_3_lut_4_lut.init = 16'h6f60;
    LUT4 i19235_3_lut_4_lut (.A(n26647), .B(index_i[2]), .C(index_i[3]), 
         .D(n29174), .Z(n21555)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;
    defparam i19235_3_lut_4_lut.init = 16'h6f60;
    LUT4 n476_bdd_3_lut_22925 (.A(n476_adj_2408), .B(n24490), .C(index_i[5]), 
         .Z(n24491)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n476_bdd_3_lut_22925.init = 16'hcaca;
    LUT4 mux_191_Mux_0_i188_3_lut (.A(n26648), .B(n931_adj_2409), .C(index_i[3]), 
         .Z(n188_adj_2410)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_0_i188_3_lut.init = 16'hcaca;
    LUT4 i18995_3_lut_3_lut_4_lut (.A(n26438), .B(index_i[3]), .C(n93_adj_2405), 
         .D(index_i[4]), .Z(n21315)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18995_3_lut_3_lut_4_lut.init = 16'h11f0;
    LUT4 i11763_2_lut_rep_793 (.A(index_q[1]), .B(index_q[2]), .C(index_q[0]), 
         .Z(n29172)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11763_2_lut_rep_793.init = 16'h7070;
    LUT4 mux_191_Mux_7_i475_3_lut_4_lut (.A(n26647), .B(index_i[2]), .C(index_i[3]), 
         .D(n29194), .Z(n475_adj_2411)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+(D)))) */ ;
    defparam mux_191_Mux_7_i475_3_lut_4_lut.init = 16'h9f90;
    PFUMX i20301 (.BLUT(n22636), .ALUT(n22637), .C0(index_i[4]), .Z(n22640));
    LUT4 i20295_3_lut (.A(n22631), .B(n22632), .C(index_q[8]), .Z(n22634)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20295_3_lut.init = 16'hcaca;
    LUT4 i20294_3_lut (.A(n22629), .B(n22630), .C(index_q[8]), .Z(n22633)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20294_3_lut.init = 16'hcaca;
    LUT4 mux_191_Mux_7_i653_3_lut_4_lut (.A(n26647), .B(index_i[2]), .C(index_i[3]), 
         .D(n70_adj_2255), .Z(n653_adj_2412)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam mux_191_Mux_7_i653_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_191_Mux_7_i891_3_lut_4_lut (.A(n26438), .B(index_i[3]), .C(index_i[4]), 
         .D(n890_adj_2378), .Z(n891_adj_2413)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_7_i891_3_lut_4_lut.init = 16'hfe0e;
    LUT4 i1_2_lut_adj_74 (.A(o_phase[11]), .B(o_phase[10]), .Z(phase_q_11__N_2233[11])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i1_2_lut_adj_74.init = 16'h9999;
    LUT4 i19009_4_lut_4_lut_4_lut (.A(n26647), .B(index_i[2]), .C(index_i[4]), 
         .D(index_i[3]), .Z(n21329)) /* synthesis lut_function=(A (B)+!A !(B (C+(D))+!B !(C+(D)))) */ ;
    defparam i19009_4_lut_4_lut_4_lut.init = 16'h999c;
    LUT4 i21730_3_lut (.A(n26845), .B(n124_adj_2414), .C(index_i[4]), 
         .Z(n22833)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21730_3_lut.init = 16'hcaca;
    PFUMX i20302 (.BLUT(n22638), .ALUT(n22639), .C0(index_i[4]), .Z(n22641));
    LUT4 i22263_3_lut (.A(n22962), .B(n22963), .C(index_i[8]), .Z(n22966)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22263_3_lut.init = 16'hcaca;
    L6MUX21 i19790 (.D0(n22117), .D1(n22118), .SD(index_q[6]), .Z(n22129));
    L6MUX21 i19791 (.D0(n22119), .D1(n22120), .SD(index_q[6]), .Z(n22130));
    LUT4 mux_191_Mux_9_i700_3_lut_4_lut (.A(n26438), .B(index_i[3]), .C(index_i[4]), 
         .D(n26485), .Z(n700_adj_2415)) /* synthesis lut_function=(!(A (C+!(D))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_9_i700_3_lut_4_lut.init = 16'h1f10;
    PFUMX i20707 (.BLUT(n557_adj_2416), .ALUT(n572_adj_2417), .C0(index_q[4]), 
          .Z(n23046));
    LUT4 mux_191_Mux_4_i158_3_lut (.A(n142_adj_2418), .B(n157_adj_2419), 
         .C(index_i[4]), .Z(n158)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_4_i158_3_lut.init = 16'hcaca;
    L6MUX21 i19792 (.D0(n22121), .D1(n22122), .SD(index_q[6]), .Z(n22131));
    CCU2D add_371_9 (.A0(quarter_wave_sample_register_i[8]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[9]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17349), .COUT(n17350), 
          .S0(o_val_pipeline_i_0__15__N_2158[8]), .S1(o_val_pipeline_i_0__15__N_2158[9]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam add_371_9.INIT0 = 16'hf555;
    defparam add_371_9.INIT1 = 16'hf555;
    defparam add_371_9.INJECT1_0 = "NO";
    defparam add_371_9.INJECT1_1 = "NO";
    PFUMX i19793 (.BLUT(n22123), .ALUT(n22124), .C0(index_q[6]), .Z(n22132));
    LUT4 n24493_bdd_3_lut (.A(n26844), .B(n444), .C(index_i[5]), .Z(n24494)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n24493_bdd_3_lut.init = 16'hcaca;
    LUT4 mux_191_Mux_2_i573_3_lut_3_lut_4_lut (.A(n26546), .B(index_i[3]), 
         .C(n557_adj_2420), .D(index_i[4]), .Z(n573_adj_2421)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_2_i573_3_lut_3_lut_4_lut.init = 16'h11f0;
    LUT4 i20157_3_lut (.A(n22492), .B(n22493), .C(index_q[8]), .Z(n22496)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20157_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_5_i700_3_lut (.A(n460_adj_2395), .B(n26727), .C(index_q[4]), 
         .Z(n700_adj_2422)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_5_i700_3_lut.init = 16'hcaca;
    LUT4 i20196_3_lut_4_lut (.A(n26546), .B(index_i[3]), .C(index_i[4]), 
         .D(n285_adj_2423), .Z(n22535)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20196_3_lut_4_lut.init = 16'hfe0e;
    LUT4 i20120_3_lut (.A(n22456), .B(n22457), .C(index_i[8]), .Z(n22459)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20120_3_lut.init = 16'hcaca;
    L6MUX21 i20730 (.D0(n23061), .D1(n23062), .SD(index_q[6]), .Z(n23069));
    LUT4 i20119_3_lut (.A(n22454), .B(n22455), .C(index_i[8]), .Z(n22458)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20119_3_lut.init = 16'hcaca;
    PFUMX i20708 (.BLUT(n589), .ALUT(n604), .C0(index_q[4]), .Z(n23047));
    LUT4 mux_191_Mux_6_i92_3_lut_4_lut_3_lut_rep_739 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26699)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_6_i92_3_lut_4_lut_3_lut_rep_739.init = 16'h6969;
    PFUMX i19218 (.BLUT(n21536), .ALUT(n21537), .C0(index_i[4]), .Z(n21538));
    LUT4 mux_191_Mux_10_i125_3_lut_4_lut_4_lut (.A(n26546), .B(index_i[3]), 
         .C(index_i[4]), .D(n26486), .Z(n125_adj_2424)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B (C (D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_10_i125_3_lut_4_lut_4_lut.init = 16'h3efe;
    L6MUX21 i20731 (.D0(n23063), .D1(n23064), .SD(index_q[6]), .Z(n23070));
    L6MUX21 i20732 (.D0(n23065), .D1(n23066), .SD(index_q[6]), .Z(n23071));
    L6MUX21 i20733 (.D0(n23067), .D1(n23068), .SD(index_q[6]), .Z(n23072));
    PFUMX i18690 (.BLUT(n21008), .ALUT(n21009), .C0(index_q[4]), .Z(n21010));
    LUT4 n699_bdd_3_lut_22837_4_lut (.A(n26546), .B(index_i[3]), .C(index_i[4]), 
         .D(n124_adj_2425), .Z(n24440)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n699_bdd_3_lut_22837_4_lut.init = 16'hf101;
    LUT4 mux_191_Mux_0_i157_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n157_adj_2426)) /* synthesis lut_function=(A (B (C+!(D))+!B !(D))+!A (B (D)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_0_i157_3_lut_4_lut.init = 16'hd4aa;
    PFUMX i20709 (.BLUT(n620_adj_2427), .ALUT(n635), .C0(index_q[4]), 
          .Z(n23048));
    LUT4 mux_192_Mux_0_i1017_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[0]), .D(index_q[3]), .Z(n1017_adj_2428)) /* synthesis lut_function=(A (B (D)+!B !((D)+!C))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_0_i1017_4_lut_4_lut_4_lut.init = 16'hdd70;
    LUT4 i20025_3_lut (.A(n22359), .B(n24311), .C(index_i[7]), .Z(n22364)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20025_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_5_i954_3_lut_4_lut_4_lut (.A(index_q[2]), .B(index_q[0]), 
         .C(index_q[3]), .D(index_q[1]), .Z(n954_adj_2429)) /* synthesis lut_function=(!(A (C)+!A (B+((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_5_i954_3_lut_4_lut_4_lut.init = 16'h0a1a;
    LUT4 i20024_3_lut (.A(n22357), .B(n22358), .C(index_i[7]), .Z(n22363)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20024_3_lut.init = 16'hcaca;
    LUT4 i22294_3_lut (.A(n22363), .B(n22364), .C(index_i[8]), .Z(n22366)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22294_3_lut.init = 16'hcaca;
    LUT4 i19980_3_lut (.A(n22315), .B(n22316), .C(index_i[8]), .Z(n22319)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19980_3_lut.init = 16'hcaca;
    PFUMX i24516 (.BLUT(n26820), .ALUT(n26821), .C0(index_i[8]), .Z(n26822));
    LUT4 mux_191_Mux_4_i573_3_lut_3_lut_4_lut_4_lut (.A(n26546), .B(index_i[3]), 
         .C(index_i[4]), .D(n26519), .Z(n573_adj_2430)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_4_i573_3_lut_3_lut_4_lut_4_lut.init = 16'h1f1c;
    CCU2D add_371_7 (.A0(quarter_wave_sample_register_i[6]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[7]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17348), .COUT(n17349), 
          .S1(o_val_pipeline_i_0__15__N_2158[7]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam add_371_7.INIT0 = 16'hf555;
    defparam add_371_7.INIT1 = 16'hf555;
    defparam add_371_7.INJECT1_0 = "NO";
    defparam add_371_7.INJECT1_1 = "NO";
    LUT4 i19481_3_lut (.A(n29163), .B(n26725), .C(index_q[3]), .Z(n21801)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19481_3_lut.init = 16'hcaca;
    LUT4 i22274_3_lut (.A(n22308), .B(n22309), .C(index_q[8]), .Z(n22312)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22274_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_0_i653_3_lut (.A(n26521), .B(n29176), .C(index_q[3]), 
         .Z(n653_adj_2431)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_0_i653_3_lut.init = 16'hcaca;
    LUT4 mux_191_Mux_3_i573_3_lut_3_lut_4_lut (.A(n26546), .B(index_i[3]), 
         .C(n397_adj_2432), .D(index_i[4]), .Z(n573_adj_2433)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_3_i573_3_lut_3_lut_4_lut.init = 16'h11f0;
    LUT4 mux_191_Mux_5_i739_rep_740 (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .Z(n26700)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_5_i739_rep_740.init = 16'h6464;
    LUT4 i19881_3_lut (.A(n22216), .B(n22217), .C(index_q[8]), .Z(n22220)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19881_3_lut.init = 16'hcaca;
    LUT4 i22280_3_lut (.A(n574_adj_2434), .B(n637), .C(index_q[6]), .Z(n21215)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22280_3_lut.init = 16'hcaca;
    LUT4 i22282_3_lut (.A(n574_adj_2435), .B(n637_adj_2296), .C(index_i[6]), 
         .Z(n21206)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22282_3_lut.init = 16'hcaca;
    PFUMX i20710 (.BLUT(n653_adj_2431), .ALUT(n668_adj_2436), .C0(index_q[4]), 
          .Z(n23049));
    PFUMX i20711 (.BLUT(n684_adj_2356), .ALUT(n699_adj_2362), .C0(index_q[4]), 
          .Z(n23050));
    PFUMX i20712 (.BLUT(n716_adj_2386), .ALUT(n731_adj_2437), .C0(index_q[4]), 
          .Z(n23051));
    LUT4 i19471_3_lut (.A(n29197), .B(n26737), .C(index_q[3]), .Z(n21791)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19471_3_lut.init = 16'hcaca;
    PFUMX i20367 (.BLUT(n732_adj_2335), .ALUT(n763_adj_2438), .C0(index_q[5]), 
          .Z(n22706));
    LUT4 i20385_3_lut (.A(n22721), .B(n22722), .C(index_q[8]), .Z(n22724)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20385_3_lut.init = 16'hcaca;
    PFUMX i19227 (.BLUT(n21545), .ALUT(n21546), .C0(index_i[4]), .Z(n21547));
    PFUMX i20713 (.BLUT(n747_adj_2299), .ALUT(n762_adj_2439), .C0(index_q[4]), 
          .Z(n23052));
    PFUMX i20714 (.BLUT(n781_adj_2285), .ALUT(n796), .C0(index_q[4]), 
          .Z(n23053));
    LUT4 i20384_3_lut (.A(n22719), .B(n22720), .C(index_q[8]), .Z(n22723)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20384_3_lut.init = 16'hcaca;
    L6MUX21 i20369 (.D0(n21388), .D1(n891_adj_2440), .SD(index_q[5]), 
            .Z(n22708));
    L6MUX21 i20372 (.D0(n22695), .D1(n22696), .SD(index_q[6]), .Z(n22711));
    L6MUX21 i20374 (.D0(n22699), .D1(n22700), .SD(index_q[6]), .Z(n22713));
    L6MUX21 i20375 (.D0(n22701), .D1(n22702), .SD(index_q[6]), .Z(n22714));
    L6MUX21 i20379 (.D0(n22709), .D1(n22710), .SD(index_q[6]), .Z(n22718));
    LUT4 i21446_3_lut (.A(n21788), .B(n21789), .C(index_q[4]), .Z(n21790)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21446_3_lut.init = 16'hcaca;
    PFUMX i20715 (.BLUT(n812_adj_2441), .ALUT(n11812), .C0(index_q[4]), 
          .Z(n23054));
    LUT4 i19296_else_4_lut (.A(index_i[2]), .B(index_i[1]), .C(index_i[4]), 
         .D(index_i[3]), .Z(n26793)) /* synthesis lut_function=(!(A (B (C)+!B (C+(D)))+!A !(B (C (D)+!C !(D))+!B (C+!(D))))) */ ;
    defparam i19296_else_4_lut.init = 16'h581f;
    PFUMX i19230 (.BLUT(n21548), .ALUT(n21549), .C0(index_i[4]), .Z(n21550));
    LUT4 i18692_3_lut (.A(n498), .B(n29173), .C(index_q[3]), .Z(n21012)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18692_3_lut.init = 16'hcaca;
    PFUMX i20717 (.BLUT(n875_adj_2442), .ALUT(n890_adj_2323), .C0(index_q[4]), 
          .Z(n23056));
    LUT4 mux_191_Mux_7_i956_3_lut_3_lut_4_lut (.A(n26437), .B(index_i[4]), 
         .C(n924_adj_2443), .D(index_i[5]), .Z(n956)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_7_i956_3_lut_3_lut_4_lut.init = 16'h11f0;
    LUT4 index_i_1__bdd_4_lut_25383 (.A(index_i[1]), .B(index_i[3]), .C(index_i[0]), 
         .D(index_i[2]), .Z(n27885)) /* synthesis lut_function=(A (B (C+(D))+!B (C (D)))+!A !(B (C)+!B !(C+(D)))) */ ;
    defparam index_i_1__bdd_4_lut_25383.init = 16'hbd94;
    CCU2D add_371_5 (.A0(quarter_wave_sample_register_i[4]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[5]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17347), .COUT(n17348));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam add_371_5.INIT0 = 16'hf555;
    defparam add_371_5.INIT1 = 16'hf555;
    defparam add_371_5.INJECT1_0 = "NO";
    defparam add_371_5.INJECT1_1 = "NO";
    LUT4 n27885_bdd_3_lut (.A(n27885), .B(index_i[1]), .C(index_i[4]), 
         .Z(n27886)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n27885_bdd_3_lut.init = 16'hcaca;
    LUT4 n77_bdd_3_lut_23888 (.A(n26727), .B(n29198), .C(index_q[3]), 
         .Z(n25591)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n77_bdd_3_lut_23888.init = 16'hacac;
    PFUMX i20718 (.BLUT(n908_adj_2444), .ALUT(n923), .C0(index_q[4]), 
          .Z(n23057));
    LUT4 mux_191_Mux_9_i763_3_lut_4_lut (.A(n26548), .B(n26601), .C(index_i[4]), 
         .D(n26472), .Z(n763_adj_2308)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;
    defparam mux_191_Mux_9_i763_3_lut_4_lut.init = 16'hf101;
    LUT4 mux_192_Mux_1_i317_3_lut (.A(n301), .B(n908_adj_2305), .C(index_q[4]), 
         .Z(n317_adj_2445)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_1_i317_3_lut.init = 16'hcaca;
    LUT4 mux_191_Mux_8_i763_3_lut_4_lut (.A(n26548), .B(n26601), .C(index_i[4]), 
         .D(n26472), .Z(n15024)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam mux_191_Mux_8_i763_3_lut_4_lut.init = 16'hfe0e;
    PFUMX i20719 (.BLUT(n939), .ALUT(n954_adj_2394), .C0(index_q[4]), 
          .Z(n23058));
    LUT4 i18709_3_lut (.A(n325), .B(n26737), .C(index_q[3]), .Z(n21029)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18709_3_lut.init = 16'hcaca;
    PFUMX i18892 (.BLUT(n318), .ALUT(n381_adj_2446), .C0(index_q[6]), 
          .Z(n21212));
    LUT4 i18707_3_lut (.A(n26724), .B(n26734), .C(index_q[3]), .Z(n21027)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18707_3_lut.init = 16'hcaca;
    LUT4 i18706_3_lut (.A(n29173), .B(n29198), .C(index_q[3]), .Z(n21026)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18706_3_lut.init = 16'hcaca;
    LUT4 i20151_3_lut (.A(n22487), .B(n22488), .C(index_i[8]), .Z(n22490)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20151_3_lut.init = 16'hcaca;
    LUT4 i20150_3_lut (.A(n22485), .B(n22486), .C(index_i[8]), .Z(n22489)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20150_3_lut.init = 16'hcaca;
    LUT4 i18704_3_lut (.A(n26740), .B(n29198), .C(index_q[3]), .Z(n21024)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18704_3_lut.init = 16'hcaca;
    PFUMX i20720 (.BLUT(n971), .ALUT(n986), .C0(index_q[4]), .Z(n23059));
    LUT4 i20089_3_lut (.A(n22425), .B(n22426), .C(index_i[8]), .Z(n22428)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20089_3_lut.init = 16'hcaca;
    LUT4 i18695_3_lut_4_lut (.A(n26569), .B(index_q[2]), .C(index_q[3]), 
         .D(n26528), .Z(n21015)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18695_3_lut_4_lut.init = 16'h6f60;
    PFUMX i18883 (.BLUT(n318_adj_2380), .ALUT(n381), .C0(index_i[6]), 
          .Z(n21203));
    LUT4 i20088_3_lut (.A(n22423), .B(n22424), .C(index_i[8]), .Z(n22427)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20088_3_lut.init = 16'hcaca;
    PFUMX i20721 (.BLUT(n1002), .ALUT(n1017_adj_2428), .C0(index_q[4]), 
          .Z(n23060));
    LUT4 i18700_3_lut (.A(n26543), .B(n29198), .C(index_q[3]), .Z(n21020)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18700_3_lut.init = 16'hcaca;
    LUT4 i19058_3_lut_4_lut_4_lut_4_lut (.A(n26569), .B(index_q[2]), .C(index_q[3]), 
         .D(index_q[4]), .Z(n21378)) /* synthesis lut_function=(A (B)+!A (B (C (D))+!B !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19058_3_lut_4_lut_4_lut_4_lut.init = 16'hc999;
    LUT4 index_i_2__bdd_4_lut_25804 (.A(index_i[2]), .B(index_i[0]), .C(index_i[4]), 
         .D(index_i[1]), .Z(n27925)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((C (D))+!B))) */ ;
    defparam index_i_2__bdd_4_lut_25804.init = 16'h0cec;
    LUT4 mux_192_Mux_2_i604_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n604_adj_2447)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)+!C !(D)))+!A (B (D)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_2_i604_3_lut_4_lut_4_lut_4_lut.init = 16'h39cf;
    LUT4 i19453_3_lut (.A(n900), .B(n29173), .C(index_q[3]), .Z(n21773)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19453_3_lut.init = 16'hcaca;
    LUT4 index_i_2__bdd_3_lut_25988 (.A(index_i[2]), .B(index_i[0]), .C(index_i[4]), 
         .Z(n27926)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B (C)+!B !(C)))) */ ;
    defparam index_i_2__bdd_3_lut_25988.init = 16'h6969;
    LUT4 i20026_3_lut (.A(n22361), .B(n22362), .C(index_i[8]), .Z(n22365)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20026_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_0_i142_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n142_adj_2448)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C))+!A !(B (C (D)+!C !(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_0_i142_3_lut_4_lut_4_lut.init = 16'ha569;
    LUT4 i19959_3_lut (.A(n22295), .B(n22296), .C(index_q[8]), .Z(n22298)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19959_3_lut.init = 16'hcaca;
    LUT4 i19958_3_lut (.A(n22293), .B(n22294), .C(index_q[8]), .Z(n22297)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19958_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_0_i762_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n762_adj_2439)) /* synthesis lut_function=(A (B+!((D)+!C))+!A !(B (D)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_0_i762_3_lut_4_lut_4_lut.init = 16'h98fc;
    LUT4 i21455_3_lut (.A(n26841), .B(n21768), .C(index_q[4]), .Z(n21769)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21455_3_lut.init = 16'hcaca;
    L6MUX21 i19961 (.D0(n21343), .D1(n21346), .SD(index_q[6]), .Z(n22300));
    LUT4 i15391_3_lut (.A(n26714), .B(n26724), .C(index_q[3]), .Z(n17541)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15391_3_lut.init = 16'hcaca;
    PFUMX i15419 (.BLUT(n17567), .ALUT(n17568), .C0(index_i[4]), .Z(n17569));
    LUT4 i15390_3_lut (.A(n26724), .B(n29171), .C(index_q[3]), .Z(n17540)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15390_3_lut.init = 16'hcaca;
    LUT4 n26603_bdd_3_lut_25604 (.A(n26486), .B(n29178), .C(index_i[4]), 
         .Z(n27928)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n26603_bdd_3_lut_25604.init = 16'hcaca;
    LUT4 mux_192_Mux_7_i475_3_lut_4_lut (.A(n26569), .B(index_q[2]), .C(index_q[3]), 
         .D(n29189), .Z(n475_adj_2449)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_7_i475_3_lut_4_lut.init = 16'h9f90;
    LUT4 i20473_3_lut (.A(n250), .B(n26528), .C(index_q[3]), .Z(n22812)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20473_3_lut.init = 16'hcaca;
    LUT4 i19277_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21597)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A (B (C (D)+!C !(D))+!B (D))) */ ;
    defparam i19277_3_lut_4_lut.init = 16'hd926;
    LUT4 i20472_3_lut (.A(n676), .B(n29187), .C(index_q[3]), .Z(n22811)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20472_3_lut.init = 16'hcaca;
    LUT4 i11407_3_lut_4_lut (.A(n26350), .B(index_i[7]), .C(index_i[8]), 
         .D(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2127[14])) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11407_3_lut_4_lut.init = 16'hffe0;
    PFUMX i20339 (.BLUT(n22674), .ALUT(n22675), .C0(index_i[4]), .Z(n22678));
    LUT4 i20471_3_lut (.A(n29181), .B(n26571), .C(index_q[3]), .Z(n22810)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20471_3_lut.init = 16'hcaca;
    LUT4 i20470_3_lut (.A(n26528), .B(n29189), .C(index_q[3]), .Z(n22809)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20470_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_2_i684_3_lut_4_lut (.A(n26569), .B(index_q[2]), .C(index_q[3]), 
         .D(n29181), .Z(n684_adj_2450)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_2_i684_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_192_Mux_3_i158_3_lut (.A(n142_adj_2451), .B(n157_adj_2452), 
         .C(index_q[4]), .Z(n158_adj_2453)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_3_i158_3_lut.init = 16'hcaca;
    PFUMX i20340 (.BLUT(n22676), .ALUT(n22677), .C0(index_i[4]), .Z(n22679));
    LUT4 mux_192_Mux_3_i125_3_lut (.A(n109_adj_2454), .B(n526_adj_2360), 
         .C(index_q[4]), .Z(n125_adj_2455)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_3_i125_3_lut.init = 16'hcaca;
    LUT4 n715_bdd_3_lut_23915_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n25632)) /* synthesis lut_function=(A (B (C+(D))+!B ((D)+!C))+!A !(B (C+(D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n715_bdd_3_lut_23915_4_lut.init = 16'haa96;
    L6MUX21 i19869 (.D0(n22192), .D1(n22193), .SD(index_q[6]), .Z(n22208));
    L6MUX21 i19870 (.D0(n22194), .D1(n22195), .SD(index_q[6]), .Z(n22209));
    L6MUX21 i19871 (.D0(n22196), .D1(n22197), .SD(index_q[6]), .Z(n22210));
    L6MUX21 i19872 (.D0(n22198), .D1(n22199), .SD(index_q[6]), .Z(n22211));
    LUT4 mux_192_Mux_7_i653_3_lut_4_lut (.A(n26569), .B(index_q[2]), .C(index_q[3]), 
         .D(n29192), .Z(n653_adj_2456)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_7_i653_3_lut_4_lut.init = 16'hf606;
    L6MUX21 i19873 (.D0(n22200), .D1(n22201), .SD(index_q[6]), .Z(n22212));
    L6MUX21 i19875 (.D0(n22204), .D1(n22205), .SD(index_q[6]), .Z(n22214));
    LUT4 i19060_4_lut_4_lut_4_lut (.A(n26569), .B(index_q[2]), .C(index_q[4]), 
         .D(index_q[3]), .Z(n21380)) /* synthesis lut_function=(A (B)+!A !(B (C+(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19060_4_lut_4_lut_4_lut.init = 16'h999c;
    LUT4 i19914_4_lut (.A(n26745), .B(n1002_adj_2457), .C(index_q[5]), 
         .D(index_q[4]), .Z(n22253)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;
    defparam i19914_4_lut.init = 16'hfaca;
    LUT4 i18913_3_lut_3_lut_4_lut (.A(n26437), .B(index_i[4]), .C(n700_adj_2415), 
         .D(index_i[5]), .Z(n21233)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18913_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 i18922_3_lut_3_lut_4_lut (.A(n26429), .B(index_q[4]), .C(n700), 
         .D(index_q[5]), .Z(n21242)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18922_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 mux_192_Mux_0_i908_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n908_adj_2444)) /* synthesis lut_function=(!(A (B (C (D))+!B !(D))+!A (B+((D)+!C)))) */ ;
    defparam mux_192_Mux_0_i908_3_lut_4_lut_4_lut.init = 16'h2a98;
    LUT4 mux_192_Mux_4_i860_3_lut (.A(n506_adj_2458), .B(n25071), .C(index_q[4]), 
         .Z(n860_adj_2459)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_4_i860_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_1_i93_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n93_adj_2460)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C+(D)))+!A !(B (C (D)+!C !(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_1_i93_3_lut_4_lut_4_lut.init = 16'h955a;
    PFUMX i24469 (.BLUT(n26746), .ALUT(n26747), .C0(index_q[2]), .Z(n26748));
    LUT4 mux_191_Mux_10_i701_4_lut_4_lut (.A(n26437), .B(index_i[4]), .C(index_i[5]), 
         .D(n26393), .Z(n701)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B (C (D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_10_i701_4_lut_4_lut.init = 16'h3efe;
    L6MUX21 i19915 (.D0(n22238), .D1(n22239), .SD(index_q[6]), .Z(n22254));
    LUT4 i21308_3_lut (.A(n21065), .B(n21066), .C(index_q[4]), .Z(n21067)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21308_3_lut.init = 16'hcaca;
    LUT4 n26462_bdd_4_lut_25711 (.A(index_q[5]), .B(index_q[2]), .C(index_q[0]), 
         .D(index_q[1]), .Z(n27992)) /* synthesis lut_function=(!(A (B (D)+!B ((D)+!C))+!A !(B (C (D)+!C !(D))+!B !(D)))) */ ;
    defparam n26462_bdd_4_lut_25711.init = 16'h40bd;
    L6MUX21 i19916 (.D0(n22240), .D1(n22241), .SD(index_q[6]), .Z(n22255));
    L6MUX21 i19917 (.D0(n22242), .D1(n22243), .SD(index_q[6]), .Z(n22256));
    LUT4 i21310_3_lut (.A(n21062), .B(n21063), .C(index_q[4]), .Z(n21064)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21310_3_lut.init = 16'hcaca;
    LUT4 n26528_bdd_3_lut_25715 (.A(index_q[2]), .B(index_q[0]), .C(index_q[4]), 
         .Z(n27995)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B (C)+!B !(C)))) */ ;
    defparam n26528_bdd_3_lut_25715.init = 16'h6969;
    PFUMX i19919 (.BLUT(n22246), .ALUT(n22247), .C0(index_q[6]), .Z(n22258));
    LUT4 mux_192_Mux_4_i700_3_lut (.A(n684_adj_2461), .B(index_q[1]), .C(index_q[4]), 
         .Z(n700_adj_2462)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_4_i700_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_4_i669_3_lut (.A(n781_adj_2303), .B(n668_adj_2336), 
         .C(index_q[4]), .Z(n669_adj_2463)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_4_i669_3_lut.init = 16'hcaca;
    PFUMX i19248 (.BLUT(n21566), .ALUT(n21567), .C0(index_q[4]), .Z(n21568));
    LUT4 mux_192_Mux_2_i189_3_lut_3_lut_4_lut (.A(index_q[1]), .B(n26539), 
         .C(n173_adj_2307), .D(index_q[4]), .Z(n189_adj_2464)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(C+(D)))) */ ;
    defparam mux_192_Mux_2_i189_3_lut_3_lut_4_lut.init = 16'h77f0;
    LUT4 mux_192_Mux_0_i851_3_lut_3_lut_rep_784 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29163)) /* synthesis lut_function=(A (B+(C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_0_i851_3_lut_3_lut_rep_784.init = 16'hadad;
    LUT4 mux_192_Mux_4_i874_3_lut_rep_785 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29164)) /* synthesis lut_function=(A (B+!(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_4_i874_3_lut_rep_785.init = 16'hdada;
    L6MUX21 i19920 (.D0(n22248), .D1(n22249), .SD(index_q[6]), .Z(n22259));
    LUT4 mux_192_Mux_4_i542_3_lut (.A(n526_adj_2360), .B(n541_adj_2288), 
         .C(index_q[4]), .Z(n542)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_4_i542_3_lut.init = 16'hcaca;
    L6MUX21 i19921 (.D0(n22250), .D1(n22251), .SD(index_q[6]), .Z(n22260));
    LUT4 i19908_4_lut (.A(n26523), .B(n26857), .C(index_q[5]), .D(index_q[4]), 
         .Z(n22247)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam i19908_4_lut.init = 16'hc5ca;
    PFUMX i19922 (.BLUT(n22252), .ALUT(n22253), .C0(index_q[6]), .Z(n22261));
    LUT4 n715_bdd_3_lut_24008 (.A(n26571), .B(n26736), .C(index_q[3]), 
         .Z(n25633)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n715_bdd_3_lut_24008.init = 16'hcaca;
    PFUMX i20346 (.BLUT(n22681), .ALUT(n22682), .C0(index_i[4]), .Z(n22685));
    L6MUX21 i20792 (.D0(n23123), .D1(n23124), .SD(index_i[6]), .Z(n23131));
    L6MUX21 i20793 (.D0(n23125), .D1(n23126), .SD(index_i[6]), .Z(n23132));
    LUT4 i11512_2_lut_3_lut_4_lut (.A(index_q[1]), .B(n26539), .C(index_q[5]), 
         .D(index_q[4]), .Z(n508)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;
    defparam i11512_2_lut_3_lut_4_lut.init = 16'hf080;
    L6MUX21 i20794 (.D0(n23127), .D1(n23128), .SD(index_i[6]), .Z(n23133));
    PFUMX i19934 (.BLUT(n286), .ALUT(n21079), .C0(index_q[5]), .Z(n22273));
    LUT4 mux_191_Mux_14_i511_4_lut_4_lut (.A(n26350), .B(index_i[7]), .C(index_i[8]), 
         .D(n254_adj_2465), .Z(n511_adj_2466)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (B (C+!(D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_14_i511_4_lut_4_lut.init = 16'h1c10;
    PFUMX i19935 (.BLUT(n349_adj_2467), .ALUT(n21082), .C0(index_q[5]), 
          .Z(n22274));
    LUT4 mux_192_Mux_4_i286_3_lut (.A(n270_adj_2468), .B(n15_adj_2469), 
         .C(index_q[4]), .Z(n286_adj_2470)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_4_i286_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_4_i94_3_lut (.A(n61), .B(n26583), .C(index_q[4]), 
         .Z(n94)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_4_i94_3_lut.init = 16'hcaca;
    LUT4 i20599_3_lut_4_lut (.A(n26451), .B(n26393), .C(index_i[4]), .D(index_i[5]), 
         .Z(n22938)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (B+((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20599_3_lut_4_lut.init = 16'hffc5;
    PFUMX i19936 (.BLUT(n413), .ALUT(n444_adj_2471), .C0(index_q[5]), 
          .Z(n22275));
    PFUMX i19937 (.BLUT(n476), .ALUT(n507), .C0(index_q[5]), .Z(n22276));
    PFUMX i19251 (.BLUT(n21569), .ALUT(n21570), .C0(index_q[4]), .Z(n21571));
    PFUMX i19938 (.BLUT(n21085), .ALUT(n573_adj_2472), .C0(index_q[5]), 
          .Z(n22277));
    PFUMX i19939 (.BLUT(n11873), .ALUT(n21088), .C0(index_q[5]), .Z(n22278));
    PFUMX i20347 (.BLUT(n22683), .ALUT(n22684), .C0(index_i[4]), .Z(n22686));
    PFUMX i19940 (.BLUT(n669), .ALUT(n700_adj_2473), .C0(index_q[5]), 
          .Z(n22279));
    L6MUX21 i19941 (.D0(n21091), .D1(n763_adj_2474), .SD(index_q[5]), 
            .Z(n22280));
    PFUMX i19943 (.BLUT(n860_adj_2475), .ALUT(n891), .C0(index_q[5]), 
          .Z(n22282));
    LUT4 mux_192_Mux_1_i620_3_lut_4_lut (.A(n26623), .B(index_q[1]), .C(index_q[3]), 
         .D(n29170), .Z(n620_adj_2476)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_1_i620_3_lut_4_lut.init = 16'hdfd0;
    PFUMX i19944 (.BLUT(n924_adj_2477), .ALUT(n21094), .C0(index_q[5]), 
          .Z(n22283));
    LUT4 index_i_1__bdd_4_lut (.A(index_i[1]), .B(index_i[0]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n29205)) /* synthesis lut_function=(A (B+(C (D)+!C !(D)))+!A !(B (C+(D))+!B !(C))) */ ;
    defparam index_i_1__bdd_4_lut.init = 16'hb89e;
    PFUMX i19945 (.BLUT(n21097), .ALUT(n1018), .C0(index_q[5]), .Z(n22284));
    LUT4 mux_192_Mux_0_i173_3_lut_4_lut (.A(n26623), .B(index_q[1]), .C(index_q[3]), 
         .D(n29171), .Z(n173_adj_2478)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_0_i173_3_lut_4_lut.init = 16'hdfd0;
    L6MUX21 i20476 (.D0(n22813), .D1(n22814), .SD(index_q[5]), .Z(n22815));
    LUT4 i18701_3_lut_4_lut (.A(n26623), .B(index_q[1]), .C(index_q[3]), 
         .D(n498), .Z(n21021)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18701_3_lut_4_lut.init = 16'hdfd0;
    PFUMX i18884 (.BLUT(n445_adj_2348), .ALUT(n508_adj_2479), .C0(index_i[6]), 
          .Z(n21204));
    PFUMX i20353 (.BLUT(n22688), .ALUT(n22689), .C0(index_i[4]), .Z(n22692));
    PFUMX i18893 (.BLUT(n445), .ALUT(n508), .C0(index_q[6]), .Z(n21213));
    PFUMX i24514 (.BLUT(n26817), .ALUT(n26818), .C0(index_q[0]), .Z(n26819));
    PFUMX i19990 (.BLUT(n956), .ALUT(n20003), .C0(index_i[6]), .Z(n22329));
    LUT4 n24537_bdd_3_lut (.A(n24537), .B(n476_adj_2408), .C(index_i[5]), 
         .Z(n24538)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n24537_bdd_3_lut.init = 16'hcaca;
    LUT4 n62_bdd_3_lut_25698 (.A(n62), .B(n125_adj_2480), .C(index_q[6]), 
         .Z(n28120)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n62_bdd_3_lut_25698.init = 16'hcaca;
    PFUMX i20354 (.BLUT(n22690), .ALUT(n22691), .C0(index_i[4]), .Z(n22693));
    PFUMX i19257 (.BLUT(n21575), .ALUT(n21576), .C0(index_q[4]), .Z(n21577));
    PFUMX i19999 (.BLUT(n94_adj_2481), .ALUT(n125_adj_2482), .C0(index_i[5]), 
          .Z(n22338));
    PFUMX i20000 (.BLUT(n17585), .ALUT(n14366), .C0(index_i[5]), .Z(n22339));
    LUT4 mux_192_Mux_0_i660_3_lut_rep_794 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29173)) /* synthesis lut_function=(A (B)+!A (B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_0_i660_3_lut_rep_794.init = 16'hc9c9;
    LUT4 i19462_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21782)) /* synthesis lut_function=(!(A (B (C (D))+!B (C (D)+!C !(D)))+!A !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19462_3_lut_4_lut_4_lut.init = 16'h5aad;
    LUT4 mux_192_Mux_9_i763_3_lut_4_lut (.A(n26567), .B(n26585), .C(index_q[4]), 
         .D(n26482), .Z(n763_adj_2329)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;
    defparam mux_192_Mux_9_i763_3_lut_4_lut.init = 16'hf101;
    L6MUX21 i20002 (.D0(n21583), .D1(n21586), .SD(index_i[5]), .Z(n22341));
    LUT4 n22825_bdd_4_lut_25695 (.A(n252_adj_2483), .B(n26429), .C(index_q[4]), 
         .D(index_q[5]), .Z(n28118)) /* synthesis lut_function=(A (B (D)+!B ((D)+!C))+!A !(B+(C+(D)))) */ ;
    defparam n22825_bdd_4_lut_25695.init = 16'haa03;
    PFUMX i19263 (.BLUT(n21581), .ALUT(n21582), .C0(index_i[4]), .Z(n21583));
    L6MUX21 i20003 (.D0(n21589), .D1(n21592), .SD(index_i[5]), .Z(n22342));
    LUT4 mux_192_Mux_8_i763_3_lut_4_lut (.A(n26567), .B(n26585), .C(index_q[4]), 
         .D(n26482), .Z(n15038)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam mux_192_Mux_8_i763_3_lut_4_lut.init = 16'hfe0e;
    LUT4 n62_bdd_4_lut_25699 (.A(n26585), .B(n26477), .C(index_q[6]), 
         .D(index_q[4]), .Z(n28121)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C+(D)))+!A (B ((D)+!C)+!B !(C)))) */ ;
    defparam n62_bdd_4_lut_25699.init = 16'h3af0;
    PFUMX i19266 (.BLUT(n21584), .ALUT(n21585), .C0(index_i[4]), .Z(n21586));
    LUT4 mux_192_Mux_3_i796_3_lut (.A(index_q[2]), .B(n781), .C(index_q[4]), 
         .Z(n796_adj_2484)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_3_i796_3_lut.init = 16'hacac;
    LUT4 i18748_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21068)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18748_3_lut_4_lut_4_lut.init = 16'hda5a;
    PFUMX i20004 (.BLUT(n413_adj_2485), .ALUT(n444_adj_2486), .C0(index_i[5]), 
          .Z(n22343));
    LUT4 mux_192_Mux_3_i781_3_lut (.A(n29182), .B(n26528), .C(index_q[3]), 
         .Z(n781)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_3_i781_3_lut.init = 16'hcaca;
    PFUMX i20005 (.BLUT(n476_adj_2487), .ALUT(n507_adj_2488), .C0(index_i[5]), 
          .Z(n22344));
    LUT4 n24541_bdd_3_lut_23046 (.A(n26837), .B(n24539), .C(index_i[5]), 
         .Z(n24542)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n24541_bdd_3_lut_23046.init = 16'hcaca;
    LUT4 n22978_bdd_4_lut_25670 (.A(n252_adj_2316), .B(n26437), .C(index_i[4]), 
         .D(index_i[5]), .Z(n28177)) /* synthesis lut_function=(A (B (D)+!B ((D)+!C))+!A !(B+(C+(D)))) */ ;
    defparam n22978_bdd_4_lut_25670.init = 16'haa03;
    LUT4 n62_bdd_3_lut_25673 (.A(n62_adj_2292), .B(n125_adj_2424), .C(index_i[6]), 
         .Z(n28179)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n62_bdd_3_lut_25673.init = 16'hcaca;
    PFUMX i20006 (.BLUT(n17575), .ALUT(n573_adj_2489), .C0(index_i[5]), 
          .Z(n22345));
    LUT4 n62_bdd_4_lut_25674 (.A(n26601), .B(n26485), .C(index_i[6]), 
         .D(index_i[4]), .Z(n28180)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C+(D)))+!A (B ((D)+!C)+!B !(C)))) */ ;
    defparam n62_bdd_4_lut_25674.init = 16'h3af0;
    LUT4 mux_192_Mux_5_i891_3_lut (.A(n875_adj_2490), .B(n890_adj_2338), 
         .C(index_q[4]), .Z(n891_adj_2491)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_5_i891_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_5_i860_3_lut (.A(n15_adj_2492), .B(n859_adj_2493), 
         .C(index_q[4]), .Z(n860_adj_2494)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_5_i860_3_lut.init = 16'hcaca;
    PFUMX i20007 (.BLUT(n605), .ALUT(n636_adj_2495), .C0(index_i[5]), 
          .Z(n22346));
    LUT4 mux_192_Mux_4_i62_4_lut (.A(n29172), .B(n61), .C(index_q[4]), 
         .D(index_q[3]), .Z(n62_adj_2496)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_4_i62_4_lut.init = 16'hc5ca;
    PFUMX i20008 (.BLUT(n21595), .ALUT(n700_adj_2497), .C0(index_i[5]), 
          .Z(n22347));
    LUT4 mux_192_Mux_4_i31_4_lut (.A(n15_adj_2469), .B(n26513), .C(index_q[4]), 
         .D(index_q[3]), .Z(n31)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_4_i31_4_lut.init = 16'h3aca;
    LUT4 i9612_3_lut_then_4_lut (.A(index_q[4]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n29207)) /* synthesis lut_function=(A (B (C)+!B !(C (D)+!C !(D)))+!A (B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9612_3_lut_then_4_lut.init = 16'hd6a5;
    LUT4 i21355_3_lut (.A(n21032), .B(n21033), .C(index_q[4]), .Z(n21034)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21355_3_lut.init = 16'hcaca;
    L6MUX21 i20009 (.D0(n732_adj_2340), .D1(n21598), .SD(index_i[5]), 
            .Z(n22348));
    PFUMX i20010 (.BLUT(n797_adj_2498), .ALUT(n828_adj_2396), .C0(index_i[5]), 
          .Z(n22349));
    LUT4 mux_192_Mux_5_i636_4_lut (.A(n157_adj_2342), .B(n26426), .C(index_q[4]), 
         .D(index_q[3]), .Z(n636_adj_2499)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_5_i636_4_lut.init = 16'h3aca;
    LUT4 i21358_3_lut (.A(n17543), .B(n17544), .C(index_q[4]), .Z(n17545)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21358_3_lut.init = 16'hcaca;
    L6MUX21 mux_192_Mux_7_i253 (.D0(n12030), .D1(n21733), .SD(index_q[5]), 
            .Z(n253)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 mux_192_Mux_9_i124_3_lut_3_lut_4_lut (.A(n26567), .B(index_q[2]), 
         .C(n26496), .D(index_q[3]), .Z(n124_adj_2500)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_9_i124_3_lut_3_lut_4_lut.init = 16'h11f0;
    LUT4 mux_192_Mux_5_i507_3_lut (.A(n491_adj_2334), .B(n506_adj_2458), 
         .C(index_q[4]), .Z(n507_adj_2501)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_5_i507_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_0_i1002_3_lut_3_lut_4_lut (.A(n26567), .B(index_q[2]), 
         .C(n1001), .D(index_q[3]), .Z(n1002)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_0_i1002_3_lut_3_lut_4_lut.init = 16'hf011;
    PFUMX i20011 (.BLUT(n860_adj_2502), .ALUT(n891_adj_2503), .C0(index_i[5]), 
          .Z(n22350));
    LUT4 mux_192_Mux_5_i476_3_lut (.A(n460_adj_2395), .B(n475), .C(index_q[4]), 
         .Z(n476_adj_2504)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_5_i476_3_lut.init = 16'hcaca;
    LUT4 i19703_2_lut (.A(index_q[3]), .B(index_q[5]), .Z(n22042)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19703_2_lut.init = 16'h8888;
    LUT4 mux_192_Mux_5_i413_3_lut (.A(n397_adj_2505), .B(n251_adj_2398), 
         .C(index_q[4]), .Z(n413_adj_2506)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_5_i413_3_lut.init = 16'hcaca;
    LUT4 i15429_3_lut (.A(n17577), .B(n17578), .C(index_q[4]), .Z(n17579)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15429_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_8_i475_3_lut_3_lut_4_lut (.A(n26567), .B(index_q[2]), 
         .C(n26496), .D(index_q[3]), .Z(n475_adj_2507)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_8_i475_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 index_i_0__bdd_4_lut_25733 (.A(index_i[0]), .B(index_i[4]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n28280)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(D))+!A !(B (D)+!B (C+!(D))))) */ ;
    defparam index_i_0__bdd_4_lut_25733.init = 16'h7e11;
    PFUMX mux_192_Mux_7_i190 (.BLUT(n21730), .ALUT(n173_adj_2508), .C0(index_q[5]), 
          .Z(n190)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 mux_192_Mux_3_i31_3_lut (.A(n781_adj_2303), .B(n30_adj_2509), .C(index_q[4]), 
         .Z(n31_adj_2510)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_3_i31_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_5_i125_3_lut (.A(n109_adj_2511), .B(n124_adj_2512), 
         .C(index_q[4]), .Z(n125_adj_2513)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_5_i125_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_5_i94_3_lut (.A(n653_adj_2514), .B(n635_adj_2515), 
         .C(index_q[4]), .Z(n94_adj_2516)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_5_i94_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_5_i31_3_lut (.A(n15_adj_2492), .B(n30_adj_2517), .C(index_q[4]), 
         .Z(n31_adj_2518)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_5_i31_3_lut.init = 16'hcaca;
    LUT4 index_i_0__bdd_2_lut (.A(index_i[0]), .B(index_i[2]), .Z(n28281)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam index_i_0__bdd_2_lut.init = 16'h6666;
    LUT4 i20639_4_lut_4_lut (.A(n26419), .B(n26506), .C(index_i[5]), .D(index_i[4]), 
         .Z(n22978)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C+(D))+!B !(C (D)+!C !(D)))) */ ;
    defparam i20639_4_lut_4_lut.init = 16'hcf50;
    LUT4 mux_191_Mux_5_i31_3_lut (.A(n15_adj_2519), .B(n30_adj_2520), .C(index_i[4]), 
         .Z(n31_adj_2521)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_5_i31_3_lut.init = 16'hcaca;
    LUT4 mux_191_Mux_4_i62_4_lut (.A(n26435), .B(n61_adj_2522), .C(index_i[4]), 
         .D(index_i[3]), .Z(n62_adj_2523)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_4_i62_4_lut.init = 16'hc5ca;
    LUT4 mux_191_Mux_4_i31_4_lut (.A(n15_adj_2524), .B(n26433), .C(index_i[4]), 
         .D(index_i[3]), .Z(n31_adj_2525)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_4_i31_4_lut.init = 16'h3aca;
    LUT4 i20421_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n22760)) /* synthesis lut_function=(A (B (C+!(D))+!B !((D)+!C))+!A !(B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20421_3_lut_4_lut_4_lut.init = 16'h81f8;
    LUT4 mux_191_Mux_3_i31_3_lut (.A(n781_adj_2526), .B(n30_adj_2527), .C(index_i[4]), 
         .Z(n31_adj_2528)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_3_i31_3_lut.init = 16'hcaca;
    LUT4 i9558_3_lut (.A(n12003), .B(n26686), .C(index_i[3]), .Z(n12004)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9558_3_lut.init = 16'hcaca;
    PFUMX i19269 (.BLUT(n21587), .ALUT(n21588), .C0(index_i[4]), .Z(n21589));
    PFUMX i20030 (.BLUT(n94_adj_2529), .ALUT(n21601), .C0(index_i[5]), 
          .Z(n22369));
    LUT4 i12213_3_lut (.A(index_i[3]), .B(index_i[1]), .C(index_i[0]), 
         .Z(n14783)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i12213_3_lut.init = 16'hecec;
    PFUMX i19272 (.BLUT(n21590), .ALUT(n21591), .C0(index_i[4]), .Z(n21592));
    PFUMX i20032 (.BLUT(n221_adj_2530), .ALUT(n252_adj_2531), .C0(index_i[5]), 
          .Z(n22371));
    LUT4 n28443_bdd_3_lut (.A(n28443), .B(index_q[1]), .C(index_q[4]), 
         .Z(n28444)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n28443_bdd_3_lut.init = 16'hcaca;
    LUT4 index_q_1__bdd_4_lut_25976 (.A(index_q[1]), .B(index_q[3]), .C(index_q[0]), 
         .D(index_q[2]), .Z(n28443)) /* synthesis lut_function=(A (B (C+(D))+!B (C (D)))+!A !(B (C)+!B !(C+(D)))) */ ;
    defparam index_q_1__bdd_4_lut_25976.init = 16'hbd94;
    PFUMX i20033 (.BLUT(n286_adj_2532), .ALUT(n21604), .C0(index_i[5]), 
          .Z(n22372));
    LUT4 i19400_3_lut_4_lut_4_lut (.A(n26647), .B(n26688), .C(index_i[3]), 
         .D(index_i[2]), .Z(n21720)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B+(C))) */ ;
    defparam i19400_3_lut_4_lut_4_lut.init = 16'hfc5c;
    LUT4 n953_bdd_3_lut_23526_4_lut_4_lut (.A(n26647), .B(n26650), .C(index_i[3]), 
         .D(index_i[2]), .Z(n25215)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B+(C))) */ ;
    defparam n953_bdd_3_lut_23526_4_lut_4_lut.init = 16'hfc5c;
    LUT4 n197_bdd_3_lut_22981 (.A(n26599), .B(index_i[3]), .C(n26703), 
         .Z(n24594)) /* synthesis lut_function=(A (B+(C))+!A !(B+!(C))) */ ;
    defparam n197_bdd_3_lut_22981.init = 16'hb8b8;
    LUT4 i19337_3_lut_4_lut (.A(n26647), .B(index_i[2]), .C(index_i[3]), 
         .D(n308), .Z(n21657)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19337_3_lut_4_lut.init = 16'hf202;
    PFUMX i20034 (.BLUT(n349_adj_2533), .ALUT(n21607), .C0(index_i[5]), 
          .Z(n22373));
    PFUMX mux_192_Mux_1_i636 (.BLUT(n620_adj_2476), .ALUT(n635_adj_2534), 
          .C0(index_q[4]), .Z(n636_adj_2535)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 n197_bdd_3_lut_23522_4_lut (.A(n26602), .B(index_i[2]), .C(index_i[3]), 
         .D(n26587), .Z(n24595)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n197_bdd_3_lut_23522_4_lut.init = 16'hf606;
    LUT4 mux_191_Mux_2_i189_3_lut_3_lut_4_lut (.A(index_i[1]), .B(n26547), 
         .C(n173_adj_2314), .D(index_i[4]), .Z(n189_adj_2536)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(C+(D)))) */ ;
    defparam mux_191_Mux_2_i189_3_lut_3_lut_4_lut.init = 16'h77f0;
    LUT4 mux_191_Mux_3_i890_3_lut_4_lut (.A(n26602), .B(index_i[2]), .C(index_i[3]), 
         .D(n396), .Z(n890_adj_2537)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_3_i890_3_lut_4_lut.init = 16'h6f60;
    LUT4 i11444_2_lut_3_lut_4_lut (.A(index_i[1]), .B(n26547), .C(index_i[5]), 
         .D(index_i[4]), .Z(n508_adj_2479)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;
    defparam i11444_2_lut_3_lut_4_lut.init = 16'hf080;
    PFUMX i19278 (.BLUT(n21596), .ALUT(n21597), .C0(index_i[4]), .Z(n21598));
    LUT4 i19214_3_lut_4_lut (.A(n26602), .B(index_i[2]), .C(index_i[3]), 
         .D(n26699), .Z(n21534)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19214_3_lut_4_lut.init = 16'hf606;
    LUT4 i1_3_lut_4_lut_adj_75 (.A(n26647), .B(n26547), .C(index_i[4]), 
         .D(n26634), .Z(n19979)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;
    defparam i1_3_lut_4_lut_adj_75.init = 16'hfff8;
    LUT4 n285_bdd_3_lut (.A(n26706), .B(n26599), .C(index_i[3]), .Z(n24597)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n285_bdd_3_lut.init = 16'hcaca;
    LUT4 mux_191_Mux_3_i796_3_lut (.A(index_i[2]), .B(n731_adj_2538), .C(index_i[4]), 
         .Z(n796_adj_2539)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_3_i796_3_lut.init = 16'hacac;
    LUT4 mux_191_Mux_6_i731_3_lut (.A(n26606), .B(n29174), .C(index_i[3]), 
         .Z(n731_adj_2538)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_6_i731_3_lut.init = 16'hcaca;
    LUT4 i19722_1_lut_2_lut (.A(index_q[2]), .B(index_q[3]), .Z(n22061)) /* synthesis lut_function=(!(A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19722_1_lut_2_lut.init = 16'h7777;
    LUT4 mux_191_Mux_5_i124_3_lut (.A(n70), .B(n26707), .C(index_i[3]), 
         .Z(n124_adj_2540)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_5_i124_3_lut.init = 16'hcaca;
    CCU2D add_371_3 (.A0(quarter_wave_sample_register_i[2]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[3]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17346), .COUT(n17347));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam add_371_3.INIT0 = 16'hf555;
    defparam add_371_3.INIT1 = 16'hf555;
    defparam add_371_3.INJECT1_0 = "NO";
    defparam add_371_3.INJECT1_1 = "NO";
    LUT4 index_i_4__bdd_4_lut_22920 (.A(index_i[4]), .B(n26437), .C(index_i[7]), 
         .D(n26485), .Z(n24245)) /* synthesis lut_function=(A (C+!(D))+!A (B+!(C))) */ ;
    defparam index_i_4__bdd_4_lut_22920.init = 16'he5ef;
    LUT4 mux_191_Mux_0_i348_3_lut_4_lut (.A(n26602), .B(index_i[2]), .C(index_i[3]), 
         .D(n26604), .Z(n348_adj_2541)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_0_i348_3_lut_4_lut.init = 16'h6f60;
    LUT4 i11640_3_lut_4_lut (.A(n26539), .B(index_q[4]), .C(index_q[5]), 
         .D(n26569), .Z(n892_adj_2542)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11640_3_lut_4_lut.init = 16'hf8f0;
    LUT4 mux_192_Mux_6_i60_3_lut_4_lut_3_lut_rep_783 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29162)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_6_i60_3_lut_4_lut_3_lut_rep_783.init = 16'hd6d6;
    LUT4 mux_192_Mux_2_i700_3_lut_4_lut (.A(index_q[1]), .B(n26585), .C(index_q[4]), 
         .D(n684_adj_2450), .Z(n700_adj_2543)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_2_i700_3_lut_4_lut.init = 16'hefe0;
    PFUMX i26216 (.BLUT(n29206), .ALUT(n29207), .C0(index_q[0]), .Z(n29208));
    LUT4 mux_192_Mux_3_i1018_3_lut_4_lut (.A(index_q[1]), .B(n26585), .C(index_q[4]), 
         .D(n19590), .Z(n1018)) /* synthesis lut_function=(A (C+!(D))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_3_i1018_3_lut_4_lut.init = 16'he0ef;
    LUT4 mux_192_Mux_1_i924_3_lut (.A(n316), .B(n923_adj_2544), .C(index_q[4]), 
         .Z(n924_adj_2545)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_1_i924_3_lut.init = 16'hcaca;
    LUT4 i11478_3_lut_4_lut (.A(n26547), .B(index_i[4]), .C(index_i[5]), 
         .D(n26647), .Z(n892_adj_2546)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11478_3_lut_4_lut.init = 16'hf8f0;
    LUT4 i20493_3_lut_3_lut_4_lut (.A(n26486), .B(index_i[3]), .C(n93_adj_2547), 
         .D(index_i[4]), .Z(n22832)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20493_3_lut_3_lut_4_lut.init = 16'hf077;
    LUT4 n254_bdd_4_lut (.A(index_q[5]), .B(index_q[3]), .C(index_q[6]), 
         .D(index_q[4]), .Z(n25806)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;
    defparam n254_bdd_4_lut.init = 16'hf8f0;
    LUT4 n404_bdd_3_lut_23498 (.A(index_i[3]), .B(n26702), .C(n26710), 
         .Z(n24637)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam n404_bdd_3_lut_23498.init = 16'he4e4;
    LUT4 mux_191_Mux_6_i251_3_lut_4_lut (.A(n26694), .B(index_i[2]), .C(index_i[3]), 
         .D(n26703), .Z(n251_adj_2548)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_6_i251_3_lut_4_lut.init = 16'hf606;
    LUT4 i9527_3_lut_4_lut (.A(n26694), .B(index_i[2]), .C(n26635), .D(n26703), 
         .Z(n444_adj_2486)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9527_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_191_Mux_4_i747_3_lut_4_lut (.A(n26694), .B(index_i[2]), .C(index_i[3]), 
         .D(n26706), .Z(n747_adj_2401)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_4_i747_3_lut_4_lut.init = 16'hf606;
    PFUMX i20039 (.BLUT(n669_adj_2549), .ALUT(n700_adj_2550), .C0(index_i[5]), 
          .Z(n22378));
    LUT4 n404_bdd_3_lut_23005 (.A(n404), .B(n26688), .C(index_i[3]), .Z(n24636)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n404_bdd_3_lut_23005.init = 16'hcaca;
    LUT4 index_q_6__bdd_4_lut_25923 (.A(index_q[6]), .B(index_q[5]), .C(index_q[1]), 
         .D(index_q[0]), .Z(n28701)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C))+!A (B (C)+!B !(C)))) */ ;
    defparam index_q_6__bdd_4_lut_25923.init = 16'h3cbc;
    LUT4 i20492_3_lut_4_lut (.A(n26486), .B(index_i[3]), .C(index_i[4]), 
         .D(n46_adj_2551), .Z(n22831)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20492_3_lut_4_lut.init = 16'h8f80;
    PFUMX i20040 (.BLUT(n21619), .ALUT(n763_adj_2402), .C0(index_i[5]), 
          .Z(n22379));
    LUT4 mux_191_Mux_3_i221_3_lut_4_lut (.A(n26486), .B(index_i[3]), .C(index_i[4]), 
         .D(n26437), .Z(n221_adj_2552)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_3_i221_3_lut_4_lut.init = 16'h08f8;
    LUT4 i21438_3_lut (.A(n21818), .B(n21819), .C(index_q[4]), .Z(n21820)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21438_3_lut.init = 16'hcaca;
    LUT4 index_q_5__bdd_3_lut (.A(index_q[5]), .B(n28702), .C(index_q[3]), 
         .Z(n28703)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam index_q_5__bdd_3_lut.init = 16'hcaca;
    LUT4 index_q_6__bdd_1_lut (.A(index_q[5]), .Z(n28700)) /* synthesis lut_function=(!(A)) */ ;
    defparam index_q_6__bdd_1_lut.init = 16'h5555;
    PFUMX i20041 (.BLUT(n21622), .ALUT(n828_adj_2553), .C0(index_i[5]), 
          .Z(n22380));
    LUT4 n470_bdd_3_lut (.A(n29177), .B(n29178), .C(index_i[3]), .Z(n24640)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n470_bdd_3_lut.init = 16'hacac;
    PFUMX i20042 (.BLUT(n860_adj_2554), .ALUT(n21625), .C0(index_i[5]), 
          .Z(n22381));
    LUT4 n26569_bdd_3_lut_26031 (.A(n26430), .B(index_q[6]), .C(index_q[5]), 
         .Z(n28704)) /* synthesis lut_function=(!(A (B)+!A (C))) */ ;
    defparam n26569_bdd_3_lut_26031.init = 16'h2727;
    LUT4 n26569_bdd_4_lut (.A(n26569), .B(index_q[6]), .C(index_q[2]), 
         .D(index_q[5]), .Z(n28705)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A !(B (C+(D))+!B (D)))) */ ;
    defparam n26569_bdd_4_lut.init = 16'h5fe0;
    LUT4 n28706_bdd_3_lut (.A(n28706), .B(n28703), .C(index_q[4]), .Z(n28707)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n28706_bdd_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_1_i349_3_lut (.A(n541_adj_2288), .B(n348_adj_2555), 
         .C(index_q[4]), .Z(n349_adj_2556)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_1_i349_3_lut.init = 16'hcaca;
    PFUMX mux_192_Mux_8_i764 (.BLUT(n716_adj_2287), .ALUT(n732_adj_2557), 
          .C0(n22040), .Z(n764)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 i21448_3_lut (.A(n21782), .B(n21783), .C(index_q[4]), .Z(n21784)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21448_3_lut.init = 16'hcaca;
    LUT4 i20633_3_lut_4_lut_4_lut (.A(n26455), .B(index_i[4]), .C(index_i[5]), 
         .D(n26470), .Z(n22972)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C)+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20633_3_lut_4_lut_4_lut.init = 16'h0434;
    LUT4 mux_191_Mux_8_i892_3_lut_4_lut (.A(n26455), .B(index_i[4]), .C(index_i[5]), 
         .D(n860_adj_2290), .Z(n892_adj_2558)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_8_i892_3_lut_4_lut.init = 16'h4f40;
    LUT4 index_i_6__bdd_4_lut_25972 (.A(index_i[6]), .B(index_i[5]), .C(index_i[1]), 
         .D(index_i[0]), .Z(n28762)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C))+!A (B (C)+!B !(C)))) */ ;
    defparam index_i_6__bdd_4_lut_25972.init = 16'h3cbc;
    LUT4 index_i_6__bdd_1_lut (.A(index_i[5]), .Z(n28761)) /* synthesis lut_function=(!(A)) */ ;
    defparam index_i_6__bdd_1_lut.init = 16'h5555;
    LUT4 index_i_5__bdd_3_lut (.A(index_i[5]), .B(n28763), .C(index_i[3]), 
         .Z(n28764)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam index_i_5__bdd_3_lut.init = 16'hcaca;
    LUT4 n26647_bdd_3_lut (.A(n26438), .B(index_i[6]), .C(index_i[5]), 
         .Z(n28765)) /* synthesis lut_function=(!(A (B)+!A (C))) */ ;
    defparam n26647_bdd_3_lut.init = 16'h2727;
    PFUMX i20061 (.BLUT(n94_adj_2559), .ALUT(n125_adj_2560), .C0(index_i[5]), 
          .Z(n22400));
    LUT4 n26647_bdd_4_lut (.A(n26647), .B(index_i[6]), .C(index_i[2]), 
         .D(index_i[5]), .Z(n28766)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A !(B (C+(D))+!B (D)))) */ ;
    defparam n26647_bdd_4_lut.init = 16'h5fe0;
    LUT4 mux_192_Mux_1_i94_3_lut (.A(index_q[0]), .B(n93_adj_2460), .C(index_q[4]), 
         .Z(n94_adj_2561)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_1_i94_3_lut.init = 16'hcaca;
    LUT4 i21570_3_lut (.A(n620_adj_2364), .B(n14450), .C(index_q[4]), 
         .Z(n21381)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21570_3_lut.init = 16'hcaca;
    LUT4 n25811_bdd_3_lut (.A(n26825), .B(n25807), .C(index_q[7]), .Z(n25812)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n25811_bdd_3_lut.init = 16'hcaca;
    LUT4 n28767_bdd_3_lut (.A(n28767), .B(n28764), .C(index_i[4]), .Z(n28768)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n28767_bdd_3_lut.init = 16'hcaca;
    PFUMX i20062 (.BLUT(n158_adj_2562), .ALUT(n189_adj_2295), .C0(index_i[5]), 
          .Z(n22401));
    LUT4 i9470_3_lut (.A(n11915), .B(n29170), .C(index_q[3]), .Z(n11916)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9470_3_lut.init = 16'hcaca;
    PFUMX i20063 (.BLUT(n221_adj_2552), .ALUT(n252_adj_2294), .C0(index_i[5]), 
          .Z(n22402));
    LUT4 mux_192_Mux_7_i892_3_lut (.A(n62_adj_2377), .B(n891_adj_2257), 
         .C(index_q[5]), .Z(n892_adj_2343)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_7_i892_3_lut.init = 16'hcaca;
    LUT4 i19238_3_lut (.A(n747_adj_2310), .B(n908_adj_2563), .C(index_q[4]), 
         .Z(n21558)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19238_3_lut.init = 16'hcaca;
    LUT4 i19237_3_lut (.A(n716_adj_2358), .B(n14848), .C(index_q[4]), 
         .Z(n21557)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19237_3_lut.init = 16'hcaca;
    PFUMX i20064 (.BLUT(n286_adj_2564), .ALUT(n21634), .C0(index_i[5]), 
          .Z(n22403));
    LUT4 n254_bdd_4_lut_adj_76 (.A(index_i[5]), .B(index_i[3]), .C(index_i[6]), 
         .D(index_i[4]), .Z(n25822)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;
    defparam n254_bdd_4_lut_adj_76.init = 16'hf8f0;
    PFUMX i20065 (.BLUT(n349_adj_2565), .ALUT(n21637), .C0(index_i[5]), 
          .Z(n22404));
    PFUMX i19293 (.BLUT(n21611), .ALUT(n21612), .C0(index_i[4]), .Z(n476_adj_2408));
    PFUMX i20066 (.BLUT(n413_adj_2566), .ALUT(n444_adj_2567), .C0(index_i[5]), 
          .Z(n22405));
    LUT4 mux_191_Mux_2_i700_3_lut_4_lut (.A(index_i[1]), .B(n26601), .C(index_i[4]), 
         .D(n684_adj_2407), .Z(n700_adj_2568)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_2_i700_3_lut_4_lut.init = 16'hefe0;
    LUT4 mux_192_Mux_10_i701_4_lut_4_lut (.A(n26429), .B(index_q[4]), .C(index_q[5]), 
         .D(n26384), .Z(n701_adj_2569)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B (C (D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_10_i701_4_lut_4_lut.init = 16'h3efe;
    PFUMX i20067 (.BLUT(n476_adj_2570), .ALUT(n507_adj_2298), .C0(index_i[5]), 
          .Z(n22406));
    LUT4 mux_192_Mux_6_i891_3_lut (.A(n875_adj_2571), .B(n890_adj_2324), 
         .C(index_q[4]), .Z(n891_adj_2572)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_6_i891_3_lut.init = 16'hcaca;
    LUT4 n25827_bdd_3_lut (.A(n26822), .B(n25823), .C(index_i[7]), .Z(n25828)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n25827_bdd_3_lut.init = 16'hcaca;
    LUT4 mux_191_Mux_3_i1018_3_lut_4_lut (.A(index_i[1]), .B(n26601), .C(index_i[4]), 
         .D(n19612), .Z(n1018_adj_2573)) /* synthesis lut_function=(A (C+!(D))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_3_i1018_3_lut_4_lut.init = 16'he0ef;
    PFUMX i20507 (.BLUT(n22830), .ALUT(n22831), .C0(index_i[5]), .Z(n22846));
    LUT4 mux_192_Mux_6_i828_4_lut (.A(n812_adj_2574), .B(n13827), .C(index_q[4]), 
         .D(index_q[2]), .Z(n828_adj_2575)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_6_i828_4_lut.init = 16'hfaca;
    PFUMX i20068 (.BLUT(n21640), .ALUT(n573_adj_2433), .C0(index_i[5]), 
          .Z(n22407));
    LUT4 mux_192_Mux_6_i797_3_lut (.A(n781_adj_2303), .B(n26356), .C(index_q[4]), 
         .Z(n797_adj_2576)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_6_i797_3_lut.init = 16'hcaca;
    PFUMX i20069 (.BLUT(n11991), .ALUT(n21643), .C0(index_i[5]), .Z(n22408));
    PFUMX i20070 (.BLUT(n669_adj_2577), .ALUT(n700_adj_2578), .C0(index_i[5]), 
          .Z(n22409));
    PFUMX i20508 (.BLUT(n22832), .ALUT(n22833), .C0(index_i[5]), .Z(n22847));
    LUT4 mux_191_Mux_8_i124_3_lut_3_lut_4_lut (.A(n26548), .B(index_i[2]), 
         .C(n26649), .D(index_i[3]), .Z(n124_adj_2387)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_8_i124_3_lut_3_lut_4_lut.init = 16'h11f0;
    LUT4 mux_192_Mux_6_i669_3_lut (.A(n653_adj_2514), .B(n668_adj_2579), 
         .C(index_q[4]), .Z(n669_adj_2580)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_6_i669_3_lut.init = 16'hcaca;
    CCU2D add_371_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(quarter_wave_sample_register_i[0]), .B1(quarter_wave_sample_register_i[1]), 
          .C1(GND_net), .D1(GND_net), .COUT(n17346));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam add_371_1.INIT0 = 16'hF000;
    defparam add_371_1.INIT1 = 16'ha666;
    defparam add_371_1.INJECT1_0 = "NO";
    defparam add_371_1.INJECT1_1 = "NO";
    L6MUX21 i20071 (.D0(n21646), .D1(n763), .SD(index_i[5]), .Z(n22410));
    L6MUX21 i20509 (.D0(n22834), .D1(n22835), .SD(index_i[5]), .Z(n22848));
    PFUMX i20073 (.BLUT(n860_adj_2581), .ALUT(n891_adj_2582), .C0(index_i[5]), 
          .Z(n22412));
    LUT4 mux_192_Mux_6_i542_3_lut (.A(n812_adj_2583), .B(n541), .C(index_q[4]), 
         .Z(n542_adj_2584)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_6_i542_3_lut.init = 16'hcaca;
    LUT4 n21206_bdd_3_lut (.A(n26352), .B(n701), .C(index_i[6]), .Z(n25853)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n21206_bdd_3_lut.init = 16'hacac;
    LUT4 index_q_4__bdd_4_lut_22960 (.A(index_q[4]), .B(n26429), .C(index_q[7]), 
         .D(n26477), .Z(n24286)) /* synthesis lut_function=(A (C+!(D))+!A (B+!(C))) */ ;
    defparam index_q_4__bdd_4_lut_22960.init = 16'he5ef;
    LUT4 mux_192_Mux_2_i955_then_4_lut (.A(index_q[4]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n26800)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B (C+!(D))+!B !(C (D)))) */ ;
    defparam mux_192_Mux_2_i955_then_4_lut.init = 16'he95d;
    LUT4 mux_192_Mux_6_i252_4_lut (.A(index_q[2]), .B(n251_adj_2398), .C(index_q[4]), 
         .D(n11010), .Z(n252_adj_2585)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_6_i252_4_lut.init = 16'hc5ca;
    LUT4 i21921_3_lut (.A(n25554), .B(n252_adj_2585), .C(index_q[5]), 
         .Z(n22112)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21921_3_lut.init = 16'hcaca;
    PFUMX mux_192_Mux_8_i574 (.BLUT(n542_adj_2371), .ALUT(n12017), .C0(index_q[5]), 
          .Z(n574)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 n25856_bdd_3_lut (.A(n28182), .B(n22975), .C(index_i[8]), .Z(n25857)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n25856_bdd_3_lut.init = 16'hcaca;
    LUT4 i19468_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21788)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (D))+!A !(B (C (D))+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19468_3_lut_3_lut_4_lut.init = 16'h4933;
    L6MUX21 i24337 (.D0(n26183), .D1(n26180), .SD(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_2142[4]));
    LUT4 mux_192_Mux_2_i955_else_4_lut (.A(index_q[4]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n26799)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+(D)))+!A !(B (C+!(D))+!B !(C+!(D))))) */ ;
    defparam mux_192_Mux_2_i955_else_4_lut.init = 16'h49c6;
    LUT4 i19223_3_lut (.A(n93_adj_2368), .B(n699), .C(index_q[4]), .Z(n21543)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19223_3_lut.init = 16'hcaca;
    LUT4 i19222_3_lut (.A(n653_adj_2456), .B(n26387), .C(index_q[4]), 
         .Z(n21542)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19222_3_lut.init = 16'hcaca;
    PFUMX i24335 (.BLUT(n26182), .ALUT(n26181), .C0(index_q[8]), .Z(n26183));
    CCU2D add_372_15 (.A0(quarter_wave_sample_register_q[14]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(\quarter_wave_sample_register_q[15] ), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17344), .S0(o_val_pipeline_q_0__15__N_2190[14]), 
          .S1(o_val_pipeline_q_0__15__N_2190[15]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(80[29:60])
    defparam add_372_15.INIT0 = 16'hf555;
    defparam add_372_15.INIT1 = 16'hf555;
    defparam add_372_15.INJECT1_0 = "NO";
    defparam add_372_15.INJECT1_1 = "NO";
    PFUMX i20074 (.BLUT(n924_adj_2586), .ALUT(n21649), .C0(index_i[5]), 
          .Z(n22413));
    LUT4 i19070_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21390)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C+(D)))+!A (B (C)+!B !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19070_3_lut_4_lut_4_lut.init = 16'hc95a;
    PFUMX i20075 (.BLUT(n21652), .ALUT(n1018_adj_2573), .C0(index_i[5]), 
          .Z(n22414));
    LUT4 mux_191_Mux_9_i124_3_lut_4_lut (.A(n26548), .B(index_i[2]), .C(index_i[3]), 
         .D(n26505), .Z(n124_adj_2425)) /* synthesis lut_function=(!(A (C+!(D))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_9_i124_3_lut_4_lut.init = 16'h1f10;
    LUT4 mux_191_Mux_3_i93_3_lut_4_lut (.A(n26548), .B(index_i[2]), .C(index_i[3]), 
         .D(n70_adj_2255), .Z(n93_adj_2587)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_3_i93_3_lut_4_lut.init = 16'hefe0;
    L6MUX21 i20512 (.D0(n22840), .D1(n22841), .SD(index_i[5]), .Z(n22851));
    L6MUX21 i20513 (.D0(n22842), .D1(n22843), .SD(index_i[5]), .Z(n22852));
    CCU2D add_372_13 (.A0(quarter_wave_sample_register_q[12]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_q[13]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17343), .COUT(n17344), 
          .S0(o_val_pipeline_q_0__15__N_2190[12]), .S1(o_val_pipeline_q_0__15__N_2190[13]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(80[29:60])
    defparam add_372_13.INIT0 = 16'hf555;
    defparam add_372_13.INIT1 = 16'hf555;
    defparam add_372_13.INJECT1_0 = "NO";
    defparam add_372_13.INJECT1_1 = "NO";
    L6MUX21 i20514 (.D0(n22844), .D1(n22845), .SD(index_i[5]), .Z(n22853));
    LUT4 mux_191_Mux_8_i475_3_lut_4_lut (.A(n26548), .B(index_i[2]), .C(index_i[3]), 
         .D(n26505), .Z(n475_adj_2588)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_8_i475_3_lut_4_lut.init = 16'hf101;
    LUT4 mux_191_Mux_0_i1002_3_lut_3_lut_4_lut (.A(n26548), .B(index_i[2]), 
         .C(n38), .D(index_i[3]), .Z(n1002_adj_2589)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_0_i1002_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 n21215_bdd_3_lut (.A(n26353), .B(n701_adj_2569), .C(index_q[6]), 
         .Z(n25863)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n21215_bdd_3_lut.init = 16'hacac;
    LUT4 mux_191_Mux_6_i890_3_lut_4_lut (.A(n26548), .B(index_i[2]), .C(index_i[3]), 
         .D(n26653), .Z(n890_adj_2590)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_6_i890_3_lut_4_lut.init = 16'hf101;
    LUT4 mux_191_Mux_8_i732_3_lut (.A(index_i[3]), .B(n15024), .C(index_i[5]), 
         .Z(n732_adj_2591)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_8_i732_3_lut.init = 16'h3a3a;
    CCU2D add_372_11 (.A0(quarter_wave_sample_register_q[10]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_q[11]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17342), .COUT(n17343), 
          .S0(o_val_pipeline_q_0__15__N_2190[10]), .S1(o_val_pipeline_q_0__15__N_2190[11]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(80[29:60])
    defparam add_372_11.INIT0 = 16'hf555;
    defparam add_372_11.INIT1 = 16'hf555;
    defparam add_372_11.INJECT1_0 = "NO";
    defparam add_372_11.INJECT1_1 = "NO";
    LUT4 n20976_bdd_3_lut_23417_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n25071)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C))+!A !(B (C+!(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n20976_bdd_3_lut_23417_4_lut_4_lut.init = 16'h5ad6;
    PFUMX i20093 (.BLUT(n158_adj_2592), .ALUT(n189_adj_2536), .C0(index_i[5]), 
          .Z(n22432));
    LUT4 n25866_bdd_3_lut (.A(n28123), .B(n22822), .C(index_q[8]), .Z(n25867)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n25866_bdd_3_lut.init = 16'hcaca;
    PFUMX i19311 (.BLUT(n21629), .ALUT(n21630), .C0(index_i[4]), .Z(n21631));
    PFUMX i24510 (.BLUT(n26811), .ALUT(n26812), .C0(index_i[1]), .Z(n26813));
    PFUMX i24332 (.BLUT(n26179), .ALUT(n22265), .C0(index_q[8]), .Z(n26180));
    PFUMX i20094 (.BLUT(n221_adj_2593), .ALUT(n21658), .C0(index_i[5]), 
          .Z(n22433));
    LUT4 i21497_3_lut (.A(n21524), .B(n21525), .C(index_i[4]), .Z(n21526)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i21497_3_lut.init = 16'hcaca;
    PFUMX i20095 (.BLUT(n286_adj_2594), .ALUT(n317_adj_2595), .C0(index_i[5]), 
          .Z(n22434));
    LUT4 i15393_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[2]), 
         .C(index_q[3]), .D(index_q[1]), .Z(n17543)) /* synthesis lut_function=(A (B (C (D))+!B !(C))+!A (B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i15393_3_lut_4_lut_4_lut_4_lut.init = 16'hd656;
    PFUMX i20096 (.BLUT(n349_adj_2596), .ALUT(n21661), .C0(index_i[5]), 
          .Z(n22435));
    LUT4 i20486_4_lut_4_lut (.A(n26410), .B(n26497), .C(index_q[5]), .D(index_q[4]), 
         .Z(n22825)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C+(D))+!B !(C (D)+!C !(D)))) */ ;
    defparam i20486_4_lut_4_lut.init = 16'hcf50;
    LUT4 mux_191_Mux_6_i60_3_lut_4_lut_4_lut_3_lut_rep_741 (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[2]), .Z(n26701)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_6_i60_3_lut_4_lut_4_lut_3_lut_rep_741.init = 16'hd6d6;
    PFUMX mux_192_Mux_2_i891 (.BLUT(n875_adj_2597), .ALUT(n890_adj_2280), 
          .C0(index_q[4]), .Z(n891_adj_2598)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 mux_191_Mux_7_i262_3_lut_rep_795 (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .Z(n29174)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_7_i262_3_lut_rep_795.init = 16'h6464;
    PFUMX i20097 (.BLUT(n413_adj_2599), .ALUT(n21664), .C0(index_i[5]), 
          .Z(n22436));
    LUT4 mux_192_Mux_5_i124_3_lut (.A(n26521), .B(n26570), .C(index_q[3]), 
         .Z(n124_adj_2512)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_5_i124_3_lut.init = 16'hcaca;
    PFUMX i18975 (.BLUT(n21293), .ALUT(n21294), .C0(index_i[5]), .Z(n21295));
    LUT4 index_i_7__bdd_4_lut_24661 (.A(index_i[7]), .B(n15074), .C(n24245), 
         .D(index_i[5]), .Z(n26340)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(B (C+(D))+!B !((D)+!C)))) */ ;
    defparam index_i_7__bdd_4_lut_24661.init = 16'h66f0;
    LUT4 i19271_3_lut_4_lut (.A(n26594), .B(index_i[2]), .C(index_i[3]), 
         .D(n26706), .Z(n21591)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19271_3_lut_4_lut.init = 16'h6f60;
    LUT4 index_i_0__bdd_4_lut_24505 (.A(index_i[0]), .B(index_i[3]), .C(index_i[1]), 
         .D(index_i[2]), .Z(n26802)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C))+!A (B (C (D)+!C !(D))+!B !(C+!(D))))) */ ;
    defparam index_i_0__bdd_4_lut_24505.init = 16'h16d3;
    LUT4 i15441_4_lut (.A(index_i[0]), .B(index_i[4]), .C(index_i[1]), 
         .D(n26601), .Z(n286_adj_2600)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i15441_4_lut.init = 16'hccc8;
    PFUMX i18978 (.BLUT(n21296), .ALUT(n21297), .C0(index_i[5]), .Z(n21298));
    LUT4 mux_191_Mux_3_i460_3_lut_4_lut (.A(n26594), .B(index_i[2]), .C(index_i[3]), 
         .D(n26709), .Z(n460_adj_2601)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_3_i460_3_lut_4_lut.init = 16'h6f60;
    PFUMX mux_192_Mux_2_i860 (.BLUT(n844_adj_2282), .ALUT(n859_adj_2602), 
          .C0(index_q[4]), .Z(n860_adj_2603)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 i21520_3_lut (.A(n716), .B(n731_adj_2604), .C(index_q[4]), .Z(n732_adj_2605)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21520_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_2_i669_3_lut (.A(n653_adj_2606), .B(n24916), .C(index_q[4]), 
         .Z(n669_adj_2607)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_2_i669_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_2_i605_3_lut (.A(n142_adj_2451), .B(n604_adj_2447), 
         .C(index_q[4]), .Z(n605_adj_2608)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_2_i605_3_lut.init = 16'hcaca;
    LUT4 i20622_3_lut_4_lut (.A(n26407), .B(n26394), .C(index_i[5]), .D(index_i[6]), 
         .Z(n22961)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (B+((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20622_3_lut_4_lut.init = 16'hffc5;
    LUT4 i21525_3_lut (.A(n26774), .B(n21114), .C(index_q[4]), .Z(n21115)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21525_3_lut.init = 16'hcaca;
    LUT4 i19968_3_lut_4_lut (.A(n26408), .B(n26386), .C(index_q[5]), .D(index_q[6]), 
         .Z(n22307)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (B+((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19968_3_lut_4_lut.init = 16'hffc5;
    PFUMX i20098 (.BLUT(n21667), .ALUT(n507_adj_2609), .C0(index_i[5]), 
          .Z(n22437));
    LUT4 i21528_3_lut (.A(n21110), .B(n21111), .C(index_q[4]), .Z(n21112)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21528_3_lut.init = 16'hcaca;
    PFUMX i24321 (.BLUT(n26166), .ALUT(n29200), .C0(index_q[3]), .Z(n26167));
    LUT4 mux_192_Mux_2_i413_3_lut (.A(n397_adj_2259), .B(n954_adj_2429), 
         .C(index_q[4]), .Z(n413_adj_2610)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_2_i413_3_lut.init = 16'hcaca;
    LUT4 i19358_3_lut_4_lut (.A(n26594), .B(index_i[2]), .C(index_i[3]), 
         .D(n26687), .Z(n21678)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19358_3_lut_4_lut.init = 16'hf606;
    LUT4 n22384_bdd_3_lut_24128 (.A(n22386), .B(n24495), .C(index_i[7]), 
         .Z(n25914)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n22384_bdd_3_lut_24128.init = 16'hcaca;
    LUT4 n187_bdd_4_lut_23712 (.A(n26486), .B(index_i[6]), .C(index_i[5]), 
         .D(n26605), .Z(n24760)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(D))+!A !(B (C+(D))+!B (D)))) */ ;
    defparam n187_bdd_4_lut_23712.init = 16'h7f40;
    LUT4 index_i_0__bdd_4_lut_24532 (.A(index_i[0]), .B(index_i[3]), .C(index_i[1]), 
         .D(index_i[2]), .Z(n26803)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C (D)))+!A !(B (C+!(D))+!B !(C+(D))))) */ ;
    defparam index_i_0__bdd_4_lut_24532.init = 16'h4ae7;
    PFUMX i20099 (.BLUT(n21670), .ALUT(n573_adj_2421), .C0(index_i[5]), 
          .Z(n22438));
    LUT4 mux_192_Mux_2_i317_3_lut (.A(n668), .B(n316_adj_2258), .C(index_q[4]), 
         .Z(n317_adj_2611)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_2_i317_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_2_i286_3_lut (.A(n270), .B(n653), .C(index_q[4]), 
         .Z(n286_adj_2612)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_2_i286_3_lut.init = 16'hcaca;
    LUT4 i20466_3_lut (.A(n26728), .B(n29189), .C(index_q[3]), .Z(n22805)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20466_3_lut.init = 16'hcaca;
    LUT4 i20465_3_lut (.A(n29181), .B(n660), .C(index_q[3]), .Z(n22804)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20465_3_lut.init = 16'hcaca;
    LUT4 i20464_3_lut (.A(n676), .B(n26571), .C(index_q[3]), .Z(n22803)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20464_3_lut.init = 16'hcaca;
    PFUMX i20100 (.BLUT(n605_adj_2613), .ALUT(n21673), .C0(index_i[5]), 
          .Z(n22439));
    LUT4 i20463_3_lut (.A(n26521), .B(n26719), .C(index_q[3]), .Z(n22802)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20463_3_lut.init = 16'hcaca;
    LUT4 i18698_3_lut (.A(n26570), .B(n29200), .C(index_q[3]), .Z(n21018)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18698_3_lut.init = 16'hcaca;
    LUT4 i21540_3_lut (.A(n142), .B(n13863), .C(index_q[4]), .Z(n158_adj_2614)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21540_3_lut.init = 16'hcaca;
    LUT4 i21374_3_lut (.A(n21017), .B(n21018), .C(index_q[4]), .Z(n21019)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21374_3_lut.init = 16'hcaca;
    LUT4 i20459_3_lut (.A(n29189), .B(n29183), .C(index_q[3]), .Z(n22798)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20459_3_lut.init = 16'hcaca;
    LUT4 i20458_3_lut (.A(n1001), .B(n26728), .C(index_q[3]), .Z(n22797)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20458_3_lut.init = 16'hcaca;
    LUT4 n22395_bdd_3_lut (.A(n22388), .B(n22389), .C(index_i[7]), .Z(n25912)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n22395_bdd_3_lut.init = 16'hcaca;
    PFUMX i20101 (.BLUT(n669_adj_2615), .ALUT(n700_adj_2568), .C0(index_i[5]), 
          .Z(n22440));
    LUT4 i20456_3_lut (.A(n29183), .B(n26521), .C(index_q[3]), .Z(n22795)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20456_3_lut.init = 16'hcaca;
    PFUMX i20102 (.BLUT(n732_adj_2616), .ALUT(n763_adj_2617), .C0(index_i[5]), 
          .Z(n22441));
    LUT4 n22384_bdd_3_lut (.A(n22384), .B(n22385), .C(index_i[7]), .Z(n25915)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n22384_bdd_3_lut.init = 16'hcaca;
    LUT4 i20267_3_lut (.A(n94_adj_2618), .B(n476_adj_2619), .C(index_q[5]), 
         .Z(n22606)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20267_3_lut.init = 16'hcaca;
    LUT4 n24763_bdd_3_lut (.A(n26813), .B(n24760), .C(index_i[4]), .Z(n24764)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n24763_bdd_3_lut.init = 16'hcaca;
    L6MUX21 i20104 (.D0(n860_adj_2268), .D1(n891_adj_2266), .SD(index_i[5]), 
            .Z(n22443));
    LUT4 i19412_3_lut (.A(n29187), .B(n250), .C(index_q[3]), .Z(n21732)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19412_3_lut.init = 16'hcaca;
    LUT4 n22942_bdd_3_lut (.A(n24599), .B(n22928), .C(index_i[6]), .Z(n25930)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n22942_bdd_3_lut.init = 16'hcaca;
    LUT4 n24950_bdd_3_lut_24141 (.A(n28283), .B(n25339), .C(index_i[6]), 
         .Z(n25932)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n24950_bdd_3_lut_24141.init = 16'hcaca;
    LUT4 i19411_3_lut (.A(n26719), .B(n29182), .C(index_q[3]), .Z(n21731)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19411_3_lut.init = 16'hcaca;
    LUT4 index_i_1__bdd_4_lut_25024 (.A(index_i[1]), .B(index_i[0]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n26804)) /* synthesis lut_function=(!(A (B (D)+!B (C+!(D)))+!A !(B (C (D)+!C !(D))+!B !((D)+!C)))) */ ;
    defparam index_i_1__bdd_4_lut_25024.init = 16'h429c;
    PFUMX i19326 (.BLUT(n21644), .ALUT(n21645), .C0(index_i[4]), .Z(n21646));
    LUT4 i19409_3_lut (.A(n29187), .B(n26521), .C(index_q[3]), .Z(n21729)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19409_3_lut.init = 16'hcaca;
    LUT4 index_q_3__bdd_3_lut_22632_3_lut_4_lut (.A(n26623), .B(index_q[1]), 
         .C(index_q[4]), .D(index_q[3]), .Z(n24165)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam index_q_3__bdd_3_lut_22632_3_lut_4_lut.init = 16'hf10f;
    LUT4 i9571_4_lut_4_lut (.A(n26623), .B(index_q[1]), .C(index_q[3]), 
         .D(n20372), .Z(n12017)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A (B (C)+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9571_4_lut_4_lut.init = 16'h0e3e;
    LUT4 i19408_3_lut (.A(n29183), .B(n250), .C(index_q[3]), .Z(n21728)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19408_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_7_i173_3_lut (.A(n26719), .B(n26521), .C(index_q[3]), 
         .Z(n173_adj_2508)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_7_i173_3_lut.init = 16'hcaca;
    LUT4 n24950_bdd_3_lut (.A(n24950), .B(n22924), .C(index_i[6]), .Z(n25933)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n24950_bdd_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_6_i70_3_lut_rep_797 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29176)) /* synthesis lut_function=(!(A (B+(C))+!A !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_6_i70_3_lut_rep_797.init = 16'h5252;
    LUT4 mux_191_Mux_6_i285_3_lut_4_lut (.A(n26594), .B(index_i[2]), .C(index_i[3]), 
         .D(n26699), .Z(n285_adj_2620)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_6_i285_3_lut_4_lut.init = 16'hf606;
    LUT4 i18756_then_4_lut (.A(index_q[0]), .B(index_q[4]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n26744)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C))+!A (B (C)+!B !(C+!(D)))) */ ;
    defparam i18756_then_4_lut.init = 16'hc34a;
    LUT4 mux_192_Mux_7_i956_3_lut_3_lut_4_lut (.A(n26429), .B(index_q[4]), 
         .C(n924_adj_2621), .D(index_q[5]), .Z(n956_adj_2622)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_7_i956_3_lut_3_lut_4_lut.init = 16'h11f0;
    LUT4 i18756_else_4_lut (.A(index_q[0]), .B(index_q[4]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n26743)) /* synthesis lut_function=(A (C)+!A !(B ((D)+!C)+!B !(C))) */ ;
    defparam i18756_else_4_lut.init = 16'hb0f0;
    LUT4 n24766_bdd_3_lut (.A(n24766), .B(n24764), .C(index_i[3]), .Z(n24767)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n24766_bdd_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_0_i572_3_lut_4_lut (.A(n26623), .B(index_q[1]), .C(index_q[3]), 
         .D(n29198), .Z(n572_adj_2417)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_0_i572_3_lut_4_lut.init = 16'hefe0;
    LUT4 i11482_2_lut_rep_389_3_lut_4_lut (.A(n26410), .B(index_q[4]), .C(index_q[6]), 
         .D(index_q[5]), .Z(n26349)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11482_2_lut_rep_389_3_lut_4_lut.init = 16'hf080;
    LUT4 mux_192_Mux_4_i158_3_lut (.A(n142_adj_2623), .B(n157_adj_2342), 
         .C(index_q[4]), .Z(n158_adj_2624)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_4_i158_3_lut.init = 16'hcaca;
    LUT4 i19405_3_lut (.A(n26592), .B(n26708), .C(index_i[3]), .Z(n21725)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19405_3_lut.init = 16'hcaca;
    LUT4 i21641_3_lut (.A(n21725), .B(n21726), .C(index_i[4]), .Z(n21727)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21641_3_lut.init = 16'hcaca;
    LUT4 i19402_3_lut (.A(n38), .B(n773), .C(index_i[3]), .Z(n21722)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19402_3_lut.init = 16'hcaca;
    LUT4 i12426_2_lut_3_lut_4_lut (.A(n26411), .B(index_q[4]), .C(index_q[6]), 
         .D(index_q[5]), .Z(n15006)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12426_2_lut_3_lut_4_lut.init = 16'hfef0;
    LUT4 i21643_3_lut (.A(n21722), .B(n21723), .C(index_i[4]), .Z(n21724)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21643_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_9_i364_3_lut_3_lut_4_lut (.A(n26623), .B(index_q[1]), 
         .C(index_q[3]), .D(n26526), .Z(n364_adj_2281)) /* synthesis lut_function=(!(A (C (D))+!A (B (C (D))+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_9_i364_3_lut_3_lut_4_lut.init = 16'h0efe;
    PFUMX i24467 (.BLUT(n26743), .ALUT(n26744), .C0(index_q[1]), .Z(n26745));
    LUT4 mux_192_Mux_5_i262_rep_583 (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .Z(n26543)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_5_i262_rep_583.init = 16'h6464;
    PFUMX i18987 (.BLUT(n21305), .ALUT(n21306), .C0(index_i[5]), .Z(n21307));
    PFUMX mux_192_Mux_3_i763 (.BLUT(n747_adj_2625), .ALUT(n762_adj_2626), 
          .C0(index_q[4]), .Z(n763_adj_2474)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    PFUMX i18990 (.BLUT(n21308), .ALUT(n21309), .C0(index_i[5]), .Z(n21310));
    PFUMX i20123 (.BLUT(n94_adj_2627), .ALUT(n21679), .C0(index_i[5]), 
          .Z(n22462));
    LUT4 i11280_3_lut (.A(index_q[3]), .B(index_q[1]), .C(index_q[0]), 
         .Z(n13839)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11280_3_lut.init = 16'hecec;
    LUT4 mux_192_Mux_6_i22_rep_584 (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .Z(n26544)) /* synthesis lut_function=(!(A (C)+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_6_i22_rep_584.init = 16'h4a4a;
    L6MUX21 i20124 (.D0(n21682), .D1(n21685), .SD(index_i[5]), .Z(n22463));
    LUT4 mux_192_Mux_3_i251_3_lut_4_lut (.A(n26623), .B(index_q[1]), .C(index_q[3]), 
         .D(n26526), .Z(n14728)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_3_i251_3_lut_4_lut.init = 16'hfe0e;
    LUT4 mux_191_Mux_0_i986_3_lut (.A(n26702), .B(n985_adj_2628), .C(index_i[3]), 
         .Z(n986_adj_2629)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_0_i986_3_lut.init = 16'hcaca;
    LUT4 mux_191_Mux_0_i971_3_lut (.A(n26710), .B(n26653), .C(index_i[3]), 
         .Z(n971_adj_2630)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_0_i971_3_lut.init = 16'hcaca;
    LUT4 i11457_2_lut_rep_415_3_lut_4_lut (.A(n26623), .B(index_q[1]), .C(index_q[4]), 
         .D(index_q[3]), .Z(n26375)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11457_2_lut_rep_415_3_lut_4_lut.init = 16'hfef0;
    LUT4 i19039_4_lut_4_lut_3_lut_4_lut (.A(n26623), .B(index_q[1]), .C(index_q[4]), 
         .D(index_q[3]), .Z(n21359)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19039_4_lut_4_lut_3_lut_4_lut.init = 16'h11ef;
    LUT4 n62_bdd_3_lut_24224_4_lut (.A(n26644), .B(index_q[3]), .C(index_q[4]), 
         .D(n30), .Z(n24458)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n62_bdd_3_lut_24224_4_lut.init = 16'hf808;
    LUT4 i19057_3_lut (.A(n526_adj_2286), .B(n15), .C(index_q[4]), .Z(n21377)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19057_3_lut.init = 16'hcaca;
    PFUMX i20126 (.BLUT(n21688), .ALUT(n317_adj_2631), .C0(index_i[5]), 
          .Z(n22465));
    LUT4 mux_191_Mux_0_i939_4_lut (.A(n773), .B(n26694), .C(index_i[3]), 
         .D(index_i[2]), .Z(n939_adj_2632)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_0_i939_4_lut.init = 16'hfaca;
    LUT4 n25073_bdd_3_lut (.A(n25073), .B(n22110), .C(index_q[6]), .Z(n25981)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n25073_bdd_3_lut.init = 16'hcaca;
    PFUMX i20127 (.BLUT(n349_adj_2633), .ALUT(n21691), .C0(index_i[5]), 
          .Z(n22466));
    LUT4 index_q_3__bdd_3_lut_24394_4_lut_4_lut (.A(n26644), .B(index_q[3]), 
         .C(index_q[4]), .D(n29190), .Z(n24166)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C))+!A !(B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam index_q_3__bdd_3_lut_24394_4_lut_4_lut.init = 16'h838f;
    LUT4 i20219_3_lut_3_lut_4_lut_4_lut (.A(n26644), .B(index_q[3]), .C(index_q[4]), 
         .D(n26526), .Z(n22558)) /* synthesis lut_function=(!(A (B (C)+!B ((D)+!C))+!A (B+((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20219_3_lut_3_lut_4_lut_4_lut.init = 16'h0838;
    LUT4 i9572_3_lut_4_lut_4_lut (.A(n26644), .B(index_q[3]), .C(index_q[5]), 
         .D(n26430), .Z(n12018)) /* synthesis lut_function=(A (B+(C (D)))+!A (B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9572_3_lut_4_lut_4_lut.init = 16'hf8c8;
    LUT4 mux_191_Mux_0_i923_3_lut (.A(n26606), .B(n29194), .C(index_i[3]), 
         .Z(n923_adj_2634)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_0_i923_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_10_i574_4_lut_4_lut (.A(n26411), .B(index_q[4]), .C(index_q[5]), 
         .D(n26401), .Z(n574_adj_2434)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_10_i574_4_lut_4_lut.init = 16'h1f1c;
    LUT4 index_q_4__bdd_4_lut_24851 (.A(index_q[4]), .B(n26411), .C(n24162), 
         .D(index_q[5]), .Z(n26346)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (B (C (D))+!B (C+!(D)))) */ ;
    defparam index_q_4__bdd_4_lut_24851.init = 16'hf099;
    PFUMX i18993 (.BLUT(n21311), .ALUT(n21312), .C0(index_i[5]), .Z(n21313));
    LUT4 i19054_3_lut (.A(n397_adj_2635), .B(n475_adj_2449), .C(index_q[4]), 
         .Z(n21374)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19054_3_lut.init = 16'hcaca;
    PFUMX i18996 (.BLUT(n21314), .ALUT(n21315), .C0(index_i[5]), .Z(n21316));
    LUT4 i19049_3_lut (.A(n348_adj_2636), .B(n443_adj_2637), .C(index_q[4]), 
         .Z(n21369)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19049_3_lut.init = 16'hcaca;
    LUT4 i19048_3_lut (.A(n397_adj_2635), .B(n781), .C(index_q[4]), .Z(n21368)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19048_3_lut.init = 16'hcaca;
    LUT4 i11298_3_lut (.A(index_q[3]), .B(index_q[1]), .C(index_q[0]), 
         .Z(n13857)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11298_3_lut.init = 16'hc8c8;
    LUT4 mux_192_Mux_3_i348_3_lut (.A(n26721), .B(n29173), .C(index_q[3]), 
         .Z(n348_adj_2638)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_3_i348_3_lut.init = 16'hcaca;
    L6MUX21 i20128 (.D0(n21694), .D1(n21697), .SD(index_i[5]), .Z(n22467));
    PFUMX i18999 (.BLUT(n21317), .ALUT(n21318), .C0(index_i[5]), .Z(n21319));
    LUT4 i19046_3_lut (.A(n364_adj_2341), .B(n890_adj_2338), .C(index_q[4]), 
         .Z(n21366)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19046_3_lut.init = 16'hcaca;
    LUT4 i19045_3_lut (.A(n333), .B(n348_adj_2636), .C(index_q[4]), .Z(n21365)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19045_3_lut.init = 16'hcaca;
    L6MUX21 i20129 (.D0(n21700), .D1(n21703), .SD(index_i[5]), .Z(n22468));
    PFUMX i19002 (.BLUT(n21320), .ALUT(n21321), .C0(index_i[5]), .Z(n21322));
    PFUMX i20769 (.BLUT(n557_adj_2639), .ALUT(n572_adj_2640), .C0(index_i[4]), 
          .Z(n23108));
    LUT4 i12402_2_lut_3_lut_4_lut (.A(n26414), .B(index_i[4]), .C(index_i[6]), 
         .D(index_i[5]), .Z(n14982)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i12402_2_lut_3_lut_4_lut.init = 16'hfef0;
    LUT4 i19394_3_lut (.A(n26709), .B(n26688), .C(index_i[3]), .Z(n21714)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19394_3_lut.init = 16'hcaca;
    PFUMX i20130 (.BLUT(n21706), .ALUT(n573_adj_2641), .C0(index_i[5]), 
          .Z(n22469));
    LUT4 i20555_3_lut_3_lut_4_lut (.A(n29190), .B(index_q[3]), .C(n93_adj_2642), 
         .D(index_q[4]), .Z(n22894)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20555_3_lut_3_lut_4_lut.init = 16'hf077;
    LUT4 mux_192_Mux_3_i908_3_lut (.A(n29167), .B(n29175), .C(index_q[3]), 
         .Z(n908_adj_2643)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_3_i908_3_lut.init = 16'hcaca;
    LUT4 n24913_bdd_3_lut_25402 (.A(n24913), .B(n22114), .C(index_q[6]), 
         .Z(n25979)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n24913_bdd_3_lut_25402.init = 16'hcaca;
    LUT4 index_i_4__bdd_4_lut (.A(index_i[4]), .B(n26414), .C(n24127), 
         .D(index_i[5]), .Z(n26347)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (B (C (D))+!B (C+!(D)))) */ ;
    defparam index_i_4__bdd_4_lut.init = 16'hf099;
    LUT4 mux_191_Mux_10_i574_4_lut_4_lut (.A(n26414), .B(index_i[4]), .C(index_i[5]), 
         .D(n26397), .Z(n574_adj_2435)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_10_i574_4_lut_4_lut.init = 16'h1f1c;
    L6MUX21 i20131 (.D0(n21709), .D1(n636), .SD(index_i[5]), .Z(n22470));
    LUT4 n24913_bdd_3_lut_24180 (.A(n22115), .B(n24919), .C(index_q[6]), 
         .Z(n25978)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n24913_bdd_3_lut_24180.init = 16'hcaca;
    PFUMX i20132 (.BLUT(n21712), .ALUT(n700_adj_2369), .C0(index_i[5]), 
          .Z(n22471));
    LUT4 mux_191_Mux_6_i653_3_lut (.A(n26689), .B(n619), .C(index_i[3]), 
         .Z(n653_adj_2644)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_6_i653_3_lut.init = 16'hcaca;
    LUT4 i19379_3_lut (.A(n26591), .B(n26703), .C(index_i[3]), .Z(n21699)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19379_3_lut.init = 16'hcaca;
    L6MUX21 i20134 (.D0(n21715), .D1(n21718), .SD(index_i[5]), .Z(n22473));
    PFUMX i20136 (.BLUT(n924_adj_2645), .ALUT(n21724), .C0(index_i[5]), 
          .Z(n22475));
    LUT4 mux_192_Mux_3_i221_3_lut_4_lut (.A(n29190), .B(index_q[3]), .C(index_q[4]), 
         .D(n26429), .Z(n221_adj_2646)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_3_i221_3_lut_4_lut.init = 16'h08f8;
    CCU2D add_372_9 (.A0(quarter_wave_sample_register_q[8]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_q[9]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17341), .COUT(n17342), 
          .S0(o_val_pipeline_q_0__15__N_2190[8]), .S1(o_val_pipeline_q_0__15__N_2190[9]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(80[29:60])
    defparam add_372_9.INIT0 = 16'hf555;
    defparam add_372_9.INIT1 = 16'hf555;
    defparam add_372_9.INJECT1_0 = "NO";
    defparam add_372_9.INJECT1_1 = "NO";
    LUT4 mux_191_Mux_5_i397_3_lut (.A(n26687), .B(n204), .C(index_i[3]), 
         .Z(n397_adj_2647)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_5_i397_3_lut.init = 16'hcaca;
    LUT4 n26603_bdd_2_lut_25991_4_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[0]), 
         .D(index_i[4]), .Z(n27929)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A !(B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n26603_bdd_2_lut_25991_4_lut.init = 16'h6400;
    PFUMX i20137 (.BLUT(n987), .ALUT(n21727), .C0(index_i[5]), .Z(n22476));
    LUT4 mux_191_Mux_0_i716_3_lut (.A(n26705), .B(n26588), .C(index_i[3]), 
         .Z(n716_adj_2648)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_0_i716_3_lut.init = 16'hcaca;
    LUT4 mux_191_Mux_6_i891_3_lut (.A(n301_adj_2256), .B(n890_adj_2590), 
         .C(index_i[4]), .Z(n891_adj_2649)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_6_i891_3_lut.init = 16'hcaca;
    LUT4 mux_191_Mux_6_i828_4_lut (.A(n812_adj_2650), .B(n14092), .C(index_i[4]), 
         .D(index_i[2]), .Z(n828_adj_2651)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_6_i828_4_lut.init = 16'hfaca;
    LUT4 mux_192_Mux_5_i491_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n491_adj_2334)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A !(B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_5_i491_3_lut_4_lut_4_lut.init = 16'ha54a;
    LUT4 mux_191_Mux_6_i797_3_lut (.A(n781_adj_2526), .B(n26358), .C(index_i[4]), 
         .Z(n797_adj_2652)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_6_i797_3_lut.init = 16'hcaca;
    LUT4 mux_191_Mux_5_i506_3_lut (.A(n26592), .B(n26591), .C(index_i[3]), 
         .Z(n506_adj_2653)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_5_i506_3_lut.init = 16'hcaca;
    LUT4 mux_191_Mux_6_i518_3_lut_3_lut_rep_742 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26702)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_6_i518_3_lut_3_lut_rep_742.init = 16'h6c6c;
    PFUMX i19005 (.BLUT(n21323), .ALUT(n21324), .C0(index_i[5]), .Z(n21325));
    PFUMX i19856 (.BLUT(n221_adj_2304), .ALUT(n252_adj_2327), .C0(index_q[5]), 
          .Z(n22195));
    LUT4 i19372_3_lut (.A(n26709), .B(n26608), .C(index_i[3]), .Z(n21692)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19372_3_lut.init = 16'hcaca;
    LUT4 mux_191_Mux_6_i669_3_lut (.A(n653_adj_2644), .B(n668_adj_2654), 
         .C(index_i[4]), .Z(n669_adj_2655)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_6_i669_3_lut.init = 16'hcaca;
    PFUMX i24508 (.BLUT(n26808), .ALUT(n26809), .C0(index_q[1]), .Z(n26810));
    LUT4 i9429_3_lut_3_lut_4_lut_4_lut (.A(index_q[2]), .B(index_q[3]), 
         .C(index_q[0]), .D(index_q[1]), .Z(n762_adj_2626)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C (D)+!C !(D)))+!A !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9429_3_lut_3_lut_4_lut_4_lut.init = 16'h700f;
    LUT4 i18742_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21062)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18742_3_lut_4_lut.init = 16'h64cc;
    LUT4 i21657_3_lut (.A(n21689), .B(n21690), .C(index_i[4]), .Z(n21691)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21657_3_lut.init = 16'hcaca;
    LUT4 mux_191_Mux_1_i317_3_lut (.A(n301_adj_2656), .B(n908_adj_2657), 
         .C(index_i[4]), .Z(n317_adj_2631)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_1_i317_3_lut.init = 16'hcaca;
    PFUMX i20569 (.BLUT(n22892), .ALUT(n22893), .C0(index_q[5]), .Z(n22908));
    LUT4 mux_191_Mux_6_i542_3_lut (.A(n526_adj_2261), .B(n541_adj_2658), 
         .C(index_i[4]), .Z(n542_adj_2659)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_6_i542_3_lut.init = 16'hcaca;
    LUT4 mux_191_Mux_5_i15_3_lut (.A(n26691), .B(n26604), .C(index_i[3]), 
         .Z(n15_adj_2519)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_5_i15_3_lut.init = 16'hcaca;
    LUT4 i19037_3_lut (.A(n491_adj_2279), .B(n541_adj_2288), .C(index_q[4]), 
         .Z(n21357)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19037_3_lut.init = 16'hcaca;
    LUT4 i19036_3_lut (.A(n557_adj_2660), .B(n475_adj_2507), .C(index_q[4]), 
         .Z(n21356)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19036_3_lut.init = 16'hcaca;
    PFUMX i20570 (.BLUT(n22894), .ALUT(n22895), .C0(index_q[5]), .Z(n22909));
    LUT4 mux_191_Mux_5_i859_3_lut (.A(n308), .B(n26691), .C(index_i[3]), 
         .Z(n859_adj_2661)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_5_i859_3_lut.init = 16'hcaca;
    LUT4 mux_191_Mux_5_i875_3_lut (.A(n70), .B(n26652), .C(index_i[3]), 
         .Z(n875_adj_2662)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_5_i875_3_lut.init = 16'hcaca;
    L6MUX21 i20571 (.D0(n22896), .D1(n22897), .SD(index_q[5]), .Z(n22910));
    PFUMX i20770 (.BLUT(n589_adj_2663), .ALUT(n604_adj_2337), .C0(index_i[4]), 
          .Z(n23109));
    LUT4 mux_192_Mux_4_i828_3_lut_4_lut (.A(index_q[4]), .B(index_q[3]), 
         .C(n812), .D(n26544), .Z(n828_adj_2664)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_4_i828_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i19028_3_lut_then_4_lut (.A(index_q[4]), .B(index_q[2]), .C(index_q[3]), 
         .D(index_q[0]), .Z(n26806)) /* synthesis lut_function=(!(A (B (C)+!B ((D)+!C))+!A !((C)+!B))) */ ;
    defparam i19028_3_lut_then_4_lut.init = 16'h5979;
    LUT4 mux_192_Mux_0_i620_3_lut (.A(n29187), .B(n29170), .C(index_q[3]), 
         .Z(n620_adj_2427)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_0_i620_3_lut.init = 16'hcaca;
    LUT4 i19034_3_lut (.A(n251), .B(n443_adj_2354), .C(index_q[4]), .Z(n21354)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19034_3_lut.init = 16'hcaca;
    LUT4 mux_191_Mux_0_i653_3_lut (.A(n70), .B(n26592), .C(index_i[3]), 
         .Z(n653_adj_2665)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_0_i653_3_lut.init = 16'hcaca;
    LUT4 mux_191_Mux_6_i250_3_lut_4_lut_3_lut_rep_743 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26703)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_6_i250_3_lut_4_lut_3_lut_rep_743.init = 16'h9696;
    LUT4 i19033_3_lut (.A(n557_adj_2660), .B(n14848), .C(index_q[4]), 
         .Z(n21353)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;
    defparam i19033_3_lut.init = 16'h3a3a;
    LUT4 mux_191_Mux_4_i61_3_lut (.A(n26709), .B(n26588), .C(index_i[3]), 
         .Z(n61_adj_2522)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_4_i61_3_lut.init = 16'hcaca;
    L6MUX21 i20574 (.D0(n22902), .D1(n22903), .SD(index_q[5]), .Z(n22913));
    LUT4 i19360_3_lut (.A(n723), .B(n26688), .C(index_i[3]), .Z(n21680)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19360_3_lut.init = 16'hcaca;
    LUT4 i19028_3_lut_else_4_lut (.A(index_q[4]), .B(index_q[2]), .C(index_q[3]), 
         .D(index_q[0]), .Z(n26805)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A !(B (C+!(D))+!B !(C)))) */ ;
    defparam i19028_3_lut_else_4_lut.init = 16'h6965;
    L6MUX21 i20575 (.D0(n22904), .D1(n22905), .SD(index_q[5]), .Z(n22914));
    LUT4 i22084_3_lut (.A(n29204), .B(n26807), .C(index_q[5]), .Z(n21349)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22084_3_lut.init = 16'hcaca;
    L6MUX21 i20576 (.D0(n22906), .D1(n22907), .SD(index_q[5]), .Z(n22915));
    LUT4 i19024_3_lut (.A(n875_adj_2571), .B(n93_adj_2368), .C(index_q[4]), 
         .Z(n21344)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19024_3_lut.init = 16'hcaca;
    PFUMX i19008 (.BLUT(n21326), .ALUT(n21327), .C0(index_i[5]), .Z(n21328));
    LUT4 i19021_3_lut (.A(n15_adj_2403), .B(n526_adj_2360), .C(index_q[4]), 
         .Z(n21341)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19021_3_lut.init = 16'hcaca;
    LUT4 i20554_3_lut_4_lut (.A(n29190), .B(index_q[3]), .C(index_q[4]), 
         .D(n46), .Z(n22893)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20554_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_192_Mux_5_i564_3_lut_3_lut_rep_796 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29175)) /* synthesis lut_function=(A (B (C))+!A !(B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_5_i564_3_lut_3_lut_rep_796.init = 16'h9595;
    PFUMX i20771 (.BLUT(n620_adj_2666), .ALUT(n635_adj_2667), .C0(index_i[4]), 
          .Z(n23110));
    LUT4 i21664_3_lut (.A(n26804), .B(n21678), .C(index_i[4]), .Z(n21679)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21664_3_lut.init = 16'hcaca;
    LUT4 mux_191_Mux_7_i892_3_lut (.A(n62_adj_2271), .B(n891_adj_2413), 
         .C(index_i[5]), .Z(n892)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_7_i892_3_lut.init = 16'hcaca;
    PFUMX i19011 (.BLUT(n21329), .ALUT(n21330), .C0(index_i[5]), .Z(n21331));
    LUT4 i19016_3_lut (.A(n747_adj_2315), .B(n762_adj_2668), .C(index_i[4]), 
         .Z(n21336)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19016_3_lut.init = 16'hcaca;
    LUT4 i19015_3_lut (.A(n716_adj_2669), .B(n14770), .C(index_i[4]), 
         .Z(n21335)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19015_3_lut.init = 16'hcaca;
    CCU2D add_372_7 (.A0(quarter_wave_sample_register_q[6]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_q[7]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17340), .COUT(n17341), 
          .S1(o_val_pipeline_q_0__15__N_2190[7]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(80[29:60])
    defparam add_372_7.INIT0 = 16'hf555;
    defparam add_372_7.INIT1 = 16'hf555;
    defparam add_372_7.INJECT1_0 = "NO";
    defparam add_372_7.INJECT1_1 = "NO";
    LUT4 mux_191_Mux_4_i270_3_lut (.A(n26686), .B(n26592), .C(index_i[3]), 
         .Z(n270_adj_2670)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_4_i270_3_lut.init = 16'hcaca;
    LUT4 mux_191_Mux_4_i15_3_lut (.A(n26591), .B(n773), .C(index_i[3]), 
         .Z(n15_adj_2524)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_4_i15_3_lut.init = 16'hcaca;
    PFUMX i24506 (.BLUT(n26805), .ALUT(n26806), .C0(index_q[1]), .Z(n26807));
    LUT4 i19013_3_lut (.A(n93_adj_2671), .B(n699_adj_2352), .C(index_i[4]), 
         .Z(n21333)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19013_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_5_i731_3_lut (.A(n26737), .B(n26734), .C(index_q[3]), 
         .Z(n731_adj_2672)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_5_i731_3_lut.init = 16'hcaca;
    PFUMX i19014 (.BLUT(n21332), .ALUT(n21333), .C0(index_i[5]), .Z(n21334));
    PFUMX mux_192_Mux_5_i732 (.BLUT(n11856), .ALUT(n731_adj_2672), .C0(index_q[4]), 
          .Z(n732_adj_2673)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 i19012_3_lut (.A(n653_adj_2412), .B(n26388), .C(index_i[4]), 
         .Z(n21332)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19012_3_lut.init = 16'hcaca;
    CCU2D add_372_5 (.A0(quarter_wave_sample_register_q[4]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_q[5]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17339), .COUT(n17340));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(80[29:60])
    defparam add_372_5.INIT0 = 16'hf555;
    defparam add_372_5.INIT1 = 16'hf555;
    defparam add_372_5.INJECT1_0 = "NO";
    defparam add_372_5.INJECT1_1 = "NO";
    LUT4 mux_191_Mux_4_i348_3_lut (.A(n26587), .B(n26697), .C(index_i[3]), 
         .Z(n348_adj_2674)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_4_i348_3_lut.init = 16'hcaca;
    LUT4 mux_191_Mux_0_i620_3_lut (.A(n26652), .B(n26686), .C(index_i[3]), 
         .Z(n620_adj_2666)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_0_i620_3_lut.init = 16'hcaca;
    PFUMX i19017 (.BLUT(n21335), .ALUT(n21336), .C0(index_i[5]), .Z(n21337));
    LUT4 i19006_3_lut (.A(n526_adj_2302), .B(n541_adj_2675), .C(index_i[4]), 
         .Z(n21326)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19006_3_lut.init = 16'hcaca;
    LUT4 i19042_3_lut_4_lut_4_lut (.A(n26430), .B(index_q[4]), .C(index_q[3]), 
         .D(n26526), .Z(n21362)) /* synthesis lut_function=(A (B (C)+!B !(C+!(D)))+!A (B (C)+!B (C+(D)))) */ ;
    defparam i19042_3_lut_4_lut_4_lut.init = 16'hd3d0;
    LUT4 mux_191_Mux_0_i589_3_lut (.A(n29194), .B(n773), .C(index_i[3]), 
         .Z(n589_adj_2663)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_0_i589_3_lut.init = 16'hcaca;
    LUT4 i21543_3_lut_then_3_lut (.A(index_q[0]), .B(index_q[4]), .C(index_q[3]), 
         .Z(n26809)) /* synthesis lut_function=(A (B)+!A (B (C)+!B !(C))) */ ;
    defparam i21543_3_lut_then_3_lut.init = 16'hc9c9;
    LUT4 mux_191_Mux_4_i684_3_lut (.A(n619), .B(n108), .C(index_i[3]), 
         .Z(n684_adj_2676)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_4_i684_3_lut.init = 16'hcaca;
    LUT4 i21543_3_lut_else_3_lut (.A(index_q[2]), .B(index_q[0]), .C(index_q[4]), 
         .D(index_q[3]), .Z(n26808)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)+!C !(D)))+!A (B (C+!(D))+!B !(C)))) */ ;
    defparam i21543_3_lut_else_3_lut.init = 16'h1e38;
    LUT4 i20553_3_lut (.A(n15), .B(n29201), .C(index_q[4]), .Z(n22892)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20553_3_lut.init = 16'hcaca;
    LUT4 i19351_3_lut (.A(n404), .B(n26599), .C(index_i[3]), .Z(n21671)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19351_3_lut.init = 16'hcaca;
    PFUMX i19362 (.BLUT(n21680), .ALUT(n21681), .C0(index_i[4]), .Z(n21682));
    LUT4 i21688_3_lut (.A(n21671), .B(n21672), .C(index_i[4]), .Z(n21673)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21688_3_lut.init = 16'hcaca;
    LUT4 i19003_3_lut (.A(n397_adj_2677), .B(n475_adj_2411), .C(index_i[4]), 
         .Z(n21323)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19003_3_lut.init = 16'hcaca;
    PFUMX i19023 (.BLUT(n21341), .ALUT(n21342), .C0(index_q[5]), .Z(n21343));
    LUT4 i23093_then_4_lut (.A(index_i[6]), .B(index_i[2]), .C(index_i[5]), 
         .D(index_i[0]), .Z(n26812)) /* synthesis lut_function=(A ((C+!(D))+!B)+!A !(B (C (D))+!B !(C+(D)))) */ ;
    defparam i23093_then_4_lut.init = 16'hb7fe;
    LUT4 i23093_else_4_lut (.A(index_i[2]), .Z(n26811)) /* synthesis lut_function=(A) */ ;
    defparam i23093_else_4_lut.init = 16'haaaa;
    LUT4 i22429_2_lut (.A(index_q[5]), .B(index_q[4]), .Z(n22040)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i22429_2_lut.init = 16'heeee;
    LUT4 i19346_3_lut (.A(n404), .B(n29177), .C(index_i[3]), .Z(n21666)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19346_3_lut.init = 16'hcaca;
    LUT4 mux_191_Mux_1_i924_3_lut (.A(n908), .B(n412_adj_2319), .C(index_i[4]), 
         .Z(n924_adj_2645)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_1_i924_3_lut.init = 16'hcaca;
    PFUMX i19026 (.BLUT(n21344), .ALUT(n21345), .C0(index_q[5]), .Z(n21346));
    L6MUX21 i20585 (.D0(n21535), .D1(n21538), .SD(index_i[5]), .Z(n22924));
    CCU2D add_372_3 (.A0(quarter_wave_sample_register_q[2]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_q[3]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17338), .COUT(n17339));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(80[29:60])
    defparam add_372_3.INIT0 = 16'hf555;
    defparam add_372_3.INIT1 = 16'hf555;
    defparam add_372_3.INJECT1_0 = "NO";
    defparam add_372_3.INJECT1_1 = "NO";
    LUT4 mux_192_Mux_6_i955_3_lut_4_lut (.A(n26496), .B(index_q[3]), .C(index_q[4]), 
         .D(n26357), .Z(n955_adj_2678)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_6_i955_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_191_Mux_5_i754_3_lut_4_lut_3_lut_rep_745 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26705)) /* synthesis lut_function=(!(A (B)+!A ((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_5_i754_3_lut_4_lut_3_lut_rep_745.init = 16'h2626;
    LUT4 i21646_3_lut (.A(n21710), .B(n21711), .C(index_i[4]), .Z(n21712)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21646_3_lut.init = 16'hcaca;
    LUT4 mux_191_Mux_5_i371_3_lut_4_lut_4_lut_3_lut_rep_746 (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[2]), .Z(n26706)) /* synthesis lut_function=(A ((C)+!B)+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_5_i371_3_lut_4_lut_4_lut_3_lut_rep_746.init = 16'hb6b6;
    LUT4 i21649_3_lut (.A(n29205), .B(n21705), .C(index_i[4]), .Z(n21706)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21649_3_lut.init = 16'hcaca;
    LUT4 i19001_3_lut (.A(n348_adj_2679), .B(n443_adj_2680), .C(index_i[4]), 
         .Z(n21321)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19001_3_lut.init = 16'hcaca;
    L6MUX21 i20589 (.D0(n21547), .D1(n17569), .SD(index_i[5]), .Z(n22928));
    L6MUX21 i20590 (.D0(n21550), .D1(n11955), .SD(index_i[5]), .Z(n22929));
    LUT4 i19000_3_lut (.A(n397_adj_2677), .B(n731_adj_2538), .C(index_i[4]), 
         .Z(n21320)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19000_3_lut.init = 16'hcaca;
    LUT4 i18998_3_lut (.A(n364_adj_2321), .B(n379_adj_2365), .C(index_i[4]), 
         .Z(n21318)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18998_3_lut.init = 16'hcaca;
    PFUMX i20772 (.BLUT(n653_adj_2665), .ALUT(n668_adj_2681), .C0(index_i[4]), 
          .Z(n23111));
    PFUMX i19035 (.BLUT(n21353), .ALUT(n21354), .C0(index_q[5]), .Z(n21355));
    LUT4 i18997_3_lut (.A(n333_adj_2682), .B(n348_adj_2679), .C(index_i[4]), 
         .Z(n21317)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18997_3_lut.init = 16'hcaca;
    LUT4 i21697_3_lut (.A(n21662), .B(n21663), .C(index_i[4]), .Z(n21664)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21697_3_lut.init = 16'hcaca;
    PFUMX i20167 (.BLUT(n956_adj_2622), .ALUT(n20006), .C0(index_q[6]), 
          .Z(n22506));
    LUT4 i19340_3_lut (.A(n29177), .B(n26707), .C(index_i[3]), .Z(n21660)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19340_3_lut.init = 16'hcaca;
    PFUMX i19365 (.BLUT(n21683), .ALUT(n21684), .C0(index_i[4]), .Z(n21685));
    LUT4 i21699_3_lut (.A(n21659), .B(n21660), .C(index_i[4]), .Z(n21661)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21699_3_lut.init = 16'hcaca;
    LUT4 i12221_3_lut (.A(index_i[3]), .B(index_i[1]), .C(index_i[0]), 
         .Z(n14791)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i12221_3_lut.init = 16'hc8c8;
    LUT4 i21702_3_lut (.A(n21656), .B(n21657), .C(index_i[4]), .Z(n21658)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21702_3_lut.init = 16'hcaca;
    PFUMX i19038 (.BLUT(n21356), .ALUT(n21357), .C0(index_q[5]), .Z(n21358));
    LUT4 mux_191_Mux_1_i349_3_lut (.A(n506_adj_2683), .B(n348), .C(index_i[4]), 
         .Z(n349_adj_2633)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_1_i349_3_lut.init = 16'hcaca;
    LUT4 mux_191_Mux_3_i348_3_lut (.A(n29178), .B(n26688), .C(index_i[3]), 
         .Z(n348_adj_2684)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_3_i348_3_lut.init = 16'hcaca;
    LUT4 i22272_3_lut (.A(n24134), .B(n22318), .C(index_i[8]), .Z(n22320)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22272_3_lut.init = 16'hcaca;
    LUT4 i21659_3_lut (.A(n21686), .B(n21687), .C(index_i[4]), .Z(n21688)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21659_3_lut.init = 16'hcaca;
    PFUMX i19041 (.BLUT(n21359), .ALUT(n21360), .C0(index_q[5]), .Z(n21361));
    LUT4 i11404_2_lut_rep_390_3_lut_4_lut (.A(n26419), .B(index_i[4]), .C(index_i[6]), 
         .D(index_i[5]), .Z(n26350)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11404_2_lut_rep_390_3_lut_4_lut.init = 16'hf080;
    PFUMX i20592 (.BLUT(n542_adj_2659), .ALUT(n573_adj_2685), .C0(index_i[5]), 
          .Z(n22931));
    LUT4 mux_191_Mux_1_i94_3_lut (.A(index_i[0]), .B(n93_adj_2686), .C(index_i[4]), 
         .Z(n94_adj_2627)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_1_i94_3_lut.init = 16'hcaca;
    LUT4 i18989_3_lut (.A(n491_adj_2687), .B(n506_adj_2683), .C(index_i[4]), 
         .Z(n21309)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18989_3_lut.init = 16'hcaca;
    LUT4 i18988_3_lut (.A(n397_adj_2432), .B(n475_adj_2588), .C(index_i[4]), 
         .Z(n21308)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18988_3_lut.init = 16'hcaca;
    PFUMX i20593 (.BLUT(n605_adj_2688), .ALUT(n636_adj_2689), .C0(index_i[5]), 
          .Z(n22932));
    LUT4 mux_191_Mux_0_i30_3_lut (.A(n26649), .B(n26605), .C(index_i[3]), 
         .Z(n30_adj_2690)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_0_i30_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_3_i747_3_lut (.A(n26543), .B(n498), .C(index_q[3]), 
         .Z(n747_adj_2625)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_3_i747_3_lut.init = 16'hcaca;
    LUT4 i18986_3_lut (.A(n251_adj_2322), .B(n443_adj_2350), .C(index_i[4]), 
         .Z(n21306)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18986_3_lut.init = 16'hcaca;
    LUT4 i19262_3_lut_4_lut (.A(n26636), .B(index_i[1]), .C(index_i[3]), 
         .D(n404), .Z(n21582)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19262_3_lut_4_lut.init = 16'hdfd0;
    LUT4 i18985_3_lut (.A(n397_adj_2432), .B(n14770), .C(index_i[4]), 
         .Z(n21305)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;
    defparam i18985_3_lut.init = 16'h3a3a;
    PFUMX i20594 (.BLUT(n669_adj_2655), .ALUT(n700_adj_2691), .C0(index_i[5]), 
          .Z(n22933));
    LUT4 i19328_3_lut (.A(n396), .B(n26688), .C(index_i[3]), .Z(n21648)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19328_3_lut.init = 16'hcaca;
    LUT4 mux_191_Mux_1_i620_3_lut_4_lut (.A(n26636), .B(index_i[1]), .C(index_i[3]), 
         .D(n26686), .Z(n620)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_1_i620_3_lut_4_lut.init = 16'hdfd0;
    LUT4 mux_191_Mux_0_i173_3_lut_4_lut (.A(n26636), .B(index_i[1]), .C(index_i[3]), 
         .D(n26697), .Z(n173_adj_2692)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_0_i173_3_lut_4_lut.init = 16'hdfd0;
    LUT4 i21723_3_lut (.A(n21647), .B(n21648), .C(index_i[4]), .Z(n21649)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21723_3_lut.init = 16'hcaca;
    PFUMX i19374 (.BLUT(n21692), .ALUT(n21693), .C0(index_i[4]), .Z(n21694));
    LUT4 i9612_3_lut_else_4_lut (.A(index_q[4]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n29206)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C+!(D)))+!A !(B (C (D)+!C !(D))+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9612_3_lut_else_4_lut.init = 16'h5295;
    LUT4 i19325_3_lut (.A(n26692), .B(n26706), .C(index_i[3]), .Z(n21645)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19325_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut (.A(index_q[0]), .B(index_q[4]), .C(index_q[2]), .Z(n20372)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_3_lut.init = 16'hfefe;
    LUT4 i21733_3_lut (.A(n21641), .B(n21642), .C(index_i[4]), .Z(n21643)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21733_3_lut.init = 16'hcaca;
    PFUMX i20595 (.BLUT(n732_adj_2693), .ALUT(n21556), .C0(index_i[5]), 
          .Z(n22934));
    LUT4 mux_191_Mux_3_i908_3_lut (.A(n26708), .B(n26588), .C(index_i[3]), 
         .Z(n908_adj_2694)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_3_i908_3_lut.init = 16'hcaca;
    PFUMX i19377 (.BLUT(n21695), .ALUT(n21696), .C0(index_i[4]), .Z(n21697));
    LUT4 i21476_3_lut (.A(n21014), .B(n21015), .C(index_q[4]), .Z(n21016)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21476_3_lut.init = 16'hcaca;
    LUT4 i21685_3_lut (.A(n716_adj_2695), .B(n731_adj_2359), .C(index_i[4]), 
         .Z(n732_adj_2616)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21685_3_lut.init = 16'hcaca;
    LUT4 mux_191_Mux_2_i669_3_lut (.A(n653_adj_2696), .B(n475_adj_2697), 
         .C(index_i[4]), .Z(n669_adj_2615)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_2_i669_3_lut.init = 16'hcaca;
    LUT4 mux_191_Mux_2_i605_3_lut (.A(n142_adj_2698), .B(n604_adj_2699), 
         .C(index_i[4]), .Z(n605_adj_2613)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_2_i605_3_lut.init = 16'hcaca;
    PFUMX i20596 (.BLUT(n797_adj_2652), .ALUT(n828_adj_2651), .C0(index_i[5]), 
          .Z(n22935));
    L6MUX21 i24185 (.D0(n25982), .D1(n25980), .SD(index_q[8]), .Z(n25983));
    PFUMX i20773 (.BLUT(n684_adj_2700), .ALUT(n699_adj_2701), .C0(index_i[4]), 
          .Z(n23112));
    PFUMX i20597 (.BLUT(n860_adj_2702), .ALUT(n891_adj_2649), .C0(index_i[5]), 
          .Z(n22936));
    LUT4 mux_191_Mux_3_i251_3_lut_4_lut (.A(n26636), .B(index_i[1]), .C(index_i[3]), 
         .D(n26519), .Z(n15026)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_3_i251_3_lut_4_lut.init = 16'hfe0e;
    LUT4 mux_191_Mux_0_i572_3_lut_4_lut (.A(n26636), .B(index_i[1]), .C(index_i[3]), 
         .D(n26710), .Z(n572_adj_2640)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_0_i572_3_lut_4_lut.init = 16'hefe0;
    LUT4 i21690_3_lut (.A(n26803), .B(n21669), .C(index_i[4]), .Z(n21670)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21690_3_lut.init = 16'hcaca;
    PFUMX i20774 (.BLUT(n716_adj_2648), .ALUT(n731_adj_2363), .C0(index_i[4]), 
          .Z(n23113));
    LUT4 i21692_3_lut (.A(n21665), .B(n21666), .C(index_i[4]), .Z(n21667)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21692_3_lut.init = 16'hcaca;
    LUT4 i9500_4_lut_4_lut (.A(n26636), .B(index_i[1]), .C(index_i[3]), 
         .D(n20376), .Z(n11946)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A (B (C)+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9500_4_lut_4_lut.init = 16'h0e3e;
    LUT4 mux_191_Mux_9_i364_3_lut_3_lut_4_lut (.A(n26636), .B(index_i[1]), 
         .C(index_i[3]), .D(n26519), .Z(n364_adj_2291)) /* synthesis lut_function=(!(A (C (D))+!A (B (C (D))+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_9_i364_3_lut_3_lut_4_lut.init = 16'h0efe;
    LUT4 i18976_3_lut (.A(n301_adj_2256), .B(n93_adj_2671), .C(index_i[4]), 
         .Z(n21296)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18976_3_lut.init = 16'hcaca;
    LUT4 index_i_3__bdd_3_lut_22608_3_lut_4_lut (.A(n26636), .B(index_i[1]), 
         .C(index_i[4]), .D(index_i[3]), .Z(n24130)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam index_i_3__bdd_3_lut_22608_3_lut_4_lut.init = 16'hf10f;
    LUT4 i11368_2_lut_rep_416_3_lut_4_lut (.A(n26636), .B(index_i[1]), .C(index_i[4]), 
         .D(index_i[3]), .Z(n26376)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11368_2_lut_rep_416_3_lut_4_lut.init = 16'hfef0;
    LUT4 i18991_4_lut_4_lut_3_lut_4_lut (.A(n26636), .B(index_i[1]), .C(index_i[4]), 
         .D(index_i[3]), .Z(n21311)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18991_4_lut_4_lut_3_lut_4_lut.init = 16'h11ef;
    LUT4 mux_191_Mux_2_i270_3_lut (.A(n26691), .B(n26607), .C(index_i[3]), 
         .Z(n270_adj_2703)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_2_i270_3_lut.init = 16'hcaca;
    PFUMX i20775 (.BLUT(n747), .ALUT(n762_adj_2704), .C0(index_i[4]), 
          .Z(n23114));
    PFUMX i24183 (.BLUT(n25981), .ALUT(n22126), .C0(index_q[7]), .Z(n25982));
    LUT4 n62_bdd_3_lut_4_lut (.A(n26637), .B(index_i[3]), .C(index_i[4]), 
         .D(n30_adj_2301), .Z(n24443)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n62_bdd_3_lut_4_lut.init = 16'hf808;
    LUT4 i20198_3_lut_3_lut_4_lut_4_lut (.A(n26637), .B(index_i[3]), .C(index_i[4]), 
         .D(n26519), .Z(n22537)) /* synthesis lut_function=(!(A (B (C)+!B ((D)+!C))+!A (B+((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20198_3_lut_3_lut_4_lut_4_lut.init = 16'h0838;
    LUT4 mux_191_Mux_2_i316_3_lut (.A(n26692), .B(n26709), .C(index_i[3]), 
         .Z(n316_adj_2705)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_2_i316_3_lut.init = 16'hcaca;
    LUT4 mux_191_Mux_2_i397_3_lut (.A(n29180), .B(n26606), .C(index_i[3]), 
         .Z(n397_adj_2706)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_2_i397_3_lut.init = 16'hcaca;
    LUT4 i19316_3_lut (.A(n26608), .B(n26592), .C(index_i[3]), .Z(n21636)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19316_3_lut.init = 16'hcaca;
    LUT4 i19315_3_lut (.A(n26710), .B(n26687), .C(index_i[3]), .Z(n21635)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19315_3_lut.init = 16'hcaca;
    LUT4 i18973_3_lut (.A(n157), .B(n30_adj_2707), .C(index_i[4]), .Z(n21293)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18973_3_lut.init = 16'hcaca;
    LUT4 mux_191_Mux_2_i413_3_lut (.A(n397_adj_2706), .B(n954_adj_2264), 
         .C(index_i[4]), .Z(n413_adj_2599)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_2_i413_3_lut.init = 16'hcaca;
    PFUMX i19044 (.BLUT(n21362), .ALUT(n21363), .C0(index_q[5]), .Z(n21364));
    LUT4 i21740_3_lut (.A(n21635), .B(n21636), .C(index_i[4]), .Z(n21637)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21740_3_lut.init = 16'hcaca;
    LUT4 index_i_3__bdd_3_lut_22640_4_lut_4_lut (.A(n26637), .B(index_i[3]), 
         .C(index_i[4]), .D(n26486), .Z(n24131)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C))+!A !(B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam index_i_3__bdd_3_lut_22640_4_lut_4_lut.init = 16'h838f;
    LUT4 mux_191_Mux_2_i317_3_lut (.A(n668_adj_2400), .B(n316_adj_2705), 
         .C(index_i[4]), .Z(n317_adj_2595)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_2_i317_3_lut.init = 16'hcaca;
    LUT4 mux_191_Mux_2_i286_3_lut (.A(n270_adj_2703), .B(n653_adj_2708), 
         .C(index_i[4]), .Z(n286_adj_2594)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_2_i286_3_lut.init = 16'hcaca;
    PFUMX i19380 (.BLUT(n21698), .ALUT(n21699), .C0(index_i[4]), .Z(n21700));
    LUT4 i9501_3_lut_4_lut_4_lut (.A(n26637), .B(index_i[3]), .C(index_i[5]), 
         .D(n26438), .Z(n11947)) /* synthesis lut_function=(A (B+(C (D)))+!A (B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9501_3_lut_4_lut_4_lut.init = 16'hf8c8;
    LUT4 i19313_3_lut (.A(n29180), .B(n26689), .C(index_i[3]), .Z(n21633)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19313_3_lut.init = 16'hcaca;
    LUT4 n25086_bdd_3_lut_25322 (.A(n22254), .B(n22255), .C(index_q[7]), 
         .Z(n26182)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n25086_bdd_3_lut_25322.init = 16'hcaca;
    LUT4 n25086_bdd_3_lut_24334 (.A(n25086), .B(n22256), .C(index_q[7]), 
         .Z(n26181)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n25086_bdd_3_lut_24334.init = 16'hacac;
    LUT4 i19312_3_lut (.A(n26650), .B(n619), .C(index_i[3]), .Z(n21632)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19312_3_lut.init = 16'hcaca;
    PFUMX i19383 (.BLUT(n21701), .ALUT(n21702), .C0(index_i[4]), .Z(n21703));
    LUT4 i21742_3_lut (.A(n21632), .B(n21633), .C(index_i[4]), .Z(n21634)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21742_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_5_i797_3_lut_4_lut (.A(index_q[4]), .B(index_q[3]), 
         .C(n26772), .D(n26543), .Z(n797_adj_2709)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_5_i797_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i21301_3_lut (.A(n21068), .B(n21069), .C(index_q[4]), .Z(n21070)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21301_3_lut.init = 16'hcaca;
    LUT4 i21707_3_lut (.A(n142_adj_2710), .B(n14127), .C(index_i[4]), 
         .Z(n158_adj_2592)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21707_3_lut.init = 16'hcaca;
    LUT4 n22265_bdd_3_lut (.A(n22258), .B(n22259), .C(index_q[7]), .Z(n26179)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n22265_bdd_3_lut.init = 16'hcaca;
    PFUMX i20200 (.BLUT(n22535), .ALUT(n22536), .C0(index_i[5]), .Z(n22539));
    PFUMX i19389 (.BLUT(n21707), .ALUT(n21708), .C0(index_i[4]), .Z(n21709));
    PFUMX i20201 (.BLUT(n22537), .ALUT(n22538), .C0(index_i[5]), .Z(n22540));
    PFUMX i20207 (.BLUT(n22542), .ALUT(n22543), .C0(index_i[5]), .Z(n22546));
    LUT4 i19304_3_lut (.A(n26706), .B(n396), .C(index_i[3]), .Z(n21624)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19304_3_lut.init = 16'hcaca;
    PFUMX i20208 (.BLUT(n22544), .ALUT(n22545), .C0(index_i[5]), .Z(n22547));
    LUT4 i21754_3_lut (.A(n21623), .B(n21624), .C(index_i[4]), .Z(n21625)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21754_3_lut.init = 16'hcaca;
    LUT4 i21721_3_lut (.A(n21650), .B(n26802), .C(index_i[4]), .Z(n21652)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21721_3_lut.init = 16'hcaca;
    PFUMX i19395 (.BLUT(n21713), .ALUT(n21714), .C0(index_i[4]), .Z(n21715));
    LUT4 mux_191_Mux_3_i924_3_lut (.A(n908_adj_2694), .B(index_i[0]), .C(index_i[4]), 
         .Z(n924_adj_2586)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_3_i924_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_6_i860_3_lut_3_lut (.A(n26387), .B(index_q[4]), .C(n844_adj_2320), 
         .Z(n860_adj_2711)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam mux_192_Mux_6_i860_3_lut_3_lut.init = 16'h7474;
    LUT4 i19022_3_lut_3_lut (.A(n26387), .B(index_q[4]), .C(n109_adj_2454), 
         .Z(n21342)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam i19022_3_lut_3_lut.init = 16'h7474;
    PFUMX i20422 (.BLUT(n22757), .ALUT(n22758), .C0(index_q[4]), .Z(n22761));
    LUT4 mux_191_Mux_3_i891_3_lut (.A(n541_adj_2658), .B(n890_adj_2537), 
         .C(index_i[4]), .Z(n891_adj_2582)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_3_i891_3_lut.init = 16'hcaca;
    LUT4 i18689_3_lut (.A(n498), .B(n26714), .C(index_q[3]), .Z(n21009)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18689_3_lut.init = 16'hcaca;
    LUT4 mux_191_Mux_3_i669_3_lut (.A(n653_adj_2708), .B(n668_adj_2400), 
         .C(index_i[4]), .Z(n669_adj_2577)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_3_i669_3_lut.init = 16'hcaca;
    PFUMX i20423 (.BLUT(n22759), .ALUT(n22760), .C0(index_q[4]), .Z(n22762));
    LUT4 i9545_4_lut (.A(n26546), .B(n26486), .C(index_i[3]), .D(index_i[4]), 
         .Z(n11991)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B ((D)+!C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9545_4_lut.init = 16'h3afa;
    LUT4 i22243_3_lut_4_lut (.A(n26495), .B(n19545), .C(index_q[8]), .D(n766), 
         .Z(n21177)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i22243_3_lut_4_lut.init = 16'hefe0;
    LUT4 i19300_3_lut (.A(n773), .B(n26709), .C(index_i[3]), .Z(n21620)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19300_3_lut.init = 16'hcaca;
    LUT4 i21735_3_lut (.A(n21638), .B(n21639), .C(index_i[4]), .Z(n21640)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21735_3_lut.init = 16'hcaca;
    LUT4 i20491_3_lut (.A(n541_adj_2675), .B(n30_adj_2690), .C(index_i[4]), 
         .Z(n22830)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20491_3_lut.init = 16'hcaca;
    LUT4 i19298_3_lut (.A(n723), .B(n396), .C(index_i[3]), .Z(n21618)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19298_3_lut.init = 16'hcaca;
    LUT4 mux_191_Mux_7_i333_3_lut (.A(n26650), .B(n70), .C(index_i[3]), 
         .Z(n333_adj_2682)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_7_i333_3_lut.init = 16'hcaca;
    LUT4 mux_191_Mux_7_i348_3_lut (.A(n26652), .B(n29194), .C(index_i[3]), 
         .Z(n348_adj_2679)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_7_i348_3_lut.init = 16'hcaca;
    LUT4 mux_191_Mux_7_i397_3_lut (.A(n26652), .B(n26650), .C(index_i[3]), 
         .Z(n397_adj_2677)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_7_i397_3_lut.init = 16'hcaca;
    PFUMX i19047 (.BLUT(n21365), .ALUT(n21366), .C0(index_q[5]), .Z(n21367));
    LUT4 mux_191_Mux_3_i476_3_lut (.A(n460_adj_2601), .B(n285_adj_2620), 
         .C(index_i[4]), .Z(n476_adj_2570)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_3_i476_3_lut.init = 16'hcaca;
    PFUMX i20776 (.BLUT(n781_adj_2379), .ALUT(n796_adj_2712), .C0(index_i[4]), 
          .Z(n23115));
    LUT4 mux_191_Mux_3_i413_3_lut (.A(n397_adj_2713), .B(n26590), .C(index_i[4]), 
         .Z(n413_adj_2566)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_3_i413_3_lut.init = 16'hcaca;
    PFUMX i24181 (.BLUT(n25979), .ALUT(n25978), .C0(index_q[7]), .Z(n25980));
    LUT4 i19291_3_lut (.A(n29180), .B(n26604), .C(index_i[3]), .Z(n21611)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19291_3_lut.init = 16'hcaca;
    LUT4 mux_191_Mux_3_i286_4_lut (.A(n93_adj_2587), .B(index_i[2]), .C(index_i[4]), 
         .D(n14791), .Z(n286_adj_2564)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_3_i286_4_lut.init = 16'h3aca;
    LUT4 mux_191_Mux_1_i986_3_lut (.A(n26652), .B(n29178), .C(index_i[3]), 
         .Z(n986_adj_2714)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_1_i986_3_lut.init = 16'hcaca;
    PFUMX i19398 (.BLUT(n21716), .ALUT(n21717), .C0(index_i[4]), .Z(n21718));
    PFUMX i20221 (.BLUT(n22556), .ALUT(n22557), .C0(index_q[5]), .Z(n22560));
    LUT4 mux_191_Mux_3_i158_3_lut (.A(n142_adj_2698), .B(n157_adj_2317), 
         .C(index_i[4]), .Z(n158_adj_2562)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_3_i158_3_lut.init = 16'hcaca;
    PFUMX i19050 (.BLUT(n21368), .ALUT(n21369), .C0(index_q[5]), .Z(n21370));
    LUT4 mux_191_Mux_3_i125_3_lut (.A(n46_adj_2715), .B(n30_adj_2707), .C(index_i[4]), 
         .Z(n125_adj_2560)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_3_i125_3_lut.init = 16'hcaca;
    PFUMX i20777 (.BLUT(n812_adj_2716), .ALUT(n12009), .C0(index_i[4]), 
          .Z(n23116));
    PFUMX i20222 (.BLUT(n22558), .ALUT(n22559), .C0(index_q[5]), .Z(n22561));
    LUT4 i19984_3_lut (.A(n190_adj_2717), .B(n25487), .C(index_i[6]), 
         .Z(n22323)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19984_3_lut.init = 16'hcaca;
    PFUMX i19056 (.BLUT(n21374), .ALUT(n21375), .C0(index_q[5]), .Z(n21376));
    LUT4 mux_192_Mux_8_i732_3_lut (.A(index_q[3]), .B(n15038), .C(index_q[5]), 
         .Z(n732_adj_2557)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_8_i732_3_lut.init = 16'h3a3a;
    LUT4 i19234_3_lut_3_lut_4_lut (.A(n26548), .B(index_i[2]), .C(n26606), 
         .D(index_i[3]), .Z(n21554)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (B (C (D))+!B (C+!(D)))) */ ;
    defparam i19234_3_lut_3_lut_4_lut.init = 16'hf099;
    LUT4 n476_bdd_3_lut_22884_4_lut (.A(n26548), .B(index_i[2]), .C(index_i[4]), 
         .D(n491_adj_2718), .Z(n24490)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+(D)))) */ ;
    defparam n476_bdd_3_lut_22884_4_lut.init = 16'h9f90;
    PFUMX i20779 (.BLUT(n875_adj_2719), .ALUT(n890_adj_2353), .C0(index_i[4]), 
          .Z(n23118));
    LUT4 i19985_3_lut (.A(n22694), .B(n21319), .C(index_i[6]), .Z(n22324)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19985_3_lut.init = 16'hcaca;
    LUT4 i20044_4_lut (.A(n21631), .B(n1002_adj_2720), .C(index_i[5]), 
         .D(index_i[4]), .Z(n22383)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;
    defparam i20044_4_lut.init = 16'hfaca;
    LUT4 mux_191_Mux_4_i860_3_lut (.A(n506_adj_2653), .B(n24948), .C(index_i[4]), 
         .Z(n860_adj_2554)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_4_i860_3_lut.init = 16'hcaca;
    PFUMX i20780 (.BLUT(n908_adj_2374), .ALUT(n923_adj_2634), .C0(index_i[4]), 
          .Z(n23119));
    PFUMX i20228 (.BLUT(n22563), .ALUT(n22564), .C0(index_q[5]), .Z(n22567));
    LUT4 i19321_3_lut_3_lut_4_lut (.A(n26548), .B(index_i[2]), .C(n70), 
         .D(index_i[3]), .Z(n21641)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (B (C (D))+!B (C+!(D)))) */ ;
    defparam i19321_3_lut_3_lut_4_lut.init = 16'hf099;
    PFUMX i20229 (.BLUT(n22565), .ALUT(n22566), .C0(index_q[5]), .Z(n22568));
    PFUMX i20781 (.BLUT(n939_adj_2632), .ALUT(n954), .C0(index_i[4]), 
          .Z(n23120));
    LUT4 i19286_3_lut (.A(n26697), .B(n26700), .C(index_i[3]), .Z(n21606)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19286_3_lut.init = 16'hcaca;
    LUT4 i19285_3_lut (.A(n26599), .B(n396), .C(index_i[3]), .Z(n21605)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19285_3_lut.init = 16'hcaca;
    LUT4 i21757_3_lut (.A(n21620), .B(n21621), .C(index_i[4]), .Z(n21622)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21757_3_lut.init = 16'hcaca;
    LUT4 i21770_3_lut (.A(n21605), .B(n21606), .C(index_i[4]), .Z(n21607)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21770_3_lut.init = 16'hcaca;
    LUT4 i19283_3_lut (.A(n26701), .B(n26592), .C(index_i[3]), .Z(n21603)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19283_3_lut.init = 16'hcaca;
    LUT4 i21759_3_lut (.A(n21617), .B(n21618), .C(index_i[4]), .Z(n21619)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21759_3_lut.init = 16'hcaca;
    LUT4 i21772_3_lut (.A(n21602), .B(n21603), .C(index_i[4]), .Z(n21604)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21772_3_lut.init = 16'hcaca;
    PFUMX i19059 (.BLUT(n21377), .ALUT(n21378), .C0(index_q[5]), .Z(n21379));
    LUT4 mux_191_Mux_3_i860_3_lut_4_lut (.A(n26548), .B(index_i[2]), .C(index_i[4]), 
         .D(n859_adj_2721), .Z(n860_adj_2581)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam mux_191_Mux_3_i860_3_lut_4_lut.init = 16'hf606;
    PFUMX i19401 (.BLUT(n21719), .ALUT(n21720), .C0(index_i[4]), .Z(n21721));
    LUT4 mux_191_Mux_4_i700_3_lut (.A(n684_adj_2676), .B(index_i[1]), .C(index_i[4]), 
         .Z(n700_adj_2550)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_4_i700_3_lut.init = 16'hcaca;
    LUT4 mux_191_Mux_4_i669_3_lut (.A(n781_adj_2526), .B(n668_adj_2373), 
         .C(index_i[4]), .Z(n669_adj_2549)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_4_i669_3_lut.init = 16'hcaca;
    LUT4 mux_191_Mux_7_i443_3_lut_4_lut (.A(n26548), .B(index_i[2]), .C(index_i[3]), 
         .D(n26606), .Z(n443_adj_2680)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;
    defparam mux_191_Mux_7_i443_3_lut_4_lut.init = 16'h6f60;
    PFUMX i19062 (.BLUT(n21380), .ALUT(n21381), .C0(index_q[5]), .Z(n21382));
    LUT4 i21776_3_lut (.A(n21599), .B(n21600), .C(index_i[4]), .Z(n21601)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21776_3_lut.init = 16'hcaca;
    LUT4 i19463_3_lut_4_lut (.A(index_q[0]), .B(n26644), .C(index_q[3]), 
         .D(n29162), .Z(n21783)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19463_3_lut_4_lut.init = 16'hfb0b;
    PFUMX i20782 (.BLUT(n971_adj_2630), .ALUT(n986_adj_2629), .C0(index_i[4]), 
          .Z(n23121));
    LUT4 mux_191_Mux_4_i542_3_lut (.A(n30_adj_2707), .B(n506_adj_2683), 
         .C(index_i[4]), .Z(n542_adj_2722)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_4_i542_3_lut.init = 16'hcaca;
    LUT4 i20038_4_lut (.A(n26451), .B(n26795), .C(index_i[5]), .D(index_i[4]), 
         .Z(n22377)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam i20038_4_lut.init = 16'hc5ca;
    LUT4 i20480_3_lut_4_lut_4_lut (.A(n26460), .B(index_q[4]), .C(index_q[5]), 
         .D(n26457), .Z(n22819)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C)+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20480_3_lut_4_lut_4_lut.init = 16'h0434;
    PFUMX i20783 (.BLUT(n1002_adj_2589), .ALUT(n1017), .C0(index_i[4]), 
          .Z(n23122));
    LUT4 mux_191_Mux_6_i668_3_lut (.A(n108), .B(n26648), .C(index_i[3]), 
         .Z(n668_adj_2654)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_6_i668_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_8_i892_3_lut_4_lut (.A(n26460), .B(index_q[4]), .C(index_q[5]), 
         .D(n860), .Z(n892_adj_2723)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_8_i892_3_lut_4_lut.init = 16'h4f40;
    LUT4 mux_191_Mux_6_i684_3_lut (.A(n70), .B(n29180), .C(index_i[3]), 
         .Z(n684_adj_2724)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_6_i684_3_lut.init = 16'hcaca;
    LUT4 i19276_3_lut (.A(n26700), .B(n26608), .C(index_i[3]), .Z(n21596)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19276_3_lut.init = 16'hcaca;
    PFUMX mux_191_Mux_1_i891 (.BLUT(n882), .ALUT(n890_adj_2725), .C0(n26562), 
          .Z(n891_adj_2328)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 mux_191_Mux_4_i286_3_lut (.A(n270_adj_2670), .B(n15_adj_2524), 
         .C(index_i[4]), .Z(n286_adj_2532)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_4_i286_3_lut.init = 16'hcaca;
    LUT4 mux_191_Mux_5_i700_3_lut (.A(n460_adj_2726), .B(n26699), .C(index_i[4]), 
         .Z(n700_adj_2497)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_5_i700_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_11_i638_4_lut_4_lut (.A(n26375), .B(index_q[5]), .C(index_q[6]), 
         .D(n26412), .Z(n638)) /* synthesis lut_function=(A (B (C (D))+!B !(C))+!A (B ((D)+!C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_11_i638_4_lut_4_lut.init = 16'hc707;
    LUT4 i19270_3_lut (.A(n396), .B(n26608), .C(index_i[3]), .Z(n21590)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19270_3_lut.init = 16'hcaca;
    LUT4 i19268_3_lut (.A(n26687), .B(n26706), .C(index_i[3]), .Z(n21588)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19268_3_lut.init = 16'hcaca;
    LUT4 mux_191_Mux_4_i94_3_lut (.A(n61_adj_2522), .B(n26593), .C(index_i[4]), 
         .Z(n94_adj_2529)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_4_i94_3_lut.init = 16'hcaca;
    LUT4 i19267_3_lut (.A(n26688), .B(n26710), .C(index_i[3]), .Z(n21587)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19267_3_lut.init = 16'hcaca;
    L6MUX21 i24144 (.D0(n25934), .D1(n25931), .SD(index_i[8]), .Z(n25935));
    LUT4 mux_192_Mux_7_i333_3_lut (.A(n26571), .B(n26521), .C(index_q[3]), 
         .Z(n333)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_7_i333_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_7_i348_3_lut (.A(n29187), .B(n29189), .C(index_q[3]), 
         .Z(n348_adj_2636)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_7_i348_3_lut.init = 16'hcaca;
    LUT4 n17750_bdd_4_lut_then_4_lut (.A(index_q[3]), .B(index_q[4]), .C(index_q[1]), 
         .D(index_q[2]), .Z(n26818)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B+(C (D)+!C !(D)))) */ ;
    defparam n17750_bdd_4_lut_then_4_lut.init = 16'hf44f;
    LUT4 mux_192_Mux_0_i731_3_lut_4_lut (.A(n26567), .B(index_q[2]), .C(index_q[3]), 
         .D(n29187), .Z(n731_adj_2437)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_0_i731_3_lut_4_lut.init = 16'h4f40;
    PFUMX i19901 (.BLUT(n158_adj_2624), .ALUT(n189_adj_2727), .C0(index_q[5]), 
          .Z(n22240));
    LUT4 i22222_3_lut_rep_392_4_lut (.A(n26478), .B(index_i[5]), .C(index_i[8]), 
         .D(n1021), .Z(n26352)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i22222_3_lut_rep_392_4_lut.init = 16'hf808;
    LUT4 i19064_3_lut_4_lut (.A(n26567), .B(index_q[2]), .C(index_q[3]), 
         .D(n29196), .Z(n21384)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19064_3_lut_4_lut.init = 16'hf404;
    LUT4 mux_192_Mux_7_i397_3_lut (.A(n29187), .B(n26571), .C(index_q[3]), 
         .Z(n397_adj_2635)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_7_i397_3_lut.init = 16'hcaca;
    LUT4 i21780_3_lut (.A(n21728), .B(n21729), .C(index_q[4]), .Z(n21730)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21780_3_lut.init = 16'hcaca;
    LUT4 i23394_then_4_lut (.A(index_q[0]), .B(index_q[4]), .C(index_q[1]), 
         .D(index_q[3]), .Z(n26747)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam i23394_then_4_lut.init = 16'h3c69;
    PFUMX i24142 (.BLUT(n25933), .ALUT(n25932), .C0(index_i[7]), .Z(n25934));
    PFUMX i23095 (.BLUT(n24765), .ALUT(n26519), .C0(index_i[4]), .Z(n24766));
    LUT4 mux_191_Mux_5_i891_3_lut (.A(n875_adj_2662), .B(n379_adj_2365), 
         .C(index_i[4]), .Z(n891_adj_2503)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_5_i891_3_lut.init = 16'hcaca;
    LUT4 mux_191_Mux_5_i860_3_lut (.A(n15_adj_2519), .B(n859_adj_2661), 
         .C(index_i[4]), .Z(n860_adj_2502)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_5_i860_3_lut.init = 16'hcaca;
    LUT4 i21788_3_lut (.A(n21593), .B(n21594), .C(index_i[4]), .Z(n21595)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21788_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_4_lut_adj_77 (.A(n26375), .B(index_q[5]), .C(index_q[8]), 
         .D(n19545), .Z(n19899)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_3_lut_4_lut_adj_77.init = 16'hfff8;
    LUT4 i23394_else_4_lut (.A(index_q[0]), .B(index_q[4]), .C(index_q[1]), 
         .D(index_q[3]), .Z(n26746)) /* synthesis lut_function=(!(A (B (C)+!B !(C (D)+!C !(D)))+!A (B ((D)+!C)+!B !((D)+!C)))) */ ;
    defparam i23394_else_4_lut.init = 16'h394b;
    LUT4 mux_191_Mux_5_i636_4_lut (.A(n157_adj_2419), .B(n26436), .C(index_i[4]), 
         .D(index_i[3]), .Z(n636_adj_2495)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_5_i636_4_lut.init = 16'h3aca;
    PFUMX i19413 (.BLUT(n21731), .ALUT(n21732), .C0(index_q[4]), .Z(n21733));
    LUT4 i21791_3_lut (.A(n17573), .B(n17574), .C(index_i[4]), .Z(n17575)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21791_3_lut.init = 16'hcaca;
    LUT4 n17750_bdd_4_lut_else_4_lut (.A(index_q[3]), .B(index_q[4]), .C(index_q[1]), 
         .D(index_q[2]), .Z(n26817)) /* synthesis lut_function=(!(A (B (D)+!B ((D)+!C))+!A !(B+!((D)+!C)))) */ ;
    defparam n17750_bdd_4_lut_else_4_lut.init = 16'h44fc;
    LUT4 i22218_3_lut_rep_393_4_lut (.A(n26476), .B(index_q[5]), .C(index_q[8]), 
         .D(n1021_adj_2728), .Z(n26353)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i22218_3_lut_rep_393_4_lut.init = 16'hf808;
    PFUMX i24139 (.BLUT(n25930), .ALUT(n22942), .C0(index_i[7]), .Z(n25931));
    LUT4 mux_191_Mux_5_i507_3_lut (.A(n491_adj_2389), .B(n506_adj_2653), 
         .C(index_i[4]), .Z(n507_adj_2488)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_5_i507_3_lut.init = 16'hcaca;
    LUT4 mux_191_Mux_5_i476_3_lut (.A(n460_adj_2726), .B(n475_adj_2399), 
         .C(index_i[4]), .Z(n476_adj_2487)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_5_i476_3_lut.init = 16'hcaca;
    LUT4 i19265_3_lut (.A(n29177), .B(n26710), .C(index_i[3]), .Z(n21585)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19265_3_lut.init = 16'hcaca;
    LUT4 mux_191_Mux_5_i413_3_lut (.A(n397_adj_2647), .B(n251_adj_2548), 
         .C(index_i[4]), .Z(n413_adj_2485)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_5_i413_3_lut.init = 16'hcaca;
    LUT4 i19261_3_lut (.A(n26700), .B(n26710), .C(index_i[3]), .Z(n21581)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19261_3_lut.init = 16'hcaca;
    L6MUX21 i24131 (.D0(n25916), .D1(n25913), .SD(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2127[4]));
    PFUMX i20460 (.BLUT(n22795), .ALUT(n22796), .C0(index_q[4]), .Z(n22799));
    LUT4 i19259_3_lut (.A(n26707), .B(n29180), .C(index_i[3]), .Z(n21579)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19259_3_lut.init = 16'hcaca;
    PFUMX i24129 (.BLUT(n25915), .ALUT(n25914), .C0(index_i[8]), .Z(n25916));
    LUT4 i20218_3_lut_3_lut_4_lut (.A(n26430), .B(index_q[3]), .C(n316_adj_2729), 
         .D(index_q[4]), .Z(n22557)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20218_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 i15435_3_lut (.A(n17583), .B(n17584), .C(index_i[4]), .Z(n17585)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15435_3_lut.init = 16'hcaca;
    LUT4 i21376_3_lut (.A(n21578), .B(n21579), .C(index_i[4]), .Z(n21580)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21376_3_lut.init = 16'hcaca;
    LUT4 mux_191_Mux_5_i125_3_lut (.A(n109_adj_2730), .B(n124_adj_2540), 
         .C(index_i[4]), .Z(n125_adj_2482)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_5_i125_3_lut.init = 16'hcaca;
    LUT4 i19256_3_lut (.A(n29171), .B(n26714), .C(index_q[3]), .Z(n21576)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19256_3_lut.init = 16'hcaca;
    LUT4 mux_191_Mux_5_i94_3_lut (.A(n653_adj_2644), .B(n635_adj_2731), 
         .C(index_i[4]), .Z(n94_adj_2481)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_5_i94_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_1_i763_3_lut_4_lut (.A(index_q[4]), .B(index_q[3]), 
         .C(n26819), .D(n26543), .Z(n763_adj_2438)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_1_i763_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i19255_3_lut (.A(n325), .B(n204_adj_2732), .C(index_q[3]), .Z(n21575)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19255_3_lut.init = 16'hcaca;
    PFUMX i20461 (.BLUT(n22797), .ALUT(n22798), .C0(index_q[4]), .Z(n22800));
    LUT4 i20352_3_lut (.A(n308), .B(n29174), .C(index_i[3]), .Z(n22691)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20352_3_lut.init = 16'hcaca;
    LUT4 i20351_3_lut (.A(n619), .B(n26652), .C(index_i[3]), .Z(n22690)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20351_3_lut.init = 16'hcaca;
    LUT4 i11947_2_lut (.A(index_q[1]), .B(index_q[3]), .Z(n541_adj_2253)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i11947_2_lut.init = 16'h1111;
    LUT4 mux_192_Mux_10_i317_3_lut_3_lut_4_lut (.A(n26430), .B(index_q[3]), 
         .C(n26457), .D(index_q[4]), .Z(n317_adj_2733)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_10_i317_3_lut_3_lut_4_lut.init = 16'hf011;
    PFUMX i20268 (.BLUT(n158_adj_2614), .ALUT(n189_adj_2464), .C0(index_q[5]), 
          .Z(n22607));
    LUT4 i20350_3_lut (.A(n26604), .B(n26650), .C(index_i[3]), .Z(n22689)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20350_3_lut.init = 16'hcaca;
    LUT4 i20349_3_lut (.A(n29174), .B(n29194), .C(index_i[3]), .Z(n22688)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20349_3_lut.init = 16'hcaca;
    PFUMX i20269 (.BLUT(n221_adj_2734), .ALUT(n21103), .C0(index_q[5]), 
          .Z(n22608));
    PFUMX i20467 (.BLUT(n22802), .ALUT(n22803), .C0(index_q[4]), .Z(n22806));
    LUT4 i15437_4_lut (.A(index_q[0]), .B(index_q[4]), .C(index_q[1]), 
         .D(n26585), .Z(n286_adj_2735)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i15437_4_lut.init = 16'hccc8;
    PFUMX i20468 (.BLUT(n22804), .ALUT(n22805), .C0(index_q[4]), .Z(n22807));
    PFUMX i20270 (.BLUT(n286_adj_2612), .ALUT(n317_adj_2611), .C0(index_q[5]), 
          .Z(n22609));
    LUT4 i21808_3_lut (.A(n21095), .B(n26768), .C(index_q[4]), .Z(n21097)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21808_3_lut.init = 16'hcaca;
    PFUMX i20271 (.BLUT(n349_adj_2736), .ALUT(n21106), .C0(index_q[5]), 
          .Z(n22610));
    PFUMX i20716 (.BLUT(n844_adj_2737), .ALUT(n11815), .C0(index_q[4]), 
          .Z(n23055));
    LUT4 i18688_3_lut (.A(n29171), .B(n325), .C(index_q[3]), .Z(n21008)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18688_3_lut.init = 16'hcaca;
    LUT4 i22339_2_lut_rep_585 (.A(index_i[1]), .B(index_i[2]), .Z(n26545)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i22339_2_lut_rep_585.init = 16'h9999;
    LUT4 n442_bdd_2_lut_23551_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[3]), 
         .Z(n25232)) /* synthesis lut_function=(A (B+(C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n442_bdd_2_lut_23551_3_lut.init = 16'hf9f9;
    LUT4 index_i_8__bdd_3_lut_24177_then_4_lut (.A(index_i[4]), .B(index_i[6]), 
         .C(index_i[5]), .D(n26419), .Z(n26821)) /* synthesis lut_function=(!(A (B (C+(D)))+!A (B (C)))) */ ;
    defparam index_i_8__bdd_3_lut_24177_then_4_lut.init = 16'h373f;
    PFUMX i24126 (.BLUT(n25912), .ALUT(n22395), .C0(index_i[8]), .Z(n25913));
    LUT4 mux_192_Mux_0_i589_3_lut (.A(n29189), .B(n931), .C(index_q[3]), 
         .Z(n589)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_0_i589_3_lut.init = 16'hcaca;
    PFUMX i20272 (.BLUT(n413_adj_2610), .ALUT(n21109), .C0(index_q[5]), 
          .Z(n22611));
    LUT4 i20631_3_lut_4_lut_4_lut (.A(n26472), .B(index_i[4]), .C(index_i[5]), 
         .D(n26419), .Z(n22970)) /* synthesis lut_function=(A ((C+!(D))+!B)+!A (B (C+!(D))+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20631_3_lut_4_lut_4_lut.init = 16'he3ef;
    LUT4 i22438_2_lut (.A(index_i[5]), .B(index_i[4]), .Z(n22013)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i22438_2_lut.init = 16'heeee;
    PFUMX i20273 (.BLUT(n21112), .ALUT(n507_adj_2738), .C0(index_q[5]), 
          .Z(n22612));
    LUT4 i18769_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21089)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A !(B (D)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18769_3_lut_3_lut_4_lut.init = 16'ha955;
    LUT4 mux_192_Mux_0_i812_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n812_adj_2441)) /* synthesis lut_function=(A (B (C+(D))+!B !(C))+!A (B (D)+!B !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_0_i812_3_lut_4_lut_4_lut_4_lut.init = 16'hcf92;
    PFUMX i20274 (.BLUT(n21115), .ALUT(n573_adj_2739), .C0(index_q[5]), 
          .Z(n22613));
    LUT4 mux_191_Mux_6_i627_3_lut_4_lut_3_lut_rep_747 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26707)) /* synthesis lut_function=(A ((C)+!B)+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_6_i627_3_lut_4_lut_3_lut_rep_747.init = 16'he6e6;
    PFUMX i20275 (.BLUT(n605_adj_2608), .ALUT(n21118), .C0(index_q[5]), 
          .Z(n22614));
    PFUMX i20778 (.BLUT(n844_adj_2740), .ALUT(n12012), .C0(index_i[4]), 
          .Z(n23117));
    LUT4 i1_3_lut_adj_78 (.A(index_i[0]), .B(index_i[4]), .C(index_i[2]), 
         .Z(n20376)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i1_3_lut_adj_78.init = 16'hfefe;
    PFUMX i20276 (.BLUT(n669_adj_2607), .ALUT(n700_adj_2543), .C0(index_q[5]), 
          .Z(n22615));
    LUT4 mux_192_Mux_3_i924_3_lut (.A(n908_adj_2643), .B(index_q[0]), .C(index_q[4]), 
         .Z(n924_adj_2477)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_3_i924_3_lut.init = 16'hcaca;
    PFUMX i20277 (.BLUT(n732_adj_2605), .ALUT(n763_adj_2741), .C0(index_q[5]), 
          .Z(n22616));
    LUT4 n315_bdd_3_lut_23235 (.A(n29195), .B(index_q[3]), .C(n26725), 
         .Z(n24908)) /* synthesis lut_function=(A (B+(C))+!A !(B+!(C))) */ ;
    defparam n315_bdd_3_lut_23235.init = 16'hb8b8;
    LUT4 mux_191_Mux_5_i683_3_lut_4_lut_4_lut_3_lut_rep_748 (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[2]), .Z(n26708)) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_5_i683_3_lut_4_lut_4_lut_3_lut_rep_748.init = 16'h6b6b;
    CCU2D add_372_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(quarter_wave_sample_register_q[0]), .B1(quarter_wave_sample_register_q[1]), 
          .C1(GND_net), .D1(GND_net), .COUT(n17338));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(80[29:60])
    defparam add_372_1.INIT0 = 16'hF000;
    defparam add_372_1.INIT1 = 16'ha666;
    defparam add_372_1.INJECT1_0 = "NO";
    defparam add_372_1.INJECT1_1 = "NO";
    LUT4 mux_191_Mux_4_i70_3_lut_3_lut_rep_749 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26709)) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_4_i70_3_lut_3_lut_rep_749.init = 16'h6a6a;
    LUT4 mux_192_Mux_0_i526_3_lut (.A(n29171), .B(n29197), .C(index_q[3]), 
         .Z(n526_adj_2252)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_0_i526_3_lut.init = 16'hcaca;
    LUT4 mux_191_Mux_0_i93_3_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .Z(n93_adj_2547)) /* synthesis lut_function=(A (B)+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_0_i93_3_lut_3_lut.init = 16'h9c9c;
    LUT4 i8238_2_lut_rep_586 (.A(index_i[1]), .B(index_i[2]), .Z(n26546)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i8238_2_lut_rep_586.init = 16'h8888;
    LUT4 i21916_3_lut (.A(n924_adj_2742), .B(n955_adj_2678), .C(index_q[5]), 
         .Z(n22123)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21916_3_lut.init = 16'hcaca;
    LUT4 i9549_2_lut_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[3]), 
         .Z(n11995)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9549_2_lut_3_lut.init = 16'h8080;
    L6MUX21 i20279 (.D0(n860_adj_2603), .D1(n891_adj_2598), .SD(index_q[5]), 
            .Z(n22618));
    LUT4 i18703_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21023)) /* synthesis lut_function=(A (B (C (D))+!B !(C (D)))+!A !(B (D)+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18703_3_lut_4_lut_4_lut.init = 16'h9366;
    LUT4 index_q_8__bdd_3_lut_then_4_lut (.A(index_q[4]), .B(index_q[6]), 
         .C(index_q[5]), .D(n26410), .Z(n26824)) /* synthesis lut_function=(!(A (B (C+(D)))+!A (B (C)))) */ ;
    defparam index_q_8__bdd_3_lut_then_4_lut.init = 16'h373f;
    LUT4 i22196_3_lut (.A(n24923), .B(n22112), .C(index_q[6]), .Z(n22126)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22196_3_lut.init = 16'hcaca;
    LUT4 mux_191_Mux_6_i467_3_lut_3_lut_3_lut_rep_750 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26710)) /* synthesis lut_function=(!(A (B)+!A (B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_6_i467_3_lut_3_lut_3_lut_rep_750.init = 16'h3636;
    LUT4 i11691_2_lut_rep_475_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[0]), 
         .Z(n26435)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11691_2_lut_rep_475_3_lut.init = 16'h7070;
    LUT4 mux_191_Mux_6_i475_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n475_adj_2697)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A !(B (C+(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_6_i475_3_lut_4_lut_4_lut.init = 16'h9936;
    LUT4 i1_3_lut_4_lut_adj_79 (.A(index_i[1]), .B(index_i[2]), .C(index_i[5]), 
         .D(n26595), .Z(n20003)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i1_3_lut_4_lut_adj_79.init = 16'hfff8;
    LUT4 i11461_2_lut_rep_491_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[3]), 
         .Z(n26451)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11461_2_lut_rep_491_3_lut.init = 16'hf8f8;
    LUT4 i20217_3_lut_4_lut (.A(n26538), .B(index_q[3]), .C(index_q[4]), 
         .D(n285_adj_2269), .Z(n22556)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20217_3_lut_4_lut.init = 16'hfe0e;
    LUT4 i11692_2_lut_rep_478_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[0]), 
         .Z(n26438)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11692_2_lut_rep_478_3_lut.init = 16'h8080;
    LUT4 i11658_3_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[3]), 
         .Z(n11010)) /* synthesis lut_function=(!((B (C))+!A)) */ ;
    defparam i11658_3_lut.init = 16'h2a2a;
    LUT4 mux_192_Mux_4_i573_3_lut_4_lut_4_lut_4_lut (.A(n26538), .B(index_q[3]), 
         .C(n26526), .D(index_q[4]), .Z(n573)) /* synthesis lut_function=(!(A (B (D)+!B ((D)+!C))+!A (B (D)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_4_i573_3_lut_4_lut_4_lut_4_lut.init = 16'h11fc;
    LUT4 n124_bdd_3_lut_22850_4_lut (.A(n26538), .B(index_q[3]), .C(index_q[4]), 
         .D(n124_adj_2500), .Z(n24455)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n124_bdd_3_lut_22850_4_lut.init = 16'hf101;
    LUT4 mux_192_Mux_10_i125_3_lut_4_lut_4_lut (.A(n26538), .B(index_q[3]), 
         .C(index_q[4]), .D(n29190), .Z(n125_adj_2480)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B (C (D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_10_i125_3_lut_4_lut_4_lut.init = 16'h3efe;
    LUT4 mux_192_Mux_2_i573_3_lut_3_lut_4_lut (.A(n26538), .B(index_q[3]), 
         .C(n557), .D(index_q[4]), .Z(n573_adj_2739)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_2_i573_3_lut_3_lut_4_lut.init = 16'h11f0;
    L6MUX21 i20303 (.D0(n22640), .D1(n22641), .SD(index_i[5]), .Z(n22642));
    LUT4 i11423_2_lut_rep_433_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n26393)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11423_2_lut_rep_433_3_lut_4_lut.init = 16'hf8f0;
    LUT4 mux_191_Mux_8_i491_3_lut_3_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n491_adj_2687)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_8_i491_3_lut_3_lut_3_lut_4_lut.init = 16'h7870;
    LUT4 mux_192_Mux_3_i573_3_lut_3_lut_4_lut (.A(n26538), .B(index_q[3]), 
         .C(n557_adj_2660), .D(index_q[4]), .Z(n573_adj_2472)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_3_i573_3_lut_3_lut_4_lut.init = 16'h11f0;
    LUT4 i11526_2_lut_rep_587 (.A(index_i[2]), .B(index_i[3]), .Z(n26547)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11526_2_lut_rep_587.init = 16'h8888;
    LUT4 i20206_3_lut_3_lut_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[4]), .D(index_i[1]), .Z(n22545)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20206_3_lut_3_lut_3_lut_4_lut.init = 16'h878f;
    LUT4 mux_192_Mux_6_i653_3_lut (.A(n26718), .B(n676), .C(index_q[3]), 
         .Z(n653_adj_2514)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_6_i653_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_6_i668_3_lut (.A(n660), .B(n29183), .C(index_q[3]), 
         .Z(n668_adj_2579)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_6_i668_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_6_i684_3_lut (.A(n26521), .B(n29200), .C(index_q[3]), 
         .Z(n684)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_6_i684_3_lut.init = 16'hcaca;
    LUT4 i11829_2_lut_rep_466_3_lut (.A(index_q[1]), .B(index_q[2]), .C(index_q[0]), 
         .Z(n26426)) /* synthesis lut_function=(A (B+!(C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11829_2_lut_rep_466_3_lut.init = 16'h8f8f;
    LUT4 i19051_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21371)) /* synthesis lut_function=(A (B (C)+!B (C (D)+!C !(D)))+!A !(B (C+!(D))+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19051_3_lut_4_lut_4_lut.init = 16'ha593;
    LUT4 i18746_3_lut_3_lut_4_lut (.A(index_q[1]), .B(index_q[2]), .C(index_q[3]), 
         .D(index_q[0]), .Z(n21066)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18746_3_lut_3_lut_4_lut.init = 16'hf80f;
    LUT4 i11734_2_lut_rep_510_3_lut (.A(index_i[2]), .B(index_i[3]), .C(index_i[1]), 
         .Z(n26470)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11734_2_lut_rep_510_3_lut.init = 16'h8080;
    LUT4 i22128_3_lut (.A(n22619), .B(n25469), .C(index_q[6]), .Z(n22628)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22128_3_lut.init = 16'hcaca;
    LUT4 i11439_2_lut_rep_434_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[4]), .D(n26548), .Z(n26394)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11439_2_lut_rep_434_3_lut_4_lut.init = 16'hf8f0;
    LUT4 index_q_8__bdd_3_lut_else_4_lut (.A(n26477), .B(index_q[4]), .C(index_q[6]), 
         .D(index_q[5]), .Z(n26823)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;
    defparam index_q_8__bdd_3_lut_else_4_lut.init = 16'hf080;
    LUT4 n572_bdd_3_lut_24005_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n25630)) /* synthesis lut_function=(A (B (C+(D)))+!A (B ((D)+!C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n572_bdd_3_lut_24005_4_lut.init = 16'hcc94;
    PFUMX i24503 (.BLUT(n26799), .ALUT(n26800), .C0(index_q[0]), .Z(n26801));
    LUT4 i11451_2_lut_3_lut_4_lut (.A(n26526), .B(n26584), .C(index_q[6]), 
         .D(index_q[5]), .Z(n254_adj_2383)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11451_2_lut_3_lut_4_lut.init = 16'hfef0;
    LUT4 i21953_3_lut (.A(n26810), .B(n62_adj_2743), .C(index_q[5]), .Z(n22605)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21953_3_lut.init = 16'hcaca;
    LUT4 i19208_3_lut (.A(n26652), .B(n308), .C(index_i[3]), .Z(n21528)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19208_3_lut.init = 16'hcaca;
    LUT4 i19205_3_lut (.A(n26652), .B(n70), .C(index_i[3]), .Z(n21525)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19205_3_lut.init = 16'hcaca;
    LUT4 i19204_3_lut (.A(n26648), .B(n308), .C(index_i[3]), .Z(n21524)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19204_3_lut.init = 16'hcaca;
    PFUMX mux_191_Mux_7_i190 (.BLUT(n21526), .ALUT(n173_adj_2744), .C0(index_i[5]), 
          .Z(n190_adj_2717)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    PFUMX i24094 (.BLUT(n25867), .ALUT(n25865), .C0(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_2142[10]));
    LUT4 mux_191_Mux_2_i491_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n491_adj_2745)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A !(B (C)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_2_i491_3_lut_4_lut_4_lut.init = 16'h6a5a;
    LUT4 i19708_1_lut_2_lut (.A(index_i[2]), .B(index_i[3]), .Z(n22047)) /* synthesis lut_function=(!(A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19708_1_lut_2_lut.init = 16'h7777;
    LUT4 mux_191_Mux_5_i460_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n460_adj_2726)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A !(B (C)+!B !(C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_5_i460_3_lut_4_lut_4_lut.init = 16'h6b5a;
    LUT4 mux_191_Mux_7_i173_3_lut (.A(n26691), .B(n70), .C(index_i[3]), 
         .Z(n173_adj_2744)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_7_i173_3_lut.init = 16'hcaca;
    LUT4 i11467_2_lut_rep_447_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[4]), .D(n26647), .Z(n26407)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11467_2_lut_rep_447_3_lut_4_lut.init = 16'hf8f0;
    LUT4 mux_191_Mux_7_i924_3_lut_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[4]), .D(n26647), .Z(n924_adj_2443)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_7_i924_3_lut_3_lut_4_lut.init = 16'h878f;
    LUT4 i11589_2_lut_rep_588 (.A(index_i[0]), .B(index_i[1]), .Z(n26548)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11589_2_lut_rep_588.init = 16'h8888;
    LUT4 mux_192_Mux_1_i986_3_lut (.A(n29187), .B(n26721), .C(index_q[3]), 
         .Z(n986_adj_2746)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_1_i986_3_lut.init = 16'hcaca;
    LUT4 mux_191_Mux_6_i635_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n635_adj_2731)) /* synthesis lut_function=(A (B (C+(D))+!B !(D))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_6_i635_3_lut_4_lut.init = 16'hcce6;
    LUT4 mux_191_Mux_1_i301_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n301_adj_2656)) /* synthesis lut_function=(A (B (C+(D))+!B !(D))+!A !(B (C+(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_1_i301_3_lut_4_lut_4_lut.init = 16'h99b6;
    LUT4 n45_bdd_3_lut_4_lut_4_lut_4_lut_adj_80 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n25263)) /* synthesis lut_function=(A (B (C+!(D))+!B ((D)+!C))+!A (B (C (D)+!C !(D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n45_bdd_3_lut_4_lut_4_lut_4_lut_adj_80.init = 16'hf38f;
    LUT4 i12485_2_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(n26635), 
         .D(index_i[2]), .Z(n15074)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i12485_2_lut_3_lut_4_lut.init = 16'hf080;
    LUT4 n301_bdd_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n25260)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+!(D)))+!A (B (D)+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n301_bdd_3_lut_4_lut_4_lut_4_lut.init = 16'h30f7;
    LUT4 mux_191_Mux_6_i812_3_lut_4_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n812_adj_2650)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(D))+!A !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_6_i812_3_lut_4_lut_3_lut_4_lut.init = 16'h7780;
    LUT4 mux_191_Mux_3_i1002_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n19612)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (D))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_3_i1002_3_lut_3_lut_4_lut.init = 16'hf708;
    LUT4 i1_3_lut_rep_518_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(n26595), .Z(n26478)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i1_3_lut_rep_518_4_lut.init = 16'hfff8;
    LUT4 mux_191_Mux_8_i526_3_lut_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n526_adj_2366)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_8_i526_3_lut_3_lut_3_lut_4_lut.init = 16'h0f70;
    PFUMX mux_191_Mux_8_i764 (.BLUT(n716_adj_2747), .ALUT(n732_adj_2591), 
          .C0(n22013), .Z(n764_adj_2390)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 mux_191_Mux_6_i781_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n781_adj_2526)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A (B (C (D)+!C !(D))+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_6_i781_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hc837;
    LUT4 i21977_3_lut (.A(n286_adj_2600), .B(n317), .C(index_i[5]), .Z(n22969)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21977_3_lut.init = 16'hcaca;
    LUT4 mux_191_Mux_6_i860_3_lut_3_lut (.A(n26388), .B(index_i[4]), .C(n844), 
         .Z(n860_adj_2702)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam mux_191_Mux_6_i860_3_lut_3_lut.init = 16'h7474;
    PFUMX mux_191_Mux_8_i574 (.BLUT(n542_adj_2367), .ALUT(n11946), .C0(index_i[5]), 
          .Z(n574_adj_2388)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 mux_192_Mux_5_i15_3_lut (.A(n26719), .B(n29181), .C(index_q[3]), 
         .Z(n15_adj_2492)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_5_i15_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_477_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n26437)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i1_2_lut_rep_477_3_lut_4_lut.init = 16'h8000;
    LUT4 mux_192_Mux_6_i875_3_lut_4_lut (.A(n26569), .B(index_q[2]), .C(index_q[3]), 
         .D(n29192), .Z(n875_adj_2571)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_6_i875_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_192_Mux_5_i397_3_lut (.A(n26724), .B(n204_adj_2732), .C(index_q[3]), 
         .Z(n397_adj_2505)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_5_i397_3_lut.init = 16'hcaca;
    LUT4 i11471_2_lut_rep_437_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n26397)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11471_2_lut_rep_437_3_lut_4_lut.init = 16'hf080;
    LUT4 mux_192_Mux_5_i506_3_lut (.A(n29176), .B(n29163), .C(index_q[3]), 
         .Z(n506_adj_2458)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_5_i506_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_4_i15_3_lut (.A(n29163), .B(n931), .C(index_q[3]), 
         .Z(n15_adj_2469)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_4_i15_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_4_i61_3_lut (.A(n29197), .B(n29175), .C(index_q[3]), 
         .Z(n61)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_4_i61_3_lut.init = 16'hcaca;
    L6MUX21 i22687 (.D0(n24249), .D1(n26340), .SD(index_i[6]), .Z(n24250));
    LUT4 mux_192_Mux_5_i939_3_lut_3_lut_4_lut (.A(n26569), .B(index_q[2]), 
         .C(n954_adj_2429), .D(index_q[4]), .Z(n939_adj_2357)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_5_i939_3_lut_3_lut_4_lut.init = 16'hf077;
    LUT4 mux_192_Mux_5_i859_3_lut (.A(n250), .B(n26719), .C(index_q[3]), 
         .Z(n859_adj_2493)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_5_i859_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_5_i875_3_lut (.A(n26521), .B(n29187), .C(index_q[3]), 
         .Z(n875_adj_2490)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_5_i875_3_lut.init = 16'hcaca;
    LUT4 mux_191_Mux_8_i172_rep_28_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n70_adj_2255)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_8_i172_rep_28_3_lut_3_lut.init = 16'h7c7c;
    LUT4 mux_191_Mux_9_i316_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n316_adj_2385)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C+(D)))+!A (B (C (D)+!C !(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_9_i316_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h3ff8;
    PFUMX i24092 (.BLUT(n21215), .ALUT(n25863), .C0(index_q[7]), .Z(n25864));
    LUT4 mux_192_Mux_4_i270_3_lut (.A(n29170), .B(n29176), .C(index_q[3]), 
         .Z(n270_adj_2468)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_4_i270_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_4_i348_3_lut (.A(n29164), .B(n29171), .C(index_q[3]), 
         .Z(n348_adj_2309)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_4_i348_3_lut.init = 16'hcaca;
    LUT4 i11499_2_lut_rep_526_3_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .Z(n26486)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11499_2_lut_rep_526_3_lut.init = 16'hf8f8;
    LUT4 mux_192_Mux_4_i684_3_lut (.A(n676), .B(n660), .C(index_q[3]), 
         .Z(n684_adj_2461)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_4_i684_3_lut.init = 16'hcaca;
    LUT4 i19956_3_lut (.A(n22289), .B(n22290), .C(index_q[7]), .Z(n22295)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19956_3_lut.init = 16'hcaca;
    PFUMX i24086 (.BLUT(n25857), .ALUT(n25855), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2127[10]));
    LUT4 i19951_3_lut (.A(n22279), .B(n22280), .C(index_q[6]), .Z(n22290)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19951_3_lut.init = 16'hcaca;
    LUT4 i20086_3_lut (.A(n22419), .B(n22420), .C(index_i[7]), .Z(n22425)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20086_3_lut.init = 16'hcaca;
    PFUMX i19224 (.BLUT(n21542), .ALUT(n21543), .C0(index_q[5]), .Z(n21544));
    L6MUX21 i19771 (.D0(n21568), .D1(n21571), .SD(index_q[5]), .Z(n22110));
    LUT4 i20081_3_lut (.A(n22409), .B(n22410), .C(index_i[6]), .Z(n22420)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20081_3_lut.init = 16'hcaca;
    LUT4 i20146_3_lut (.A(n22477), .B(n22478), .C(index_i[7]), .Z(n22485)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20146_3_lut.init = 16'hcaca;
    LUT4 i20139_3_lut (.A(n22463), .B(n25276), .C(index_i[6]), .Z(n22478)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20139_3_lut.init = 16'hcaca;
    LUT4 mux_191_Mux_4_i1002_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n1002_adj_2720)) /* synthesis lut_function=(A (B (C (D))+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_4_i1002_3_lut_3_lut_4_lut.init = 16'hf007;
    LUT4 n285_bdd_3_lut_adj_81 (.A(n29195), .B(n26734), .C(index_q[3]), 
         .Z(n24911)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n285_bdd_3_lut_adj_81.init = 16'hacac;
    L6MUX21 i19775 (.D0(n21577), .D1(n17542), .SD(index_q[5]), .Z(n22114));
    L6MUX21 i19776 (.D0(n21010), .D1(n11827), .SD(index_q[5]), .Z(n22115));
    LUT4 i19498_3_lut_3_lut_4_lut (.A(n26569), .B(index_q[2]), .C(n1001), 
         .D(index_q[3]), .Z(n21818)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19498_3_lut_3_lut_4_lut.init = 16'hf077;
    LUT4 i21989_3_lut (.A(n924_adj_2748), .B(n955), .C(index_i[5]), .Z(n22937)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21989_3_lut.init = 16'hcaca;
    PFUMX i19778 (.BLUT(n542_adj_2584), .ALUT(n573_adj_2749), .C0(index_q[5]), 
          .Z(n22117));
    LUT4 i20148_3_lut (.A(n22481), .B(n22482), .C(index_i[7]), .Z(n22487)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20148_3_lut.init = 16'hcaca;
    LUT4 i20142_3_lut (.A(n22469), .B(n22470), .C(index_i[6]), .Z(n22481)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20142_3_lut.init = 16'hcaca;
    PFUMX i24084 (.BLUT(n21206), .ALUT(n25853), .C0(index_i[7]), .Z(n25854));
    PFUMX i19779 (.BLUT(n605_adj_2750), .ALUT(n636_adj_2751), .C0(index_q[5]), 
          .Z(n22118));
    PFUMX i19780 (.BLUT(n669_adj_2580), .ALUT(n700_adj_2270), .C0(index_q[5]), 
          .Z(n22119));
    LUT4 i20380_3_lut (.A(n22711), .B(n22712), .C(index_q[7]), .Z(n22719)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20380_3_lut.init = 16'hcaca;
    LUT4 i20373_3_lut (.A(n22697), .B(n25596), .C(index_q[6]), .Z(n22712)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20373_3_lut.init = 16'hcaca;
    LUT4 i20382_3_lut (.A(n22715), .B(n22716), .C(index_q[7]), .Z(n22721)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20382_3_lut.init = 16'hcaca;
    LUT4 i20376_3_lut (.A(n25635), .B(n22704), .C(index_q[6]), .Z(n22715)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20376_3_lut.init = 16'hcaca;
    PFUMX i19781 (.BLUT(n732), .ALUT(n21016), .C0(index_q[5]), .Z(n22120));
    LUT4 mux_192_Mux_2_i731_3_lut_3_lut_4_lut (.A(index_q[2]), .B(index_q[3]), 
         .C(index_q[1]), .D(index_q[0]), .Z(n731_adj_2604)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(B (C)+!B !(C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_2_i731_3_lut_3_lut_4_lut.init = 16'h69f0;
    LUT4 i19330_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21650)) /* synthesis lut_function=(!(A (B)+!A (B (C+(D))+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19330_3_lut_3_lut_4_lut.init = 16'h3326;
    LUT4 i22427_2_lut (.A(index_q[3]), .B(index_q[2]), .Z(n22054)) /* synthesis lut_function=(A+!(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i22427_2_lut.init = 16'hbbbb;
    PFUMX i19782 (.BLUT(n797_adj_2576), .ALUT(n828_adj_2575), .C0(index_q[5]), 
          .Z(n22121));
    PFUMX i24071 (.BLUT(n25828), .ALUT(n1022_adj_2382), .C0(index_i[9]), 
          .Z(quarter_wave_sample_register_i_15__N_2127[12]));
    PFUMX i19783 (.BLUT(n860_adj_2711), .ALUT(n891_adj_2572), .C0(index_q[5]), 
          .Z(n22122));
    LUT4 i19976_3_lut (.A(n24445), .B(n28768), .C(index_i[7]), .Z(n22315)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19976_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_2_i653_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n653_adj_2606)) /* synthesis lut_function=(A (B (C+!(D))+!B !(D))+!A !(B (C+!(D))+!B !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_2_i653_3_lut_4_lut.init = 16'h94aa;
    LUT4 i20019_3_lut (.A(n22347), .B(n22348), .C(index_i[6]), .Z(n22358)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20019_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_6_i924_3_lut_4_lut (.A(index_q[2]), .B(index_q[3]), 
         .C(index_q[4]), .D(n908_adj_2563), .Z(n924_adj_2742)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_6_i924_3_lut_4_lut.init = 16'h6f60;
    LUT4 i12082_2_lut_rep_590 (.A(index_q[2]), .B(index_q[0]), .Z(n26550)) /* synthesis lut_function=(A (B)) */ ;
    defparam i12082_2_lut_rep_590.init = 16'h8888;
    L6MUX21 i20722 (.D0(n23045), .D1(n23046), .SD(index_q[5]), .Z(n23061));
    LUT4 i20115_3_lut (.A(n24543), .B(n22447), .C(index_i[7]), .Z(n22454)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20115_3_lut.init = 16'hcaca;
    LUT4 i20153_3_lut (.A(n24460), .B(n28707), .C(index_q[7]), .Z(n22492)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20153_3_lut.init = 16'hcaca;
    L6MUX21 i20723 (.D0(n23047), .D1(n23048), .SD(index_q[5]), .Z(n23062));
    LUT4 i20290_3_lut (.A(n22621), .B(n22622), .C(index_q[7]), .Z(n22629)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20290_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_3_i700_3_lut_4_lut (.A(index_q[4]), .B(index_q[3]), 
         .C(n684_adj_2752), .D(n26544), .Z(n700_adj_2473)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_3_i700_3_lut_4_lut.init = 16'hf4b0;
    PFUMX i24066 (.BLUT(n254), .ALUT(n25822), .C0(index_i[8]), .Z(n25823));
    L6MUX21 i20724 (.D0(n23049), .D1(n23050), .SD(index_q[5]), .Z(n23063));
    LUT4 n21012_bdd_3_lut (.A(n29196), .B(n29198), .C(index_q[3]), .Z(n24914)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n21012_bdd_3_lut.init = 16'hcaca;
    L6MUX21 i20725 (.D0(n23051), .D1(n23052), .SD(index_q[5]), .Z(n23064));
    L6MUX21 i20341 (.D0(n22678), .D1(n22679), .SD(index_i[5]), .Z(n22680));
    PFUMX i19239 (.BLUT(n21557), .ALUT(n21558), .C0(index_q[5]), .Z(n21559));
    L6MUX21 i20726 (.D0(n23053), .D1(n23054), .SD(index_q[5]), .Z(n23065));
    L6MUX21 i20727 (.D0(n23055), .D1(n23056), .SD(index_q[5]), .Z(n23066));
    L6MUX21 i20348 (.D0(n22685), .D1(n22686), .SD(index_i[5]), .Z(n22687));
    L6MUX21 i20728 (.D0(n23057), .D1(n23058), .SD(index_q[5]), .Z(n23067));
    L6MUX21 i20729 (.D0(n23059), .D1(n23060), .SD(index_q[5]), .Z(n23068));
    PFUMX i24061 (.BLUT(n25812), .ALUT(n1022), .C0(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_2142[12]));
    L6MUX21 i20355 (.D0(n22692), .D1(n22693), .SD(index_i[5]), .Z(n22694));
    PFUMX i20356 (.BLUT(n11916), .ALUT(n62_adj_2278), .C0(index_q[5]), 
          .Z(n22695));
    PFUMX i20357 (.BLUT(n94_adj_2561), .ALUT(n21769), .C0(index_q[5]), 
          .Z(n22696));
    LUT4 mux_191_Mux_5_i30_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n30_adj_2520)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A (B+!(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_5_i30_3_lut_4_lut.init = 16'hcc67;
    PFUMX i25959 (.BLUT(n28766), .ALUT(n28765), .C0(index_i[3]), .Z(n28767));
    L6MUX21 i20358 (.D0(n21775), .D1(n21781), .SD(index_q[5]), .Z(n22697));
    LUT4 i18974_3_lut_3_lut (.A(n26388), .B(index_i[4]), .C(n46_adj_2715), 
         .Z(n21294)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam i18974_3_lut_3_lut.init = 16'h7474;
    LUT4 n308_bdd_3_lut (.A(n26740), .B(n26721), .C(index_q[3]), .Z(n24917)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n308_bdd_3_lut.init = 16'hacac;
    LUT4 i19874_3_lut (.A(n22202), .B(n22203), .C(index_q[6]), .Z(n22213)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19874_3_lut.init = 16'hcaca;
    PFUMX mux_192_Mux_1_i891 (.BLUT(n882_adj_2262), .ALUT(n890_adj_2753), 
          .C0(n26565), .Z(n891_adj_2440)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    PFUMX i25956 (.BLUT(n28762), .ALUT(n28761), .C0(index_i[2]), .Z(n28763));
    LUT4 i11616_4_lut_4_lut (.A(index_i[3]), .B(index_i[2]), .C(index_i[0]), 
         .D(index_i[1]), .Z(n875_adj_2719)) /* synthesis lut_function=((B (C)+!B (D))+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11616_4_lut_4_lut.init = 16'hf7d5;
    PFUMX i20360 (.BLUT(n21784), .ALUT(n317_adj_2445), .C0(index_q[5]), 
          .Z(n22699));
    LUT4 mux_191_Mux_1_i987_3_lut_4_lut_4_lut (.A(index_i[3]), .B(n986_adj_2714), 
         .C(index_i[4]), .D(n29174), .Z(n987)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_1_i987_3_lut_4_lut_4_lut.init = 16'hc5c0;
    LUT4 i20204_3_lut_4_lut_3_lut (.A(index_i[3]), .B(index_i[4]), .C(n26486), 
         .Z(n22543)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20204_3_lut_4_lut_3_lut.init = 16'h6464;
    PFUMX i22685 (.BLUT(n26354), .ALUT(n26373), .C0(index_i[7]), .Z(n24249));
    LUT4 n24921_bdd_3_lut (.A(n24921), .B(n157_adj_2754), .C(index_q[4]), 
         .Z(n24922)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n24921_bdd_3_lut.init = 16'hcaca;
    LUT4 i9533_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n11979)) /* synthesis lut_function=(!(A (B (D)+!B (C+!(D)))+!A !(B (D)+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9533_3_lut_4_lut_4_lut.init = 16'h4699;
    LUT4 i19963_3_lut (.A(n25357), .B(n22763), .C(index_q[6]), .Z(n22302)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19963_3_lut.init = 16'hcaca;
    LUT4 n20971_bdd_3_lut_23276 (.A(n26598), .B(n26699), .C(index_i[3]), 
         .Z(n24947)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n20971_bdd_3_lut_23276.init = 16'hcaca;
    LUT4 mux_191_Mux_1_i573_3_lut_4_lut_4_lut (.A(index_i[3]), .B(n557_adj_2755), 
         .C(index_i[4]), .D(n29174), .Z(n573_adj_2641)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B ((D)+!C)+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_1_i573_3_lut_4_lut_4_lut.init = 16'h5c0c;
    LUT4 i20478_3_lut_4_lut_4_lut (.A(n26482), .B(index_q[4]), .C(index_q[5]), 
         .D(n26410), .Z(n22817)) /* synthesis lut_function=(A ((C+!(D))+!B)+!A (B (C+!(D))+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20478_3_lut_4_lut_4_lut.init = 16'he3ef;
    PFUMX i20361 (.BLUT(n349_adj_2556), .ALUT(n21790), .C0(index_q[5]), 
          .Z(n22700));
    LUT4 i11532_2_lut_3_lut_3_lut (.A(index_i[3]), .B(index_i[1]), .C(index_i[0]), 
         .Z(n14092)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11532_2_lut_3_lut_3_lut.init = 16'h4040;
    LUT4 mux_192_Mux_3_i684_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[4]), .Z(n684_adj_2752)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A !(B ((D)+!C)+!B (C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_3_i684_3_lut_3_lut_4_lut.init = 16'h5594;
    L6MUX21 i23011 (.D0(n24641), .D1(n24638), .SD(index_i[5]), .Z(n24642));
    L6MUX21 i20362 (.D0(n21793), .D1(n21799), .SD(index_q[5]), .Z(n22701));
    PFUMX i25914 (.BLUT(n28705), .ALUT(n28704), .C0(index_q[3]), .Z(n28706));
    L6MUX21 i20363 (.D0(n21802), .D1(n21808), .SD(index_q[5]), .Z(n22702));
    PFUMX i23009 (.BLUT(n24640), .ALUT(n475_adj_2697), .C0(index_i[4]), 
          .Z(n24641));
    LUT4 i8820_4_lut_4_lut (.A(index_i[3]), .B(index_i[0]), .C(index_i[1]), 
         .D(index_i[2]), .Z(n11225)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (D)+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i8820_4_lut_4_lut.init = 16'h0bf4;
    L6MUX21 i20365 (.D0(n21817), .D1(n636_adj_2535), .SD(index_q[5]), 
            .Z(n22704));
    LUT4 i22522_2_lut_rep_412_3_lut_4_lut (.A(n26569), .B(index_q[2]), .C(index_q[5]), 
         .D(n26584), .Z(n26372)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i22522_2_lut_rep_412_3_lut_4_lut.init = 16'h0f7f;
    PFUMX i23006 (.BLUT(n24637), .ALUT(n24636), .C0(index_i[4]), .Z(n24638));
    PFUMX i20366 (.BLUT(n21820), .ALUT(n700_adj_2361), .C0(index_q[5]), 
          .Z(n22705));
    L6MUX21 i20368 (.D0(n21373), .D1(n21385), .SD(index_q[5]), .Z(n22707));
    LUT4 i19246_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21566)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C))+!A !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19246_3_lut_4_lut_4_lut.init = 16'h5a52;
    PFUMX i25911 (.BLUT(n28701), .ALUT(n28700), .C0(index_q[2]), .Z(n28702));
    LUT4 i19385_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21705)) /* synthesis lut_function=(A (B (C+(D))+!B ((D)+!C))+!A !(B (C+(D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19385_3_lut_4_lut.init = 16'haa96;
    LUT4 mux_191_Mux_0_i124_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n124_adj_2414)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A !(B (D)+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_0_i124_3_lut_4_lut_4_lut.init = 16'h6c99;
    LUT4 i19019_4_lut_3_lut (.A(index_i[3]), .B(index_i[4]), .C(n26438), 
         .Z(n21339)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19019_4_lut_3_lut.init = 16'h6565;
    LUT4 mux_191_Mux_2_i221_4_lut_4_lut (.A(index_i[3]), .B(index_i[4]), 
         .C(n26438), .D(n26397), .Z(n221_adj_2593)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (B+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_2_i221_4_lut_4_lut.init = 16'hf7c4;
    PFUMX i20370 (.BLUT(n924_adj_2545), .ALUT(n21391), .C0(index_q[5]), 
          .Z(n22709));
    PFUMX i24057 (.BLUT(n254_adj_2274), .ALUT(n25806), .C0(index_q[8]), 
          .Z(n25807));
    PFUMX i20371 (.BLUT(n987_adj_2756), .ALUT(n21394), .C0(index_q[5]), 
          .Z(n22710));
    LUT4 i9502_3_lut_3_lut (.A(index_i[3]), .B(index_i[4]), .C(n11947), 
         .Z(n11948)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9502_3_lut_3_lut.init = 16'h7474;
    LUT4 mux_191_Mux_6_i459_rep_798 (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .Z(n29177)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_6_i459_rep_798.init = 16'h4d4d;
    LUT4 mux_191_Mux_11_i638_4_lut_4_lut (.A(n26376), .B(index_i[5]), .C(index_i[6]), 
         .D(n26415), .Z(n638_adj_2757)) /* synthesis lut_function=(A (B (C (D))+!B !(C))+!A (B ((D)+!C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_11_i638_4_lut_4_lut.init = 16'hc707;
    LUT4 mux_191_Mux_6_i732_3_lut_4_lut (.A(n26650), .B(index_i[3]), .C(index_i[4]), 
         .D(n731_adj_2538), .Z(n732_adj_2693)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_6_i732_3_lut_4_lut.init = 16'hf909;
    LUT4 i11630_2_lut_rep_448_3_lut_4_lut (.A(index_q[2]), .B(index_q[3]), 
         .C(index_q[4]), .D(n26569), .Z(n26408)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11630_2_lut_rep_448_3_lut_4_lut.init = 16'hf8f0;
    LUT4 mux_191_Mux_6_i700_3_lut_4_lut (.A(n26650), .B(index_i[3]), .C(index_i[4]), 
         .D(n684_adj_2724), .Z(n700_adj_2691)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_6_i700_3_lut_4_lut.init = 16'h9f90;
    LUT4 i11357_2_lut_3_lut_4_lut (.A(n26519), .B(n26595), .C(index_i[6]), 
         .D(index_i[5]), .Z(n254_adj_2465)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i11357_2_lut_3_lut_4_lut.init = 16'hfef0;
    LUT4 mux_192_Mux_3_i859_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n859_adj_2758)) /* synthesis lut_function=(!(A (B (D)+!B !(D))+!A (B (C+(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_3_i859_3_lut_3_lut_4_lut.init = 16'h339c;
    LUT4 i18697_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21017)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(D))+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18697_3_lut_3_lut_4_lut.init = 16'h3319;
    L6MUX21 i22986 (.D0(n24598), .D1(n24596), .SD(index_i[5]), .Z(n24599));
    LUT4 index_i_5__bdd_3_lut_4_lut (.A(index_i[0]), .B(index_i[2]), .C(n251_adj_2548), 
         .D(index_i[5]), .Z(n25335)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam index_i_5__bdd_3_lut_4_lut.init = 16'hf066;
    LUT4 i15424_3_lut_3_lut (.A(index_i[0]), .B(index_i[2]), .C(index_i[3]), 
         .Z(n17574)) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i15424_3_lut_3_lut.init = 16'h6a6a;
    LUT4 n20971_bdd_3_lut_23642_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n24948)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C))+!A !(B (C+!(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n20971_bdd_3_lut_23642_4_lut_4_lut.init = 16'h5ad6;
    PFUMX i22984 (.BLUT(n24597), .ALUT(n285_adj_2620), .C0(index_i[4]), 
          .Z(n24598));
    LUT4 mux_191_Mux_4_i349_3_lut_4_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[4]), .D(n348_adj_2674), .Z(n349_adj_2533)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_4_i349_3_lut_4_lut.init = 16'hf606;
    LUT4 i19496_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[2]), .C(index_q[3]), 
         .D(index_q[1]), .Z(n21816)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+!(D)))+!A !(B+!(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19496_3_lut_4_lut_4_lut.init = 16'h6c67;
    LUT4 mux_191_Mux_4_i828_3_lut_4_lut (.A(index_i[4]), .B(index_i[3]), 
         .C(n812_adj_2293), .D(n26598), .Z(n828_adj_2553)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_4_i828_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_191_Mux_5_i797_3_lut_4_lut (.A(index_i[4]), .B(index_i[3]), 
         .C(n26757), .D(n26700), .Z(n797_adj_2498)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_5_i797_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_191_Mux_1_i763_3_lut_4_lut (.A(index_i[4]), .B(index_i[3]), 
         .C(n26834), .D(n26700), .Z(n763_adj_2326)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_1_i763_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12222_2_lut_rep_601 (.A(index_i[2]), .B(index_i[0]), .Z(n26561)) /* synthesis lut_function=(A (B)) */ ;
    defparam i12222_2_lut_rep_601.init = 16'h8888;
    LUT4 i20105_4_lut_4_lut (.A(index_i[4]), .B(index_i[5]), .C(n26763), 
         .D(n908_adj_2657), .Z(n22444)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam i20105_4_lut_4_lut.init = 16'hd1c0;
    LUT4 i22432_2_lut_rep_602 (.A(index_i[4]), .B(index_i[3]), .Z(n26562)) /* synthesis lut_function=((B)+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i22432_2_lut_rep_602.init = 16'hdddd;
    LUT4 i19274_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21594)) /* synthesis lut_function=(A (B (C)+!B !(C (D)+!C !(D)))+!A (B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19274_3_lut_4_lut_4_lut.init = 16'hd6a5;
    LUT4 mux_191_Mux_3_i797_3_lut_4_lut (.A(index_i[4]), .B(index_i[3]), 
         .C(n796_adj_2539), .D(n70_adj_2255), .Z(n797_adj_2311)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_3_i797_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i18766_3_lut_3_lut_4_lut (.A(index_q[2]), .B(n26567), .C(n26521), 
         .D(index_q[3]), .Z(n21086)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (B (C (D))+!B (C+!(D)))) */ ;
    defparam i18766_3_lut_3_lut_4_lut.init = 16'hf099;
    LUT4 mux_191_Mux_3_i700_3_lut_4_lut (.A(index_i[4]), .B(index_i[3]), 
         .C(n684_adj_2759), .D(n26598), .Z(n700_adj_2578)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_3_i700_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i11459_2_lut_rep_641 (.A(index_i[2]), .B(index_i[3]), .Z(n26601)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11459_2_lut_rep_641.init = 16'heeee;
    LUT4 i22000_3_lut (.A(n25585), .B(n21561), .C(index_q[5]), .Z(n21562)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22000_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_7_i443_3_lut_4_lut (.A(index_q[2]), .B(n26567), .C(index_q[3]), 
         .D(n29182), .Z(n443_adj_2637)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;
    defparam mux_192_Mux_7_i443_3_lut_4_lut.init = 16'h6f60;
    LUT4 i20225_3_lut_4_lut_3_lut (.A(index_q[3]), .B(index_q[4]), .C(n29190), 
         .Z(n22564)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20225_3_lut_4_lut_3_lut.init = 16'h6464;
    LUT4 mux_192_Mux_1_i987_3_lut_4_lut_4_lut (.A(index_q[3]), .B(n986_adj_2746), 
         .C(index_q[4]), .D(n26528), .Z(n987_adj_2756)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_1_i987_3_lut_4_lut_4_lut.init = 16'hc5c0;
    LUT4 i8841_4_lut_4_lut (.A(index_q[3]), .B(index_q[0]), .C(index_q[1]), 
         .D(index_q[2]), .Z(n11249)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (D)+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i8841_4_lut_4_lut.init = 16'h0bf4;
    LUT4 i11107_4_lut_4_lut (.A(index_q[3]), .B(index_q[2]), .C(index_q[0]), 
         .D(index_q[1]), .Z(n875_adj_2442)) /* synthesis lut_function=((B (C)+!B (D))+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11107_4_lut_4_lut.init = 16'hf7d5;
    LUT4 i19241_4_lut_3_lut (.A(index_q[3]), .B(index_q[4]), .C(n26430), 
         .Z(n21561)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19241_4_lut_3_lut.init = 16'h6565;
    LUT4 mux_192_Mux_2_i221_4_lut_4_lut (.A(index_q[3]), .B(index_q[4]), 
         .C(n26430), .D(n26401), .Z(n221_adj_2734)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (B+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_2_i221_4_lut_4_lut.init = 16'hf7c4;
    LUT4 i9573_3_lut_3_lut (.A(index_q[3]), .B(index_q[4]), .C(n12018), 
         .Z(n12019)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9573_3_lut_3_lut.init = 16'h7474;
    LUT4 i18694_3_lut_3_lut_4_lut (.A(index_q[2]), .B(n26567), .C(n29182), 
         .D(index_q[3]), .Z(n21014)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (B (C (D))+!B (C+!(D)))) */ ;
    defparam i18694_3_lut_3_lut_4_lut.init = 16'hf099;
    LUT4 i19297_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21617)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19297_3_lut_4_lut.init = 16'h64cc;
    LUT4 i9568_4_lut_4_lut (.A(index_q[4]), .B(n22042), .C(n29208), .D(n29192), 
         .Z(n12014)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam i9568_4_lut_4_lut.init = 16'hf4b0;
    LUT4 i20280_4_lut_4_lut (.A(index_q[4]), .B(index_q[5]), .C(n26801), 
         .D(n908_adj_2305), .Z(n22619)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam i20280_4_lut_4_lut.init = 16'hd1c0;
    LUT4 i22453_2_lut_rep_605 (.A(index_q[4]), .B(index_q[3]), .Z(n26565)) /* synthesis lut_function=((B)+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i22453_2_lut_rep_605.init = 16'hdddd;
    LUT4 mux_192_Mux_3_i797_3_lut_4_lut (.A(index_q[4]), .B(index_q[3]), 
         .C(n796_adj_2484), .D(n29192), .Z(n797)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_3_i797_3_lut_4_lut.init = 16'hf2d0;
    LUT4 mux_191_Mux_5_i731_3_lut (.A(n26608), .B(n26706), .C(index_i[3]), 
         .Z(n731)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_5_i731_3_lut.init = 16'hcaca;
    LUT4 mux_191_Mux_0_i142_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n142_adj_2760)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C))+!A !(B (C (D)+!C !(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_0_i142_3_lut_4_lut_4_lut.init = 16'ha569;
    LUT4 n627_bdd_3_lut_23766_4_lut_4_lut (.A(index_q[2]), .B(n676), .C(index_q[3]), 
         .D(n26569), .Z(n25449)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B ((D)+!C)+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n627_bdd_3_lut_23766_4_lut_4_lut.init = 16'h5c0c;
    LUT4 i11267_2_lut_rep_607 (.A(index_q[0]), .B(index_q[1]), .Z(n26567)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11267_2_lut_rep_607.init = 16'h8888;
    LUT4 mux_192_Mux_3_i1002_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n19590)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (D))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_3_i1002_3_lut_3_lut_4_lut.init = 16'hf708;
    LUT4 mux_192_Mux_4_i491_3_lut_4_lut_4_lut (.A(index_q[2]), .B(n29187), 
         .C(index_q[3]), .D(n26567), .Z(n491_adj_2761)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_4_i491_3_lut_4_lut_4_lut.init = 16'hfc5c;
    LUT4 mux_192_Mux_3_i860_3_lut_4_lut (.A(index_q[2]), .B(n26567), .C(index_q[4]), 
         .D(n859_adj_2758), .Z(n860_adj_2475)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam mux_192_Mux_3_i860_3_lut_4_lut.init = 16'hf606;
    LUT4 i11318_2_lut_rep_425_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n26385)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A (B+((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11318_2_lut_rep_425_4_lut_4_lut_4_lut.init = 16'h0038;
    LUT4 mux_192_Mux_3_i93_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n93_adj_2254)) /* synthesis lut_function=(A (B (C+!(D))+!B (D))+!A (B ((D)+!C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_3_i93_3_lut_4_lut_4_lut_4_lut.init = 16'hf78c;
    LUT4 n10961_bdd_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n25355)) /* synthesis lut_function=(A (B (C+!(D))+!B ((D)+!C))+!A (B (C (D)+!C !(D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n10961_bdd_3_lut_4_lut_4_lut_4_lut.init = 16'hf38f;
    LUT4 i1_4_lut_adj_82 (.A(index_q[6]), .B(n26482), .C(index_q[5]), 
         .D(index_q[4]), .Z(n19975)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_4_lut_adj_82.init = 16'hfffe;
    PFUMX i20122 (.BLUT(n12004), .ALUT(n62_adj_2762), .C0(index_i[5]), 
          .Z(n22461));
    LUT4 n476_bdd_3_lut_23393_3_lut_4_lut (.A(index_q[2]), .B(n26567), .C(n491_adj_2761), 
         .D(index_q[4]), .Z(n25081)) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))+!A !(B ((D)+!C)+!B !(C+(D)))) */ ;
    defparam n476_bdd_3_lut_23393_3_lut_4_lut.init = 16'h99f0;
    LUT4 mux_192_Mux_5_i781_3_lut_4_lut_4_lut_else_4_lut (.A(index_q[3]), 
         .B(index_q[0]), .C(index_q[4]), .Z(n26770)) /* synthesis lut_function=(!(A (C)+!A (B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_5_i781_3_lut_4_lut_4_lut_else_4_lut.init = 16'h1f1f;
    LUT4 i17442_4_lut (.A(n26622), .B(n892_adj_2542), .C(index_q[6]), 
         .D(index_q[5]), .Z(n19624)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D))))) */ ;
    defparam i17442_4_lut.init = 16'h3a35;
    PFUMX i20060 (.BLUT(n31_adj_2528), .ALUT(n62_adj_2763), .C0(index_i[5]), 
          .Z(n22399));
    LUT4 i22211_3_lut (.A(n19624), .B(n19975), .C(index_q[7]), .Z(n22495)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22211_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_7_i924_3_lut_3_lut_4_lut (.A(index_q[2]), .B(index_q[3]), 
         .C(index_q[4]), .D(n26569), .Z(n924_adj_2621)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_7_i924_3_lut_3_lut_4_lut.init = 16'h878f;
    LUT4 i18782_3_lut_4_lut_4_lut (.A(index_q[2]), .B(n250), .C(index_q[3]), 
         .D(n26569), .Z(n21102)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18782_3_lut_4_lut_4_lut.init = 16'hc5c0;
    PFUMX i20029 (.BLUT(n31_adj_2525), .ALUT(n62_adj_2523), .C0(index_i[5]), 
          .Z(n22368));
    PFUMX i25613 (.BLUT(n28281), .ALUT(n28280), .C0(index_i[1]), .Z(n28282));
    PFUMX i19998 (.BLUT(n31_adj_2521), .ALUT(n21580), .C0(index_i[5]), 
          .Z(n22337));
    PFUMX i19853 (.BLUT(n31_adj_2518), .ALUT(n21019), .C0(index_q[5]), 
          .Z(n22192));
    PFUMX i22982 (.BLUT(n24595), .ALUT(n24594), .C0(index_i[4]), .Z(n24596));
    LUT4 mux_191_Mux_1_i732_3_lut (.A(n716_adj_2347), .B(n491_adj_2389), 
         .C(index_i[4]), .Z(n732_adj_2325)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_1_i732_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_rep_516_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(n26584), .Z(n26476)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_3_lut_rep_516_4_lut.init = 16'hfff8;
    PFUMX i19854 (.BLUT(n94_adj_2516), .ALUT(n125_adj_2513), .C0(index_q[5]), 
          .Z(n22193));
    LUT4 i19486_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n21806)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A (B (C)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19486_3_lut_4_lut_4_lut.init = 16'h3c8c;
    LUT4 i11685_2_lut_rep_497_3_lut (.A(index_q[2]), .B(index_q[3]), .C(index_q[1]), 
         .Z(n26457)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11685_2_lut_rep_497_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_rep_674 (.A(index_i[5]), .B(index_i[6]), .Z(n26634)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i1_2_lut_rep_674.init = 16'heeee;
    LUT4 i1_3_lut_4_lut_adj_83 (.A(index_i[5]), .B(index_i[6]), .C(index_i[7]), 
         .D(n26635), .Z(n20065)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i1_3_lut_4_lut_adj_83.init = 16'hfffe;
    LUT4 i11449_2_lut_rep_675 (.A(index_i[3]), .B(index_i[4]), .Z(n26635)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11449_2_lut_rep_675.init = 16'h8888;
    LUT4 i20632_3_lut_3_lut_4_lut (.A(index_i[3]), .B(index_i[4]), .C(n413_adj_2318), 
         .D(index_i[5]), .Z(n22971)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20632_3_lut_3_lut_4_lut.init = 16'h77f0;
    LUT4 i12188_2_lut_3_lut (.A(index_i[3]), .B(index_i[4]), .C(index_i[5]), 
         .Z(n14756)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i12188_2_lut_3_lut.init = 16'hf8f8;
    LUT4 i22145_3_lut (.A(n22444), .B(n25237), .C(index_i[6]), .Z(n22453)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22145_3_lut.init = 16'hcaca;
    PFUMX i19930 (.BLUT(n31_adj_2510), .ALUT(n62_adj_2764), .C0(index_q[5]), 
          .Z(n22269));
    LUT4 mux_192_Mux_4_i1002_3_lut_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n1002_adj_2457)) /* synthesis lut_function=(A (B (C (D))+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_4_i1002_3_lut_3_lut_3_lut_4_lut.init = 16'hf007;
    LUT4 i1_2_lut_3_lut_adj_84 (.A(index_i[3]), .B(index_i[4]), .C(index_i[5]), 
         .Z(n20230)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i1_2_lut_3_lut_adj_84.init = 16'h8080;
    LUT4 i12214_2_lut_rep_676 (.A(index_i[2]), .B(index_i[0]), .Z(n26636)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i12214_2_lut_rep_676.init = 16'heeee;
    LUT4 i19067_3_lut_4_lut (.A(n26569), .B(index_q[2]), .C(index_q[3]), 
         .D(n29173), .Z(n21387)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19067_3_lut_4_lut.init = 16'hdfd0;
    PFUMX i19855 (.BLUT(n17579), .ALUT(n14391), .C0(index_q[5]), .Z(n22194));
    LUT4 i20418_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n22757)) /* synthesis lut_function=(A (B (D)+!B !(C (D)+!C !(D)))+!A !(B (C+!(D))+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20418_3_lut_4_lut_4_lut.init = 16'h8f30;
    L6MUX21 i19857 (.D0(n21022), .D1(n21025), .SD(index_q[5]), .Z(n22196));
    LUT4 i1_2_lut_rep_545_3_lut (.A(index_i[2]), .B(index_i[0]), .C(index_i[1]), 
         .Z(n26505)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_545_3_lut.init = 16'hfefe;
    L6MUX21 i19858 (.D0(n21028), .D1(n21031), .SD(index_q[5]), .Z(n22197));
    LUT4 i11268_2_lut_2_lut_3_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[3]), 
         .Z(n13827)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11268_2_lut_2_lut_3_lut.init = 16'h0808;
    LUT4 i11091_2_lut_rep_441_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n26401)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11091_2_lut_rep_441_3_lut_4_lut.init = 16'hf080;
    LUT4 mux_191_Mux_9_i285_3_lut_3_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[1]), .Z(n285_adj_2423)) /* synthesis lut_function=(A (C)+!A !(B+(C+(D)))) */ ;
    defparam mux_191_Mux_9_i285_3_lut_3_lut_4_lut_4_lut.init = 16'ha0a1;
    LUT4 mux_192_Mux_6_i812_3_lut_4_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n812_adj_2574)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(D))+!A !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_6_i812_3_lut_4_lut_3_lut_4_lut.init = 16'h7780;
    LUT4 mux_191_Mux_5_i954_3_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[1]), .Z(n954_adj_2264)) /* synthesis lut_function=(!(A (C)+!A (B+((D)+!C)))) */ ;
    defparam mux_191_Mux_5_i954_3_lut_4_lut_4_lut.init = 16'h0a1a;
    PFUMX i19859 (.BLUT(n413_adj_2506), .ALUT(n444_adj_2397), .C0(index_q[5]), 
          .Z(n22198));
    LUT4 i1_2_lut_rep_469_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n26429)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_2_lut_rep_469_3_lut_4_lut.init = 16'h8000;
    LUT4 i11724_2_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(n26622), 
         .D(index_q[2]), .Z(n125)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11724_2_lut_3_lut_4_lut.init = 16'hf080;
    PFUMX i19860 (.BLUT(n476_adj_2504), .ALUT(n507_adj_2501), .C0(index_q[5]), 
          .Z(n22199));
    LUT4 mux_191_Mux_0_i46_3_lut_4_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[1]), .D(index_i[3]), .Z(n46_adj_2551)) /* synthesis lut_function=(A (D)+!A (B+(C+!(D)))) */ ;
    defparam mux_191_Mux_0_i46_3_lut_4_lut_4_lut_4_lut.init = 16'hfe55;
    LUT4 mux_191_Mux_8_i716_3_lut_4_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[1]), .D(index_i[3]), .Z(n716_adj_2747)) /* synthesis lut_function=(!(A (D)+!A !(B+(C+(D))))) */ ;
    defparam mux_191_Mux_8_i716_3_lut_4_lut_4_lut_4_lut.init = 16'h55fe;
    LUT4 mux_192_Mux_6_i730_3_lut_rep_568_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n26528)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_6_i730_3_lut_rep_568_3_lut.init = 16'h3838;
    LUT4 mux_192_Mux_8_i526_3_lut_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n526_adj_2370)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_8_i526_3_lut_3_lut_3_lut_4_lut.init = 16'h0f70;
    LUT4 mux_192_Mux_7_i491_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n491_adj_2765)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(D))+!A (B (C+!(D))+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_7_i491_3_lut_4_lut_4_lut_4_lut.init = 16'h3780;
    LUT4 i11367_2_lut_rep_454_3_lut_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[1]), .Z(n26414)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;
    defparam i11367_2_lut_rep_454_3_lut_4_lut.init = 16'hf0e0;
    LUT4 n45_bdd_2_lut_3_lut_3_lut_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[1]), .D(index_i[3]), .Z(n25327)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B ((D)+!C)))) */ ;
    defparam n45_bdd_2_lut_3_lut_3_lut_4_lut.init = 16'h00fe;
    LUT4 n875_bdd_3_lut_24339_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n25352)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+!(D)))+!A (B (D)+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n875_bdd_3_lut_24339_4_lut_4_lut_4_lut.init = 16'h30f7;
    PFUMX i19861 (.BLUT(n17545), .ALUT(n573_adj_2766), .C0(index_q[5]), 
          .Z(n22200));
    LUT4 i11599_2_lut_rep_677 (.A(index_i[1]), .B(index_i[2]), .Z(n26637)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11599_2_lut_rep_677.init = 16'heeee;
    LUT4 mux_192_Mux_1_i348_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n348_adj_2555)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A (B (C+!(D))+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_1_i348_3_lut_4_lut_4_lut.init = 16'h3f80;
    PFUMX i19862 (.BLUT(n605_adj_2767), .ALUT(n636_adj_2499), .C0(index_q[5]), 
          .Z(n22201));
    LUT4 mux_192_Mux_9_i316_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), 
         .B(index_q[1]), .C(index_q[3]), .D(index_q[2]), .Z(n316_adj_2729)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C+(D)))+!A (B (C (D)+!C !(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_9_i316_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h3ff8;
    LUT4 mux_192_Mux_5_i30_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n30_adj_2517)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A (B+!(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_5_i30_3_lut_4_lut.init = 16'hcc67;
    PFUMX i19863 (.BLUT(n21034), .ALUT(n700_adj_2422), .C0(index_q[5]), 
          .Z(n22202));
    LUT4 i11278_2_lut_rep_609 (.A(index_q[0]), .B(index_q[1]), .Z(n26569)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11278_2_lut_rep_609.init = 16'heeee;
    PFUMX i19899 (.BLUT(n31), .ALUT(n62_adj_2496), .C0(index_q[5]), .Z(n22238));
    LUT4 mux_191_Mux_5_i781_3_lut_4_lut_4_lut_then_4_lut (.A(index_i[3]), 
         .B(index_i[0]), .C(index_i[4]), .D(index_i[2]), .Z(n26756)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_5_i781_3_lut_4_lut_4_lut_then_4_lut.init = 16'hece0;
    LUT4 i11445_2_lut_rep_546_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[3]), 
         .Z(n26506)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11445_2_lut_rep_546_3_lut.init = 16'he0e0;
    LUT4 mux_191_Mux_9_i93_3_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .Z(n93_adj_2405)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_9_i93_3_lut_3_lut.init = 16'hc1c1;
    LUT4 i11694_2_lut_rep_473_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[0]), 
         .Z(n26433)) /* synthesis lut_function=(A (C)+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11694_2_lut_rep_473_3_lut.init = 16'hf1f1;
    LUT4 mux_191_Mux_8_i412_3_lut_4_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .Z(n14770)) /* synthesis lut_function=(A (B+!(C))+!A !((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_8_i412_3_lut_4_lut_3_lut.init = 16'h8e8e;
    LUT4 i19279_3_lut_4_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n21599)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19279_3_lut_4_lut_3_lut_4_lut.init = 16'h0fe0;
    LUT4 i22037_3_lut (.A(n27886), .B(n25217), .C(index_i[5]), .Z(n22382)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22037_3_lut.init = 16'hcaca;
    L6MUX21 i19864 (.D0(n732_adj_2673), .D1(n21037), .SD(index_q[5]), 
            .Z(n22203));
    PFUMX i19865 (.BLUT(n797_adj_2709), .ALUT(n828), .C0(index_q[5]), 
          .Z(n22204));
    LUT4 i11270_2_lut_rep_566_3_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .Z(n26526)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11270_2_lut_rep_566_3_lut.init = 16'he0e0;
    LUT4 mux_192_Mux_0_i333_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n333_adj_2768)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_0_i333_3_lut_3_lut_4_lut.init = 16'hf10e;
    PFUMX i19866 (.BLUT(n860_adj_2494), .ALUT(n891_adj_2491), .C0(index_q[5]), 
          .Z(n22205));
    LUT4 n10365_bdd_3_lut_22614_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[4]), .D(index_i[3]), .Z(n24127)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C+(D)))+!A (B (C (D)+!C !(D))+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n10365_bdd_3_lut_22614_4_lut_4_lut_4_lut.init = 16'hc10f;
    L6MUX21 i25532 (.D0(n28181), .D1(n28178), .SD(index_i[7]), .Z(n28182));
    LUT4 i11319_2_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n635_adj_2534)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A (B (C+!(D))+!B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11319_2_lut_4_lut_4_lut.init = 16'hf1fc;
    PFUMX i25530 (.BLUT(n28180), .ALUT(n28179), .C0(index_i[5]), .Z(n28181));
    LUT4 mux_191_Mux_9_i412_3_lut_3_lut_4_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .Z(n412_adj_2319)) /* synthesis lut_function=(!(A (B (C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_9_i412_3_lut_3_lut_4_lut_3_lut.init = 16'h7e7e;
    PFUMX i22928 (.BLUT(n24542), .ALUT(n24538), .C0(index_i[6]), .Z(n24543));
    PFUMX i25528 (.BLUT(n22978), .ALUT(n28177), .C0(index_i[6]), .Z(n28178));
    LUT4 n17762_bdd_4_lut_then_4_lut (.A(index_i[3]), .B(index_i[4]), .C(index_i[1]), 
         .D(index_i[2]), .Z(n26833)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B+(C (D)+!C !(D)))) */ ;
    defparam n17762_bdd_4_lut_then_4_lut.init = 16'hf44f;
    LUT4 mux_191_Mux_4_i236_3_lut_4_lut_3_lut_rep_630_4_lut (.A(index_i[1]), 
         .B(index_i[2]), .C(index_i[3]), .D(index_i[0]), .Z(n26590)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_4_i236_3_lut_4_lut_3_lut_rep_630_4_lut.init = 16'hf01f;
    LUT4 n17762_bdd_4_lut_else_4_lut (.A(index_i[3]), .B(index_i[4]), .C(index_i[1]), 
         .D(index_i[2]), .Z(n26832)) /* synthesis lut_function=(!(A (B (D)+!B ((D)+!C))+!A !(B+!((D)+!C)))) */ ;
    defparam n17762_bdd_4_lut_else_4_lut.init = 16'h44fc;
    LUT4 i11290_2_lut_rep_450_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n26410)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11290_2_lut_rep_450_3_lut_4_lut.init = 16'hfef0;
    LUT4 i11446_2_lut_rep_455_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[4]), .D(index_i[3]), .Z(n26415)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11446_2_lut_rep_455_3_lut_4_lut.init = 16'hfef0;
    LUT4 i19406_3_lut_3_lut_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[3]), 
         .Z(n21726)) /* synthesis lut_function=(A (C)+!A (B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19406_3_lut_3_lut_3_lut.init = 16'he5e5;
    LUT4 n903_bdd_3_lut_4_lut_3_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .Z(n26166)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n903_bdd_3_lut_4_lut_3_lut.init = 16'h6161;
    LUT4 i18781_3_lut_3_lut_4_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n21101)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18781_3_lut_3_lut_4_lut_3_lut_4_lut.init = 16'h11ef;
    LUT4 mux_192_Mux_3_i30_3_lut_3_lut_4_lut_3_lut_4_lut (.A(index_q[0]), 
         .B(index_q[1]), .C(index_q[3]), .D(index_q[2]), .Z(n30_adj_2509)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_3_i30_3_lut_3_lut_4_lut_3_lut_4_lut.init = 16'hfe11;
    LUT4 mux_192_Mux_6_i796_3_lut_rep_396_3_lut_3_lut_4_lut (.A(index_q[0]), 
         .B(index_q[1]), .C(index_q[3]), .D(index_q[2]), .Z(n26356)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_6_i796_3_lut_rep_396_3_lut_3_lut_4_lut.init = 16'hfe01;
    LUT4 mux_192_Mux_3_i557_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n557_adj_2660)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_3_i557_3_lut_3_lut_4_lut.init = 16'hf10f;
    LUT4 i12169_1_lut_rep_410_2_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n26370)) /* synthesis lut_function=(!(A (C+(D))+!A (B (C+(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12169_1_lut_rep_410_2_lut_3_lut_4_lut.init = 16'h010f;
    LUT4 i18796_3_lut (.A(n498), .B(n29195), .C(index_q[3]), .Z(n21116)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18796_3_lut.init = 16'hcaca;
    LUT4 i22041_3_lut (.A(n542_adj_2722), .B(n573_adj_2430), .C(index_i[5]), 
         .Z(n22376)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22041_3_lut.init = 16'hcaca;
    LUT4 i22926_then_3_lut (.A(index_i[0]), .B(index_i[4]), .C(index_i[3]), 
         .Z(n26836)) /* synthesis lut_function=(A (B)+!A (B (C)+!B !(C))) */ ;
    defparam i22926_then_3_lut.init = 16'hc9c9;
    L6MUX21 i20424 (.D0(n22761), .D1(n22762), .SD(index_q[5]), .Z(n22763));
    LUT4 i22926_else_3_lut (.A(index_i[2]), .B(index_i[0]), .C(index_i[4]), 
         .D(index_i[3]), .Z(n26835)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)+!C !(D)))+!A (B (C+!(D))+!B !(C)))) */ ;
    defparam i22926_else_3_lut.init = 16'h1e38;
    LUT4 i19459_3_lut_4_lut (.A(n26569), .B(index_q[2]), .C(index_q[3]), 
         .D(n29182), .Z(n21779)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19459_3_lut_4_lut.init = 16'hdfd0;
    LUT4 i21523_3_lut (.A(n21116), .B(n21117), .C(index_q[4]), .Z(n21118)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21523_3_lut.init = 16'hcaca;
    LUT4 i19460_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n21780)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C+(D)))+!A (B (C (D)+!C !(D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19460_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h3ef0;
    L6MUX21 i25492 (.D0(n28122), .D1(n28119), .SD(index_q[7]), .Z(n28123));
    LUT4 mux_192_Mux_6_i908_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), 
         .B(index_q[1]), .C(index_q[3]), .D(index_q[2]), .Z(n908_adj_2563)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A (B (C (D)+!C !(D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_6_i908_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h1cf0;
    PFUMX i25490 (.BLUT(n28121), .ALUT(n28120), .C0(index_q[5]), .Z(n28122));
    LUT4 i11679_2_lut_rep_522_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n26482)) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11679_2_lut_rep_522_3_lut_4_lut.init = 16'he000;
    LUT4 mux_192_Mux_3_i157_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n157_adj_2452)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_3_i157_3_lut_3_lut_4_lut.init = 16'h1ff0;
    PFUMX i25488 (.BLUT(n22825), .ALUT(n28118), .C0(index_q[6]), .Z(n28119));
    LUT4 i22485_2_lut_rep_495_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n26455)) /* synthesis lut_function=(!(A+(B+(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i22485_2_lut_rep_495_3_lut_4_lut.init = 16'h0111;
    LUT4 i20224_3_lut_3_lut_4_lut (.A(n26526), .B(index_q[3]), .C(n923_adj_2544), 
         .D(index_q[4]), .Z(n22563)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20224_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 i19472_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n21792)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B ((D)+!C)+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19472_3_lut_4_lut_4_lut.init = 16'hfc1c;
    LUT4 mux_192_Mux_3_i109_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n109_adj_2454)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (D)+!B !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_3_i109_3_lut_4_lut_4_lut.init = 16'hcf10;
    LUT4 mux_191_Mux_5_i781_3_lut_4_lut_4_lut_else_4_lut (.A(index_i[3]), 
         .B(index_i[0]), .C(index_i[4]), .Z(n26755)) /* synthesis lut_function=(!(A (C)+!A (B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_5_i781_3_lut_4_lut_4_lut_else_4_lut.init = 16'h1f1f;
    LUT4 i11700_2_lut_rep_525_3_lut (.A(index_i[2]), .B(index_i[3]), .C(index_i[1]), 
         .Z(n26485)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11700_2_lut_rep_525_3_lut.init = 16'hfefe;
    LUT4 mux_192_Mux_2_i250_3_lut_3_lut_4_lut_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n250)) /* synthesis lut_function=(A ((C)+!B)+!A (B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_2_i250_3_lut_3_lut_4_lut_3_lut.init = 16'he7e7;
    LUT4 mux_192_Mux_5_i53_3_lut_4_lut_3_lut_rep_610 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n26570)) /* synthesis lut_function=(A ((C)+!B)+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_5_i53_3_lut_4_lut_3_lut_rep_610.init = 16'he6e6;
    LUT4 mux_192_Mux_7_i506_3_lut_4_lut_4_lut (.A(index_q[2]), .B(n29187), 
         .C(index_q[3]), .D(n26569), .Z(n506_adj_2769)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B ((D)+!C)+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_7_i506_3_lut_4_lut_4_lut.init = 16'h5c0c;
    LUT4 mux_192_Mux_6_i691_3_lut_rep_611 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n26571)) /* synthesis lut_function=(A (B+!(C))+!A !((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_6_i691_3_lut_rep_611.init = 16'h8e8e;
    LUT4 i11890_3_lut_3_lut_4_lut_4_lut (.A(index_q[2]), .B(index_q[3]), 
         .C(index_q[1]), .D(index_q[0]), .Z(n14450)) /* synthesis lut_function=(!(A+!(B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11890_3_lut_3_lut_4_lut_4_lut.init = 16'h4555;
    LUT4 mux_192_Mux_0_i557_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n557_adj_2416)) /* synthesis lut_function=(A ((D)+!C)+!A !((D)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_0_i557_3_lut_4_lut.init = 16'haa4e;
    LUT4 i19454_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21774)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A (B (D)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19454_3_lut_4_lut.init = 16'h18cc;
    LUT4 i18763_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21083)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)))+!A !(B (C+!(D))+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18763_3_lut_3_lut_4_lut.init = 16'h71cc;
    LUT4 mux_192_Mux_6_i635_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n635_adj_2515)) /* synthesis lut_function=(A (B (C+(D))+!B !(D))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_6_i635_3_lut_4_lut.init = 16'hcce6;
    LUT4 mux_192_Mux_3_i142_3_lut_4_lut_3_lut (.A(index_q[2]), .B(index_q[3]), 
         .C(index_q[1]), .Z(n142_adj_2451)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_3_i142_3_lut_4_lut_3_lut.init = 16'h6464;
    LUT4 mux_192_Mux_11_i766_3_lut (.A(n638), .B(n765), .C(index_q[7]), 
         .Z(n766)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_11_i766_3_lut.init = 16'h3a3a;
    LUT4 i7157_2_lut_rep_684 (.A(index_q[1]), .B(index_q[2]), .Z(n26644)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i7157_2_lut_rep_684.init = 16'heeee;
    L6MUX21 i20784 (.D0(n23107), .D1(n23108), .SD(index_i[5]), .Z(n23123));
    LUT4 mux_192_Mux_8_i412_3_lut_4_lut_3_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .Z(n14848)) /* synthesis lut_function=(A (B+!(C))+!A !((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_8_i412_3_lut_4_lut_3_lut.init = 16'h8e8e;
    LUT4 i18791_3_lut (.A(n498), .B(n26740), .C(index_q[3]), .Z(n21111)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18791_3_lut.init = 16'hcaca;
    PFUMX i19900 (.BLUT(n94), .ALUT(n21046), .C0(index_q[5]), .Z(n22239));
    LUT4 i11513_2_lut_rep_537_3_lut (.A(index_q[1]), .B(index_q[2]), .C(index_q[3]), 
         .Z(n26497)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11513_2_lut_rep_537_3_lut.init = 16'he0e0;
    L6MUX21 i20785 (.D0(n23109), .D1(n23110), .SD(index_i[5]), .Z(n23124));
    PFUMX i19902 (.BLUT(n221_adj_2770), .ALUT(n252_adj_2771), .C0(index_q[5]), 
          .Z(n22241));
    LUT4 n10831_bdd_3_lut_24390_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[4]), .D(index_q[3]), .Z(n24162)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C+(D)))+!A (B (C (D)+!C !(D))+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n10831_bdd_3_lut_24390_4_lut_4_lut_4_lut.init = 16'hc10f;
    LUT4 mux_192_Mux_9_i93_3_lut_3_lut_3_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .Z(n93)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_9_i93_3_lut_3_lut_3_lut.init = 16'hc1c1;
    PFUMX i19903 (.BLUT(n286_adj_2470), .ALUT(n21049), .C0(index_q[5]), 
          .Z(n22242));
    LUT4 mux_192_Mux_4_i236_3_lut_4_lut_3_lut_rep_622_4_lut (.A(index_q[1]), 
         .B(index_q[2]), .C(index_q[3]), .D(index_q[0]), .Z(n26582)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_4_i236_3_lut_4_lut_3_lut_rep_622_4_lut.init = 16'hf01f;
    L6MUX21 i23918 (.D0(n25634), .D1(n25631), .SD(index_q[5]), .Z(n25635));
    LUT4 index_q_1__bdd_4_lut_25534 (.A(index_q[1]), .B(index_q[0]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n26841)) /* synthesis lut_function=(!(A (B (D)+!B (C+!(D)))+!A !(B (C (D)+!C !(D))+!B !((D)+!C)))) */ ;
    defparam index_q_1__bdd_4_lut_25534.init = 16'h429c;
    PFUMX i19904 (.BLUT(n349), .ALUT(n21052), .C0(index_q[5]), .Z(n22243));
    LUT4 i22885_then_4_lut (.A(index_i[0]), .B(index_i[4]), .C(index_i[1]), 
         .D(index_i[3]), .Z(n26843)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam i22885_then_4_lut.init = 16'h3c69;
    LUT4 mux_192_Mux_1_i923_3_lut_3_lut_4_lut_3_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .Z(n923_adj_2544)) /* synthesis lut_function=(!(A (B (C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_1_i923_3_lut_3_lut_4_lut_3_lut.init = 16'h7e7e;
    PFUMX i24499 (.BLUT(n26793), .ALUT(n26794), .C0(index_i[0]), .Z(n26795));
    LUT4 i12102_3_lut_3_lut (.A(index_q[2]), .B(index_q[0]), .C(index_q[1]), 
         .Z(n1001)) /* synthesis lut_function=(A (C)+!A (B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12102_3_lut_3_lut.init = 16'hf4f4;
    PFUMX i23916 (.BLUT(n25633), .ALUT(n25632), .C0(index_q[4]), .Z(n25634));
    LUT4 i22885_else_4_lut (.A(index_i[0]), .B(index_i[4]), .C(index_i[1]), 
         .D(index_i[3]), .Z(n26842)) /* synthesis lut_function=(!(A (B (C)+!B !(C (D)+!C !(D)))+!A (B ((D)+!C)+!B !((D)+!C)))) */ ;
    defparam i22885_else_4_lut.init = 16'h394b;
    LUT4 i11514_2_lut_rep_452_3_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[4]), .D(index_q[3]), .Z(n26412)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11514_2_lut_rep_452_3_lut_4_lut.init = 16'hfef0;
    LUT4 i11764_2_lut_rep_553_3_lut (.A(index_q[1]), .B(index_q[2]), .C(index_q[0]), 
         .Z(n26513)) /* synthesis lut_function=(A (C)+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11764_2_lut_rep_553_3_lut.init = 16'hf1f1;
    LUT4 i18724_3_lut_4_lut_3_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .D(index_q[0]), .Z(n21044)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18724_3_lut_4_lut_3_lut_4_lut.init = 16'h0fe0;
    L6MUX21 i25379 (.D0(n29161), .D1(n27994), .SD(index_q[3]), .Z(n27998));
    PFUMX i19909 (.BLUT(n669_adj_2463), .ALUT(n700_adj_2462), .C0(index_q[5]), 
          .Z(n22248));
    PFUMX i19910 (.BLUT(n21064), .ALUT(n763_adj_2392), .C0(index_q[5]), 
          .Z(n22249));
    PFUMX i25375 (.BLUT(n27993), .ALUT(n27992), .C0(index_q[4]), .Z(n27994));
    PFUMX i19911 (.BLUT(n21067), .ALUT(n828_adj_2664), .C0(index_q[5]), 
          .Z(n22250));
    LUT4 i11303_3_lut_3_lut_4_lut_4_lut (.A(index_q[2]), .B(index_q[3]), 
         .C(index_q[1]), .D(index_q[0]), .Z(n13863)) /* synthesis lut_function=(!(A ((C+(D))+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11303_3_lut_3_lut_4_lut_4_lut.init = 16'h555d;
    LUT4 i21530_3_lut (.A(n21107), .B(n21108), .C(index_q[4]), .Z(n21109)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21530_3_lut.init = 16'hcaca;
    LUT4 i18785_3_lut (.A(n26740), .B(n26570), .C(index_q[3]), .Z(n21105)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18785_3_lut.init = 16'hcaca;
    LUT4 index_i_0__bdd_4_lut_25253 (.A(index_i[0]), .B(index_i[3]), .C(index_i[1]), 
         .D(index_i[2]), .Z(n26845)) /* synthesis lut_function=(A (B (C)+!B !(C+!(D)))+!A !(B ((D)+!C)+!B !(C (D)+!C !(D)))) */ ;
    defparam index_i_0__bdd_4_lut_25253.init = 16'h92c1;
    LUT4 i21534_3_lut (.A(n21104), .B(n21105), .C(index_q[4]), .Z(n21106)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21534_3_lut.init = 16'hcaca;
    PFUMX i19912 (.BLUT(n860_adj_2459), .ALUT(n21070), .C0(index_q[5]), 
          .Z(n22251));
    LUT4 mux_192_Mux_2_i931_3_lut_4_lut_3_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[0]), .Z(n931_adj_2372)) /* synthesis lut_function=(!(A (B)+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_2_i931_3_lut_4_lut_3_lut.init = 16'h7676;
    LUT4 mux_192_Mux_6_i636_4_lut_4_lut (.A(index_q[1]), .B(index_q[4]), 
         .C(n635_adj_2515), .D(n14395), .Z(n636_adj_2751)) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_6_i636_4_lut_4_lut.init = 16'hf3d1;
    LUT4 mux_191_Mux_3_i349_3_lut_3_lut (.A(index_i[1]), .B(index_i[4]), 
         .C(n348_adj_2684), .Z(n349_adj_2565)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_3_i349_3_lut_3_lut.init = 16'hd1d1;
    LUT4 i21538_3_lut (.A(n21101), .B(n21102), .C(index_q[4]), .Z(n21103)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21538_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_2_i62_3_lut_3_lut (.A(index_q[1]), .B(index_q[4]), 
         .C(n812_adj_2583), .Z(n62_adj_2743)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_2_i62_3_lut_3_lut.init = 16'h7474;
    L6MUX21 i20786 (.D0(n23111), .D1(n23112), .SD(index_i[5]), .Z(n23125));
    L6MUX21 i20787 (.D0(n23113), .D1(n23114), .SD(index_i[5]), .Z(n23126));
    L6MUX21 i20788 (.D0(n23115), .D1(n23116), .SD(index_i[5]), .Z(n23127));
    PFUMX i23913 (.BLUT(n25630), .ALUT(n26385), .C0(index_q[4]), .Z(n25631));
    LUT4 i22626_then_4_lut (.A(index_q[0]), .B(index_q[4]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n26850)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)+!C !(D))+!B (C (D)))) */ ;
    defparam i22626_then_4_lut.init = 16'hda0e;
    LUT4 mux_192_Mux_2_i94_3_lut_3_lut (.A(index_q[1]), .B(index_q[4]), 
         .C(n124_adj_2512), .Z(n94_adj_2618)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_2_i94_3_lut_3_lut.init = 16'hd1d1;
    L6MUX21 i20789 (.D0(n23117), .D1(n23118), .SD(index_i[5]), .Z(n23128));
    L6MUX21 i20790 (.D0(n23119), .D1(n23120), .SD(index_i[5]), .Z(n23129));
    L6MUX21 i20791 (.D0(n23121), .D1(n23122), .SD(index_i[5]), .Z(n23130));
    LUT4 i19073_3_lut_4_lut_3_lut (.A(index_q[1]), .B(index_q[3]), .C(index_q[2]), 
         .Z(n21393)) /* synthesis lut_function=(A (B)+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19073_3_lut_4_lut_3_lut.init = 16'hd9d9;
    L6MUX21 i20462 (.D0(n22799), .D1(n22800), .SD(index_q[5]), .Z(n22801));
    LUT4 i22626_else_4_lut (.A(index_q[0]), .B(index_q[4]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n26849)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C))+!A (B (C)+!B (C+(D)))) */ ;
    defparam i22626_else_4_lut.init = 16'hf178;
    PFUMX i19931 (.BLUT(n94_adj_2772), .ALUT(n125_adj_2455), .C0(index_q[5]), 
          .Z(n22270));
    LUT4 mux_192_Mux_3_i349_3_lut_3_lut (.A(index_q[1]), .B(index_q[4]), 
         .C(n348_adj_2638), .Z(n349_adj_2467)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_3_i349_3_lut_3_lut.init = 16'hd1d1;
    LUT4 mux_192_Mux_5_i924_4_lut_3_lut (.A(index_q[2]), .B(n13839), .C(index_q[4]), 
         .Z(n924_adj_2773)) /* synthesis lut_function=(!(A (B+(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_5_i924_4_lut_3_lut.init = 16'h5656;
    LUT4 i22065_3_lut (.A(n286_adj_2735), .B(n317_adj_2733), .C(index_q[5]), 
         .Z(n22816)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22065_3_lut.init = 16'hcaca;
    LUT4 i11831_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), .B(n26539), .C(index_q[4]), 
         .D(index_q[0]), .Z(n14391)) /* synthesis lut_function=(!(A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11831_3_lut_4_lut_4_lut_4_lut.init = 16'h55d5;
    L6MUX21 i20469 (.D0(n22806), .D1(n22807), .SD(index_q[5]), .Z(n22808));
    PFUMX i19932 (.BLUT(n158_adj_2453), .ALUT(n189), .C0(index_q[5]), 
          .Z(n22271));
    PFUMX i19933 (.BLUT(n221_adj_2646), .ALUT(n252), .C0(index_q[5]), 
          .Z(n22272));
    LUT4 i19352_3_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[3]), .C(index_i[2]), 
         .D(index_i[0]), .Z(n21672)) /* synthesis lut_function=(A (B (D)+!B (C (D)+!C !(D)))+!A (B (D)+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19352_3_lut_4_lut_4_lut.init = 16'hfc13;
    LUT4 i19495_3_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[2]), .C(index_q[0]), 
         .D(index_q[3]), .Z(n21815)) /* synthesis lut_function=(!(A ((D)+!B)+!A !(B (D)+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19495_3_lut_4_lut_4_lut.init = 16'h4588;
    PFUMX i20474 (.BLUT(n22809), .ALUT(n22810), .C0(index_q[4]), .Z(n22813));
    L6MUX21 i25317 (.D0(n27930), .D1(n27927), .SD(index_i[5]), .Z(n27931));
    PFUMX i20475 (.BLUT(n22811), .ALUT(n22812), .C0(index_q[4]), .Z(n22814));
    PFUMX i25315 (.BLUT(n27929), .ALUT(n27928), .C0(index_i[3]), .Z(n27930));
    PFUMX i26214 (.BLUT(n29202), .ALUT(n29203), .C0(index_q[0]), .Z(n29204));
    PFUMX i15392 (.BLUT(n17540), .ALUT(n17541), .C0(index_q[4]), .Z(n17542));
    PFUMX i19960 (.BLUT(n22297), .ALUT(n22298), .C0(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_2142[3]));
    LUT4 i22317_2_lut_rep_686 (.A(index_q[1]), .B(index_q[2]), .Z(n26646)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i22317_2_lut_rep_686.init = 16'h9999;
    PFUMX i25312 (.BLUT(n27926), .ALUT(n27925), .C0(index_i[3]), .Z(n27927));
    PFUMX i20028 (.BLUT(n22365), .ALUT(n22366), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2127[5]));
    PFUMX i19455 (.BLUT(n21773), .ALUT(n21774), .C0(index_q[4]), .Z(n21775));
    PFUMX i20090 (.BLUT(n22427), .ALUT(n22428), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2127[3]));
    LUT4 i11324_2_lut_rep_772 (.A(index_q[0]), .B(index_q[1]), .Z(n26732)) /* synthesis lut_function=(A+!(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11324_2_lut_rep_772.init = 16'hbbbb;
    L6MUX21 i23893 (.D0(n25595), .D1(n25593), .SD(index_q[4]), .Z(n25596));
    LUT4 i11323_2_lut_rep_751 (.A(index_q[0]), .B(index_q[1]), .Z(n26711)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11323_2_lut_rep_751.init = 16'h2222;
    PFUMX i18702 (.BLUT(n21020), .ALUT(n21021), .C0(index_q[4]), .Z(n21022));
    LUT4 n378_bdd_2_lut_23790_3_lut (.A(index_q[1]), .B(index_q[2]), .C(index_q[3]), 
         .Z(n25464)) /* synthesis lut_function=(A (B+(C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n378_bdd_2_lut_23790_3_lut.init = 16'hf9f9;
    PFUMX i18705 (.BLUT(n21023), .ALUT(n21024), .C0(index_q[4]), .Z(n21025));
    LUT4 mux_192_Mux_0_i93_3_lut_3_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .Z(n93_adj_2642)) /* synthesis lut_function=(A (B)+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_0_i93_3_lut_3_lut.init = 16'h9c9c;
    LUT4 i12244_2_lut_rep_687 (.A(index_i[0]), .B(index_i[1]), .Z(n26647)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i12244_2_lut_rep_687.init = 16'heeee;
    LUT4 i22073_3_lut (.A(n25329), .B(n21339), .C(index_i[5]), .Z(n21340)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22073_3_lut.init = 16'hcaca;
    PFUMX i23891 (.BLUT(n26401), .ALUT(n25594), .C0(index_q[5]), .Z(n25595));
    PFUMX i20152 (.BLUT(n22489), .ALUT(n22490), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2127[1]));
    LUT4 i17428_4_lut (.A(n26635), .B(n892_adj_2546), .C(index_i[6]), 
         .D(index_i[5]), .Z(n19605)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D))))) */ ;
    defparam i17428_4_lut.init = 16'h3a35;
    PFUMX i19461 (.BLUT(n21779), .ALUT(n21780), .C0(index_q[4]), .Z(n21781));
    LUT4 i22224_3_lut (.A(n19605), .B(n19979), .C(index_i[7]), .Z(n22318)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22224_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_6_i157_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n157_adj_2754)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (D))+!A !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_6_i157_3_lut_4_lut_4_lut_4_lut.init = 16'h5d22;
    LUT4 mux_191_Mux_3_i142_3_lut_4_lut_3_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[1]), .Z(n142_adj_2698)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_3_i142_3_lut_4_lut_3_lut.init = 16'h6464;
    LUT4 mux_191_Mux_8_i397_3_lut_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n397_adj_2432)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B ((D)+!C))) */ ;
    defparam mux_191_Mux_8_i397_3_lut_3_lut_3_lut_4_lut.init = 16'hf10f;
    LUT4 mux_192_Mux_4_i205_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n205)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_4_i205_3_lut_4_lut_4_lut.init = 16'h5a2a;
    PFUMX i23889 (.BLUT(n25592), .ALUT(n25591), .C0(index_q[5]), .Z(n25593));
    LUT4 mux_191_Mux_0_i333_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n333_adj_2774)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B (D))) */ ;
    defparam mux_191_Mux_0_i333_3_lut_3_lut_4_lut.init = 16'hf10e;
    PFUMX i18708 (.BLUT(n21026), .ALUT(n21027), .C0(index_q[4]), .Z(n21028));
    LUT4 mux_191_Mux_2_i716_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n716_adj_2695)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)+!C !(D)))+!A (B (D)+!B !((D)+!C)))) */ ;
    defparam mux_191_Mux_2_i716_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h31cf;
    LUT4 i19382_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n21702)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)+!C !(D)))+!A (B (C+!(D))+!B ((D)+!C)))) */ ;
    defparam i19382_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h0e30;
    LUT4 mux_191_Mux_3_i157_3_lut_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n157_adj_2317)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B !(C+(D))))) */ ;
    defparam mux_191_Mux_3_i157_3_lut_3_lut_3_lut_4_lut.init = 16'h1ff0;
    PFUMX i18711 (.BLUT(n21029), .ALUT(n21030), .C0(index_q[4]), .Z(n21031));
    LUT4 mux_191_Mux_4_i491_3_lut_4_lut_4_lut (.A(index_i[2]), .B(n26652), 
         .C(index_i[3]), .D(n26548), .Z(n491_adj_2718)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_4_i491_3_lut_4_lut_4_lut.init = 16'hfc5c;
    LUT4 n476_bdd_3_lut_23045_3_lut (.A(index_i[1]), .B(index_i[4]), .C(n124_adj_2540), 
         .Z(n24537)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n476_bdd_3_lut_23045_3_lut.init = 16'hd1d1;
    LUT4 i11401_2_lut_rep_459_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n26419)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i11401_2_lut_rep_459_3_lut_4_lut.init = 16'hfef0;
    PFUMX i20001 (.BLUT(n221), .ALUT(n252_adj_2345), .C0(index_i[5]), 
          .Z(n22340));
    LUT4 mux_191_Mux_7_i308_3_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n308)) /* synthesis lut_function=(A ((C)+!B)+!A (B+!(C))) */ ;
    defparam mux_191_Mux_7_i308_3_lut_4_lut_3_lut.init = 16'he7e7;
    LUT4 i19373_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n21693)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (B (C+!(D))+!B (D))) */ ;
    defparam i19373_3_lut_4_lut_4_lut_4_lut.init = 16'hf1cc;
    LUT4 i12207_3_lut_3_lut (.A(index_i[2]), .B(index_i[0]), .C(index_i[1]), 
         .Z(n38)) /* synthesis lut_function=(A (C)+!A (B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i12207_3_lut_3_lut.init = 16'hf4f4;
    LUT4 mux_191_Mux_8_i46_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n46_adj_2715)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (B (C)+!B !(C (D)+!C !(D)))) */ ;
    defparam mux_191_Mux_8_i46_3_lut_4_lut_4_lut_4_lut.init = 16'hc1f0;
    LUT4 i11525_3_lut_3_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n14085)) /* synthesis lut_function=(!(A+!(B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11525_3_lut_3_lut_4_lut_4_lut.init = 16'h4555;
    LUT4 i12409_1_lut_rep_407_2_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n26367)) /* synthesis lut_function=(!(A (C+(D))+!A (B (C+(D))+!B (C)))) */ ;
    defparam i12409_1_lut_rep_407_2_lut_3_lut_4_lut.init = 16'h010f;
    LUT4 mux_191_Mux_5_i924_4_lut_3_lut (.A(index_i[2]), .B(n14783), .C(index_i[4]), 
         .Z(n924)) /* synthesis lut_function=(!(A (B+(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_5_i924_4_lut_3_lut.init = 16'h5656;
    PFUMX i23881 (.BLUT(n25584), .ALUT(n25583), .C0(index_q[4]), .Z(n25585));
    LUT4 index_i_6__bdd_4_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[6]), 
         .C(index_i[5]), .D(n26519), .Z(n24765)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (D))+!A (B (C (D))+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam index_i_6__bdd_4_lut_4_lut_4_lut.init = 16'h04f7;
    PFUMX i20386 (.BLUT(n22723), .ALUT(n22724), .C0(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_2142[1]));
    LUT4 mux_191_Mux_2_i142_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n142_adj_2710)) /* synthesis lut_function=(!(A (B (D)+!B (C (D)+!C !(D)))+!A (B (D)+!B (C+!(D))))) */ ;
    defparam mux_191_Mux_2_i142_3_lut_4_lut_4_lut_4_lut.init = 16'h03ec;
    LUT4 i18741_then_4_lut (.A(index_q[1]), .B(index_q[2]), .C(index_q[4]), 
         .D(index_q[3]), .Z(n26856)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+(D)))+!A !(B (C)+!B !(C+!(D)))) */ ;
    defparam i18741_then_4_lut.init = 16'h9c97;
    LUT4 mux_191_Mux_7_i506_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n506)) /* synthesis lut_function=(!(A (B (D)+!B ((D)+!C))+!A (B (D)+!B (C+!(D))))) */ ;
    defparam mux_191_Mux_7_i506_3_lut_4_lut_4_lut_4_lut.init = 16'h01ec;
    LUT4 mux_191_Mux_8_i506_3_lut_4_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n506_adj_2683)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B ((D)+!C)))) */ ;
    defparam mux_191_Mux_8_i506_3_lut_4_lut_3_lut_4_lut.init = 16'h0ef0;
    LUT4 index_i_5__bdd_3_lut_23647_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n25226)) /* synthesis lut_function=(A (B (C)+!B (C+(D)))+!A (B (C)+!B !(C (D)+!C !(D)))) */ ;
    defparam index_i_5__bdd_3_lut_23647_4_lut_4_lut_4_lut.init = 16'he3f0;
    PFUMX i19473 (.BLUT(n21791), .ALUT(n21792), .C0(index_q[4]), .Z(n21793));
    LUT4 i11567_3_lut_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n14127)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B !(C+!(D))))) */ ;
    defparam i11567_3_lut_3_lut_3_lut_4_lut.init = 16'h10ff;
    LUT4 i19336_3_lut_3_lut_4_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n21656)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B !((D)+!C)))) */ ;
    defparam i19336_3_lut_3_lut_4_lut_3_lut_4_lut.init = 16'h11ef;
    PFUMX i9381 (.BLUT(n12046), .ALUT(n12047), .C0(n22061), .Z(n11827));
    LUT4 i11728_2_lut_rep_512_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n26472)) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;
    defparam i11728_2_lut_rep_512_3_lut_4_lut.init = 16'he000;
    LUT4 mux_191_Mux_3_i747_3_lut (.A(n26700), .B(n404), .C(index_i[3]), 
         .Z(n747_adj_2276)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_3_i747_3_lut.init = 16'hcaca;
    LUT4 mux_191_Mux_2_i931_3_lut_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n931_adj_2409)) /* synthesis lut_function=(!(A (B (C))+!A (B (C)+!B !(C)))) */ ;
    defparam mux_191_Mux_2_i931_3_lut_3_lut_3_lut.init = 16'h3e3e;
    LUT4 mux_191_Mux_7_i572_3_lut_rep_398_3_lut_3_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n26358)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)+!C !(D)))) */ ;
    defparam mux_191_Mux_7_i572_3_lut_rep_398_3_lut_3_lut_4_lut.init = 16'hfe01;
    LUT4 i11503_2_lut_rep_559_3_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .Z(n26519)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i11503_2_lut_rep_559_3_lut.init = 16'he0e0;
    LUT4 i11595_2_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n635_adj_2260)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A (B (C+!(D))+!B (C+(D)))) */ ;
    defparam i11595_2_lut_4_lut_4_lut.init = 16'hf1fc;
    LUT4 mux_191_Mux_3_i30_3_lut_3_lut_4_lut_4_lut_3_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[2]), .D(index_i[3]), .Z(n30_adj_2527)) /* synthesis lut_function=(A (C)+!A (B (C)+!B ((D)+!C))) */ ;
    defparam mux_191_Mux_3_i30_3_lut_3_lut_4_lut_4_lut_3_lut_4_lut.init = 16'hf1e1;
    LUT4 mux_191_Mux_7_i235_3_lut_rep_646_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26606)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C)+!B !(C))) */ ;
    defparam mux_191_Mux_7_i235_3_lut_rep_646_3_lut.init = 16'he3e3;
    LUT4 mux_191_Mux_7_i762_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n762_adj_2668)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A (B (C (D)+!C !(D))+!B !(C)))) */ ;
    defparam mux_191_Mux_7_i762_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h1cf0;
    LUT4 i19364_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n21684)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C+(D)))+!A (B (C (D)+!C !(D))+!B !(C)))) */ ;
    defparam i19364_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h3ef0;
    LUT4 mux_191_Mux_7_i541_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n541_adj_2675)) /* synthesis lut_function=(A (B (D)+!B (C+!(D)))+!A (B (D)+!B !(D))) */ ;
    defparam mux_191_Mux_7_i541_3_lut_4_lut_4_lut_4_lut.init = 16'hec33;
    LUT4 i19363_3_lut_4_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n21683)) /* synthesis lut_function=(A (B (D)+!B ((D)+!C))+!A (B (D)+!B (C+!(D)))) */ ;
    defparam i19363_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'hfe13;
    LUT4 mux_191_Mux_7_i60_3_lut_3_lut_4_lut_3_lut_rep_688 (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[2]), .Z(n26648)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B+!(C)))) */ ;
    defparam mux_191_Mux_7_i60_3_lut_3_lut_4_lut_3_lut_rep_688.init = 16'h1818;
    LUT4 i9596_3_lut_4_lut_3_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[4]), 
         .Z(n12046)) /* synthesis lut_function=(!(A (B)+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9596_3_lut_4_lut_3_lut.init = 16'h6262;
    LUT4 mux_191_Mux_8_i116_3_lut_rep_689 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26649)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B !(C))) */ ;
    defparam mux_191_Mux_8_i116_3_lut_rep_689.init = 16'hc1c1;
    LUT4 mux_191_Mux_7_i29_3_lut_rep_690 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26650)) /* synthesis lut_function=(A (B+!(C))+!A !((C)+!B)) */ ;
    defparam mux_191_Mux_7_i29_3_lut_rep_690.init = 16'h8e8e;
    PFUMX i9583 (.BLUT(n12064), .ALUT(n12065), .C0(n22054), .Z(n12030));
    PFUMX i19883 (.BLUT(n22220), .ALUT(n22221), .C0(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_2142[5]));
    LUT4 mux_192_Mux_0_i985_3_lut_3_lut_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n985)) /* synthesis lut_function=(!(A (B+!(C))+!A (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_0_i985_3_lut_3_lut_3_lut.init = 16'h2525;
    PFUMX i9509 (.BLUT(n12058), .ALUT(n12059), .C0(n22047), .Z(n11955));
    LUT4 mux_191_Mux_7_i340_3_lut_rep_692 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26652)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B (C)+!B !(C)))) */ ;
    defparam mux_191_Mux_7_i340_3_lut_rep_692.init = 16'h1c1c;
    LUT4 mux_192_Mux_0_i708_3_lut_4_lut_3_lut_rep_752 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n26712)) /* synthesis lut_function=(!(A (B)+!A ((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_0_i708_3_lut_4_lut_3_lut_rep_752.init = 16'h2626;
    LUT4 mux_191_Mux_7_i691_3_lut_rep_693 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26653)) /* synthesis lut_function=(!(A (B (C))+!A !(B+(C)))) */ ;
    defparam mux_191_Mux_7_i691_3_lut_rep_693.init = 16'h7e7e;
    PFUMX i19479 (.BLUT(n21797), .ALUT(n21798), .C0(index_q[4]), .Z(n21799));
    LUT4 mux_192_Mux_6_i347_3_lut_4_lut_3_lut_rep_754 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n26714)) /* synthesis lut_function=(!(A (B+!(C))+!A ((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_6_i347_3_lut_4_lut_3_lut_rep_754.init = 16'h2424;
    PFUMX i19975 (.BLUT(n22312), .ALUT(n22313), .C0(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_2142[8]));
    LUT4 mux_191_Mux_8_i30_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n30_adj_2707)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A !(B ((D)+!C)+!B (C (D)+!C !(D))))) */ ;
    defparam mux_191_Mux_8_i30_3_lut_3_lut_4_lut.init = 16'h7e0f;
    PFUMX i19482 (.BLUT(n21800), .ALUT(n21801), .C0(index_q[4]), .Z(n21802));
    LUT4 mux_191_Mux_0_i699_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n699_adj_2701)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (D))+!A (B (C+!(D))+!B !(C+!(D))))) */ ;
    defparam mux_191_Mux_0_i699_3_lut_3_lut_4_lut.init = 16'h1c33;
    PFUMX i19982 (.BLUT(n22319), .ALUT(n22320), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2127[9]));
    PFUMX i19488 (.BLUT(n21806), .ALUT(n21807), .C0(index_q[4]), .Z(n21808));
    PFUMX i22887 (.BLUT(n24494), .ALUT(n24491), .C0(index_i[6]), .Z(n24495));
    LUT4 i19319_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21639)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B (C (D)+!C !(D))))) */ ;
    defparam i19319_3_lut_3_lut_4_lut.init = 16'h0f1c;
    PFUMX i19497 (.BLUT(n21815), .ALUT(n21816), .C0(index_q[4]), .Z(n21817));
    LUT4 mux_192_Mux_4_i221_3_lut_3_lut (.A(index_q[0]), .B(index_q[4]), 
         .C(n205), .Z(n221_adj_2770)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_4_i221_3_lut_3_lut.init = 16'h7474;
    LUT4 i18741_else_4_lut (.A(index_q[1]), .B(index_q[2]), .C(index_q[4]), 
         .D(index_q[3]), .Z(n26855)) /* synthesis lut_function=(!(A (B (C)+!B !(C (D)+!C !(D)))+!A (B (C+(D))+!B !(C+!(D))))) */ ;
    defparam i18741_else_4_lut.init = 16'h381f;
    LUT4 mux_191_Mux_2_i955_then_4_lut (.A(index_i[4]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n26762)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B (C+!(D))+!B !(C (D)))) */ ;
    defparam mux_191_Mux_2_i955_then_4_lut.init = 16'he95d;
    PFUMX i20121 (.BLUT(n22458), .ALUT(n22459), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2127[2]));
    LUT4 mux_192_Mux_1_i890_4_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[3]), 
         .C(n26521), .D(index_q[4]), .Z(n890_adj_2753)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (D))+!A !((C+(D))+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_1_i890_4_lut_4_lut_4_lut_4_lut.init = 16'h55f3;
    LUT4 mux_192_Mux_0_i491_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n491_adj_2775)) /* synthesis lut_function=(!(A (B (D)+!B !(C+!(D)))+!A ((C+!(D))+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_0_i491_3_lut_4_lut.init = 16'h24aa;
    LUT4 mux_192_Mux_2_i859_3_lut_4_lut_4_lut (.A(index_q[0]), .B(n29195), 
         .C(index_q[3]), .D(n26644), .Z(n859_adj_2602)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B ((D)+!C)+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_2_i859_3_lut_4_lut_4_lut.init = 16'h5c0c;
    PFUMX i20159 (.BLUT(n22496), .ALUT(n22497), .C0(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_2142[9]));
    LUT4 i19396_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21716)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C (D)))+!A (B (C+(D))+!B !(C)))) */ ;
    defparam i19396_4_lut_4_lut_4_lut.init = 16'h301c;
    LUT4 mux_191_Mux_3_i653_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n653_adj_2708)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A !(B (D)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_3_i653_3_lut_4_lut_4_lut.init = 16'h4d99;
    LUT4 mux_191_Mux_7_i716_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n716_adj_2669)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C+!(D))+!B (C)))) */ ;
    defparam mux_191_Mux_7_i716_3_lut_3_lut_4_lut.init = 16'h0f81;
    LUT4 n476_bdd_3_lut_24561 (.A(n476_adj_2619), .B(n25081), .C(index_q[5]), 
         .Z(n25082)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n476_bdd_3_lut_24561.init = 16'hcaca;
    LUT4 mux_191_Mux_0_i557_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n557_adj_2639)) /* synthesis lut_function=(A ((D)+!C)+!A !((D)+!B)) */ ;
    defparam mux_191_Mux_0_i557_3_lut_4_lut.init = 16'haa4e;
    LUT4 i19318_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21638)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)))+!A !(B (C+!(D))+!B (D)))) */ ;
    defparam i19318_3_lut_3_lut_4_lut.init = 16'h71cc;
    LUT4 n316_bdd_3_lut_24380_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n25307)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A !(B ((D)+!C)+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n316_bdd_3_lut_24380_3_lut_4_lut.init = 16'h552c;
    LUT4 mux_192_Mux_2_i348_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n348_adj_2776)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_2_i348_3_lut_4_lut_4_lut.init = 16'h52a5;
    LUT4 n45_bdd_3_lut_23576_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n25262)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C (D)+!C !(D))+!B (C)))) */ ;
    defparam n45_bdd_3_lut_23576_3_lut_4_lut.init = 16'h0fc1;
    LUT4 mux_191_Mux_2_i557_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n557_adj_2420)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C+!(D))+!B (C (D)+!C !(D))))) */ ;
    defparam mux_191_Mux_2_i557_3_lut_3_lut_4_lut.init = 16'h0f18;
    LUT4 i19361_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21681)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A (B (D)+!B !(C (D))))) */ ;
    defparam i19361_3_lut_4_lut.init = 16'h18cc;
    LUT4 mux_192_Mux_5_i573_3_lut_3_lut (.A(index_q[0]), .B(index_q[4]), 
         .C(n572_adj_2777), .Z(n573_adj_2766)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_5_i573_3_lut_3_lut.init = 16'hd1d1;
    PFUMX i20031 (.BLUT(n158), .ALUT(n189_adj_2778), .C0(index_i[5]), 
          .Z(n22370));
    LUT4 mux_192_Mux_2_i507_3_lut_3_lut (.A(index_q[0]), .B(index_q[4]), 
         .C(n491_adj_2384), .Z(n507_adj_2738)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_2_i507_3_lut_3_lut.init = 16'h7474;
    PFUMX i20629 (.BLUT(n22966), .ALUT(n22967), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2127[8]));
    LUT4 index_q_0__bdd_4_lut_24486 (.A(index_q[0]), .B(index_q[3]), .C(index_q[1]), 
         .D(index_q[2]), .Z(n26768)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C))+!A (B (C (D)+!C !(D))+!B !(C+!(D))))) */ ;
    defparam index_q_0__bdd_4_lut_24486.init = 16'h16d3;
    LUT4 mux_191_Mux_4_i389_3_lut_3_lut_3_lut_rep_799 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29178)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_4_i389_3_lut_3_lut_3_lut_rep_799.init = 16'h9393;
    LUT4 i18775_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21095)) /* synthesis lut_function=(!(A (B)+!A (B (C+(D))+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18775_3_lut_3_lut_4_lut.init = 16'h3326;
    PFUMX i23856 (.BLUT(n25553), .ALUT(n26741), .C0(index_q[4]), .Z(n25554));
    PFUMX i20296 (.BLUT(n22633), .ALUT(n22634), .C0(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_2142[2]));
    LUT4 i11835_2_lut_3_lut_3_lut (.A(index_q[0]), .B(index_q[3]), .C(index_q[2]), 
         .Z(n14395)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11835_2_lut_3_lut_3_lut.init = 16'h4040;
    LUT4 mux_192_Mux_2_i349_3_lut_3_lut (.A(index_q[0]), .B(index_q[4]), 
         .C(n348_adj_2776), .Z(n349_adj_2736)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_2_i349_3_lut_3_lut.init = 16'hd1d1;
    LUT4 i9469_3_lut_4_lut_4_lut (.A(index_q[0]), .B(n931), .C(index_q[4]), 
         .D(n26644), .Z(n11915)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B ((D)+!C)+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9469_3_lut_4_lut_4_lut.init = 16'h5c0c;
    PFUMX i20495 (.BLUT(n142_adj_2760), .ALUT(n157_adj_2426), .C0(index_i[4]), 
          .Z(n22834));
    LUT4 mux_191_Mux_2_i955_else_4_lut (.A(index_i[4]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n26761)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+(D)))+!A !(B (C+!(D))+!B !(C+!(D))))) */ ;
    defparam mux_191_Mux_2_i955_else_4_lut.init = 16'h49c6;
    LUT4 mux_192_Mux_2_i763_4_lut_4_lut (.A(index_q[0]), .B(n11877), .C(index_q[4]), 
         .D(n157_adj_2754), .Z(n763_adj_2741)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_2_i763_4_lut_4_lut.init = 16'hdfd0;
    PFUMX i20496 (.BLUT(n173_adj_2692), .ALUT(n188_adj_2410), .C0(index_i[4]), 
          .Z(n22835));
    PFUMX i18717 (.BLUT(n21035), .ALUT(n21036), .C0(index_q[4]), .Z(n21037));
    LUT4 i18772_3_lut_4_lut_4_lut (.A(index_q[0]), .B(n29167), .C(index_q[3]), 
         .D(n26644), .Z(n21092)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18772_3_lut_4_lut_4_lut.init = 16'hc5c0;
    LUT4 i18773_3_lut (.A(n325), .B(n29173), .C(index_q[3]), .Z(n21093)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18773_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_4_i142_3_lut_4_lut_3_lut (.A(index_q[0]), .B(index_q[3]), 
         .C(index_q[2]), .Z(n142_adj_2623)) /* synthesis lut_function=(A (B (C))+!A !(B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_4_i142_3_lut_4_lut_3_lut.init = 16'h9595;
    LUT4 i21810_3_lut (.A(n21092), .B(n21093), .C(index_q[4]), .Z(n21094)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21810_3_lut.init = 16'hcaca;
    LUT4 i19072_3_lut (.A(n29176), .B(n29167), .C(index_q[3]), .Z(n21392)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19072_3_lut.init = 16'hcaca;
    PFUMX mux_192_Mux_14_i1023 (.BLUT(n511), .ALUT(n19899), .C0(index_q[9]), 
          .Z(quarter_wave_sample_register_q_15__N_2142[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 mux_192_Mux_3_i444_3_lut_4_lut (.A(index_q[0]), .B(index_q[3]), 
         .C(n26538), .D(index_q[4]), .Z(n444_adj_2471)) /* synthesis lut_function=(!(A (B (D)+!B (C (D)))+!A !(B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_3_i444_3_lut_4_lut.init = 16'h46aa;
    LUT4 mux_192_Mux_4_i252_4_lut_4_lut (.A(index_q[0]), .B(index_q[3]), 
         .C(n26644), .D(index_q[4]), .Z(n252_adj_2771)) /* synthesis lut_function=(!(A (B (D)+!B !(D))+!A !(B ((D)+!C)+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_4_i252_4_lut_4_lut.init = 16'h669d;
    LUT4 mux_191_Mux_11_i766_3_lut (.A(n638_adj_2757), .B(n765_adj_2381), 
         .C(index_i[7]), .Z(n766_adj_2779)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_11_i766_3_lut.init = 16'h3a3a;
    LUT4 i22245_3_lut (.A(n766_adj_2779), .B(n20065), .C(index_i[8]), 
         .Z(n21171)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22245_3_lut.init = 16'hcaca;
    LUT4 i21427_3_lut (.A(n21392), .B(n21393), .C(index_q[4]), .Z(n21394)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21427_3_lut.init = 16'hcaca;
    PFUMX i20501 (.BLUT(n333_adj_2774), .ALUT(n348_adj_2541), .C0(index_i[4]), 
          .Z(n22840));
    LUT4 mux_192_Mux_3_i62_3_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[4]), .D(n812_adj_2574), .Z(n62_adj_2764)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_3_i62_3_lut_4_lut.init = 16'h6f60;
    PFUMX i20502 (.BLUT(n364_adj_2780), .ALUT(n379), .C0(index_i[4]), 
          .Z(n22841));
    L6MUX21 i12939362_i1 (.D0(n22922), .D1(n23075), .SD(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_2142[0]));
    LUT4 i19027_3_lut_then_4_lut (.A(index_q[4]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n29203)) /* synthesis lut_function=(A (B (C)+!B !(C (D)+!C !(D)))+!A !(B (C)+!B !(C (D)+!C !(D)))) */ ;
    defparam i19027_3_lut_then_4_lut.init = 16'h96a5;
    L6MUX21 i12927356_i1 (.D0(n22860), .D1(n23137), .SD(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2127[0]));
    PFUMX mux_191_Mux_14_i1023 (.BLUT(n511_adj_2466), .ALUT(n20039), .C0(index_i[9]), 
          .Z(quarter_wave_sample_register_i_15__N_2127[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    PFUMX i20503 (.BLUT(n397_adj_2404), .ALUT(n412_adj_2351), .C0(index_i[4]), 
          .Z(n22842));
    LUT4 i18797_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n21117)) /* synthesis lut_function=(A (C+(D))+!A !(B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18797_3_lut_4_lut_4_lut.init = 16'haba5;
    PFUMX i20504 (.BLUT(n428_adj_2346), .ALUT(n443), .C0(index_i[4]), 
          .Z(n22843));
    LUT4 index_q_4__bdd_3_lut_22718_4_lut (.A(n26496), .B(index_q[3]), .C(index_q[5]), 
         .D(index_q[4]), .Z(n24289)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam index_q_4__bdd_3_lut_22718_4_lut.init = 16'hf080;
    PFUMX i20505 (.BLUT(n460_adj_2331), .ALUT(n475_adj_2406), .C0(index_i[4]), 
          .Z(n22844));
    LUT4 i21578_3_lut (.A(n491_adj_2765), .B(n506_adj_2769), .C(index_q[4]), 
         .Z(n21375)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21578_3_lut.init = 16'hcaca;
    LUT4 i20288_3_lut (.A(n25452), .B(n22618), .C(index_q[6]), .Z(n22627)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20288_3_lut.init = 16'hcaca;
    LUT4 i19052_3_lut (.A(n29197), .B(n29173), .C(index_q[3]), .Z(n21372)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19052_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_3_i94_3_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[4]), .D(n93_adj_2254), .Z(n94_adj_2772)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_3_i94_3_lut_4_lut.init = 16'hf606;
    LUT4 i20624_3_lut (.A(n22956), .B(n22957), .C(index_i[7]), .Z(n22963)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20624_3_lut.init = 16'hcaca;
    LUT4 i20623_3_lut (.A(n22954), .B(n24767), .C(index_i[7]), .Z(n22962)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20623_3_lut.init = 16'hcaca;
    L6MUX21 i23808 (.D0(n25486), .D1(n25484), .SD(index_i[5]), .Z(n25487));
    LUT4 i22319_2_lut_rep_757 (.A(index_q[0]), .B(index_q[1]), .Z(n26717)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i22319_2_lut_rep_757.init = 16'h9999;
    PFUMX i20506 (.BLUT(n491_adj_2781), .ALUT(n11225), .C0(index_i[4]), 
          .Z(n22845));
    PFUMX i23806 (.BLUT(n25485), .ALUT(n70), .C0(index_i[3]), .Z(n25486));
    LUT4 i15428_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n17578)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i15428_3_lut_4_lut_4_lut_4_lut.init = 16'h3999;
    LUT4 i22135_3_lut (.A(n11948), .B(n892_adj_2558), .C(index_i[6]), 
         .Z(n22960)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22135_3_lut.init = 16'hcaca;
    PFUMX i23804 (.BLUT(n25483), .ALUT(n21528), .C0(index_i[4]), .Z(n25484));
    LUT4 n25864_bdd_3_lut_3_lut (.A(n1021_adj_2728), .B(index_q[8]), .C(n25864), 
         .Z(n25865)) /* synthesis lut_function=(A (B+(C))+!A !(B+!(C))) */ ;
    defparam n25864_bdd_3_lut_3_lut.init = 16'hb8b8;
    L6MUX21 i22855 (.D0(n24459), .D1(n24457), .SD(index_q[6]), .Z(n24460));
    PFUMX i18852 (.BLUT(n21170), .ALUT(n21171), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2127[11]));
    LUT4 i18770_3_lut (.A(n26720), .B(n26734), .C(index_q[3]), .Z(n21090)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18770_3_lut.init = 16'hcaca;
    PFUMX i22853 (.BLUT(n24458), .ALUT(n62_adj_2377), .C0(index_q[5]), 
          .Z(n24459));
    LUT4 i7662_2_lut_rep_624 (.A(index_q[3]), .B(index_q[4]), .Z(n26584)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i7662_2_lut_rep_624.init = 16'heeee;
    LUT4 i9385_3_lut_4_lut (.A(index_q[3]), .B(index_q[4]), .C(n26717), 
         .D(n29200), .Z(n605_adj_2750)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9385_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i18858 (.BLUT(n21176), .ALUT(n21177), .C0(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_2142[11]));
    LUT4 i20628_3_lut (.A(n22964), .B(n22965), .C(index_i[8]), .Z(n22967)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20628_3_lut.init = 16'hcaca;
    LUT4 i9406_3_lut_3_lut_4_lut (.A(index_q[3]), .B(index_q[4]), .C(n29197), 
         .D(index_q[0]), .Z(n605_adj_2767)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9406_3_lut_3_lut_4_lut.init = 16'h10fe;
    LUT4 i9436_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n875_adj_2597)) /* synthesis lut_function=(A (C (D))+!A !(B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9436_3_lut_4_lut_4_lut_4_lut.init = 16'hb555;
    LUT4 i9614_3_lut_4_lut_3_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[4]), 
         .Z(n12064)) /* synthesis lut_function=(A (B)+!A !(B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9614_3_lut_4_lut_3_lut.init = 16'h9898;
    LUT4 i20611_3_lut (.A(n22945), .B(n22946), .C(index_i[7]), .Z(n22950)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20611_3_lut.init = 16'hcaca;
    PFUMX i22851 (.BLUT(n24456), .ALUT(n24455), .C0(index_q[5]), .Z(n24457));
    LUT4 i11806_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(n26547), .C(index_i[4]), 
         .D(index_i[0]), .Z(n14366)) /* synthesis lut_function=(!(A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11806_3_lut_4_lut_4_lut_4_lut.init = 16'h55d5;
    LUT4 i1_2_lut_rep_625 (.A(index_q[3]), .B(index_q[2]), .Z(n26585)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_2_lut_rep_625.init = 16'heeee;
    LUT4 mux_192_Mux_6_i204_3_lut_3_lut_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n204_adj_2732)) /* synthesis lut_function=(!(A (C)+!A !((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_6_i204_3_lut_3_lut_3_lut.init = 16'h5b5b;
    LUT4 mux_192_Mux_6_i498_3_lut_4_lut_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n498)) /* synthesis lut_function=(A (B+!(C))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_6_i498_3_lut_4_lut_3_lut.init = 16'h9b9b;
    LUT4 i22497_2_lut_rep_500_3_lut_4_lut (.A(index_q[3]), .B(index_q[2]), 
         .C(index_q[1]), .D(index_q[0]), .Z(n26460)) /* synthesis lut_function=(!(A+(B+(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i22497_2_lut_rep_500_3_lut_4_lut.init = 16'h0111;
    L6MUX21 i23788 (.D0(n25468), .D1(n25466), .SD(index_q[5]), .Z(n25469));
    LUT4 i11732_2_lut_rep_517_3_lut (.A(index_q[3]), .B(index_q[2]), .C(index_q[1]), 
         .Z(n26477)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11732_2_lut_rep_517_3_lut.init = 16'hfefe;
    LUT4 i20735_3_lut (.A(n23071), .B(n23072), .C(index_q[7]), .Z(n23074)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20735_3_lut.init = 16'hcaca;
    LUT4 i9412_3_lut_3_lut_4_lut (.A(index_q[3]), .B(index_q[2]), .C(index_q[1]), 
         .D(index_q[0]), .Z(n812_adj_2583)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9412_3_lut_3_lut_4_lut.init = 16'h1ef0;
    PFUMX i23786 (.BLUT(n572_adj_2777), .ALUT(n25467), .C0(index_q[4]), 
          .Z(n25468));
    LUT4 i20603_3_lut (.A(n22929), .B(n24642), .C(index_i[6]), .Z(n22942)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20603_3_lut.init = 16'hcaca;
    LUT4 i9431_2_lut_3_lut (.A(index_q[1]), .B(index_q[2]), .C(index_q[3]), 
         .Z(n11877)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9431_2_lut_3_lut.init = 16'h8080;
    LUT4 mux_191_Mux_6_i924_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[4]), .D(n762_adj_2668), .Z(n924_adj_2748)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_6_i924_3_lut_4_lut.init = 16'h6f60;
    PFUMX i23783 (.BLUT(n25465), .ALUT(n25464), .C0(index_q[4]), .Z(n25466));
    LUT4 mux_191_Mux_3_i94_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[4]), .D(n93_adj_2587), .Z(n94_adj_2559)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_3_i94_3_lut_4_lut.init = 16'hf606;
    LUT4 i20734_3_lut (.A(n23069), .B(n23070), .C(index_q[7]), .Z(n23073)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20734_3_lut.init = 16'hcaca;
    LUT4 mux_191_Mux_3_i62_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[4]), .D(n812_adj_2650), .Z(n62_adj_2763)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_3_i62_3_lut_4_lut.init = 16'h6f60;
    L6MUX21 i22842 (.D0(n24444), .D1(n24442), .SD(index_i[6]), .Z(n24445));
    PFUMX i22840 (.BLUT(n24443), .ALUT(n62_adj_2271), .C0(index_i[5]), 
          .Z(n24444));
    LUT4 i20113_3_lut (.A(n25231), .B(n22443), .C(index_i[6]), .Z(n22452)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20113_3_lut.init = 16'hcaca;
    LUT4 n25854_bdd_3_lut_3_lut (.A(n1021), .B(index_i[8]), .C(n25854), 
         .Z(n25855)) /* synthesis lut_function=(A (B+(C))+!A !(B+!(C))) */ ;
    defparam n25854_bdd_3_lut_3_lut.init = 16'hb8b8;
    PFUMX i22838 (.BLUT(n24441), .ALUT(n24440), .C0(index_i[5]), .Z(n24442));
    L6MUX21 i23769 (.D0(n25451), .D1(n25448), .SD(index_q[5]), .Z(n25452));
    PFUMX i23767 (.BLUT(n25450), .ALUT(n25449), .C0(index_q[4]), .Z(n25451));
    LUT4 mux_191_Mux_4_i221_3_lut_3_lut (.A(index_i[0]), .B(index_i[4]), 
         .C(n205_adj_2782), .Z(n221_adj_2530)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_4_i221_3_lut_3_lut.init = 16'h7474;
    LUT4 i9557_3_lut_4_lut_4_lut (.A(index_i[0]), .B(n773), .C(index_i[4]), 
         .D(n26637), .Z(n12003)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B ((D)+!C)+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9557_3_lut_4_lut_4_lut.init = 16'h5c0c;
    LUT4 index_q_0__bdd_4_lut_24853 (.A(index_q[0]), .B(index_q[3]), .C(index_q[1]), 
         .D(index_q[2]), .Z(n26774)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C (D)))+!A !(B (C+!(D))+!B !(C+(D))))) */ ;
    defparam index_q_0__bdd_4_lut_24853.init = 16'h4ae7;
    LUT4 i19797_3_lut (.A(n22131), .B(n22132), .C(index_q[7]), .Z(n22136)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19797_3_lut.init = 16'hcaca;
    PFUMX i23764 (.BLUT(n26370), .ALUT(n25447), .C0(index_q[4]), .Z(n25448));
    LUT4 i19069_3_lut (.A(n1001), .B(n931), .C(index_q[3]), .Z(n21389)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19069_3_lut.init = 16'hcaca;
    LUT4 i19327_3_lut_4_lut_4_lut (.A(index_i[0]), .B(n26708), .C(index_i[3]), 
         .D(n26637), .Z(n21647)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19327_3_lut_4_lut_4_lut.init = 16'hc5c0;
    LUT4 i11804_2_lut_rep_476_3_lut_3_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[1]), .Z(n26436)) /* synthesis lut_function=((B (C))+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11804_2_lut_rep_476_3_lut_3_lut.init = 16'hd5d5;
    LUT4 i11103_2_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n844_adj_2737)) /* synthesis lut_function=(A (B+!(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11103_2_lut_3_lut_4_lut.init = 16'h9ff9;
    LUT4 i21429_3_lut (.A(n21389), .B(n21390), .C(index_q[4]), .Z(n21391)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21429_3_lut.init = 16'hcaca;
    LUT4 i9383_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n541)) /* synthesis lut_function=(A (B (C (D))+!B !(C (D)))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9383_3_lut_4_lut_4_lut_4_lut.init = 16'h9333;
    LUT4 mux_191_Mux_9_i62_3_lut_4_lut_then_4_lut (.A(index_i[4]), .B(index_i[2]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n26862)) /* synthesis lut_function=(!(A (B (C+(D)))+!A (B+(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_9_i62_3_lut_4_lut_then_4_lut.init = 16'h222b;
    LUT4 i11508_2_lut_rep_426_3_lut_4_lut (.A(index_q[2]), .B(index_q[3]), 
         .C(index_q[4]), .D(n26567), .Z(n26386)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11508_2_lut_rep_426_3_lut_4_lut.init = 16'hf8f0;
    LUT4 mux_191_Mux_9_i62_3_lut_4_lut_else_4_lut (.A(index_i[4]), .B(index_i[2]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n26861)) /* synthesis lut_function=((B+(C (D)))+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_9_i62_3_lut_4_lut_else_4_lut.init = 16'hfddd;
    LUT4 mux_191_Mux_6_i204_3_lut_4_lut_3_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .Z(n204)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_6_i204_3_lut_4_lut_3_lut_3_lut.init = 16'h3d3d;
    LUT4 n21654_bdd_3_lut_3_lut (.A(index_i[1]), .B(n526_adj_2261), .C(index_i[4]), 
         .Z(n24539)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n21654_bdd_3_lut_3_lut.init = 16'h5c5c;
    LUT4 mux_191_Mux_1_i890_4_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[3]), 
         .C(n70), .D(index_i[4]), .Z(n890_adj_2725)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (D))+!A !((C+(D))+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_1_i890_4_lut_4_lut_4_lut_4_lut.init = 16'h55f3;
    LUT4 mux_191_Mux_6_i636_4_lut_4_lut (.A(index_i[1]), .B(index_i[4]), 
         .C(n635_adj_2731), .D(n14367), .Z(n636_adj_2689)) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_6_i636_4_lut_4_lut.init = 16'hf3d1;
    LUT4 i12193_1_lut_2_lut_3_lut_4_lut (.A(n26526), .B(index_q[3]), .C(index_q[5]), 
         .D(index_q[4]), .Z(n381_adj_2446)) /* synthesis lut_function=(!(A (C+(D))+!A (B (C+(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12193_1_lut_2_lut_3_lut_4_lut.init = 16'h010f;
    LUT4 i19264_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21584)) /* synthesis lut_function=(A (B (C (D))+!B !(C (D)))+!A !(B (D)+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19264_3_lut_4_lut_4_lut.init = 16'h9366;
    LUT4 i11530_3_lut_3_lut_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[0]), 
         .Z(n619)) /* synthesis lut_function=(!(A ((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11530_3_lut_3_lut_3_lut.init = 16'h5d5d;
    LUT4 i11669_4_lut (.A(n26495), .B(index_q[7]), .C(n892_adj_2542), 
         .D(index_q[6]), .Z(n1021_adj_2728)) /* synthesis lut_function=(A (B+(C (D)))+!A (B+(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11669_4_lut.init = 16'hfcdd;
    LUT4 i11582_2_lut_rep_642 (.A(index_i[1]), .B(index_i[0]), .Z(n26602)) /* synthesis lut_function=((B)+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11582_2_lut_rep_642.init = 16'hdddd;
    LUT4 mux_191_Mux_2_i349_3_lut_3_lut (.A(index_i[0]), .B(index_i[4]), 
         .C(n348_adj_2783), .Z(n349_adj_2596)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_2_i349_3_lut_3_lut.init = 16'hd1d1;
    LUT4 i19273_3_lut_4_lut_4_lut (.A(index_i[0]), .B(n26709), .C(index_i[3]), 
         .D(n26546), .Z(n21593)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19273_3_lut_4_lut_4_lut.init = 16'hcfc5;
    LUT4 i11479_4_lut (.A(n14756), .B(index_i[7]), .C(n892_adj_2546), 
         .D(index_i[6]), .Z(n1021)) /* synthesis lut_function=(A (B+(C (D)))+!A (B+(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11479_4_lut.init = 16'hfcdd;
    LUT4 i11522_3_lut_3_lut_3_lut_rep_644 (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .Z(n26604)) /* synthesis lut_function=(!(A+!(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11522_3_lut_3_lut_3_lut_rep_644.init = 16'h4545;
    LUT4 mux_191_Mux_2_i507_3_lut_3_lut (.A(index_i[0]), .B(index_i[4]), 
         .C(n491_adj_2745), .Z(n507_adj_2609)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_2_i507_3_lut_3_lut.init = 16'h7474;
    LUT4 mux_191_Mux_5_i573_3_lut_3_lut (.A(index_i[0]), .B(index_i[4]), 
         .C(n572_adj_2784), .Z(n573_adj_2489)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_5_i573_3_lut_3_lut.init = 16'hd1d1;
    LUT4 mux_191_Mux_2_i763_4_lut_4_lut (.A(index_i[0]), .B(n11995), .C(index_i[4]), 
         .D(n157_adj_2785), .Z(n763_adj_2617)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_2_i763_4_lut_4_lut.init = 16'hdfd0;
    LUT4 mux_191_Mux_0_i684_3_lut_4_lut_4_lut (.A(index_i[0]), .B(n26685), 
         .C(index_i[3]), .D(n26637), .Z(n684_adj_2700)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B ((D)+!C)+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_0_i684_3_lut_4_lut_4_lut.init = 16'h5c0c;
    LUT4 mux_191_Mux_8_i85_3_lut_rep_645 (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .Z(n26605)) /* synthesis lut_function=(A (B (C))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_8_i85_3_lut_rep_645.init = 16'h9191;
    LUT4 i11807_2_lut_3_lut_3_lut (.A(index_i[0]), .B(index_i[3]), .C(index_i[2]), 
         .Z(n14367)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11807_2_lut_3_lut_3_lut.init = 16'h4040;
    LUT4 mux_192_Mux_10_i252_3_lut_4_lut_4_lut (.A(n26526), .B(index_q[3]), 
         .C(index_q[4]), .D(n29190), .Z(n252_adj_2483)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B (C (D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_10_i252_3_lut_4_lut_4_lut.init = 16'h3efe;
    LUT4 mux_191_Mux_2_i859_3_lut_4_lut_4_lut (.A(index_i[0]), .B(n26599), 
         .C(index_i[3]), .D(n26637), .Z(n859)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B ((D)+!C)+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_2_i859_3_lut_4_lut_4_lut.init = 16'h5c0c;
    LUT4 i22335_2_lut_rep_724 (.A(index_i[0]), .B(index_i[1]), .Z(n26684)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i22335_2_lut_rep_724.init = 16'h9999;
    LUT4 mux_191_Mux_6_i573_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[4]), .D(n572_adj_2786), .Z(n573_adj_2685)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_6_i573_3_lut_4_lut.init = 16'hf909;
    LUT4 mux_191_Mux_7_i45_3_lut_3_lut_rep_647_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26607)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_7_i45_3_lut_3_lut_rep_647_3_lut.init = 16'h3939;
    LUT4 mux_191_Mux_4_i77_3_lut_3_lut_rep_628_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26588)) /* synthesis lut_function=(A (B (C))+!A !(B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_4_i77_3_lut_3_lut_rep_628_3_lut.init = 16'h9595;
    LUT4 mux_191_Mux_6_i498_3_lut_4_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n404)) /* synthesis lut_function=(A (B+!(C))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_6_i498_3_lut_4_lut_4_lut_3_lut.init = 16'h9b9b;
    LUT4 i15433_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n17583)) /* synthesis lut_function=(A (B)+!A !(B (C (D))+!B !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i15433_3_lut_4_lut_4_lut.init = 16'h9ccc;
    LUT4 mux_191_Mux_4_i142_3_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[3]), 
         .C(index_i[2]), .Z(n142_adj_2418)) /* synthesis lut_function=(A (B (C))+!A !(B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_4_i142_3_lut_4_lut_3_lut.init = 16'h9595;
    LUT4 mux_191_Mux_4_i340_3_lut_rep_627 (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[1]), .Z(n26587)) /* synthesis lut_function=(A ((C)+!B)+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_4_i340_3_lut_rep_627.init = 16'he6e6;
    LUT4 mux_191_Mux_8_i93_3_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .D(index_i[3]), .Z(n93_adj_2671)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(D))+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_8_i93_3_lut_3_lut_4_lut.init = 16'h3391;
    LUT4 i9513_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n541_adj_2658)) /* synthesis lut_function=(A (B (C (D))+!B !(C (D)))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9513_3_lut_4_lut_4_lut_4_lut.init = 16'h9333;
    LUT4 mux_191_Mux_5_i505_3_lut_4_lut_3_lut_rep_631 (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[1]), .Z(n26591)) /* synthesis lut_function=(A (B+(C))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_5_i505_3_lut_4_lut_3_lut_rep_631.init = 16'hb9b9;
    LUT4 i19378_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n21698)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !(B (C+!(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19378_3_lut_4_lut_4_lut.init = 16'ha5a9;
    LUT4 mux_191_Mux_5_i572_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n572_adj_2784)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A !(B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_5_i572_3_lut_4_lut_4_lut.init = 16'ha9a5;
    LUT4 i11527_2_lut_rep_634 (.A(index_i[0]), .B(index_i[1]), .Z(n26594)) /* synthesis lut_function=((B)+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11527_2_lut_rep_634.init = 16'hdddd;
    LUT4 mux_191_Mux_0_i635_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n635_adj_2667)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_0_i635_3_lut_4_lut_4_lut.init = 16'hfd0a;
    LUT4 i19216_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n21536)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (D))+!A !(D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19216_3_lut_4_lut_4_lut_4_lut.init = 16'ha25d;
    LUT4 mux_191_Mux_3_i444_3_lut_4_lut (.A(index_i[0]), .B(index_i[3]), 
         .C(n26546), .D(index_i[4]), .Z(n444_adj_2567)) /* synthesis lut_function=(!(A (B (D)+!B (C (D)))+!A !(B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_3_i444_3_lut_4_lut.init = 16'h46aa;
    LUT4 mux_191_Mux_1_i93_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n93_adj_2686)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C+(D)))+!A !(B (C (D)+!C !(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_1_i93_3_lut_4_lut_4_lut_4_lut.init = 16'h955a;
    LUT4 i11615_2_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n844_adj_2740)) /* synthesis lut_function=(A (B+!(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11615_2_lut_3_lut_4_lut.init = 16'h9ff9;
    LUT4 mux_191_Mux_7_i620_3_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .D(index_i[3]), .Z(n620_adj_2284)) /* synthesis lut_function=(A (B (C+!(D)))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_7_i620_3_lut_4_lut_4_lut.init = 16'h9199;
    LUT4 mux_191_Mux_2_i908_3_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .D(index_i[3]), .Z(n908_adj_2657)) /* synthesis lut_function=(!(A (B+!(D))+!A !(B+!(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_2_i908_3_lut_4_lut_4_lut.init = 16'h6645;
    LUT4 n53_bdd_3_lut_4_lut_4_lut_adj_85 (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[1]), .D(index_i[3]), .Z(n24945)) /* synthesis lut_function=(A (B+!((D)+!C))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n53_bdd_3_lut_4_lut_4_lut_adj_85.init = 16'h99b9;
    LUT4 i19366_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[2]), .C(index_i[1]), 
         .D(index_i[3]), .Z(n21686)) /* synthesis lut_function=(!(A (B (D)+!B !(C+(D)))+!A !(B (D)+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19366_3_lut_4_lut_4_lut.init = 16'h66b9;
    LUT4 mux_191_Mux_0_i796_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[1]), .D(index_i[3]), .Z(n796_adj_2712)) /* synthesis lut_function=(A (B (C+(D))+!B (C (D)))+!A !(B ((D)+!C)+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_0_i796_3_lut_4_lut_4_lut.init = 16'hb9c0;
    LUT4 i9541_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(n26547), .D(index_i[4]), .Z(n189_adj_2778)) /* synthesis lut_function=(A (B (C (D)))+!A !(B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9541_3_lut_4_lut_4_lut_4_lut.init = 16'h9555;
    LUT4 mux_191_Mux_4_i252_4_lut_4_lut (.A(index_i[0]), .B(index_i[3]), 
         .C(n26637), .D(index_i[4]), .Z(n252_adj_2531)) /* synthesis lut_function=(!(A (B (D)+!B !(D))+!A !(B ((D)+!C)+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_4_i252_4_lut_4_lut.init = 16'h669d;
    LUT4 mux_191_Mux_1_i62_3_lut_4_lut (.A(index_i[0]), .B(index_i[3]), 
         .C(index_i[2]), .D(index_i[4]), .Z(n62_adj_2762)) /* synthesis lut_function=(A (B (D)+!B ((D)+!C))+!A !(B (D)+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_1_i62_3_lut_4_lut.init = 16'haa56;
    LUT4 i19387_3_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[0]), 
         .D(index_i[3]), .Z(n21707)) /* synthesis lut_function=(!(A ((D)+!B)+!A !(B (D)+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19387_3_lut_4_lut_4_lut.init = 16'h4588;
    LUT4 i19303_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[2]), .C(index_i[1]), 
         .D(index_i[3]), .Z(n21623)) /* synthesis lut_function=(A ((C (D))+!B)+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19303_3_lut_4_lut_4_lut.init = 16'he666;
    LUT4 i7509_2_lut_rep_635 (.A(index_i[3]), .B(index_i[4]), .Z(n26595)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i7509_2_lut_rep_635.init = 16'heeee;
    LUT4 i9529_3_lut_3_lut_4_lut (.A(index_i[3]), .B(index_i[4]), .C(n26709), 
         .D(index_i[0]), .Z(n605)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9529_3_lut_3_lut_4_lut.init = 16'h10fe;
    LUT4 i9515_3_lut_4_lut (.A(index_i[3]), .B(index_i[4]), .C(n26684), 
         .D(n29180), .Z(n605_adj_2688)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9515_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i19381_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[0]), 
         .D(index_i[3]), .Z(n21701)) /* synthesis lut_function=(!(A (B (D)+!B !(C+!(D)))+!A !(B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19381_3_lut_4_lut.init = 16'h64aa;
    LUT4 mux_191_Mux_2_i604_3_lut_4_lut_4_lut_4_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n604_adj_2699)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)+!C !(D)))+!A (B (C)+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_2_i604_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'h3c9f;
    PFUMX i20557 (.BLUT(n142_adj_2448), .ALUT(n157_adj_2263), .C0(index_q[4]), 
          .Z(n22896));
    LUT4 i19309_3_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[0]), 
         .D(index_i[3]), .Z(n21629)) /* synthesis lut_function=(!(A (B+!(C+(D)))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19309_3_lut_4_lut_4_lut.init = 16'h6664;
    LUT4 i22171_3_lut (.A(n12019), .B(n892_adj_2723), .C(index_q[6]), 
         .Z(n22306)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22171_3_lut.init = 16'hcaca;
    LUT4 index_i_5__bdd_4_lut_24068_4_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n25337)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B (C)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam index_i_5__bdd_4_lut_24068_4_lut_4_lut.init = 16'h3d2d;
    LUT4 mux_192_Mux_5_i109_3_lut_3_lut_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .Z(n109_adj_2511)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_5_i109_3_lut_3_lut_3_lut.init = 16'h3939;
    LUT4 i11603_2_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n668_adj_2681)) /* synthesis lut_function=(!(A ((D)+!B)+!A (B ((D)+!C)+!B (C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11603_2_lut_4_lut_4_lut_4_lut.init = 16'h00c9;
    L6MUX21 i23673 (.D0(n25356), .D1(n25353), .SD(index_q[5]), .Z(n25357));
    PFUMX i23671 (.BLUT(n25355), .ALUT(n25354), .C0(index_q[4]), .Z(n25356));
    LUT4 mux_191_Mux_6_i435_3_lut_4_lut_4_lut_3_lut_rep_648 (.A(index_i[1]), 
         .B(index_i[0]), .C(index_i[2]), .Z(n26608)) /* synthesis lut_function=(A (B+(C))+!A !(B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_6_i435_3_lut_4_lut_4_lut_3_lut_rep_648.init = 16'hbdbd;
    LUT4 mux_191_Mux_5_i109_3_lut_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .Z(n109_adj_2730)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_5_i109_3_lut_3_lut_3_lut.init = 16'h3939;
    PFUMX i20558 (.BLUT(n173_adj_2478), .ALUT(n188), .C0(index_q[4]), 
          .Z(n22897));
    LUT4 i11295_2_lut_rep_578 (.A(index_q[1]), .B(index_q[2]), .Z(n26538)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11295_2_lut_rep_578.init = 16'h8888;
    LUT4 i19349_3_lut_4_lut (.A(index_i[1]), .B(index_i[0]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21669)) /* synthesis lut_function=(A (B+(C+(D)))+!A !(B (C+(D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19349_3_lut_4_lut.init = 16'haabd;
    PFUMX i23668 (.BLUT(n875_adj_2571), .ALUT(n25352), .C0(index_q[4]), 
          .Z(n25353));
    LUT4 i9609_3_lut_3_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n12059)) /* synthesis lut_function=(!(A (B (D)+!B !(C+(D)))+!A (B (C+(D))+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9609_3_lut_3_lut_4_lut_4_lut.init = 16'h22bd;
    LUT4 i9423_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(n26539), .D(index_q[4]), .Z(n189_adj_2727)) /* synthesis lut_function=(A (B (C (D)))+!A !(B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9423_3_lut_4_lut_4_lut_4_lut.init = 16'h9555;
    LUT4 mux_191_Mux_0_i364_3_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n364_adj_2780)) /* synthesis lut_function=(A (B (D)+!B (C+!(D)))+!A !(B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_0_i364_3_lut_3_lut_4_lut.init = 16'hbd33;
    LUT4 i19388_3_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[0]), 
         .D(index_i[3]), .Z(n21708)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A (B (C)+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19388_3_lut_4_lut_4_lut.init = 16'h3c9d;
    PFUMX i20563 (.BLUT(n333_adj_2768), .ALUT(n348_adj_2376), .C0(index_q[4]), 
          .Z(n22902));
    LUT4 i15434_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n17584)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i15434_3_lut_4_lut_4_lut_4_lut.init = 16'h3999;
    PFUMX i23654 (.BLUT(n25337), .ALUT(n25336), .C0(index_i[5]), .Z(n25338));
    LUT4 mux_191_Mux_2_i836_3_lut_4_lut_3_lut_rep_725 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26685)) /* synthesis lut_function=(A (B)+!A !(B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_2_i836_3_lut_4_lut_3_lut_rep_725.init = 16'h9898;
    LUT4 mux_191_Mux_4_i262_3_lut_3_lut_rep_726 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26686)) /* synthesis lut_function=(A (B+(C))+!A !(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_4_i262_3_lut_3_lut_rep_726.init = 16'ha9a9;
    LUT4 mux_191_Mux_6_i378_3_lut_4_lut_3_lut_rep_727 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26687)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_6_i378_3_lut_4_lut_3_lut_rep_727.init = 16'h4949;
    L6MUX21 i19957 (.D0(n22291), .D1(n22292), .SD(index_q[7]), .Z(n22296));
    LUT4 i11273_2_lut_rep_424_3_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .D(index_q[0]), .Z(n26384)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11273_2_lut_rep_424_3_lut_4_lut.init = 16'hf8f0;
    PFUMX i23645 (.BLUT(n25328), .ALUT(n25327), .C0(index_i[4]), .Z(n25329));
    LUT4 mux_191_Mux_6_i505_3_lut_rep_728 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26688)) /* synthesis lut_function=(A (B)+!A (B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_6_i505_3_lut_rep_728.init = 16'hc9c9;
    LUT4 i11099_2_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n668_adj_2436)) /* synthesis lut_function=(!(A ((D)+!B)+!A (B ((D)+!C)+!B (C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11099_2_lut_4_lut_4_lut_4_lut.init = 16'h00c9;
    LUT4 mux_191_Mux_5_i38_3_lut_3_lut_4_lut_3_lut_rep_729 (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[2]), .Z(n26689)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_5_i38_3_lut_3_lut_4_lut_3_lut_rep_729.init = 16'h1919;
    LUT4 mux_191_Mux_7_i77_3_lut_3_lut_rep_731 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26691)) /* synthesis lut_function=(A (B)+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_7_i77_3_lut_3_lut_rep_731.init = 16'h9c9c;
    LUT4 mux_191_Mux_3_i676_3_lut_4_lut_3_lut_rep_732 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26692)) /* synthesis lut_function=(A (B (C))+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_3_i676_3_lut_4_lut_3_lut_rep_732.init = 16'h9494;
    LUT4 i19393_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21713)) /* synthesis lut_function=(A (B (C)+!B (C (D)+!C !(D)))+!A !(B (C+!(D))+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19393_3_lut_4_lut_4_lut.init = 16'ha593;
    LUT4 n20976_bdd_3_lut_23380 (.A(n26544), .B(n26727), .C(index_q[3]), 
         .Z(n25070)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n20976_bdd_3_lut_23380.init = 16'hcaca;
    LUT4 mux_192_Mux_5_i781_3_lut_4_lut_4_lut_then_4_lut (.A(index_q[3]), 
         .B(index_q[0]), .C(index_q[4]), .D(index_q[2]), .Z(n26771)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_5_i781_3_lut_4_lut_4_lut_then_4_lut.init = 16'hece0;
    LUT4 mux_191_Mux_3_i684_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[4]), .Z(n684_adj_2759)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A !(B ((D)+!C)+!B (C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_3_i684_3_lut_3_lut_4_lut.init = 16'h5594;
    LUT4 mux_192_Mux_5_i572_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n572_adj_2777)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A !(B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_5_i572_3_lut_4_lut_4_lut.init = 16'ha9a5;
    LUT4 mux_191_Mux_2_i653_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n653_adj_2696)) /* synthesis lut_function=(A (B (C+!(D))+!B !(D))+!A !(B (C+!(D))+!B !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_2_i653_3_lut_4_lut.init = 16'h94aa;
    LUT4 mux_191_Mux_1_i557_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n557_adj_2755)) /* synthesis lut_function=(A (B (C+(D)))+!A (B ((D)+!C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_1_i557_3_lut_4_lut.init = 16'hcc94;
    LUT4 mux_191_Mux_3_i859_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n859_adj_2721)) /* synthesis lut_function=(!(A (B (D)+!B !(D))+!A (B (C+(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_3_i859_3_lut_3_lut_4_lut.init = 16'h339c;
    LUT4 mux_191_Mux_6_i572_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n572_adj_2786)) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_6_i572_3_lut_4_lut.init = 16'hccd9;
    LUT4 i19258_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21578)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(D))+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19258_3_lut_3_lut_4_lut.init = 16'h3319;
    LUT4 n12055_bdd_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[4]), 
         .D(index_i[2]), .Z(n25485)) /* synthesis lut_function=(A (B)+!A !(B (D)+!B !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n12055_bdd_3_lut_4_lut.init = 16'h98cc;
    LUT4 i19403_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21723)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C+(D)))+!A (B (C)+!B !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19403_3_lut_4_lut_4_lut.init = 16'hc95a;
    LUT4 i20797_3_lut (.A(n23133), .B(n23134), .C(index_i[7]), .Z(n23136)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20797_3_lut.init = 16'hcaca;
    L6MUX21 i22776 (.D0(n24361), .D1(n24359), .SD(index_q[6]), .Z(n24362));
    LUT4 i19369_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21689)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (D))+!A !(B (C (D))+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19369_3_lut_3_lut_4_lut.init = 16'h4933;
    LUT4 i19324_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21644)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A !(B (D)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19324_3_lut_3_lut_4_lut.init = 16'ha955;
    LUT4 i19480_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n21800)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !(B (C+!(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19480_3_lut_4_lut_4_lut.init = 16'ha5a9;
    L6MUX21 i23628 (.D0(n25311), .D1(n25308), .SD(index_q[5]), .Z(n25312));
    LUT4 mux_191_Mux_3_i397_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n397_adj_2713)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !(B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_3_i397_3_lut_4_lut_4_lut.init = 16'ha95a;
    LUT4 mux_191_Mux_0_i762_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n762_adj_2704)) /* synthesis lut_function=(A (B+!((D)+!C))+!A !(B (D)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_0_i762_3_lut_4_lut_4_lut.init = 16'h98fc;
    LUT4 i20796_3_lut (.A(n23131), .B(n23132), .C(index_i[7]), .Z(n23135)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20796_3_lut.init = 16'hcaca;
    PFUMX i23626 (.BLUT(n25310), .ALUT(n25309), .C0(index_q[4]), .Z(n25311));
    LUT4 i11569_2_lut_rep_734 (.A(index_i[0]), .B(index_i[1]), .Z(n26694)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11569_2_lut_rep_734.init = 16'h2222;
    PFUMX i22774 (.BLUT(n924_adj_2773), .ALUT(n24360), .C0(index_q[5]), 
          .Z(n24361));
    LUT4 mux_191_Mux_4_i723_3_lut_4_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n723)) /* synthesis lut_function=(A ((C)+!B)+!A !(B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_4_i723_3_lut_4_lut_4_lut_3_lut.init = 16'hb2b2;
    LUT4 i20226_3_lut_4_lut (.A(n26526), .B(index_q[3]), .C(index_q[4]), 
         .D(n26460), .Z(n22565)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20226_3_lut_4_lut.init = 16'hfe0e;
    PFUMX i23623 (.BLUT(n25307), .ALUT(n316), .C0(index_q[4]), .Z(n25308));
    LUT4 i11528_2_lut_rep_637 (.A(index_i[0]), .B(index_i[1]), .Z(n26597)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11528_2_lut_rep_637.init = 16'h4444;
    LUT4 i15427_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n17577)) /* synthesis lut_function=(A (B)+!A !(B (C (D))+!B !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i15427_3_lut_4_lut_4_lut.init = 16'h9ccc;
    L6MUX21 i22635 (.D0(n24167), .D1(n26346), .SD(index_q[6]), .Z(n24168));
    LUT4 i19926_3_lut (.A(n22260), .B(n22261), .C(index_q[7]), .Z(n22265)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19926_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_3_i828_3_lut_3_lut_4_lut (.A(n26526), .B(index_q[3]), 
         .C(n157_adj_2452), .D(index_q[4]), .Z(n828_adj_2277)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_3_i828_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 mux_191_Mux_2_i348_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n348_adj_2783)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)+!C !(D)))+!A !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_2_i348_3_lut_4_lut_4_lut_4_lut.init = 16'h5a25;
    PFUMX i22633 (.BLUT(n24166), .ALUT(n24165), .C0(index_q[5]), .Z(n24167));
    LUT4 mux_191_Mux_4_i205_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n205_adj_2782)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_4_i205_3_lut_4_lut_4_lut.init = 16'h5a2a;
    L6MUX21 i23591 (.D0(n25275), .D1(n25273), .SD(index_i[4]), .Z(n25276));
    LUT4 mux_192_Mux_6_i573_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[4]), .D(n572), .Z(n573_adj_2749)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_6_i573_3_lut_4_lut.init = 16'hf909;
    LUT4 mux_191_Mux_4_i204_3_lut_3_lut_rep_632_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26592)) /* synthesis lut_function=(!(A (B+(C))+!A !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_4_i204_3_lut_3_lut_rep_632_3_lut.init = 16'h5252;
    LUT4 i19213_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n21533)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (D))+!A !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19213_3_lut_4_lut_4_lut_4_lut.init = 16'h55a2;
    PFUMX i23589 (.BLUT(n26397), .ALUT(n25274), .C0(index_i[5]), .Z(n25275));
    PFUMX i23587 (.BLUT(n25272), .ALUT(n25271), .C0(index_i[5]), .Z(n25273));
    PFUMX i20564 (.BLUT(n364), .ALUT(n379_adj_2355), .C0(index_q[4]), 
          .Z(n22903));
    LUT4 mux_191_Mux_6_i157_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n157_adj_2785)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (D))+!A !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_6_i157_3_lut_4_lut_4_lut_4_lut.init = 16'h5d22;
    L6MUX21 i23579 (.D0(n25264), .D1(n25261), .SD(index_i[5]), .Z(n25265));
    PFUMX i23577 (.BLUT(n25263), .ALUT(n25262), .C0(index_i[4]), .Z(n25264));
    PFUMX i20565 (.BLUT(n397_adj_2344), .ALUT(n412), .C0(index_q[4]), 
          .Z(n22904));
    PFUMX i23574 (.BLUT(n301_adj_2256), .ALUT(n25260), .C0(index_i[4]), 
          .Z(n25261));
    PFUMX i20566 (.BLUT(n428), .ALUT(n443_adj_2306), .C0(index_q[4]), 
          .Z(n22905));
    LUT4 mux_191_Mux_0_i985_3_lut_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n985_adj_2628)) /* synthesis lut_function=(!(A (B+!(C))+!A (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_0_i985_3_lut_3_lut_3_lut.init = 16'h2525;
    PFUMX i20567 (.BLUT(n460_adj_2339), .ALUT(n475_adj_2393), .C0(index_q[4]), 
          .Z(n22906));
    PFUMX i22772 (.BLUT(n24358), .ALUT(n26476), .C0(index_q[5]), .Z(n24359));
    L6MUX21 i23549 (.D0(n25236), .D1(n25234), .SD(index_i[5]), .Z(n25237));
    PFUMX i23547 (.BLUT(n572_adj_2784), .ALUT(n25235), .C0(index_i[4]), 
          .Z(n25236));
    PFUMX i22628 (.BLUT(n21242), .ALUT(n24160), .C0(index_q[6]), .Z(n24161));
    L6MUX21 i22611 (.D0(n24132), .D1(n26347), .SD(index_i[6]), .Z(n24133));
    PFUMX i22609 (.BLUT(n24131), .ALUT(n24130), .C0(index_i[5]), .Z(n24132));
    LUT4 mux_191_Mux_6_i371_3_lut_4_lut_3_lut_rep_735 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26695)) /* synthesis lut_function=(!(A (B+!(C))+!A ((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_6_i371_3_lut_4_lut_3_lut_rep_735.init = 16'h2424;
    PFUMX i23544 (.BLUT(n25233), .ALUT(n25232), .C0(index_i[4]), .Z(n25234));
    L6MUX21 i23542 (.D0(n25230), .D1(n25228), .SD(index_i[4]), .Z(n25231));
    PFUMX i23540 (.BLUT(n25229), .ALUT(n26367), .C0(index_i[5]), .Z(n25230));
    PFUMX i23538 (.BLUT(n25227), .ALUT(n25226), .C0(index_i[5]), .Z(n25228));
    PFUMX i23527 (.BLUT(n25216), .ALUT(n25215), .C0(index_i[4]), .Z(n25217));
    L6MUX21 i23518 (.D0(n25208), .D1(n25205), .SD(index_i[5]), .Z(n25209));
    PFUMX i22604 (.BLUT(n21233), .ALUT(n24125), .C0(index_i[6]), .Z(n24126));
    LUT4 mux_191_Mux_6_i389_3_lut_4_lut_3_lut_rep_737 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26697)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_6_i389_3_lut_4_lut_3_lut_rep_737.init = 16'h9292;
    PFUMX i23516 (.BLUT(n25207), .ALUT(n25206), .C0(index_i[4]), .Z(n25208));
    PFUMX i20568 (.BLUT(n491_adj_2775), .ALUT(n11249), .C0(index_q[4]), 
          .Z(n22907));
    PFUMX i18738 (.BLUT(n21056), .ALUT(n21057), .C0(index_q[4]), .Z(n476_adj_2619));
    LUT4 mux_191_Mux_0_i812_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n812_adj_2716)) /* synthesis lut_function=(A (B (C+(D))+!B !(C))+!A (B (D)+!B !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_0_i812_3_lut_4_lut_4_lut_4_lut.init = 16'hcf92;
    LUT4 mux_192_Mux_5_i38_3_lut_4_lut_3_lut_rep_758 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n26718)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_5_i38_3_lut_4_lut_3_lut_rep_758.init = 16'h1919;
    PFUMX i23513 (.BLUT(n25204), .ALUT(n908), .C0(index_i[4]), .Z(n25205));
    LUT4 i19339_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21659)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C))+!A !(B ((D)+!C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19339_3_lut_4_lut_4_lut.init = 16'h925a;
    LUT4 i8009_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n157_adj_2419)) /* synthesis lut_function=(!(A (C (D))+!A !(B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i8009_3_lut_4_lut_4_lut.init = 16'h4aaa;
    LUT4 mux_192_Mux_2_i262_3_lut_3_lut_rep_759 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n26719)) /* synthesis lut_function=(A (B)+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_2_i262_3_lut_3_lut_rep_759.init = 16'h9c9c;
    LUT4 i19282_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21602)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A !(B (C+!(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19282_3_lut_4_lut_4_lut.init = 16'ha52b;
    LUT4 mux_192_Mux_10_i413_3_lut_3_lut_4_lut (.A(n26526), .B(index_q[3]), 
         .C(n26457), .D(index_q[4]), .Z(n413_adj_2313)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_192_Mux_10_i413_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 i19992_3_lut (.A(n22324), .B(n22325), .C(index_i[7]), .Z(n22331)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19992_3_lut.init = 16'hcaca;
    LUT4 n908_bdd_3_lut_24451_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n25204)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A !(B ((D)+!C)+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n908_bdd_3_lut_24451_3_lut_4_lut.init = 16'h552c;
    LUT4 mux_191_Mux_0_i491_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n491_adj_2781)) /* synthesis lut_function=(!(A (B (D)+!B !(C+!(D)))+!A ((C+!(D))+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_191_Mux_0_i491_3_lut_4_lut.init = 16'h24aa;
    
endmodule
//
// Verilog Description of module \nco(OW=12)_U1 
//

module \nco(OW=12)_U1  (increment, GND_net, o_phase, dac_clk_p_c, n26683) /* synthesis syn_module_defined=1 */ ;
    input [30:0]increment;
    input GND_net;
    output [11:0]o_phase;
    input dac_clk_p_c;
    input n26683;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(29[49:58])
    
    wire n17470;
    wire [31:0]n233;
    wire [31:0]n133;
    
    wire n17471, n17469, n17468, n17467, n17481, n17480, n17479, 
        n17478, n17477, n17476, n17475, n17474, n17473, n17472;
    
    CCU2D phase_register_545_add_4_10 (.A0(increment[8]), .B0(n233[8]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[9]), .B1(n233[9]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17470), .COUT(n17471), .S0(n133[8]), 
          .S1(n133[9]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_545_add_4_10.INIT0 = 16'h5666;
    defparam phase_register_545_add_4_10.INIT1 = 16'h5666;
    defparam phase_register_545_add_4_10.INJECT1_0 = "NO";
    defparam phase_register_545_add_4_10.INJECT1_1 = "NO";
    CCU2D phase_register_545_add_4_8 (.A0(increment[6]), .B0(n233[6]), .C0(GND_net), 
          .D0(GND_net), .A1(increment[7]), .B1(n233[7]), .C1(GND_net), 
          .D1(GND_net), .CIN(n17469), .COUT(n17470), .S0(n133[6]), .S1(n133[7]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_545_add_4_8.INIT0 = 16'h5666;
    defparam phase_register_545_add_4_8.INIT1 = 16'h5666;
    defparam phase_register_545_add_4_8.INJECT1_0 = "NO";
    defparam phase_register_545_add_4_8.INJECT1_1 = "NO";
    CCU2D phase_register_545_add_4_6 (.A0(increment[4]), .B0(n233[4]), .C0(GND_net), 
          .D0(GND_net), .A1(increment[5]), .B1(n233[5]), .C1(GND_net), 
          .D1(GND_net), .CIN(n17468), .COUT(n17469), .S0(n133[4]), .S1(n133[5]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_545_add_4_6.INIT0 = 16'h5666;
    defparam phase_register_545_add_4_6.INIT1 = 16'h5666;
    defparam phase_register_545_add_4_6.INJECT1_0 = "NO";
    defparam phase_register_545_add_4_6.INJECT1_1 = "NO";
    CCU2D phase_register_545_add_4_4 (.A0(increment[2]), .B0(n233[2]), .C0(GND_net), 
          .D0(GND_net), .A1(increment[3]), .B1(n233[3]), .C1(GND_net), 
          .D1(GND_net), .CIN(n17467), .COUT(n17468), .S0(n133[2]), .S1(n133[3]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_545_add_4_4.INIT0 = 16'h5666;
    defparam phase_register_545_add_4_4.INIT1 = 16'h5666;
    defparam phase_register_545_add_4_4.INJECT1_0 = "NO";
    defparam phase_register_545_add_4_4.INJECT1_1 = "NO";
    CCU2D phase_register_545_add_4_2 (.A0(increment[0]), .B0(n233[0]), .C0(GND_net), 
          .D0(GND_net), .A1(increment[1]), .B1(n233[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n17467), .S1(n133[1]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_545_add_4_2.INIT0 = 16'h7000;
    defparam phase_register_545_add_4_2.INIT1 = 16'h5666;
    defparam phase_register_545_add_4_2.INJECT1_0 = "NO";
    defparam phase_register_545_add_4_2.INJECT1_1 = "NO";
    LUT4 i15351_2_lut (.A(increment[0]), .B(n233[0]), .Z(n133[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i15351_2_lut.init = 16'h6666;
    CCU2D phase_register_545_add_4_32 (.A0(increment[30]), .B0(o_phase[10]), 
          .C0(GND_net), .D0(GND_net), .A1(o_phase[11]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n17481), .S0(n133[30]), .S1(n133[31]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_545_add_4_32.INIT0 = 16'h5666;
    defparam phase_register_545_add_4_32.INIT1 = 16'hfaaa;
    defparam phase_register_545_add_4_32.INJECT1_0 = "NO";
    defparam phase_register_545_add_4_32.INJECT1_1 = "NO";
    FD1S3DX phase_register_545__i31 (.D(n133[31]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(o_phase[11])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_545__i31.GSR = "DISABLED";
    FD1S3DX phase_register_545__i30 (.D(n133[30]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(o_phase[10])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_545__i30.GSR = "DISABLED";
    FD1S3DX phase_register_545__i29 (.D(n133[29]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(o_phase[9])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_545__i29.GSR = "DISABLED";
    FD1S3DX phase_register_545__i28 (.D(n133[28]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(o_phase[8])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_545__i28.GSR = "DISABLED";
    FD1S3DX phase_register_545__i27 (.D(n133[27]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(o_phase[7])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_545__i27.GSR = "DISABLED";
    FD1S3DX phase_register_545__i26 (.D(n133[26]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(o_phase[6])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_545__i26.GSR = "DISABLED";
    FD1S3DX phase_register_545__i25 (.D(n133[25]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(o_phase[5])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_545__i25.GSR = "DISABLED";
    FD1S3DX phase_register_545__i24 (.D(n133[24]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(o_phase[4])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_545__i24.GSR = "DISABLED";
    FD1S3DX phase_register_545__i23 (.D(n133[23]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(o_phase[3])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_545__i23.GSR = "DISABLED";
    FD1S3DX phase_register_545__i22 (.D(n133[22]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(o_phase[2])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_545__i22.GSR = "DISABLED";
    FD1S3DX phase_register_545__i21 (.D(n133[21]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(o_phase[1])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_545__i21.GSR = "DISABLED";
    FD1S3DX phase_register_545__i20 (.D(n133[20]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(o_phase[0])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_545__i20.GSR = "DISABLED";
    FD1S3DX phase_register_545__i19 (.D(n133[19]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(n233[19])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_545__i19.GSR = "DISABLED";
    FD1S3DX phase_register_545__i18 (.D(n133[18]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(n233[18])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_545__i18.GSR = "DISABLED";
    FD1S3DX phase_register_545__i17 (.D(n133[17]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(n233[17])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_545__i17.GSR = "DISABLED";
    FD1S3DX phase_register_545__i16 (.D(n133[16]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(n233[16])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_545__i16.GSR = "DISABLED";
    FD1S3DX phase_register_545__i15 (.D(n133[15]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(n233[15])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_545__i15.GSR = "DISABLED";
    FD1S3DX phase_register_545__i14 (.D(n133[14]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(n233[14])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_545__i14.GSR = "DISABLED";
    FD1S3DX phase_register_545__i13 (.D(n133[13]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(n233[13])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_545__i13.GSR = "DISABLED";
    FD1S3DX phase_register_545__i12 (.D(n133[12]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(n233[12])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_545__i12.GSR = "DISABLED";
    FD1S3DX phase_register_545__i11 (.D(n133[11]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(n233[11])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_545__i11.GSR = "DISABLED";
    FD1S3DX phase_register_545__i10 (.D(n133[10]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(n233[10])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_545__i10.GSR = "DISABLED";
    FD1S3DX phase_register_545__i9 (.D(n133[9]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(n233[9])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_545__i9.GSR = "DISABLED";
    FD1S3DX phase_register_545__i8 (.D(n133[8]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(n233[8])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_545__i8.GSR = "DISABLED";
    FD1S3DX phase_register_545__i7 (.D(n133[7]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(n233[7])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_545__i7.GSR = "DISABLED";
    FD1S3DX phase_register_545__i6 (.D(n133[6]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(n233[6])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_545__i6.GSR = "DISABLED";
    FD1S3DX phase_register_545__i5 (.D(n133[5]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(n233[5])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_545__i5.GSR = "DISABLED";
    FD1S3DX phase_register_545__i4 (.D(n133[4]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(n233[4])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_545__i4.GSR = "DISABLED";
    FD1S3DX phase_register_545__i3 (.D(n133[3]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(n233[3])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_545__i3.GSR = "DISABLED";
    FD1S3DX phase_register_545__i2 (.D(n133[2]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(n233[2])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_545__i2.GSR = "DISABLED";
    FD1S3DX phase_register_545__i1 (.D(n133[1]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(n233[1])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_545__i1.GSR = "DISABLED";
    FD1S3DX phase_register_545__i0 (.D(n133[0]), .CK(dac_clk_p_c), .CD(n26683), 
            .Q(n233[0])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_545__i0.GSR = "DISABLED";
    CCU2D phase_register_545_add_4_30 (.A0(increment[28]), .B0(o_phase[8]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[29]), .B1(o_phase[9]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17480), .COUT(n17481), .S0(n133[28]), 
          .S1(n133[29]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_545_add_4_30.INIT0 = 16'h5666;
    defparam phase_register_545_add_4_30.INIT1 = 16'h5666;
    defparam phase_register_545_add_4_30.INJECT1_0 = "NO";
    defparam phase_register_545_add_4_30.INJECT1_1 = "NO";
    CCU2D phase_register_545_add_4_28 (.A0(increment[26]), .B0(o_phase[6]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[27]), .B1(o_phase[7]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17479), .COUT(n17480), .S0(n133[26]), 
          .S1(n133[27]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_545_add_4_28.INIT0 = 16'h5666;
    defparam phase_register_545_add_4_28.INIT1 = 16'h5666;
    defparam phase_register_545_add_4_28.INJECT1_0 = "NO";
    defparam phase_register_545_add_4_28.INJECT1_1 = "NO";
    CCU2D phase_register_545_add_4_26 (.A0(increment[24]), .B0(o_phase[4]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[25]), .B1(o_phase[5]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17478), .COUT(n17479), .S0(n133[24]), 
          .S1(n133[25]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_545_add_4_26.INIT0 = 16'h5666;
    defparam phase_register_545_add_4_26.INIT1 = 16'h5666;
    defparam phase_register_545_add_4_26.INJECT1_0 = "NO";
    defparam phase_register_545_add_4_26.INJECT1_1 = "NO";
    CCU2D phase_register_545_add_4_24 (.A0(increment[22]), .B0(o_phase[2]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[23]), .B1(o_phase[3]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17477), .COUT(n17478), .S0(n133[22]), 
          .S1(n133[23]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_545_add_4_24.INIT0 = 16'h5666;
    defparam phase_register_545_add_4_24.INIT1 = 16'h5666;
    defparam phase_register_545_add_4_24.INJECT1_0 = "NO";
    defparam phase_register_545_add_4_24.INJECT1_1 = "NO";
    CCU2D phase_register_545_add_4_22 (.A0(increment[20]), .B0(o_phase[0]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[21]), .B1(o_phase[1]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17476), .COUT(n17477), .S0(n133[20]), 
          .S1(n133[21]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_545_add_4_22.INIT0 = 16'h5666;
    defparam phase_register_545_add_4_22.INIT1 = 16'h5666;
    defparam phase_register_545_add_4_22.INJECT1_0 = "NO";
    defparam phase_register_545_add_4_22.INJECT1_1 = "NO";
    CCU2D phase_register_545_add_4_20 (.A0(increment[18]), .B0(n233[18]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[19]), .B1(n233[19]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17475), .COUT(n17476), .S0(n133[18]), 
          .S1(n133[19]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_545_add_4_20.INIT0 = 16'h5666;
    defparam phase_register_545_add_4_20.INIT1 = 16'h5666;
    defparam phase_register_545_add_4_20.INJECT1_0 = "NO";
    defparam phase_register_545_add_4_20.INJECT1_1 = "NO";
    CCU2D phase_register_545_add_4_18 (.A0(increment[16]), .B0(n233[16]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[17]), .B1(n233[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17474), .COUT(n17475), .S0(n133[16]), 
          .S1(n133[17]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_545_add_4_18.INIT0 = 16'h5666;
    defparam phase_register_545_add_4_18.INIT1 = 16'h5666;
    defparam phase_register_545_add_4_18.INJECT1_0 = "NO";
    defparam phase_register_545_add_4_18.INJECT1_1 = "NO";
    CCU2D phase_register_545_add_4_16 (.A0(increment[14]), .B0(n233[14]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[15]), .B1(n233[15]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17473), .COUT(n17474), .S0(n133[14]), 
          .S1(n133[15]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_545_add_4_16.INIT0 = 16'h5666;
    defparam phase_register_545_add_4_16.INIT1 = 16'h5666;
    defparam phase_register_545_add_4_16.INJECT1_0 = "NO";
    defparam phase_register_545_add_4_16.INJECT1_1 = "NO";
    CCU2D phase_register_545_add_4_14 (.A0(increment[12]), .B0(n233[12]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[13]), .B1(n233[13]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17472), .COUT(n17473), .S0(n133[12]), 
          .S1(n133[13]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_545_add_4_14.INIT0 = 16'h5666;
    defparam phase_register_545_add_4_14.INIT1 = 16'h5666;
    defparam phase_register_545_add_4_14.INJECT1_0 = "NO";
    defparam phase_register_545_add_4_14.INJECT1_1 = "NO";
    CCU2D phase_register_545_add_4_12 (.A0(increment[10]), .B0(n233[10]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[11]), .B1(n233[11]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17471), .COUT(n17472), .S0(n133[10]), 
          .S1(n133[11]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_545_add_4_12.INIT0 = 16'h5666;
    defparam phase_register_545_add_4_12.INIT1 = 16'h5666;
    defparam phase_register_545_add_4_12.INJECT1_0 = "NO";
    defparam phase_register_545_add_4_12.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module dynamic_pll
//

module dynamic_pll (i_clk_2f_N_2250, lo_pll_out, i_ref_clk_c, pll_clk, 
            pll_rst, pll_stb, pll_we, pll_data_i, pll_addr, pll_data_o, 
            pll_ack, GND_net) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;
    output i_clk_2f_N_2250;
    output lo_pll_out;
    input i_ref_clk_c;
    input pll_clk;
    input pll_rst;
    input pll_stb;
    input pll_we;
    input [7:0]pll_data_i;
    input [4:0]pll_addr;
    output [7:0]pll_data_o;
    output pll_ack;
    input GND_net;
    
    wire i_clk_2f_N_2250 /* synthesis is_inv_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/clock_phase_shifter.v(11[21:28])
    wire lo_pll_out /* synthesis is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(157[6:16])
    wire i_ref_clk_c /* synthesis is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(23[12:21])
    
    INV i26296 (.A(lo_pll_out), .Z(i_clk_2f_N_2250));
    EHXPLLJ PLLInst_0 (.CLKI(i_ref_clk_c), .CLKFB(lo_pll_out), .PHASESEL0(GND_net), 
            .PHASESEL1(GND_net), .PHASEDIR(GND_net), .PHASESTEP(GND_net), 
            .LOADREG(GND_net), .STDBY(GND_net), .PLLWAKESYNC(GND_net), 
            .RST(GND_net), .RESETC(GND_net), .RESETD(GND_net), .RESETM(GND_net), 
            .ENCLKOP(GND_net), .ENCLKOS(GND_net), .ENCLKOS2(GND_net), 
            .ENCLKOS3(GND_net), .PLLCLK(pll_clk), .PLLRST(pll_rst), .PLLSTB(pll_stb), 
            .PLLWE(pll_we), .PLLDATI0(pll_data_i[0]), .PLLDATI1(pll_data_i[1]), 
            .PLLDATI2(pll_data_i[2]), .PLLDATI3(pll_data_i[3]), .PLLDATI4(pll_data_i[4]), 
            .PLLDATI5(pll_data_i[5]), .PLLDATI6(pll_data_i[6]), .PLLDATI7(pll_data_i[7]), 
            .PLLADDR0(pll_addr[0]), .PLLADDR1(pll_addr[1]), .PLLADDR2(pll_addr[2]), 
            .PLLADDR3(pll_addr[3]), .PLLADDR4(pll_addr[4]), .CLKOP(lo_pll_out), 
            .PLLDATO0(pll_data_o[0]), .PLLDATO1(pll_data_o[1]), .PLLDATO2(pll_data_o[2]), 
            .PLLDATO3(pll_data_o[3]), .PLLDATO4(pll_data_o[4]), .PLLDATO5(pll_data_o[5]), 
            .PLLDATO6(pll_data_o[6]), .PLLDATO7(pll_data_o[7]), .PLLACK(pll_ack)) /* synthesis FREQUENCY_PIN_CLKOP="420.000000", FREQUENCY_PIN_CLKI="12.000000", ICP_CURRENT="6", LPF_RESISTOR="8", syn_instantiated=1, LSE_LINE_FILE_ID=8, LSE_LCOL=13, LSE_RCOL=5, LSE_LLINE=164, LSE_RLINE=175 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(164[13] 175[5])
    defparam PLLInst_0.CLKI_DIV = 1;
    defparam PLLInst_0.CLKFB_DIV = 35;
    defparam PLLInst_0.CLKOP_DIV = 1;
    defparam PLLInst_0.CLKOS_DIV = 1;
    defparam PLLInst_0.CLKOS2_DIV = 1;
    defparam PLLInst_0.CLKOS3_DIV = 1;
    defparam PLLInst_0.CLKOP_ENABLE = "ENABLED";
    defparam PLLInst_0.CLKOS_ENABLE = "DISABLED";
    defparam PLLInst_0.CLKOS2_ENABLE = "DISABLED";
    defparam PLLInst_0.CLKOS3_ENABLE = "DISABLED";
    defparam PLLInst_0.VCO_BYPASS_A0 = "DISABLED";
    defparam PLLInst_0.VCO_BYPASS_B0 = "DISABLED";
    defparam PLLInst_0.VCO_BYPASS_C0 = "DISABLED";
    defparam PLLInst_0.VCO_BYPASS_D0 = "DISABLED";
    defparam PLLInst_0.CLKOP_CPHASE = 0;
    defparam PLLInst_0.CLKOS_CPHASE = 0;
    defparam PLLInst_0.CLKOS2_CPHASE = 0;
    defparam PLLInst_0.CLKOS3_CPHASE = 0;
    defparam PLLInst_0.CLKOP_FPHASE = 0;
    defparam PLLInst_0.CLKOS_FPHASE = 0;
    defparam PLLInst_0.CLKOS2_FPHASE = 0;
    defparam PLLInst_0.CLKOS3_FPHASE = 0;
    defparam PLLInst_0.FEEDBK_PATH = "CLKOP";
    defparam PLLInst_0.FRACN_ENABLE = "ENABLED";
    defparam PLLInst_0.FRACN_DIV = 2731;
    defparam PLLInst_0.CLKOP_TRIM_POL = "RISING";
    defparam PLLInst_0.CLKOP_TRIM_DELAY = 0;
    defparam PLLInst_0.CLKOS_TRIM_POL = "FALLING";
    defparam PLLInst_0.CLKOS_TRIM_DELAY = 0;
    defparam PLLInst_0.PLL_USE_WB = "ENABLED";
    defparam PLLInst_0.PREDIVIDER_MUXA1 = 0;
    defparam PLLInst_0.PREDIVIDER_MUXB1 = 0;
    defparam PLLInst_0.PREDIVIDER_MUXC1 = 0;
    defparam PLLInst_0.PREDIVIDER_MUXD1 = 0;
    defparam PLLInst_0.OUTDIVIDER_MUXA2 = "DIVA";
    defparam PLLInst_0.OUTDIVIDER_MUXB2 = "DIVB";
    defparam PLLInst_0.OUTDIVIDER_MUXC2 = "DIVC";
    defparam PLLInst_0.OUTDIVIDER_MUXD2 = "DIVD";
    defparam PLLInst_0.PLL_LOCK_MODE = 0;
    defparam PLLInst_0.STDBY_ENABLE = "DISABLED";
    defparam PLLInst_0.DPHASE_SOURCE = "DISABLED";
    defparam PLLInst_0.PLLRST_ENA = "DISABLED";
    defparam PLLInst_0.MRST_ENA = "DISABLED";
    defparam PLLInst_0.DCRST_ENA = "DISABLED";
    defparam PLLInst_0.DDRST_ENA = "DISABLED";
    defparam PLLInst_0.INTFB_WAKE = "DISABLED";
    
endmodule
