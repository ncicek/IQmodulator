// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.11.3.469
// Netlist written on Wed Jan 13 20:58:38 2021
//
// Verilog Description of module top
//

module top (i_ref_clk, i_resetb, i_wbu_uart_rx, o_wbu_uart_tx, o_baseband_i, 
            o_baseband_q, dac_clk_p, dac_clk_n, i_clk_p, i_clk_n, 
            q_clk_p, q_clk_n) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(4[8:11])
    input i_ref_clk;   // d:/documents/git_local/fm_modulator/rtl/top.v(22[12:21])
    input i_resetb;   // d:/documents/git_local/fm_modulator/rtl/top.v(22[23:31])
    input i_wbu_uart_rx;   // d:/documents/git_local/fm_modulator/rtl/top.v(24[12:25])
    output o_wbu_uart_tx;   // d:/documents/git_local/fm_modulator/rtl/top.v(25[13:26])
    output [9:0]o_baseband_i;   // d:/documents/git_local/fm_modulator/rtl/top.v(27[38:50])
    output [9:0]o_baseband_q;   // d:/documents/git_local/fm_modulator/rtl/top.v(27[52:64])
    output dac_clk_p;   // d:/documents/git_local/fm_modulator/rtl/top.v(28[49:58])
    output dac_clk_n;   // d:/documents/git_local/fm_modulator/rtl/top.v(28[60:69])
    output i_clk_p;   // d:/documents/git_local/fm_modulator/rtl/top.v(28[13:20])
    output i_clk_n;   // d:/documents/git_local/fm_modulator/rtl/top.v(28[22:29])
    output q_clk_p;   // d:/documents/git_local/fm_modulator/rtl/top.v(28[31:38])
    output q_clk_n;   // d:/documents/git_local/fm_modulator/rtl/top.v(28[40:47])
    
    wire i_ref_clk_c /* synthesis SET_AS_NETWORK=i_ref_clk_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(22[12:21])
    wire o_baseband_i_c_15 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[37:47])
    wire o_baseband_i_c_14 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[37:47])
    wire o_baseband_i_c_13 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[37:47])
    wire o_baseband_i_c_12 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[37:47])
    wire o_baseband_i_c_11 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[37:47])
    wire o_baseband_i_c_10 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[37:47])
    wire n3607 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[37:47])
    wire o_baseband_i_c_8 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[37:47])
    wire o_baseband_i_c_7 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[37:47])
    wire o_baseband_q_c_15 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[49:59])
    wire o_baseband_q_c_14 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[49:59])
    wire o_baseband_q_c_13 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[49:59])
    wire o_baseband_q_c_12 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[49:59])
    wire o_baseband_q_c_11 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[49:59])
    wire o_baseband_q_c_10 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[49:59])
    wire n3608 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[49:59])
    wire o_baseband_q_c_8 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[49:59])
    wire o_baseband_q_c_7 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[49:59])
    wire lo_pll_out /* synthesis is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(159[6:16])
    wire i_clk_2f_N_2249 /* synthesis is_inv_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/clock_phase_shifter.v(11[21:28])
    
    wire GND_net, VCC_net, i_resetb_c, i_wbu_uart_rx_c, o_wbu_uart_tx_c, 
        o_baseband_i_c_9, o_baseband_q_c_9, i_clk_p_c, q_clk_p_c, i_resetb_N_301, 
        rx_stb;
    wire [7:0]rx_data;   // d:/documents/git_local/fm_modulator/rtl/top.v(50[12:19])
    
    wire tx_busy, wb_stb, wb_we;
    wire [29:0]wb_addr;   // d:/documents/git_local/fm_modulator/rtl/top.v(67[13:20])
    wire [31:0]wb_odata;   // d:/documents/git_local/fm_modulator/rtl/top.v(68[13:21])
    
    wire wb_ack, wb_err;
    wire [31:0]wb_idata;   // d:/documents/git_local/fm_modulator/rtl/top.v(73[12:20])
    wire [29:0]bus_err_address;   // d:/documents/git_local/fm_modulator/rtl/top.v(97[12:27])
    
    wire wb_fm_ack;
    wire [31:0]wb_fm_data;   // d:/documents/git_local/fm_modulator/rtl/top.v(101[13:23])
    wire [31:0]wb_smpl_data;   // d:/documents/git_local/fm_modulator/rtl/top.v(104[12:24])
    
    wire wb_smpl_ack;
    wire [23:0]chg_counter;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(97[17:28])
    wire [7:0]wb_lo_data;   // d:/documents/git_local/fm_modulator/rtl/top.v(137[12:22])
    
    wire wb_lo_ack, pll_clk, pll_rst, pll_stb, pll_we, pll_ack;
    wire [7:0]pll_data_i;   // d:/documents/git_local/fm_modulator/rtl/top.v(143[12:22])
    wire [7:0]pll_data_o;   // d:/documents/git_local/fm_modulator/rtl/top.v(143[24:34])
    wire [4:0]pll_addr;   // d:/documents/git_local/fm_modulator/rtl/top.v(144[12:20])
    wire [31:0]smpl_register;   // d:/documents/git_local/fm_modulator/rtl/top.v(197[13:26])
    wire [31:0]power_counter;   // d:/documents/git_local/fm_modulator/rtl/top.v(197[28:41])
    
    wire smpl_interrupt, none_sel, wb_fm_data_31__N_63, wb_lo_data_7__N_96;
    wire [31:0]wb_smpl_data_31__N_64;
    wire [31:0]power_counter_31__N_232;
    wire [30:0]power_counter_31__N_201;
    wire [31:0]power_counter_31__N_129;
    wire [31:0]wb_idata_31__N_266;
    wire [31:0]wb_idata_31__N_1;
    
    wire chg_counter_23__N_406, n19615, n19739, n19731;
    wire [3:0]state_adj_3110;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(83[12:17])
    wire [7:0]lcl_data;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(84[12:20])
    
    wire zero_baud_counter, o_busy_N_536;
    wire [7:0]lcl_data_7__N_511;
    
    wire zero_baud_counter_N_526, zero_baud_counter_N_525, i_clk_n_c, 
        q_clk_n_c, i_ref_clk_c_enable_278, n19695, n19691, n19689, 
        n19456, n25134, n19685, n2139, n2138, n2137, n2136, n24789, 
        n2134, n2133, n2132, n24790, n24791, n2129, n2128, n2127, 
        n2126, n2125, n24792, n24793, n24794, n2121, n24795, n2119, 
        n2118, n2117, n2116, n2115, n2114, n2113, n2112, n2110, 
        n2109, i_ref_clk_c_enable_180, n2, n19627, n19625, n9456, 
        n17288, n17568, n17268, n17287, n17269, n17286, n17274, 
        n17285, n17282, n17272, n17284, n17281, n17267, n17280, 
        n17297, n17279, n17296, n17278, n17295, n17277, n17294, 
        n17276, n17293, n12729, n24992, n17283, n17275, n17292, 
        n4, n17273, n17291, n24890, n17271, n38, n36, n34, n24788, 
        i_ref_clk_c_enable_98, n32, n11785, n30, i_ref_clk_c_enable_193, 
        i_ref_clk_c_enable_66, i_ref_clk_c_enable_106, n26, n25, n17290, 
        n22, n27585, i_ref_clk_c_enable_329, n17270, n2_adj_3058, 
        n1, n2_adj_3059, n1_adj_3060, n2_adj_3061, n2_adj_3062, n1_adj_3063, 
        n2_adj_3064, n1_adj_3065, n2_adj_3066, n1_adj_3067, n2_adj_3068, 
        n1_adj_3069, n2_adj_3070, n1_adj_3071, n2_adj_3072, n1_adj_3073, 
        n2_adj_3074, n1_adj_3075, n2_adj_3076, n1_adj_3077, n2_adj_3078, 
        n24809, n2_adj_3079, n1_adj_3080, n2_adj_3081, n25213, n24808, 
        n17289, n2_adj_3082, n2_adj_3083, n24806, n2_adj_3084, n1_adj_3085, 
        n2_adj_3086, n1_adj_3087, n2_adj_3088, n1_adj_3089, n2_adj_3090, 
        n1_adj_3091, n2_adj_3092, n1_adj_3093, n2_adj_3094, n2_adj_3095, 
        n2_adj_3096, n1_adj_3097, n2_adj_3098, n1_adj_3099, n2_adj_3100, 
        n1_adj_3101, n2_adj_3102, n24803, n27530, n2_adj_3103, n1_adj_3104, 
        n2_adj_3105, n1_adj_3106, n2_adj_3107, n1_adj_3108, n27529;
    
    VHI i2 (.Z(VCC_net));
    GSR GSR_INST (.GSR(i_resetb_N_301)) /* synthesis syn_instantiated=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(38[5:28])
    FD1S3AX wb_smpl_data_i0 (.D(wb_smpl_data_31__N_64[0]), .CK(i_ref_clk_c), 
            .Q(wb_smpl_data[0]));   // d:/documents/git_local/fm_modulator/rtl/top.v(214[9] 222[10])
    defparam wb_smpl_data_i0.GSR = "DISABLED";
    hbbus genbus (.i_ref_clk_c(i_ref_clk_c), .wb_odata({wb_odata}), .n27585(n27585), 
          .wb_addr({wb_addr}), .wb_we(wb_we), .wb_stb(wb_stb), .n27530(n27530), 
          .GND_net(GND_net), .wb_err(wb_err), .wb_ack(wb_ack), .\wb_idata[0] (wb_idata[0]), 
          .\wb_idata[2] (wb_idata[2]), .\wb_idata[3] (wb_idata[3]), .\wb_idata[4] (wb_idata[4]), 
          .\wb_idata[5] (wb_idata[5]), .\wb_idata[6] (wb_idata[6]), .\wb_idata[7] (wb_idata[7]), 
          .\wb_idata[8] (wb_idata[8]), .\wb_idata[9] (wb_idata[9]), .\wb_idata[10] (wb_idata[10]), 
          .\wb_idata[11] (wb_idata[11]), .\wb_idata[12] (wb_idata[12]), 
          .\wb_idata[13] (wb_idata[13]), .\wb_idata[14] (wb_idata[14]), 
          .\wb_idata[15] (wb_idata[15]), .\wb_idata[16] (wb_idata[16]), 
          .\wb_idata[17] (wb_idata[17]), .\wb_idata[18] (wb_idata[18]), 
          .\wb_idata[19] (wb_idata[19]), .\wb_idata[20] (wb_idata[20]), 
          .\wb_idata[21] (wb_idata[21]), .\wb_idata[22] (wb_idata[22]), 
          .\wb_idata[23] (wb_idata[23]), .\wb_idata[24] (wb_idata[24]), 
          .\wb_idata[25] (wb_idata[25]), .\wb_idata[26] (wb_idata[26]), 
          .\wb_idata[27] (wb_idata[27]), .\wb_idata[28] (wb_idata[28]), 
          .\wb_idata[29] (wb_idata[29]), .\wb_idata[30] (wb_idata[30]), 
          .\wb_idata[31] (wb_idata[31]), .n2(n2), .n12729(n12729), .VCC_net(VCC_net), 
          .\rx_data[6] (rx_data[6]), .\rx_data[0] (rx_data[0]), .\rx_data[5] (rx_data[5]), 
          .\rx_data[1] (rx_data[1]), .\rx_data[2] (rx_data[2]), .rx_stb(rx_stb), 
          .\rx_data[3] (rx_data[3]), .\rx_data[4] (rx_data[4]), .tx_busy(tx_busy), 
          .n24992(n24992), .\lcl_data[1] (lcl_data[1]), .\lcl_data_7__N_511[0] (lcl_data_7__N_511[0]), 
          .\lcl_data[2] (lcl_data[2]), .\lcl_data_7__N_511[1] (lcl_data_7__N_511[1]), 
          .\lcl_data[3] (lcl_data[3]), .\lcl_data_7__N_511[2] (lcl_data_7__N_511[2]), 
          .\lcl_data[4] (lcl_data[4]), .\lcl_data_7__N_511[3] (lcl_data_7__N_511[3]), 
          .\lcl_data[5] (lcl_data[5]), .\lcl_data_7__N_511[4] (lcl_data_7__N_511[4]), 
          .\lcl_data[6] (lcl_data[6]), .\lcl_data_7__N_511[5] (lcl_data_7__N_511[5]), 
          .\lcl_data[7] (lcl_data[7]), .\lcl_data_7__N_511[6] (lcl_data_7__N_511[6]), 
          .n24890(n24890), .zero_baud_counter_N_526(zero_baud_counter_N_526), 
          .zero_baud_counter_N_525(zero_baud_counter_N_525), .zero_baud_counter(zero_baud_counter), 
          .i_ref_clk_c_enable_329(i_ref_clk_c_enable_329), .o_busy_N_536(o_busy_N_536), 
          .\state[0] (state_adj_3110[0]), .n17568(n17568)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(76[7] 92[22])
    FD1S3AX power_counter_i0 (.D(power_counter_31__N_129[0]), .CK(i_ref_clk_c), 
            .Q(power_counter[0])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(226[9] 231[54])
    defparam power_counter_i0.GSR = "DISABLED";
    FD1S3AX wb_idata_i0 (.D(wb_idata_31__N_1[0]), .CK(i_ref_clk_c), .Q(wb_idata[0]));   // d:/documents/git_local/fm_modulator/rtl/top.v(267[9] 275[22])
    defparam wb_idata_i0.GSR = "DISABLED";
    FD1S3JX wb_ack_70 (.D(n4), .CK(i_ref_clk_c), .PD(wb_smpl_ack), .Q(wb_ack)) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(264[9] 265[57])
    defparam wb_ack_70.GSR = "DISABLED";
    PUR PUR_INST (.PUR(i_resetb_N_301)) /* synthesis syn_instantiated=1 */ ;
    defparam PUR_INST.RST_PULSE = 1;
    FD1S3IX wb_smpl_ack_63 (.D(wb_stb), .CK(i_ref_clk_c), .CD(n24809), 
            .Q(wb_smpl_ack)) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(200[9] 201[44])
    defparam wb_smpl_ack_63.GSR = "DISABLED";
    fm_generator_wb_slave wb_fm_data_31__I_0 (.i_ref_clk_c(i_ref_clk_c), .i_ref_clk_c_enable_106(i_ref_clk_c_enable_106), 
            .i_resetb_N_301(i_resetb_N_301), .wb_odata({wb_odata}), .i_ref_clk_c_enable_66(i_ref_clk_c_enable_66), 
            .i_ref_clk_c_enable_98(i_ref_clk_c_enable_98), .wb_fm_data({wb_fm_data}), 
            .wb_fm_ack(wb_fm_ack), .wb_fm_data_31__N_63(wb_fm_data_31__N_63), 
            .GND_net(GND_net), .\wb_addr[1] (wb_addr[1]), .\wb_addr[0] (wb_addr[0]), 
            .\power_counter[1] (power_counter[1]), .\smpl_register[1] (smpl_register[1]), 
            .n2139(n2139), .i_resetb_c(i_resetb_c), .n24803(n24803), .n2(n2_adj_3102), 
            .\smpl_register[5] (smpl_register[5]), .n24788(n24788), .n2_adj_1(n2_adj_3061), 
            .\smpl_register[29] (smpl_register[29]), .n24795(n24795), .n2_adj_2(n2_adj_3078), 
            .\smpl_register[20] (smpl_register[20]), .n24794(n24794), .n2_adj_3(n2_adj_3081), 
            .\smpl_register[18] (smpl_register[18]), .n24793(n24793), .n2_adj_4(n2_adj_3082), 
            .\smpl_register[17] (smpl_register[17]), .n24792(n24792), .n2_adj_5(n2_adj_3083), 
            .\smpl_register[16] (smpl_register[16]), .n24791(n24791), .n2_adj_6(n2_adj_3094), 
            .\smpl_register[10] (smpl_register[10]), .n24790(n24790), .n2_adj_7(n2_adj_3095), 
            .\smpl_register[9] (smpl_register[9]), .n24789(n24789), .o_baseband_i_c_15(o_baseband_i_c_15), 
            .o_baseband_i_c_14(o_baseband_i_c_14), .o_baseband_i_c_13(o_baseband_i_c_13), 
            .o_baseband_i_c_12(o_baseband_i_c_12), .o_baseband_i_c_11(o_baseband_i_c_11), 
            .o_baseband_i_c_10(o_baseband_i_c_10), .n3607(n3607), .o_baseband_q_c_7(o_baseband_q_c_7), 
            .o_baseband_i_c_7(o_baseband_i_c_7), .o_baseband_i_c_8(o_baseband_i_c_8), 
            .n27529(n27529), .o_baseband_q_c_15(o_baseband_q_c_15), .o_baseband_q_c_14(o_baseband_q_c_14), 
            .o_baseband_q_c_13(o_baseband_q_c_13), .o_baseband_q_c_12(o_baseband_q_c_12), 
            .o_baseband_q_c_11(o_baseband_q_c_11), .o_baseband_q_c_10(o_baseband_q_c_10), 
            .n3608(n3608), .o_baseband_q_c_8(o_baseband_q_c_8)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(123[2] 134[2])
    FD1P3AX smpl_register_i0_i0 (.D(wb_odata[0]), .SP(i_ref_clk_c_enable_278), 
            .CK(i_ref_clk_c), .Q(smpl_register[0]));   // d:/documents/git_local/fm_modulator/rtl/top.v(204[9] 212[6])
    defparam smpl_register_i0_i0.GSR = "DISABLED";
    FD1S3IX wb_err_68 (.D(none_sel), .CK(i_ref_clk_c), .CD(n2), .Q(wb_err));   // d:/documents/git_local/fm_modulator/rtl/top.v(253[9] 254[34])
    defparam wb_err_68.GSR = "DISABLED";
    OB o_baseband_i_pad_7 (.I(o_baseband_i_c_14), .O(o_baseband_i[7]));   // d:/documents/git_local/fm_modulator/rtl/top.v(27[38:50])
    OB o_baseband_i_pad_8 (.I(o_baseband_i_c_15), .O(o_baseband_i[8]));   // d:/documents/git_local/fm_modulator/rtl/top.v(27[38:50])
    OB o_baseband_i_pad_9 (.I(o_baseband_i_c_9), .O(o_baseband_i[9]));   // d:/documents/git_local/fm_modulator/rtl/top.v(27[38:50])
    OB o_wbu_uart_tx_pad (.I(o_wbu_uart_tx_c), .O(o_wbu_uart_tx));   // d:/documents/git_local/fm_modulator/rtl/top.v(25[13:26])
    FD1P3AX bus_err_address_i0_i0 (.D(wb_addr[0]), .SP(wb_err), .CK(i_ref_clk_c), 
            .Q(bus_err_address[0])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(257[9] 259[31])
    defparam bus_err_address_i0_i0.GSR = "DISABLED";
    CCU2D add_35_31 (.A0(power_counter[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17297), .S0(power_counter_31__N_201[29]), 
          .S1(power_counter_31__N_201[30]));   // d:/documents/git_local/fm_modulator/rtl/top.v(231[27:53])
    defparam add_35_31.INIT0 = 16'h5aaa;
    defparam add_35_31.INIT1 = 16'h5aaa;
    defparam add_35_31.INJECT1_0 = "NO";
    defparam add_35_31.INJECT1_1 = "NO";
    CCU2D add_35_29 (.A0(power_counter[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17296), .COUT(n17297), .S0(power_counter_31__N_201[27]), 
          .S1(power_counter_31__N_201[28]));   // d:/documents/git_local/fm_modulator/rtl/top.v(231[27:53])
    defparam add_35_29.INIT0 = 16'h5aaa;
    defparam add_35_29.INIT1 = 16'h5aaa;
    defparam add_35_29.INJECT1_0 = "NO";
    defparam add_35_29.INJECT1_1 = "NO";
    CCU2D add_34_25 (.A0(power_counter[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17278), .COUT(n17279), .S0(power_counter_31__N_232[23]), 
          .S1(power_counter_31__N_232[24]));   // d:/documents/git_local/fm_modulator/rtl/top.v(229[21:41])
    defparam add_34_25.INIT0 = 16'h5aaa;
    defparam add_34_25.INIT1 = 16'h5aaa;
    defparam add_34_25.INJECT1_0 = "NO";
    defparam add_34_25.INJECT1_1 = "NO";
    FD1P3AX smpl_interrupt_65 (.D(wb_odata[0]), .SP(i_ref_clk_c_enable_193), 
            .CK(i_ref_clk_c), .Q(smpl_interrupt)) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(204[9] 212[6])
    defparam smpl_interrupt_65.GSR = "DISABLED";
    CCU2D add_35_27 (.A0(power_counter[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17295), .COUT(n17296), .S0(power_counter_31__N_201[25]), 
          .S1(power_counter_31__N_201[26]));   // d:/documents/git_local/fm_modulator/rtl/top.v(231[27:53])
    defparam add_35_27.INIT0 = 16'h5aaa;
    defparam add_35_27.INIT1 = 16'h5aaa;
    defparam add_35_27.INJECT1_0 = "NO";
    defparam add_35_27.INJECT1_1 = "NO";
    CCU2D add_34_23 (.A0(power_counter[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17277), .COUT(n17278), .S0(power_counter_31__N_232[21]), 
          .S1(power_counter_31__N_232[22]));   // d:/documents/git_local/fm_modulator/rtl/top.v(229[21:41])
    defparam add_34_23.INIT0 = 16'h5aaa;
    defparam add_34_23.INIT1 = 16'h5aaa;
    defparam add_34_23.INJECT1_0 = "NO";
    defparam add_34_23.INJECT1_1 = "NO";
    CCU2D add_35_25 (.A0(power_counter[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17294), .COUT(n17295), .S0(power_counter_31__N_201[23]), 
          .S1(power_counter_31__N_201[24]));   // d:/documents/git_local/fm_modulator/rtl/top.v(231[27:53])
    defparam add_35_25.INIT0 = 16'h5aaa;
    defparam add_35_25.INIT1 = 16'h5aaa;
    defparam add_35_25.INJECT1_0 = "NO";
    defparam add_35_25.INJECT1_1 = "NO";
    CCU2D add_34_21 (.A0(power_counter[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17276), .COUT(n17277), .S0(power_counter_31__N_232[19]), 
          .S1(power_counter_31__N_232[20]));   // d:/documents/git_local/fm_modulator/rtl/top.v(229[21:41])
    defparam add_34_21.INIT0 = 16'h5aaa;
    defparam add_34_21.INIT1 = 16'h5aaa;
    defparam add_34_21.INJECT1_0 = "NO";
    defparam add_34_21.INJECT1_1 = "NO";
    CCU2D add_35_23 (.A0(power_counter[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17293), .COUT(n17294), .S0(power_counter_31__N_201[21]), 
          .S1(power_counter_31__N_201[22]));   // d:/documents/git_local/fm_modulator/rtl/top.v(231[27:53])
    defparam add_35_23.INIT0 = 16'h5aaa;
    defparam add_35_23.INIT1 = 16'h5aaa;
    defparam add_35_23.INJECT1_0 = "NO";
    defparam add_35_23.INJECT1_1 = "NO";
    LUT4 o_clk_q_I_0_1_lut (.A(q_clk_p_c), .Z(q_clk_n_c)) /* synthesis lut_function=(!(A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/clock_phase_shifter.v(18[16:24])
    defparam o_clk_q_I_0_1_lut.init = 16'h5555;
    LUT4 o_clk_i_I_0_1_lut (.A(i_clk_p_c), .Z(i_clk_n_c)) /* synthesis lut_function=(!(A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/clock_phase_shifter.v(14[16:24])
    defparam o_clk_i_I_0_1_lut.init = 16'h5555;
    FD1P3AX smpl_register_i0_i31 (.D(wb_odata[31]), .SP(i_ref_clk_c_enable_278), 
            .CK(i_ref_clk_c), .Q(smpl_register[31]));   // d:/documents/git_local/fm_modulator/rtl/top.v(204[9] 212[6])
    defparam smpl_register_i0_i31.GSR = "DISABLED";
    LUT4 i3_4_lut (.A(wb_addr[1]), .B(wb_addr[0]), .C(n24806), .D(n9456), 
         .Z(i_ref_clk_c_enable_278)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i3_4_lut.init = 16'h0040;
    LUT4 equal_371_i3_2_lut (.A(wb_addr[2]), .B(wb_addr[3]), .Z(n9456)) /* synthesis lut_function=(A+(B)) */ ;
    defparam equal_371_i3_2_lut.init = 16'heeee;
    FD1P3AX smpl_register_i0_i30 (.D(wb_odata[30]), .SP(i_ref_clk_c_enable_278), 
            .CK(i_ref_clk_c), .Q(smpl_register[30]));   // d:/documents/git_local/fm_modulator/rtl/top.v(204[9] 212[6])
    defparam smpl_register_i0_i30.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i29 (.D(wb_odata[29]), .SP(i_ref_clk_c_enable_278), 
            .CK(i_ref_clk_c), .Q(smpl_register[29]));   // d:/documents/git_local/fm_modulator/rtl/top.v(204[9] 212[6])
    defparam smpl_register_i0_i29.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i28 (.D(wb_odata[28]), .SP(i_ref_clk_c_enable_278), 
            .CK(i_ref_clk_c), .Q(smpl_register[28]));   // d:/documents/git_local/fm_modulator/rtl/top.v(204[9] 212[6])
    defparam smpl_register_i0_i28.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i27 (.D(wb_odata[27]), .SP(i_ref_clk_c_enable_278), 
            .CK(i_ref_clk_c), .Q(smpl_register[27]));   // d:/documents/git_local/fm_modulator/rtl/top.v(204[9] 212[6])
    defparam smpl_register_i0_i27.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i26 (.D(wb_odata[26]), .SP(i_ref_clk_c_enable_278), 
            .CK(i_ref_clk_c), .Q(smpl_register[26]));   // d:/documents/git_local/fm_modulator/rtl/top.v(204[9] 212[6])
    defparam smpl_register_i0_i26.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i25 (.D(wb_odata[25]), .SP(i_ref_clk_c_enable_278), 
            .CK(i_ref_clk_c), .Q(smpl_register[25]));   // d:/documents/git_local/fm_modulator/rtl/top.v(204[9] 212[6])
    defparam smpl_register_i0_i25.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i24 (.D(wb_odata[24]), .SP(i_ref_clk_c_enable_278), 
            .CK(i_ref_clk_c), .Q(smpl_register[24]));   // d:/documents/git_local/fm_modulator/rtl/top.v(204[9] 212[6])
    defparam smpl_register_i0_i24.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i23 (.D(wb_odata[23]), .SP(i_ref_clk_c_enable_278), 
            .CK(i_ref_clk_c), .Q(smpl_register[23]));   // d:/documents/git_local/fm_modulator/rtl/top.v(204[9] 212[6])
    defparam smpl_register_i0_i23.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i22 (.D(wb_odata[22]), .SP(i_ref_clk_c_enable_278), 
            .CK(i_ref_clk_c), .Q(smpl_register[22]));   // d:/documents/git_local/fm_modulator/rtl/top.v(204[9] 212[6])
    defparam smpl_register_i0_i22.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i21 (.D(wb_odata[21]), .SP(i_ref_clk_c_enable_278), 
            .CK(i_ref_clk_c), .Q(smpl_register[21]));   // d:/documents/git_local/fm_modulator/rtl/top.v(204[9] 212[6])
    defparam smpl_register_i0_i21.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i20 (.D(wb_odata[20]), .SP(i_ref_clk_c_enable_278), 
            .CK(i_ref_clk_c), .Q(smpl_register[20]));   // d:/documents/git_local/fm_modulator/rtl/top.v(204[9] 212[6])
    defparam smpl_register_i0_i20.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i19 (.D(wb_odata[19]), .SP(i_ref_clk_c_enable_278), 
            .CK(i_ref_clk_c), .Q(smpl_register[19]));   // d:/documents/git_local/fm_modulator/rtl/top.v(204[9] 212[6])
    defparam smpl_register_i0_i19.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i18 (.D(wb_odata[18]), .SP(i_ref_clk_c_enable_278), 
            .CK(i_ref_clk_c), .Q(smpl_register[18]));   // d:/documents/git_local/fm_modulator/rtl/top.v(204[9] 212[6])
    defparam smpl_register_i0_i18.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i17 (.D(wb_odata[17]), .SP(i_ref_clk_c_enable_278), 
            .CK(i_ref_clk_c), .Q(smpl_register[17]));   // d:/documents/git_local/fm_modulator/rtl/top.v(204[9] 212[6])
    defparam smpl_register_i0_i17.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i16 (.D(wb_odata[16]), .SP(i_ref_clk_c_enable_278), 
            .CK(i_ref_clk_c), .Q(smpl_register[16]));   // d:/documents/git_local/fm_modulator/rtl/top.v(204[9] 212[6])
    defparam smpl_register_i0_i16.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i15 (.D(wb_odata[15]), .SP(i_ref_clk_c_enable_278), 
            .CK(i_ref_clk_c), .Q(smpl_register[15]));   // d:/documents/git_local/fm_modulator/rtl/top.v(204[9] 212[6])
    defparam smpl_register_i0_i15.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i14 (.D(wb_odata[14]), .SP(i_ref_clk_c_enable_278), 
            .CK(i_ref_clk_c), .Q(smpl_register[14]));   // d:/documents/git_local/fm_modulator/rtl/top.v(204[9] 212[6])
    defparam smpl_register_i0_i14.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i13 (.D(wb_odata[13]), .SP(i_ref_clk_c_enable_278), 
            .CK(i_ref_clk_c), .Q(smpl_register[13]));   // d:/documents/git_local/fm_modulator/rtl/top.v(204[9] 212[6])
    defparam smpl_register_i0_i13.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i12 (.D(wb_odata[12]), .SP(i_ref_clk_c_enable_278), 
            .CK(i_ref_clk_c), .Q(smpl_register[12]));   // d:/documents/git_local/fm_modulator/rtl/top.v(204[9] 212[6])
    defparam smpl_register_i0_i12.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i11 (.D(wb_odata[11]), .SP(i_ref_clk_c_enable_278), 
            .CK(i_ref_clk_c), .Q(smpl_register[11]));   // d:/documents/git_local/fm_modulator/rtl/top.v(204[9] 212[6])
    defparam smpl_register_i0_i11.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i10 (.D(wb_odata[10]), .SP(i_ref_clk_c_enable_278), 
            .CK(i_ref_clk_c), .Q(smpl_register[10]));   // d:/documents/git_local/fm_modulator/rtl/top.v(204[9] 212[6])
    defparam smpl_register_i0_i10.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i9 (.D(wb_odata[9]), .SP(i_ref_clk_c_enable_278), 
            .CK(i_ref_clk_c), .Q(smpl_register[9]));   // d:/documents/git_local/fm_modulator/rtl/top.v(204[9] 212[6])
    defparam smpl_register_i0_i9.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i8 (.D(wb_odata[8]), .SP(i_ref_clk_c_enable_278), 
            .CK(i_ref_clk_c), .Q(smpl_register[8]));   // d:/documents/git_local/fm_modulator/rtl/top.v(204[9] 212[6])
    defparam smpl_register_i0_i8.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i7 (.D(wb_odata[7]), .SP(i_ref_clk_c_enable_278), 
            .CK(i_ref_clk_c), .Q(smpl_register[7]));   // d:/documents/git_local/fm_modulator/rtl/top.v(204[9] 212[6])
    defparam smpl_register_i0_i7.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i6 (.D(wb_odata[6]), .SP(i_ref_clk_c_enable_278), 
            .CK(i_ref_clk_c), .Q(smpl_register[6]));   // d:/documents/git_local/fm_modulator/rtl/top.v(204[9] 212[6])
    defparam smpl_register_i0_i6.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i5 (.D(wb_odata[5]), .SP(i_ref_clk_c_enable_278), 
            .CK(i_ref_clk_c), .Q(smpl_register[5]));   // d:/documents/git_local/fm_modulator/rtl/top.v(204[9] 212[6])
    defparam smpl_register_i0_i5.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i4 (.D(wb_odata[4]), .SP(i_ref_clk_c_enable_278), 
            .CK(i_ref_clk_c), .Q(smpl_register[4]));   // d:/documents/git_local/fm_modulator/rtl/top.v(204[9] 212[6])
    defparam smpl_register_i0_i4.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i3 (.D(wb_odata[3]), .SP(i_ref_clk_c_enable_278), 
            .CK(i_ref_clk_c), .Q(smpl_register[3]));   // d:/documents/git_local/fm_modulator/rtl/top.v(204[9] 212[6])
    defparam smpl_register_i0_i3.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i2 (.D(wb_odata[2]), .SP(i_ref_clk_c_enable_278), 
            .CK(i_ref_clk_c), .Q(smpl_register[2]));   // d:/documents/git_local/fm_modulator/rtl/top.v(204[9] 212[6])
    defparam smpl_register_i0_i2.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i1 (.D(wb_odata[1]), .SP(i_ref_clk_c_enable_278), 
            .CK(i_ref_clk_c), .Q(smpl_register[1]));   // d:/documents/git_local/fm_modulator/rtl/top.v(204[9] 212[6])
    defparam smpl_register_i0_i1.GSR = "DISABLED";
    CCU2D add_34_19 (.A0(power_counter[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17275), .COUT(n17276), .S0(power_counter_31__N_232[17]), 
          .S1(power_counter_31__N_232[18]));   // d:/documents/git_local/fm_modulator/rtl/top.v(229[21:41])
    defparam add_34_19.INIT0 = 16'h5aaa;
    defparam add_34_19.INIT1 = 16'h5aaa;
    defparam add_34_19.INJECT1_0 = "NO";
    defparam add_34_19.INJECT1_1 = "NO";
    LUT4 i1_4_lut (.A(chg_counter_23__N_406), .B(n19689), .C(n19739), 
         .D(n19685), .Z(i_ref_clk_c_enable_180)) /* synthesis lut_function=(A+!(B (C (D)))) */ ;
    defparam i1_4_lut.init = 16'hbfff;
    LUT4 i17378_4_lut (.A(chg_counter[18]), .B(chg_counter[23]), .C(chg_counter[3]), 
         .D(chg_counter[16]), .Z(n19689)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i17378_4_lut.init = 16'h8000;
    LUT4 i17427_4_lut (.A(n19627), .B(n19731), .C(n19695), .D(n19625), 
         .Z(n19739)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i17427_4_lut.init = 16'h8000;
    LUT4 i17374_4_lut (.A(chg_counter[19]), .B(chg_counter[13]), .C(chg_counter[2]), 
         .D(chg_counter[14]), .Z(n19685)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i17374_4_lut.init = 16'h8000;
    LUT4 i17326_2_lut (.A(chg_counter[10]), .B(chg_counter[0]), .Z(n19627)) /* synthesis lut_function=(A (B)) */ ;
    defparam i17326_2_lut.init = 16'h8888;
    LUT4 i17419_4_lut (.A(chg_counter[12]), .B(n19691), .C(n19615), .D(chg_counter[11]), 
         .Z(n19731)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i17419_4_lut.init = 16'h8000;
    LUT4 i17384_4_lut (.A(chg_counter[8]), .B(chg_counter[1]), .C(chg_counter[9]), 
         .D(chg_counter[6]), .Z(n19695)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i17384_4_lut.init = 16'h8000;
    LUT4 i17324_2_lut (.A(chg_counter[20]), .B(chg_counter[5]), .Z(n19625)) /* synthesis lut_function=(A (B)) */ ;
    defparam i17324_2_lut.init = 16'h8888;
    LUT4 i17380_4_lut (.A(chg_counter[21]), .B(chg_counter[7]), .C(chg_counter[4]), 
         .D(chg_counter[15]), .Z(n19691)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i17380_4_lut.init = 16'h8000;
    LUT4 i17314_2_lut (.A(chg_counter[17]), .B(chg_counter[22]), .Z(n19615)) /* synthesis lut_function=(A (B)) */ ;
    defparam i17314_2_lut.init = 16'h8888;
    LUT4 i2_3_lut_4_lut (.A(wb_addr[9]), .B(n11785), .C(wb_addr[8]), .D(n27585), 
         .Z(wb_lo_data_7__N_96)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[21:47])
    defparam i2_3_lut_4_lut.init = 16'h2000;
    LUT4 i17398_3_lut (.A(n11785), .B(wb_addr[8]), .C(wb_addr[9]), .Z(none_sel)) /* synthesis lut_function=(A+!(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(249[20:68])
    defparam i17398_3_lut.init = 16'habab;
    LUT4 i_resetb_I_0_1_lut (.A(i_resetb_c), .Z(i_resetb_N_301)) /* synthesis lut_function=(!(A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(36[16:25])
    defparam i_resetb_I_0_1_lut.init = 16'h5555;
    LUT4 mux_373_i1_4_lut (.A(smpl_interrupt), .B(wb_addr[0]), .C(n25134), 
         .D(n19456), .Z(wb_smpl_data_31__N_64[0])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(215[3] 222[10])
    defparam mux_373_i1_4_lut.init = 16'hca0a;
    LUT4 i1_4_lut_adj_106 (.A(smpl_register[0]), .B(n9456), .C(power_counter[0]), 
         .D(wb_addr[1]), .Z(n19456)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(215[3] 222[10])
    defparam i1_4_lut_adj_106.init = 16'h3022;
    LUT4 i1_2_lut_rep_248_3_lut (.A(wb_addr[9]), .B(n11785), .C(wb_addr[8]), 
         .Z(n24808)) /* synthesis lut_function=((B+(C))+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[21:47])
    defparam i1_2_lut_rep_248_3_lut.init = 16'hfdfd;
    LUT4 wb_stb_I_0_72_2_lut_3_lut_4_lut (.A(wb_addr[9]), .B(n11785), .C(wb_stb), 
         .D(wb_addr[8]), .Z(wb_fm_data_31__N_63)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[21:47])
    defparam wb_stb_I_0_72_2_lut_3_lut_4_lut.init = 16'h0020;
    LUT4 i1_2_lut_rep_243_3_lut_4_lut (.A(wb_addr[9]), .B(n11785), .C(n25213), 
         .D(wb_addr[8]), .Z(n24803)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[21:47])
    defparam i1_2_lut_rep_243_3_lut_4_lut.init = 16'h0020;
    LUT4 power_counter_31__I_0_77_i1_3_lut (.A(power_counter_31__N_232[0]), 
         .B(power_counter_31__N_201[0]), .C(power_counter[31]), .Z(power_counter_31__N_129[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(231[4:54])
    defparam power_counter_31__I_0_77_i1_3_lut.init = 16'hcaca;
    LUT4 i719_1_lut (.A(o_baseband_i_c_15), .Z(o_baseband_i_c_9)) /* synthesis lut_function=(!(A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(112[31:66])
    defparam i719_1_lut.init = 16'h5555;
    LUT4 wb_idata_31__I_0_i1_3_lut (.A(wb_idata_31__N_266[0]), .B(wb_fm_data[0]), 
         .C(wb_fm_ack), .Z(wb_idata_31__N_1[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[8] 275[22])
    defparam wb_idata_31__I_0_i1_3_lut.init = 16'hcaca;
    LUT4 mux_59_i1_4_lut (.A(wb_lo_data[0]), .B(wb_smpl_data[0]), .C(wb_smpl_ack), 
         .D(wb_lo_ack), .Z(wb_idata_31__N_266[0])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(272[8] 275[22])
    defparam mux_59_i1_4_lut.init = 16'hcac0;
    LUT4 i1_2_lut (.A(wb_fm_ack), .B(wb_lo_ack), .Z(n4)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(265[13:56])
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i19_4_lut (.A(n25), .B(n38), .C(n34), .D(n26), .Z(n11785)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[21:47])
    defparam i19_4_lut.init = 16'hfffe;
    LUT4 i5_2_lut (.A(wb_addr[12]), .B(wb_addr[15]), .Z(n25)) /* synthesis lut_function=(A+!(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[21:47])
    defparam i5_2_lut.init = 16'hbbbb;
    LUT4 i18_4_lut (.A(wb_addr[20]), .B(n36), .C(n30), .D(wb_addr[21]), 
         .Z(n38)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[21:47])
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i14_4_lut (.A(wb_addr[13]), .B(wb_addr[29]), .C(wb_addr[19]), 
         .D(wb_addr[28]), .Z(n34)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[21:47])
    defparam i14_4_lut.init = 16'hfffe;
    LUT4 i6_2_lut (.A(wb_addr[22]), .B(wb_addr[24]), .Z(n26)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[21:47])
    defparam i6_2_lut.init = 16'heeee;
    LUT4 i16_4_lut (.A(wb_addr[14]), .B(n32), .C(n22), .D(wb_addr[26]), 
         .Z(n36)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[21:47])
    defparam i16_4_lut.init = 16'hfffe;
    LUT4 i10_2_lut (.A(wb_addr[10]), .B(wb_addr[16]), .Z(n30)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[21:47])
    defparam i10_2_lut.init = 16'heeee;
    LUT4 i12_4_lut (.A(wb_addr[11]), .B(wb_addr[18]), .C(wb_addr[27]), 
         .D(wb_addr[23]), .Z(n32)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[21:47])
    defparam i12_4_lut.init = 16'hfffe;
    LUT4 i2_2_lut (.A(wb_addr[17]), .B(wb_addr[25]), .Z(n22)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[21:47])
    defparam i2_2_lut.init = 16'heeee;
    LUT4 mux_374_Mux_31_i2_3_lut (.A(bus_err_address[29]), .B(power_counter[31]), 
         .C(wb_addr[0]), .Z(n2_adj_3058)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(215[3] 222[10])
    defparam mux_374_Mux_31_i2_3_lut.init = 16'hcaca;
    LUT4 i11097_2_lut (.A(smpl_register[31]), .B(wb_addr[0]), .Z(n1)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(215[3] 222[10])
    defparam i11097_2_lut.init = 16'h8888;
    LUT4 mux_374_Mux_30_i2_3_lut (.A(bus_err_address[28]), .B(power_counter[30]), 
         .C(wb_addr[0]), .Z(n2_adj_3059)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(215[3] 222[10])
    defparam mux_374_Mux_30_i2_3_lut.init = 16'hcaca;
    LUT4 i11096_2_lut (.A(smpl_register[30]), .B(wb_addr[0]), .Z(n1_adj_3060)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(215[3] 222[10])
    defparam i11096_2_lut.init = 16'h8888;
    LUT4 mux_374_Mux_29_i2_3_lut (.A(bus_err_address[27]), .B(power_counter[29]), 
         .C(wb_addr[0]), .Z(n2_adj_3061)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(215[3] 222[10])
    defparam mux_374_Mux_29_i2_3_lut.init = 16'hcaca;
    LUT4 wb_idata_31__I_0_i32_4_lut (.A(wb_smpl_data[31]), .B(wb_fm_data[31]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_1[31])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[8] 275[22])
    defparam wb_idata_31__I_0_i32_4_lut.init = 16'hcac0;
    LUT4 mux_374_Mux_28_i2_3_lut (.A(bus_err_address[26]), .B(power_counter[28]), 
         .C(wb_addr[0]), .Z(n2_adj_3062)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(215[3] 222[10])
    defparam mux_374_Mux_28_i2_3_lut.init = 16'hcaca;
    LUT4 i11094_2_lut (.A(smpl_register[28]), .B(wb_addr[0]), .Z(n1_adj_3063)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(215[3] 222[10])
    defparam i11094_2_lut.init = 16'h8888;
    LUT4 mux_374_Mux_27_i2_3_lut (.A(bus_err_address[25]), .B(power_counter[27]), 
         .C(wb_addr[0]), .Z(n2_adj_3064)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(215[3] 222[10])
    defparam mux_374_Mux_27_i2_3_lut.init = 16'hcaca;
    LUT4 i11093_2_lut (.A(smpl_register[27]), .B(wb_addr[0]), .Z(n1_adj_3065)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(215[3] 222[10])
    defparam i11093_2_lut.init = 16'h8888;
    LUT4 mux_374_Mux_26_i2_3_lut (.A(bus_err_address[24]), .B(power_counter[26]), 
         .C(wb_addr[0]), .Z(n2_adj_3066)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(215[3] 222[10])
    defparam mux_374_Mux_26_i2_3_lut.init = 16'hcaca;
    LUT4 i11092_2_lut (.A(smpl_register[26]), .B(wb_addr[0]), .Z(n1_adj_3067)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(215[3] 222[10])
    defparam i11092_2_lut.init = 16'h8888;
    LUT4 mux_374_Mux_25_i2_3_lut (.A(bus_err_address[23]), .B(power_counter[25]), 
         .C(wb_addr[0]), .Z(n2_adj_3068)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(215[3] 222[10])
    defparam mux_374_Mux_25_i2_3_lut.init = 16'hcaca;
    LUT4 i11091_2_lut (.A(smpl_register[25]), .B(wb_addr[0]), .Z(n1_adj_3069)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(215[3] 222[10])
    defparam i11091_2_lut.init = 16'h8888;
    LUT4 mux_374_Mux_24_i2_3_lut (.A(bus_err_address[22]), .B(power_counter[24]), 
         .C(wb_addr[0]), .Z(n2_adj_3070)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(215[3] 222[10])
    defparam mux_374_Mux_24_i2_3_lut.init = 16'hcaca;
    LUT4 i11090_2_lut (.A(smpl_register[24]), .B(wb_addr[0]), .Z(n1_adj_3071)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(215[3] 222[10])
    defparam i11090_2_lut.init = 16'h8888;
    LUT4 mux_374_Mux_23_i2_3_lut (.A(bus_err_address[21]), .B(power_counter[23]), 
         .C(wb_addr[0]), .Z(n2_adj_3072)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(215[3] 222[10])
    defparam mux_374_Mux_23_i2_3_lut.init = 16'hcaca;
    LUT4 i11089_2_lut (.A(smpl_register[23]), .B(wb_addr[0]), .Z(n1_adj_3073)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(215[3] 222[10])
    defparam i11089_2_lut.init = 16'h8888;
    LUT4 mux_374_Mux_22_i2_3_lut (.A(bus_err_address[20]), .B(power_counter[22]), 
         .C(wb_addr[0]), .Z(n2_adj_3074)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(215[3] 222[10])
    defparam mux_374_Mux_22_i2_3_lut.init = 16'hcaca;
    LUT4 i11088_2_lut (.A(smpl_register[22]), .B(wb_addr[0]), .Z(n1_adj_3075)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(215[3] 222[10])
    defparam i11088_2_lut.init = 16'h8888;
    LUT4 mux_374_Mux_21_i2_3_lut (.A(bus_err_address[19]), .B(power_counter[21]), 
         .C(wb_addr[0]), .Z(n2_adj_3076)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(215[3] 222[10])
    defparam mux_374_Mux_21_i2_3_lut.init = 16'hcaca;
    LUT4 i11087_2_lut (.A(smpl_register[21]), .B(wb_addr[0]), .Z(n1_adj_3077)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(215[3] 222[10])
    defparam i11087_2_lut.init = 16'h8888;
    LUT4 mux_374_Mux_20_i2_3_lut (.A(bus_err_address[18]), .B(power_counter[20]), 
         .C(wb_addr[0]), .Z(n2_adj_3078)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(215[3] 222[10])
    defparam mux_374_Mux_20_i2_3_lut.init = 16'hcaca;
    LUT4 mux_374_Mux_19_i2_3_lut (.A(bus_err_address[17]), .B(power_counter[19]), 
         .C(wb_addr[0]), .Z(n2_adj_3079)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(215[3] 222[10])
    defparam mux_374_Mux_19_i2_3_lut.init = 16'hcaca;
    LUT4 i11085_2_lut (.A(smpl_register[19]), .B(wb_addr[0]), .Z(n1_adj_3080)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(215[3] 222[10])
    defparam i11085_2_lut.init = 16'h8888;
    LUT4 mux_374_Mux_18_i2_3_lut (.A(bus_err_address[16]), .B(power_counter[18]), 
         .C(wb_addr[0]), .Z(n2_adj_3081)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(215[3] 222[10])
    defparam mux_374_Mux_18_i2_3_lut.init = 16'hcaca;
    LUT4 i21100_2_lut_3_lut_4_lut (.A(n24808), .B(n25213), .C(wb_addr[0]), 
         .D(wb_addr[1]), .Z(i_ref_clk_c_enable_106)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(125[39:58])
    defparam i21100_2_lut_3_lut_4_lut.init = 16'h0004;
    LUT4 mux_374_Mux_17_i2_3_lut (.A(bus_err_address[15]), .B(power_counter[17]), 
         .C(wb_addr[0]), .Z(n2_adj_3082)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(215[3] 222[10])
    defparam mux_374_Mux_17_i2_3_lut.init = 16'hcaca;
    LUT4 i21096_2_lut_3_lut_4_lut (.A(n24808), .B(n25213), .C(wb_addr[0]), 
         .D(wb_addr[1]), .Z(i_ref_clk_c_enable_66)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(125[39:58])
    defparam i21096_2_lut_3_lut_4_lut.init = 16'h0040;
    LUT4 mux_374_Mux_16_i2_3_lut (.A(bus_err_address[14]), .B(power_counter[16]), 
         .C(wb_addr[0]), .Z(n2_adj_3083)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(215[3] 222[10])
    defparam mux_374_Mux_16_i2_3_lut.init = 16'hcaca;
    LUT4 mux_374_Mux_15_i2_3_lut (.A(bus_err_address[13]), .B(power_counter[15]), 
         .C(wb_addr[0]), .Z(n2_adj_3084)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(215[3] 222[10])
    defparam mux_374_Mux_15_i2_3_lut.init = 16'hcaca;
    LUT4 i11081_2_lut (.A(smpl_register[15]), .B(wb_addr[0]), .Z(n1_adj_3085)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(215[3] 222[10])
    defparam i11081_2_lut.init = 16'h8888;
    LUT4 mux_374_Mux_14_i2_3_lut (.A(bus_err_address[12]), .B(power_counter[14]), 
         .C(wb_addr[0]), .Z(n2_adj_3086)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(215[3] 222[10])
    defparam mux_374_Mux_14_i2_3_lut.init = 16'hcaca;
    LUT4 i11080_2_lut (.A(smpl_register[14]), .B(wb_addr[0]), .Z(n1_adj_3087)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(215[3] 222[10])
    defparam i11080_2_lut.init = 16'h8888;
    LUT4 mux_374_Mux_13_i2_3_lut (.A(bus_err_address[11]), .B(power_counter[13]), 
         .C(wb_addr[0]), .Z(n2_adj_3088)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(215[3] 222[10])
    defparam mux_374_Mux_13_i2_3_lut.init = 16'hcaca;
    LUT4 i11079_2_lut (.A(smpl_register[13]), .B(wb_addr[0]), .Z(n1_adj_3089)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(215[3] 222[10])
    defparam i11079_2_lut.init = 16'h8888;
    LUT4 mux_374_Mux_12_i2_3_lut (.A(bus_err_address[10]), .B(power_counter[12]), 
         .C(wb_addr[0]), .Z(n2_adj_3090)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(215[3] 222[10])
    defparam mux_374_Mux_12_i2_3_lut.init = 16'hcaca;
    LUT4 i11078_2_lut (.A(smpl_register[12]), .B(wb_addr[0]), .Z(n1_adj_3091)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(215[3] 222[10])
    defparam i11078_2_lut.init = 16'h8888;
    LUT4 mux_374_Mux_11_i2_3_lut (.A(bus_err_address[9]), .B(power_counter[11]), 
         .C(wb_addr[0]), .Z(n2_adj_3092)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(215[3] 222[10])
    defparam mux_374_Mux_11_i2_3_lut.init = 16'hcaca;
    LUT4 i11077_2_lut (.A(smpl_register[11]), .B(wb_addr[0]), .Z(n1_adj_3093)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(215[3] 222[10])
    defparam i11077_2_lut.init = 16'h8888;
    LUT4 mux_374_Mux_10_i2_3_lut (.A(bus_err_address[8]), .B(power_counter[10]), 
         .C(wb_addr[0]), .Z(n2_adj_3094)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(215[3] 222[10])
    defparam mux_374_Mux_10_i2_3_lut.init = 16'hcaca;
    LUT4 i21094_3_lut_4_lut (.A(n24808), .B(n25213), .C(wb_addr[0]), .D(wb_addr[1]), 
         .Z(i_ref_clk_c_enable_98)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(125[39:58])
    defparam i21094_3_lut_4_lut.init = 16'h0400;
    LUT4 mux_374_Mux_9_i2_3_lut (.A(bus_err_address[7]), .B(power_counter[9]), 
         .C(wb_addr[0]), .Z(n2_adj_3095)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(215[3] 222[10])
    defparam mux_374_Mux_9_i2_3_lut.init = 16'hcaca;
    LUT4 mux_374_Mux_8_i2_3_lut (.A(bus_err_address[6]), .B(power_counter[8]), 
         .C(wb_addr[0]), .Z(n2_adj_3096)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(215[3] 222[10])
    defparam mux_374_Mux_8_i2_3_lut.init = 16'hcaca;
    LUT4 i11074_2_lut (.A(smpl_register[8]), .B(wb_addr[0]), .Z(n1_adj_3097)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(215[3] 222[10])
    defparam i11074_2_lut.init = 16'h8888;
    LUT4 mux_374_Mux_7_i2_3_lut (.A(bus_err_address[5]), .B(power_counter[7]), 
         .C(wb_addr[0]), .Z(n2_adj_3098)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(215[3] 222[10])
    defparam mux_374_Mux_7_i2_3_lut.init = 16'hcaca;
    LUT4 i11073_2_lut (.A(smpl_register[7]), .B(wb_addr[0]), .Z(n1_adj_3099)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(215[3] 222[10])
    defparam i11073_2_lut.init = 16'h8888;
    LUT4 mux_374_Mux_6_i2_3_lut (.A(bus_err_address[4]), .B(power_counter[6]), 
         .C(wb_addr[0]), .Z(n2_adj_3100)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(215[3] 222[10])
    defparam mux_374_Mux_6_i2_3_lut.init = 16'hcaca;
    LUT4 i11072_2_lut (.A(smpl_register[6]), .B(wb_addr[0]), .Z(n1_adj_3101)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(215[3] 222[10])
    defparam i11072_2_lut.init = 16'h8888;
    LUT4 mux_374_Mux_5_i2_3_lut (.A(bus_err_address[3]), .B(power_counter[5]), 
         .C(wb_addr[0]), .Z(n2_adj_3102)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(215[3] 222[10])
    defparam mux_374_Mux_5_i2_3_lut.init = 16'hcaca;
    LUT4 mux_374_Mux_4_i2_3_lut (.A(bus_err_address[2]), .B(power_counter[4]), 
         .C(wb_addr[0]), .Z(n2_adj_3103)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(215[3] 222[10])
    defparam mux_374_Mux_4_i2_3_lut.init = 16'hcaca;
    LUT4 i11070_2_lut (.A(smpl_register[4]), .B(wb_addr[0]), .Z(n1_adj_3104)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(215[3] 222[10])
    defparam i11070_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_rep_653 (.A(wb_stb), .B(wb_we), .Z(n25213)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(205[7:30])
    defparam i1_2_lut_rep_653.init = 16'h8888;
    LUT4 i21063_2_lut_3_lut_3_lut_4_lut (.A(wb_stb), .B(wb_we), .C(n24809), 
         .D(n25134), .Z(i_ref_clk_c_enable_193)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(205[7:30])
    defparam i21063_2_lut_3_lut_3_lut_4_lut.init = 16'h0008;
    LUT4 mux_374_Mux_3_i2_3_lut (.A(bus_err_address[1]), .B(power_counter[3]), 
         .C(wb_addr[0]), .Z(n2_adj_3105)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(215[3] 222[10])
    defparam mux_374_Mux_3_i2_3_lut.init = 16'hcaca;
    LUT4 i11069_2_lut (.A(smpl_register[3]), .B(wb_addr[0]), .Z(n1_adj_3106)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(215[3] 222[10])
    defparam i11069_2_lut.init = 16'h8888;
    LUT4 mux_374_Mux_2_i2_3_lut (.A(bus_err_address[0]), .B(power_counter[2]), 
         .C(wb_addr[0]), .Z(n2_adj_3107)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(215[3] 222[10])
    defparam mux_374_Mux_2_i2_3_lut.init = 16'hcaca;
    LUT4 i11068_2_lut (.A(smpl_register[2]), .B(wb_addr[0]), .Z(n1_adj_3108)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(215[3] 222[10])
    defparam i11068_2_lut.init = 16'h8888;
    LUT4 i2_3_lut_rep_249 (.A(n11785), .B(wb_addr[9]), .C(wb_addr[8]), 
         .Z(n24809)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(243[23:49])
    defparam i2_3_lut_rep_249.init = 16'hefef;
    LUT4 i1_2_lut_rep_246_4_lut (.A(n11785), .B(wb_addr[9]), .C(wb_addr[8]), 
         .D(n25213), .Z(n24806)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(243[23:49])
    defparam i1_2_lut_rep_246_4_lut.init = 16'h1000;
    PFUMX mux_374_Mux_2_i3 (.BLUT(n1_adj_3108), .ALUT(n2_adj_3107), .C0(wb_addr[1]), 
          .Z(n2138));
    PFUMX mux_374_Mux_3_i3 (.BLUT(n1_adj_3106), .ALUT(n2_adj_3105), .C0(wb_addr[1]), 
          .Z(n2137));
    PFUMX mux_374_Mux_4_i3 (.BLUT(n1_adj_3104), .ALUT(n2_adj_3103), .C0(wb_addr[1]), 
          .Z(n2136));
    PFUMX mux_374_Mux_6_i3 (.BLUT(n1_adj_3101), .ALUT(n2_adj_3100), .C0(wb_addr[1]), 
          .Z(n2134));
    PFUMX mux_374_Mux_7_i3 (.BLUT(n1_adj_3099), .ALUT(n2_adj_3098), .C0(wb_addr[1]), 
          .Z(n2133));
    PFUMX mux_374_Mux_8_i3 (.BLUT(n1_adj_3097), .ALUT(n2_adj_3096), .C0(wb_addr[1]), 
          .Z(n2132));
    PFUMX mux_374_Mux_11_i3 (.BLUT(n1_adj_3093), .ALUT(n2_adj_3092), .C0(wb_addr[1]), 
          .Z(n2129));
    PFUMX mux_374_Mux_12_i3 (.BLUT(n1_adj_3091), .ALUT(n2_adj_3090), .C0(wb_addr[1]), 
          .Z(n2128));
    PFUMX mux_374_Mux_13_i3 (.BLUT(n1_adj_3089), .ALUT(n2_adj_3088), .C0(wb_addr[1]), 
          .Z(n2127));
    PFUMX mux_374_Mux_14_i3 (.BLUT(n1_adj_3087), .ALUT(n2_adj_3086), .C0(wb_addr[1]), 
          .Z(n2126));
    PFUMX mux_374_Mux_15_i3 (.BLUT(n1_adj_3085), .ALUT(n2_adj_3084), .C0(wb_addr[1]), 
          .Z(n2125));
    PFUMX mux_374_Mux_19_i3 (.BLUT(n1_adj_3080), .ALUT(n2_adj_3079), .C0(wb_addr[1]), 
          .Z(n2121));
    PFUMX mux_374_Mux_21_i3 (.BLUT(n1_adj_3077), .ALUT(n2_adj_3076), .C0(wb_addr[1]), 
          .Z(n2119));
    PFUMX mux_374_Mux_22_i3 (.BLUT(n1_adj_3075), .ALUT(n2_adj_3074), .C0(wb_addr[1]), 
          .Z(n2118));
    PFUMX mux_374_Mux_23_i3 (.BLUT(n1_adj_3073), .ALUT(n2_adj_3072), .C0(wb_addr[1]), 
          .Z(n2117));
    PFUMX mux_374_Mux_24_i3 (.BLUT(n1_adj_3071), .ALUT(n2_adj_3070), .C0(wb_addr[1]), 
          .Z(n2116));
    PFUMX mux_374_Mux_25_i3 (.BLUT(n1_adj_3069), .ALUT(n2_adj_3068), .C0(wb_addr[1]), 
          .Z(n2115));
    PFUMX mux_374_Mux_26_i3 (.BLUT(n1_adj_3067), .ALUT(n2_adj_3066), .C0(wb_addr[1]), 
          .Z(n2114));
    PFUMX mux_374_Mux_27_i3 (.BLUT(n1_adj_3065), .ALUT(n2_adj_3064), .C0(wb_addr[1]), 
          .Z(n2113));
    PFUMX mux_374_Mux_28_i3 (.BLUT(n1_adj_3063), .ALUT(n2_adj_3062), .C0(wb_addr[1]), 
          .Z(n2112));
    PFUMX mux_374_Mux_30_i3 (.BLUT(n1_adj_3060), .ALUT(n2_adj_3059), .C0(wb_addr[1]), 
          .Z(n2110));
    PFUMX mux_374_Mux_31_i3 (.BLUT(n1), .ALUT(n2_adj_3058), .C0(wb_addr[1]), 
          .Z(n2109));
    FD1S3AX wb_idata_i31 (.D(wb_idata_31__N_1[31]), .CK(i_ref_clk_c), .Q(wb_idata[31]));   // d:/documents/git_local/fm_modulator/rtl/top.v(267[9] 275[22])
    defparam wb_idata_i31.GSR = "DISABLED";
    LUT4 wb_idata_31__I_0_i31_4_lut (.A(wb_smpl_data[30]), .B(wb_fm_data[30]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_1[30])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[8] 275[22])
    defparam wb_idata_31__I_0_i31_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i30_4_lut (.A(wb_smpl_data[29]), .B(wb_fm_data[29]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_1[29])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[8] 275[22])
    defparam wb_idata_31__I_0_i30_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i29_4_lut (.A(wb_smpl_data[28]), .B(wb_fm_data[28]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_1[28])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[8] 275[22])
    defparam wb_idata_31__I_0_i29_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i28_4_lut (.A(wb_smpl_data[27]), .B(wb_fm_data[27]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_1[27])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[8] 275[22])
    defparam wb_idata_31__I_0_i28_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i27_4_lut (.A(wb_smpl_data[26]), .B(wb_fm_data[26]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_1[26])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[8] 275[22])
    defparam wb_idata_31__I_0_i27_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i26_4_lut (.A(wb_smpl_data[25]), .B(wb_fm_data[25]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_1[25])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[8] 275[22])
    defparam wb_idata_31__I_0_i26_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i25_4_lut (.A(wb_smpl_data[24]), .B(wb_fm_data[24]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_1[24])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[8] 275[22])
    defparam wb_idata_31__I_0_i25_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i24_4_lut (.A(wb_smpl_data[23]), .B(wb_fm_data[23]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_1[23])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[8] 275[22])
    defparam wb_idata_31__I_0_i24_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i23_4_lut (.A(wb_smpl_data[22]), .B(wb_fm_data[22]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_1[22])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[8] 275[22])
    defparam wb_idata_31__I_0_i23_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i22_4_lut (.A(wb_smpl_data[21]), .B(wb_fm_data[21]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_1[21])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[8] 275[22])
    defparam wb_idata_31__I_0_i22_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i21_4_lut (.A(wb_smpl_data[20]), .B(wb_fm_data[20]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_1[20])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[8] 275[22])
    defparam wb_idata_31__I_0_i21_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i20_4_lut (.A(wb_smpl_data[19]), .B(wb_fm_data[19]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_1[19])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[8] 275[22])
    defparam wb_idata_31__I_0_i20_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i19_4_lut (.A(wb_smpl_data[18]), .B(wb_fm_data[18]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_1[18])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[8] 275[22])
    defparam wb_idata_31__I_0_i19_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i18_4_lut (.A(wb_smpl_data[17]), .B(wb_fm_data[17]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_1[17])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[8] 275[22])
    defparam wb_idata_31__I_0_i18_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i17_4_lut (.A(wb_smpl_data[16]), .B(wb_fm_data[16]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_1[16])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[8] 275[22])
    defparam wb_idata_31__I_0_i17_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i16_4_lut (.A(wb_smpl_data[15]), .B(wb_fm_data[15]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_1[15])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[8] 275[22])
    defparam wb_idata_31__I_0_i16_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i15_4_lut (.A(wb_smpl_data[14]), .B(wb_fm_data[14]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_1[14])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[8] 275[22])
    defparam wb_idata_31__I_0_i15_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i14_4_lut (.A(wb_smpl_data[13]), .B(wb_fm_data[13]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_1[13])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[8] 275[22])
    defparam wb_idata_31__I_0_i14_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i13_4_lut (.A(wb_smpl_data[12]), .B(wb_fm_data[12]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_1[12])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[8] 275[22])
    defparam wb_idata_31__I_0_i13_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i12_4_lut (.A(wb_smpl_data[11]), .B(wb_fm_data[11]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_1[11])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[8] 275[22])
    defparam wb_idata_31__I_0_i12_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i11_4_lut (.A(wb_smpl_data[10]), .B(wb_fm_data[10]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_1[10])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[8] 275[22])
    defparam wb_idata_31__I_0_i11_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i10_4_lut (.A(wb_smpl_data[9]), .B(wb_fm_data[9]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_1[9])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[8] 275[22])
    defparam wb_idata_31__I_0_i10_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i9_4_lut (.A(wb_smpl_data[8]), .B(wb_fm_data[8]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_1[8])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[8] 275[22])
    defparam wb_idata_31__I_0_i9_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i8_3_lut (.A(wb_idata_31__N_266[7]), .B(wb_fm_data[7]), 
         .C(wb_fm_ack), .Z(wb_idata_31__N_1[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[8] 275[22])
    defparam wb_idata_31__I_0_i8_3_lut.init = 16'hcaca;
    LUT4 mux_59_i8_4_lut (.A(wb_lo_data[7]), .B(wb_smpl_data[7]), .C(wb_smpl_ack), 
         .D(wb_lo_ack), .Z(wb_idata_31__N_266[7])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(272[8] 275[22])
    defparam mux_59_i8_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i7_3_lut (.A(wb_idata_31__N_266[6]), .B(wb_fm_data[6]), 
         .C(wb_fm_ack), .Z(wb_idata_31__N_1[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[8] 275[22])
    defparam wb_idata_31__I_0_i7_3_lut.init = 16'hcaca;
    LUT4 mux_59_i7_4_lut (.A(wb_lo_data[6]), .B(wb_smpl_data[6]), .C(wb_smpl_ack), 
         .D(wb_lo_ack), .Z(wb_idata_31__N_266[6])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(272[8] 275[22])
    defparam mux_59_i7_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i6_3_lut (.A(wb_idata_31__N_266[5]), .B(wb_fm_data[5]), 
         .C(wb_fm_ack), .Z(wb_idata_31__N_1[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[8] 275[22])
    defparam wb_idata_31__I_0_i6_3_lut.init = 16'hcaca;
    LUT4 mux_59_i6_4_lut (.A(wb_lo_data[5]), .B(wb_smpl_data[5]), .C(wb_smpl_ack), 
         .D(wb_lo_ack), .Z(wb_idata_31__N_266[5])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(272[8] 275[22])
    defparam mux_59_i6_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i5_3_lut (.A(wb_idata_31__N_266[4]), .B(wb_fm_data[4]), 
         .C(wb_fm_ack), .Z(wb_idata_31__N_1[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[8] 275[22])
    defparam wb_idata_31__I_0_i5_3_lut.init = 16'hcaca;
    LUT4 mux_59_i5_4_lut (.A(wb_lo_data[4]), .B(wb_smpl_data[4]), .C(wb_smpl_ack), 
         .D(wb_lo_ack), .Z(wb_idata_31__N_266[4])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(272[8] 275[22])
    defparam mux_59_i5_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i4_3_lut (.A(wb_idata_31__N_266[3]), .B(wb_fm_data[3]), 
         .C(wb_fm_ack), .Z(wb_idata_31__N_1[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[8] 275[22])
    defparam wb_idata_31__I_0_i4_3_lut.init = 16'hcaca;
    LUT4 mux_59_i4_4_lut (.A(wb_lo_data[3]), .B(wb_smpl_data[3]), .C(wb_smpl_ack), 
         .D(wb_lo_ack), .Z(wb_idata_31__N_266[3])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(272[8] 275[22])
    defparam mux_59_i4_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i3_3_lut (.A(wb_idata_31__N_266[2]), .B(wb_fm_data[2]), 
         .C(wb_fm_ack), .Z(wb_idata_31__N_1[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[8] 275[22])
    defparam wb_idata_31__I_0_i3_3_lut.init = 16'hcaca;
    LUT4 mux_59_i3_4_lut (.A(wb_lo_data[2]), .B(wb_smpl_data[2]), .C(wb_smpl_ack), 
         .D(wb_lo_ack), .Z(wb_idata_31__N_266[2])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(272[8] 275[22])
    defparam mux_59_i3_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i2_3_lut (.A(wb_idata_31__N_266[1]), .B(wb_fm_data[1]), 
         .C(wb_fm_ack), .Z(wb_idata_31__N_1[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(270[8] 275[22])
    defparam wb_idata_31__I_0_i2_3_lut.init = 16'hcaca;
    LUT4 mux_59_i2_4_lut (.A(wb_lo_data[1]), .B(wb_smpl_data[1]), .C(wb_smpl_ack), 
         .D(wb_lo_ack), .Z(wb_idata_31__N_266[1])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(272[8] 275[22])
    defparam mux_59_i2_4_lut.init = 16'hcac0;
    LUT4 i10086_1_lut (.A(wb_idata[1]), .Z(n12729)) /* synthesis lut_function=(!(A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(267[9] 275[22])
    defparam i10086_1_lut.init = 16'h5555;
    FD1S3AX wb_idata_i30 (.D(wb_idata_31__N_1[30]), .CK(i_ref_clk_c), .Q(wb_idata[30]));   // d:/documents/git_local/fm_modulator/rtl/top.v(267[9] 275[22])
    defparam wb_idata_i30.GSR = "DISABLED";
    FD1S3AX wb_idata_i29 (.D(wb_idata_31__N_1[29]), .CK(i_ref_clk_c), .Q(wb_idata[29]));   // d:/documents/git_local/fm_modulator/rtl/top.v(267[9] 275[22])
    defparam wb_idata_i29.GSR = "DISABLED";
    FD1S3AX wb_idata_i28 (.D(wb_idata_31__N_1[28]), .CK(i_ref_clk_c), .Q(wb_idata[28]));   // d:/documents/git_local/fm_modulator/rtl/top.v(267[9] 275[22])
    defparam wb_idata_i28.GSR = "DISABLED";
    FD1S3AX wb_idata_i27 (.D(wb_idata_31__N_1[27]), .CK(i_ref_clk_c), .Q(wb_idata[27]));   // d:/documents/git_local/fm_modulator/rtl/top.v(267[9] 275[22])
    defparam wb_idata_i27.GSR = "DISABLED";
    FD1S3AX wb_idata_i26 (.D(wb_idata_31__N_1[26]), .CK(i_ref_clk_c), .Q(wb_idata[26]));   // d:/documents/git_local/fm_modulator/rtl/top.v(267[9] 275[22])
    defparam wb_idata_i26.GSR = "DISABLED";
    FD1S3AX wb_idata_i25 (.D(wb_idata_31__N_1[25]), .CK(i_ref_clk_c), .Q(wb_idata[25]));   // d:/documents/git_local/fm_modulator/rtl/top.v(267[9] 275[22])
    defparam wb_idata_i25.GSR = "DISABLED";
    FD1S3AX wb_idata_i24 (.D(wb_idata_31__N_1[24]), .CK(i_ref_clk_c), .Q(wb_idata[24]));   // d:/documents/git_local/fm_modulator/rtl/top.v(267[9] 275[22])
    defparam wb_idata_i24.GSR = "DISABLED";
    FD1S3AX wb_idata_i23 (.D(wb_idata_31__N_1[23]), .CK(i_ref_clk_c), .Q(wb_idata[23]));   // d:/documents/git_local/fm_modulator/rtl/top.v(267[9] 275[22])
    defparam wb_idata_i23.GSR = "DISABLED";
    FD1S3AX wb_idata_i22 (.D(wb_idata_31__N_1[22]), .CK(i_ref_clk_c), .Q(wb_idata[22]));   // d:/documents/git_local/fm_modulator/rtl/top.v(267[9] 275[22])
    defparam wb_idata_i22.GSR = "DISABLED";
    FD1S3AX wb_idata_i21 (.D(wb_idata_31__N_1[21]), .CK(i_ref_clk_c), .Q(wb_idata[21]));   // d:/documents/git_local/fm_modulator/rtl/top.v(267[9] 275[22])
    defparam wb_idata_i21.GSR = "DISABLED";
    FD1S3AX wb_idata_i20 (.D(wb_idata_31__N_1[20]), .CK(i_ref_clk_c), .Q(wb_idata[20]));   // d:/documents/git_local/fm_modulator/rtl/top.v(267[9] 275[22])
    defparam wb_idata_i20.GSR = "DISABLED";
    FD1S3AX wb_idata_i19 (.D(wb_idata_31__N_1[19]), .CK(i_ref_clk_c), .Q(wb_idata[19]));   // d:/documents/git_local/fm_modulator/rtl/top.v(267[9] 275[22])
    defparam wb_idata_i19.GSR = "DISABLED";
    LUT4 power_counter_31__I_0_77_i31_3_lut (.A(power_counter_31__N_232[30]), 
         .B(power_counter_31__N_201[30]), .C(power_counter[31]), .Z(power_counter_31__N_129[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(231[4:54])
    defparam power_counter_31__I_0_77_i31_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_77_i30_3_lut (.A(power_counter_31__N_232[29]), 
         .B(power_counter_31__N_201[29]), .C(power_counter[31]), .Z(power_counter_31__N_129[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(231[4:54])
    defparam power_counter_31__I_0_77_i30_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_77_i29_3_lut (.A(power_counter_31__N_232[28]), 
         .B(power_counter_31__N_201[28]), .C(power_counter[31]), .Z(power_counter_31__N_129[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(231[4:54])
    defparam power_counter_31__I_0_77_i29_3_lut.init = 16'hcaca;
    FD1S3AX wb_idata_i18 (.D(wb_idata_31__N_1[18]), .CK(i_ref_clk_c), .Q(wb_idata[18]));   // d:/documents/git_local/fm_modulator/rtl/top.v(267[9] 275[22])
    defparam wb_idata_i18.GSR = "DISABLED";
    LUT4 power_counter_31__I_0_77_i28_3_lut (.A(power_counter_31__N_232[27]), 
         .B(power_counter_31__N_201[27]), .C(power_counter[31]), .Z(power_counter_31__N_129[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(231[4:54])
    defparam power_counter_31__I_0_77_i28_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_77_i27_3_lut (.A(power_counter_31__N_232[26]), 
         .B(power_counter_31__N_201[26]), .C(power_counter[31]), .Z(power_counter_31__N_129[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(231[4:54])
    defparam power_counter_31__I_0_77_i27_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_77_i26_3_lut (.A(power_counter_31__N_232[25]), 
         .B(power_counter_31__N_201[25]), .C(power_counter[31]), .Z(power_counter_31__N_129[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(231[4:54])
    defparam power_counter_31__I_0_77_i26_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_77_i25_3_lut (.A(power_counter_31__N_232[24]), 
         .B(power_counter_31__N_201[24]), .C(power_counter[31]), .Z(power_counter_31__N_129[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(231[4:54])
    defparam power_counter_31__I_0_77_i25_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_77_i24_3_lut (.A(power_counter_31__N_232[23]), 
         .B(power_counter_31__N_201[23]), .C(power_counter[31]), .Z(power_counter_31__N_129[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(231[4:54])
    defparam power_counter_31__I_0_77_i24_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_77_i23_3_lut (.A(power_counter_31__N_232[22]), 
         .B(power_counter_31__N_201[22]), .C(power_counter[31]), .Z(power_counter_31__N_129[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(231[4:54])
    defparam power_counter_31__I_0_77_i23_3_lut.init = 16'hcaca;
    FD1S3AX wb_idata_i17 (.D(wb_idata_31__N_1[17]), .CK(i_ref_clk_c), .Q(wb_idata[17]));   // d:/documents/git_local/fm_modulator/rtl/top.v(267[9] 275[22])
    defparam wb_idata_i17.GSR = "DISABLED";
    LUT4 power_counter_31__I_0_77_i22_3_lut (.A(power_counter_31__N_232[21]), 
         .B(power_counter_31__N_201[21]), .C(power_counter[31]), .Z(power_counter_31__N_129[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(231[4:54])
    defparam power_counter_31__I_0_77_i22_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_77_i21_3_lut (.A(power_counter_31__N_232[20]), 
         .B(power_counter_31__N_201[20]), .C(power_counter[31]), .Z(power_counter_31__N_129[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(231[4:54])
    defparam power_counter_31__I_0_77_i21_3_lut.init = 16'hcaca;
    FD1S3AX wb_idata_i16 (.D(wb_idata_31__N_1[16]), .CK(i_ref_clk_c), .Q(wb_idata[16]));   // d:/documents/git_local/fm_modulator/rtl/top.v(267[9] 275[22])
    defparam wb_idata_i16.GSR = "DISABLED";
    FD1S3AX wb_idata_i15 (.D(wb_idata_31__N_1[15]), .CK(i_ref_clk_c), .Q(wb_idata[15]));   // d:/documents/git_local/fm_modulator/rtl/top.v(267[9] 275[22])
    defparam wb_idata_i15.GSR = "DISABLED";
    LUT4 power_counter_31__I_0_77_i20_3_lut (.A(power_counter_31__N_232[19]), 
         .B(power_counter_31__N_201[19]), .C(power_counter[31]), .Z(power_counter_31__N_129[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(231[4:54])
    defparam power_counter_31__I_0_77_i20_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_77_i19_3_lut (.A(power_counter_31__N_232[18]), 
         .B(power_counter_31__N_201[18]), .C(power_counter[31]), .Z(power_counter_31__N_129[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(231[4:54])
    defparam power_counter_31__I_0_77_i19_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_77_i18_3_lut (.A(power_counter_31__N_232[17]), 
         .B(power_counter_31__N_201[17]), .C(power_counter[31]), .Z(power_counter_31__N_129[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(231[4:54])
    defparam power_counter_31__I_0_77_i18_3_lut.init = 16'hcaca;
    FD1S3AX wb_idata_i14 (.D(wb_idata_31__N_1[14]), .CK(i_ref_clk_c), .Q(wb_idata[14]));   // d:/documents/git_local/fm_modulator/rtl/top.v(267[9] 275[22])
    defparam wb_idata_i14.GSR = "DISABLED";
    FD1S3AX wb_idata_i13 (.D(wb_idata_31__N_1[13]), .CK(i_ref_clk_c), .Q(wb_idata[13]));   // d:/documents/git_local/fm_modulator/rtl/top.v(267[9] 275[22])
    defparam wb_idata_i13.GSR = "DISABLED";
    LUT4 power_counter_31__I_0_77_i17_3_lut (.A(power_counter_31__N_232[16]), 
         .B(power_counter_31__N_201[16]), .C(power_counter[31]), .Z(power_counter_31__N_129[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(231[4:54])
    defparam power_counter_31__I_0_77_i17_3_lut.init = 16'hcaca;
    FD1S3AX wb_idata_i12 (.D(wb_idata_31__N_1[12]), .CK(i_ref_clk_c), .Q(wb_idata[12]));   // d:/documents/git_local/fm_modulator/rtl/top.v(267[9] 275[22])
    defparam wb_idata_i12.GSR = "DISABLED";
    LUT4 power_counter_31__I_0_77_i16_3_lut (.A(power_counter_31__N_232[15]), 
         .B(power_counter_31__N_201[15]), .C(power_counter[31]), .Z(power_counter_31__N_129[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(231[4:54])
    defparam power_counter_31__I_0_77_i16_3_lut.init = 16'hcaca;
    FD1S3AX wb_idata_i11 (.D(wb_idata_31__N_1[11]), .CK(i_ref_clk_c), .Q(wb_idata[11]));   // d:/documents/git_local/fm_modulator/rtl/top.v(267[9] 275[22])
    defparam wb_idata_i11.GSR = "DISABLED";
    FD1S3AX wb_idata_i10 (.D(wb_idata_31__N_1[10]), .CK(i_ref_clk_c), .Q(wb_idata[10]));   // d:/documents/git_local/fm_modulator/rtl/top.v(267[9] 275[22])
    defparam wb_idata_i10.GSR = "DISABLED";
    FD1S3AX wb_idata_i9 (.D(wb_idata_31__N_1[9]), .CK(i_ref_clk_c), .Q(wb_idata[9]));   // d:/documents/git_local/fm_modulator/rtl/top.v(267[9] 275[22])
    defparam wb_idata_i9.GSR = "DISABLED";
    LUT4 power_counter_31__I_0_77_i15_3_lut (.A(power_counter_31__N_232[14]), 
         .B(power_counter_31__N_201[14]), .C(power_counter[31]), .Z(power_counter_31__N_129[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(231[4:54])
    defparam power_counter_31__I_0_77_i15_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_77_i14_3_lut (.A(power_counter_31__N_232[13]), 
         .B(power_counter_31__N_201[13]), .C(power_counter[31]), .Z(power_counter_31__N_129[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(231[4:54])
    defparam power_counter_31__I_0_77_i14_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_77_i13_3_lut (.A(power_counter_31__N_232[12]), 
         .B(power_counter_31__N_201[12]), .C(power_counter[31]), .Z(power_counter_31__N_129[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(231[4:54])
    defparam power_counter_31__I_0_77_i13_3_lut.init = 16'hcaca;
    FD1S3AX wb_idata_i8 (.D(wb_idata_31__N_1[8]), .CK(i_ref_clk_c), .Q(wb_idata[8]));   // d:/documents/git_local/fm_modulator/rtl/top.v(267[9] 275[22])
    defparam wb_idata_i8.GSR = "DISABLED";
    LUT4 power_counter_31__I_0_77_i12_3_lut (.A(power_counter_31__N_232[11]), 
         .B(power_counter_31__N_201[11]), .C(power_counter[31]), .Z(power_counter_31__N_129[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(231[4:54])
    defparam power_counter_31__I_0_77_i12_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_77_i11_3_lut (.A(power_counter_31__N_232[10]), 
         .B(power_counter_31__N_201[10]), .C(power_counter[31]), .Z(power_counter_31__N_129[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(231[4:54])
    defparam power_counter_31__I_0_77_i11_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_77_i10_3_lut (.A(power_counter_31__N_232[9]), 
         .B(power_counter_31__N_201[9]), .C(power_counter[31]), .Z(power_counter_31__N_129[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(231[4:54])
    defparam power_counter_31__I_0_77_i10_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_77_i9_3_lut (.A(power_counter_31__N_232[8]), 
         .B(power_counter_31__N_201[8]), .C(power_counter[31]), .Z(power_counter_31__N_129[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(231[4:54])
    defparam power_counter_31__I_0_77_i9_3_lut.init = 16'hcaca;
    FD1S3AX wb_idata_i7 (.D(wb_idata_31__N_1[7]), .CK(i_ref_clk_c), .Q(wb_idata[7]));   // d:/documents/git_local/fm_modulator/rtl/top.v(267[9] 275[22])
    defparam wb_idata_i7.GSR = "DISABLED";
    LUT4 power_counter_31__I_0_77_i8_3_lut (.A(power_counter_31__N_232[7]), 
         .B(power_counter_31__N_201[7]), .C(power_counter[31]), .Z(power_counter_31__N_129[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(231[4:54])
    defparam power_counter_31__I_0_77_i8_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_77_i7_3_lut (.A(power_counter_31__N_232[6]), 
         .B(power_counter_31__N_201[6]), .C(power_counter[31]), .Z(power_counter_31__N_129[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(231[4:54])
    defparam power_counter_31__I_0_77_i7_3_lut.init = 16'hcaca;
    FD1S3AX wb_idata_i6 (.D(wb_idata_31__N_1[6]), .CK(i_ref_clk_c), .Q(wb_idata[6]));   // d:/documents/git_local/fm_modulator/rtl/top.v(267[9] 275[22])
    defparam wb_idata_i6.GSR = "DISABLED";
    FD1S3AX wb_idata_i5 (.D(wb_idata_31__N_1[5]), .CK(i_ref_clk_c), .Q(wb_idata[5]));   // d:/documents/git_local/fm_modulator/rtl/top.v(267[9] 275[22])
    defparam wb_idata_i5.GSR = "DISABLED";
    LUT4 power_counter_31__I_0_77_i6_3_lut (.A(power_counter_31__N_232[5]), 
         .B(power_counter_31__N_201[5]), .C(power_counter[31]), .Z(power_counter_31__N_129[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(231[4:54])
    defparam power_counter_31__I_0_77_i6_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_77_i5_3_lut (.A(power_counter_31__N_232[4]), 
         .B(power_counter_31__N_201[4]), .C(power_counter[31]), .Z(power_counter_31__N_129[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(231[4:54])
    defparam power_counter_31__I_0_77_i5_3_lut.init = 16'hcaca;
    FD1S3AX wb_idata_i4 (.D(wb_idata_31__N_1[4]), .CK(i_ref_clk_c), .Q(wb_idata[4]));   // d:/documents/git_local/fm_modulator/rtl/top.v(267[9] 275[22])
    defparam wb_idata_i4.GSR = "DISABLED";
    LUT4 power_counter_31__I_0_77_i4_3_lut (.A(power_counter_31__N_232[3]), 
         .B(power_counter_31__N_201[3]), .C(power_counter[31]), .Z(power_counter_31__N_129[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(231[4:54])
    defparam power_counter_31__I_0_77_i4_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_77_i3_3_lut (.A(power_counter_31__N_232[2]), 
         .B(power_counter_31__N_201[2]), .C(power_counter[31]), .Z(power_counter_31__N_129[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(231[4:54])
    defparam power_counter_31__I_0_77_i3_3_lut.init = 16'hcaca;
    FD1S3AX wb_idata_i3 (.D(wb_idata_31__N_1[3]), .CK(i_ref_clk_c), .Q(wb_idata[3]));   // d:/documents/git_local/fm_modulator/rtl/top.v(267[9] 275[22])
    defparam wb_idata_i3.GSR = "DISABLED";
    FD1S3AX wb_idata_i2 (.D(wb_idata_31__N_1[2]), .CK(i_ref_clk_c), .Q(wb_idata[2]));   // d:/documents/git_local/fm_modulator/rtl/top.v(267[9] 275[22])
    defparam wb_idata_i2.GSR = "DISABLED";
    LUT4 power_counter_31__I_0_77_i2_3_lut (.A(power_counter_31__N_232[1]), 
         .B(power_counter_31__N_201[1]), .C(power_counter[31]), .Z(power_counter_31__N_129[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(231[4:54])
    defparam power_counter_31__I_0_77_i2_3_lut.init = 16'hcaca;
    FD1S3AX wb_idata_i1 (.D(wb_idata_31__N_1[1]), .CK(i_ref_clk_c), .Q(wb_idata[1]));   // d:/documents/git_local/fm_modulator/rtl/top.v(267[9] 275[22])
    defparam wb_idata_i1.GSR = "DISABLED";
    LUT4 i755_1_lut (.A(o_baseband_q_c_15), .Z(o_baseband_q_c_9)) /* synthesis lut_function=(!(A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(113[31:66])
    defparam i755_1_lut.init = 16'h5555;
    LUT4 i3_4_lut_rep_574 (.A(wb_addr[3]), .B(wb_addr[2]), .C(wb_addr[0]), 
         .D(wb_addr[1]), .Z(n25134)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(209[4:8])
    defparam i3_4_lut_rep_574.init = 16'hfffb;
    efb_inst wb_lo_data_7__I_0 (.i_ref_clk_c(i_ref_clk_c), .i_resetb_N_301(i_resetb_N_301), 
            .n27585(n27585), .wb_lo_data_7__N_96(wb_lo_data_7__N_96), .wb_we(wb_we), 
            .\wb_addr[7] (wb_addr[7]), .\wb_addr[6] (wb_addr[6]), .\wb_addr[5] (wb_addr[5]), 
            .\wb_addr[4] (wb_addr[4]), .\wb_addr[3] (wb_addr[3]), .\wb_addr[2] (wb_addr[2]), 
            .\wb_addr[1] (wb_addr[1]), .\wb_addr[0] (wb_addr[0]), .\wb_odata[7] (wb_odata[7]), 
            .\wb_odata[6] (wb_odata[6]), .\wb_odata[5] (wb_odata[5]), .\wb_odata[4] (wb_odata[4]), 
            .\wb_odata[3] (wb_odata[3]), .\wb_odata[2] (wb_odata[2]), .\wb_odata[1] (wb_odata[1]), 
            .\wb_odata[0] (wb_odata[0]), .pll_data_o({pll_data_o}), .pll_ack(pll_ack), 
            .wb_lo_data({wb_lo_data}), .wb_lo_ack(wb_lo_ack), .pll_clk(pll_clk), 
            .pll_rst(pll_rst), .pll_stb(pll_stb), .pll_we(pll_we), .pll_addr({pll_addr}), 
            .pll_data_i({pll_data_i}), .GND_net(GND_net), .VCC_net(VCC_net)) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(179[10] 191[3])
    VLO i1 (.Z(GND_net));
    clock_phase_shifter clock_phase_shifter_inst (.q_clk_p_c(q_clk_p_c), .i_clk_2f_N_2249(i_clk_2f_N_2249), 
            .q_clk_n_c(q_clk_n_c), .i_clk_p_c(i_clk_p_c), .lo_pll_out(lo_pll_out), 
            .i_clk_n_c(i_clk_n_c)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(160[21] 164[2])
    CCU2D add_35_21 (.A0(power_counter[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17292), .COUT(n17293), .S0(power_counter_31__N_201[19]), 
          .S1(power_counter_31__N_201[20]));   // d:/documents/git_local/fm_modulator/rtl/top.v(231[27:53])
    defparam add_35_21.INIT0 = 16'h5aaa;
    defparam add_35_21.INIT1 = 16'h5aaa;
    defparam add_35_21.INJECT1_0 = "NO";
    defparam add_35_21.INJECT1_1 = "NO";
    CCU2D add_34_17 (.A0(power_counter[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17274), .COUT(n17275), .S0(power_counter_31__N_232[15]), 
          .S1(power_counter_31__N_232[16]));   // d:/documents/git_local/fm_modulator/rtl/top.v(229[21:41])
    defparam add_34_17.INIT0 = 16'h5aaa;
    defparam add_34_17.INIT1 = 16'h5aaa;
    defparam add_34_17.INJECT1_0 = "NO";
    defparam add_34_17.INJECT1_1 = "NO";
    CCU2D add_35_19 (.A0(power_counter[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17291), .COUT(n17292), .S0(power_counter_31__N_201[17]), 
          .S1(power_counter_31__N_201[18]));   // d:/documents/git_local/fm_modulator/rtl/top.v(231[27:53])
    defparam add_35_19.INIT0 = 16'h5aaa;
    defparam add_35_19.INIT1 = 16'h5aaa;
    defparam add_35_19.INJECT1_0 = "NO";
    defparam add_35_19.INJECT1_1 = "NO";
    CCU2D add_34_15 (.A0(power_counter[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17273), .COUT(n17274), .S0(power_counter_31__N_232[13]), 
          .S1(power_counter_31__N_232[14]));   // d:/documents/git_local/fm_modulator/rtl/top.v(229[21:41])
    defparam add_34_15.INIT0 = 16'h5aaa;
    defparam add_34_15.INIT1 = 16'h5aaa;
    defparam add_34_15.INJECT1_0 = "NO";
    defparam add_34_15.INJECT1_1 = "NO";
    CCU2D add_35_17 (.A0(power_counter[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17290), .COUT(n17291), .S0(power_counter_31__N_201[15]), 
          .S1(power_counter_31__N_201[16]));   // d:/documents/git_local/fm_modulator/rtl/top.v(231[27:53])
    defparam add_35_17.INIT0 = 16'h5aaa;
    defparam add_35_17.INIT1 = 16'h5aaa;
    defparam add_35_17.INJECT1_0 = "NO";
    defparam add_35_17.INJECT1_1 = "NO";
    CCU2D add_34_5 (.A0(power_counter[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17268), .COUT(n17269), .S0(power_counter_31__N_232[3]), 
          .S1(power_counter_31__N_232[4]));   // d:/documents/git_local/fm_modulator/rtl/top.v(229[21:41])
    defparam add_34_5.INIT0 = 16'h5aaa;
    defparam add_34_5.INIT1 = 16'h5aaa;
    defparam add_34_5.INJECT1_0 = "NO";
    defparam add_34_5.INJECT1_1 = "NO";
    CCU2D add_35_15 (.A0(power_counter[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17289), .COUT(n17290), .S0(power_counter_31__N_201[13]), 
          .S1(power_counter_31__N_201[14]));   // d:/documents/git_local/fm_modulator/rtl/top.v(231[27:53])
    defparam add_35_15.INIT0 = 16'h5aaa;
    defparam add_35_15.INIT1 = 16'h5aaa;
    defparam add_35_15.INJECT1_0 = "NO";
    defparam add_35_15.INJECT1_1 = "NO";
    OB o_baseband_i_pad_6 (.I(o_baseband_i_c_13), .O(o_baseband_i[6]));   // d:/documents/git_local/fm_modulator/rtl/top.v(27[38:50])
    FD1P3AX power_counter_i31 (.D(n27530), .SP(power_counter_31__N_232[31]), 
            .CK(i_ref_clk_c), .Q(power_counter[31])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(226[9] 231[54])
    defparam power_counter_i31.GSR = "DISABLED";
    FD1S3AX power_counter_i30 (.D(power_counter_31__N_129[30]), .CK(i_ref_clk_c), 
            .Q(power_counter[30])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(226[9] 231[54])
    defparam power_counter_i30.GSR = "DISABLED";
    FD1S3AX power_counter_i29 (.D(power_counter_31__N_129[29]), .CK(i_ref_clk_c), 
            .Q(power_counter[29])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(226[9] 231[54])
    defparam power_counter_i29.GSR = "DISABLED";
    FD1S3AX power_counter_i28 (.D(power_counter_31__N_129[28]), .CK(i_ref_clk_c), 
            .Q(power_counter[28])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(226[9] 231[54])
    defparam power_counter_i28.GSR = "DISABLED";
    FD1S3AX power_counter_i27 (.D(power_counter_31__N_129[27]), .CK(i_ref_clk_c), 
            .Q(power_counter[27])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(226[9] 231[54])
    defparam power_counter_i27.GSR = "DISABLED";
    FD1S3AX power_counter_i26 (.D(power_counter_31__N_129[26]), .CK(i_ref_clk_c), 
            .Q(power_counter[26])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(226[9] 231[54])
    defparam power_counter_i26.GSR = "DISABLED";
    FD1S3AX power_counter_i25 (.D(power_counter_31__N_129[25]), .CK(i_ref_clk_c), 
            .Q(power_counter[25])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(226[9] 231[54])
    defparam power_counter_i25.GSR = "DISABLED";
    FD1S3AX power_counter_i24 (.D(power_counter_31__N_129[24]), .CK(i_ref_clk_c), 
            .Q(power_counter[24])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(226[9] 231[54])
    defparam power_counter_i24.GSR = "DISABLED";
    FD1S3AX power_counter_i23 (.D(power_counter_31__N_129[23]), .CK(i_ref_clk_c), 
            .Q(power_counter[23])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(226[9] 231[54])
    defparam power_counter_i23.GSR = "DISABLED";
    FD1S3AX power_counter_i22 (.D(power_counter_31__N_129[22]), .CK(i_ref_clk_c), 
            .Q(power_counter[22])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(226[9] 231[54])
    defparam power_counter_i22.GSR = "DISABLED";
    FD1S3AX power_counter_i21 (.D(power_counter_31__N_129[21]), .CK(i_ref_clk_c), 
            .Q(power_counter[21])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(226[9] 231[54])
    defparam power_counter_i21.GSR = "DISABLED";
    FD1S3AX power_counter_i20 (.D(power_counter_31__N_129[20]), .CK(i_ref_clk_c), 
            .Q(power_counter[20])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(226[9] 231[54])
    defparam power_counter_i20.GSR = "DISABLED";
    FD1S3AX power_counter_i19 (.D(power_counter_31__N_129[19]), .CK(i_ref_clk_c), 
            .Q(power_counter[19])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(226[9] 231[54])
    defparam power_counter_i19.GSR = "DISABLED";
    FD1S3AX power_counter_i18 (.D(power_counter_31__N_129[18]), .CK(i_ref_clk_c), 
            .Q(power_counter[18])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(226[9] 231[54])
    defparam power_counter_i18.GSR = "DISABLED";
    FD1S3AX power_counter_i17 (.D(power_counter_31__N_129[17]), .CK(i_ref_clk_c), 
            .Q(power_counter[17])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(226[9] 231[54])
    defparam power_counter_i17.GSR = "DISABLED";
    CCU2D add_35_13 (.A0(power_counter[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17288), .COUT(n17289), .S0(power_counter_31__N_201[11]), 
          .S1(power_counter_31__N_201[12]));   // d:/documents/git_local/fm_modulator/rtl/top.v(231[27:53])
    defparam add_35_13.INIT0 = 16'h5aaa;
    defparam add_35_13.INIT1 = 16'h5aaa;
    defparam add_35_13.INJECT1_0 = "NO";
    defparam add_35_13.INJECT1_1 = "NO";
    CCU2D add_35_11 (.A0(power_counter[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17287), .COUT(n17288), .S0(power_counter_31__N_201[9]), 
          .S1(power_counter_31__N_201[10]));   // d:/documents/git_local/fm_modulator/rtl/top.v(231[27:53])
    defparam add_35_11.INIT0 = 16'h5aaa;
    defparam add_35_11.INIT1 = 16'h5aaa;
    defparam add_35_11.INJECT1_0 = "NO";
    defparam add_35_11.INJECT1_1 = "NO";
    CCU2D add_35_9 (.A0(power_counter[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17286), .COUT(n17287), .S0(power_counter_31__N_201[7]), 
          .S1(power_counter_31__N_201[8]));   // d:/documents/git_local/fm_modulator/rtl/top.v(231[27:53])
    defparam add_35_9.INIT0 = 16'h5aaa;
    defparam add_35_9.INIT1 = 16'h5aaa;
    defparam add_35_9.INJECT1_0 = "NO";
    defparam add_35_9.INJECT1_1 = "NO";
    CCU2D add_34_9 (.A0(power_counter[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17270), .COUT(n17271), .S0(power_counter_31__N_232[7]), 
          .S1(power_counter_31__N_232[8]));   // d:/documents/git_local/fm_modulator/rtl/top.v(229[21:41])
    defparam add_34_9.INIT0 = 16'h5aaa;
    defparam add_34_9.INIT1 = 16'h5aaa;
    defparam add_34_9.INJECT1_0 = "NO";
    defparam add_34_9.INJECT1_1 = "NO";
    CCU2D add_35_7 (.A0(power_counter[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17285), .COUT(n17286), .S0(power_counter_31__N_201[5]), 
          .S1(power_counter_31__N_201[6]));   // d:/documents/git_local/fm_modulator/rtl/top.v(231[27:53])
    defparam add_35_7.INIT0 = 16'h5aaa;
    defparam add_35_7.INIT1 = 16'h5aaa;
    defparam add_35_7.INJECT1_0 = "NO";
    defparam add_35_7.INJECT1_1 = "NO";
    CCU2D add_35_5 (.A0(power_counter[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17284), .COUT(n17285), .S0(power_counter_31__N_201[3]), 
          .S1(power_counter_31__N_201[4]));   // d:/documents/git_local/fm_modulator/rtl/top.v(231[27:53])
    defparam add_35_5.INIT0 = 16'h5aaa;
    defparam add_35_5.INIT1 = 16'h5aaa;
    defparam add_35_5.INJECT1_0 = "NO";
    defparam add_35_5.INJECT1_1 = "NO";
    CCU2D add_34_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(power_counter[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n17267), .S1(power_counter_31__N_232[0]));   // d:/documents/git_local/fm_modulator/rtl/top.v(229[21:41])
    defparam add_34_1.INIT0 = 16'hF000;
    defparam add_34_1.INIT1 = 16'h5555;
    defparam add_34_1.INJECT1_0 = "NO";
    defparam add_34_1.INJECT1_1 = "NO";
    CCU2D add_35_3 (.A0(power_counter[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17283), .COUT(n17284), .S0(power_counter_31__N_201[1]), 
          .S1(power_counter_31__N_201[2]));   // d:/documents/git_local/fm_modulator/rtl/top.v(231[27:53])
    defparam add_35_3.INIT0 = 16'h5aaa;
    defparam add_35_3.INIT1 = 16'h5aaa;
    defparam add_35_3.INJECT1_0 = "NO";
    defparam add_35_3.INJECT1_1 = "NO";
    CCU2D add_35_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(power_counter[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n17283), .S1(power_counter_31__N_201[0]));   // d:/documents/git_local/fm_modulator/rtl/top.v(231[27:53])
    defparam add_35_1.INIT0 = 16'hF000;
    defparam add_35_1.INIT1 = 16'h5555;
    defparam add_35_1.INJECT1_0 = "NO";
    defparam add_35_1.INJECT1_1 = "NO";
    CCU2D add_34_3 (.A0(power_counter[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17267), .COUT(n17268), .S0(power_counter_31__N_232[1]), 
          .S1(power_counter_31__N_232[2]));   // d:/documents/git_local/fm_modulator/rtl/top.v(229[21:41])
    defparam add_34_3.INIT0 = 16'h5aaa;
    defparam add_34_3.INIT1 = 16'h5aaa;
    defparam add_34_3.INJECT1_0 = "NO";
    defparam add_34_3.INJECT1_1 = "NO";
    CCU2D add_34_33 (.A0(power_counter[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n17282), .S0(power_counter_31__N_232[31]));   // d:/documents/git_local/fm_modulator/rtl/top.v(229[21:41])
    defparam add_34_33.INIT0 = 16'h5aaa;
    defparam add_34_33.INIT1 = 16'h0000;
    defparam add_34_33.INJECT1_0 = "NO";
    defparam add_34_33.INJECT1_1 = "NO";
    CCU2D add_34_13 (.A0(power_counter[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17272), .COUT(n17273), .S0(power_counter_31__N_232[11]), 
          .S1(power_counter_31__N_232[12]));   // d:/documents/git_local/fm_modulator/rtl/top.v(229[21:41])
    defparam add_34_13.INIT0 = 16'h5aaa;
    defparam add_34_13.INIT1 = 16'h5aaa;
    defparam add_34_13.INJECT1_0 = "NO";
    defparam add_34_13.INJECT1_1 = "NO";
    CCU2D add_34_31 (.A0(power_counter[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17281), .COUT(n17282), .S0(power_counter_31__N_232[29]), 
          .S1(power_counter_31__N_232[30]));   // d:/documents/git_local/fm_modulator/rtl/top.v(229[21:41])
    defparam add_34_31.INIT0 = 16'h5aaa;
    defparam add_34_31.INIT1 = 16'h5aaa;
    defparam add_34_31.INJECT1_0 = "NO";
    defparam add_34_31.INJECT1_1 = "NO";
    CCU2D add_34_7 (.A0(power_counter[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17269), .COUT(n17270), .S0(power_counter_31__N_232[5]), 
          .S1(power_counter_31__N_232[6]));   // d:/documents/git_local/fm_modulator/rtl/top.v(229[21:41])
    defparam add_34_7.INIT0 = 16'h5aaa;
    defparam add_34_7.INIT1 = 16'h5aaa;
    defparam add_34_7.INJECT1_0 = "NO";
    defparam add_34_7.INJECT1_1 = "NO";
    CCU2D add_34_29 (.A0(power_counter[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17280), .COUT(n17281), .S0(power_counter_31__N_232[27]), 
          .S1(power_counter_31__N_232[28]));   // d:/documents/git_local/fm_modulator/rtl/top.v(229[21:41])
    defparam add_34_29.INIT0 = 16'h5aaa;
    defparam add_34_29.INIT1 = 16'h5aaa;
    defparam add_34_29.INJECT1_0 = "NO";
    defparam add_34_29.INJECT1_1 = "NO";
    CCU2D add_34_11 (.A0(power_counter[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17271), .COUT(n17272), .S0(power_counter_31__N_232[9]), 
          .S1(power_counter_31__N_232[10]));   // d:/documents/git_local/fm_modulator/rtl/top.v(229[21:41])
    defparam add_34_11.INIT0 = 16'h5aaa;
    defparam add_34_11.INIT1 = 16'h5aaa;
    defparam add_34_11.INJECT1_0 = "NO";
    defparam add_34_11.INJECT1_1 = "NO";
    CCU2D add_34_27 (.A0(power_counter[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17279), .COUT(n17280), .S0(power_counter_31__N_232[25]), 
          .S1(power_counter_31__N_232[26]));   // d:/documents/git_local/fm_modulator/rtl/top.v(229[21:41])
    defparam add_34_27.INIT0 = 16'h5aaa;
    defparam add_34_27.INIT1 = 16'h5aaa;
    defparam add_34_27.INJECT1_0 = "NO";
    defparam add_34_27.INJECT1_1 = "NO";
    FD1S3AX power_counter_i16 (.D(power_counter_31__N_129[16]), .CK(i_ref_clk_c), 
            .Q(power_counter[16])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(226[9] 231[54])
    defparam power_counter_i16.GSR = "DISABLED";
    TSALL TSALL_INST (.TSALL(GND_net));
    LUT4 m1_lut (.Z(n27530)) /* synthesis lut_function=1, syn_instantiated=1 */ ;
    defparam m1_lut.init = 16'hffff;
    FD1S3AX power_counter_i15 (.D(power_counter_31__N_129[15]), .CK(i_ref_clk_c), 
            .Q(power_counter[15])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(226[9] 231[54])
    defparam power_counter_i15.GSR = "DISABLED";
    FD1S3AX power_counter_i14 (.D(power_counter_31__N_129[14]), .CK(i_ref_clk_c), 
            .Q(power_counter[14])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(226[9] 231[54])
    defparam power_counter_i14.GSR = "DISABLED";
    FD1S3AX power_counter_i13 (.D(power_counter_31__N_129[13]), .CK(i_ref_clk_c), 
            .Q(power_counter[13])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(226[9] 231[54])
    defparam power_counter_i13.GSR = "DISABLED";
    FD1S3AX power_counter_i12 (.D(power_counter_31__N_129[12]), .CK(i_ref_clk_c), 
            .Q(power_counter[12])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(226[9] 231[54])
    defparam power_counter_i12.GSR = "DISABLED";
    FD1S3AX power_counter_i11 (.D(power_counter_31__N_129[11]), .CK(i_ref_clk_c), 
            .Q(power_counter[11])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(226[9] 231[54])
    defparam power_counter_i11.GSR = "DISABLED";
    FD1S3AX power_counter_i10 (.D(power_counter_31__N_129[10]), .CK(i_ref_clk_c), 
            .Q(power_counter[10])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(226[9] 231[54])
    defparam power_counter_i10.GSR = "DISABLED";
    FD1S3AX power_counter_i9 (.D(power_counter_31__N_129[9]), .CK(i_ref_clk_c), 
            .Q(power_counter[9])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(226[9] 231[54])
    defparam power_counter_i9.GSR = "DISABLED";
    FD1S3AX power_counter_i8 (.D(power_counter_31__N_129[8]), .CK(i_ref_clk_c), 
            .Q(power_counter[8])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(226[9] 231[54])
    defparam power_counter_i8.GSR = "DISABLED";
    FD1S3AX power_counter_i7 (.D(power_counter_31__N_129[7]), .CK(i_ref_clk_c), 
            .Q(power_counter[7])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(226[9] 231[54])
    defparam power_counter_i7.GSR = "DISABLED";
    FD1S3AX power_counter_i6 (.D(power_counter_31__N_129[6]), .CK(i_ref_clk_c), 
            .Q(power_counter[6])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(226[9] 231[54])
    defparam power_counter_i6.GSR = "DISABLED";
    FD1S3AX power_counter_i5 (.D(power_counter_31__N_129[5]), .CK(i_ref_clk_c), 
            .Q(power_counter[5])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(226[9] 231[54])
    defparam power_counter_i5.GSR = "DISABLED";
    FD1S3AX power_counter_i4 (.D(power_counter_31__N_129[4]), .CK(i_ref_clk_c), 
            .Q(power_counter[4])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(226[9] 231[54])
    defparam power_counter_i4.GSR = "DISABLED";
    FD1S3AX power_counter_i3 (.D(power_counter_31__N_129[3]), .CK(i_ref_clk_c), 
            .Q(power_counter[3])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(226[9] 231[54])
    defparam power_counter_i3.GSR = "DISABLED";
    FD1S3AX power_counter_i2 (.D(power_counter_31__N_129[2]), .CK(i_ref_clk_c), 
            .Q(power_counter[2])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(226[9] 231[54])
    defparam power_counter_i2.GSR = "DISABLED";
    FD1S3AX power_counter_i1 (.D(power_counter_31__N_129[1]), .CK(i_ref_clk_c), 
            .Q(power_counter[1])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(226[9] 231[54])
    defparam power_counter_i1.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i31 (.D(n2109), .CK(i_ref_clk_c), .CD(n9456), 
            .Q(wb_smpl_data[31]));   // d:/documents/git_local/fm_modulator/rtl/top.v(214[9] 222[10])
    defparam wb_smpl_data_i31.GSR = "DISABLED";
    \rxuartlite(CLOCKS_PER_BAUD=20)  rxtransport (.i_ref_clk_c(i_ref_clk_c), 
            .\rx_data[0] (rx_data[0]), .rx_stb(rx_stb), .i_wbu_uart_rx_c(i_wbu_uart_rx_c), 
            .chg_counter({chg_counter}), .i_ref_clk_c_enable_180(i_ref_clk_c_enable_180), 
            .chg_counter_23__N_406(chg_counter_23__N_406), .GND_net(GND_net), 
            .\rx_data[6] (rx_data[6]), .\rx_data[5] (rx_data[5]), .\rx_data[4] (rx_data[4]), 
            .\rx_data[3] (rx_data[3]), .\rx_data[2] (rx_data[2]), .\rx_data[1] (rx_data[1])) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(54[54:102])
    FD1S3IX wb_smpl_data_i30 (.D(n2110), .CK(i_ref_clk_c), .CD(n9456), 
            .Q(wb_smpl_data[30]));   // d:/documents/git_local/fm_modulator/rtl/top.v(214[9] 222[10])
    defparam wb_smpl_data_i30.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i29 (.D(n24795), .CK(i_ref_clk_c), .CD(n9456), 
            .Q(wb_smpl_data[29]));   // d:/documents/git_local/fm_modulator/rtl/top.v(214[9] 222[10])
    defparam wb_smpl_data_i29.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i28 (.D(n2112), .CK(i_ref_clk_c), .CD(n9456), 
            .Q(wb_smpl_data[28]));   // d:/documents/git_local/fm_modulator/rtl/top.v(214[9] 222[10])
    defparam wb_smpl_data_i28.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i27 (.D(n2113), .CK(i_ref_clk_c), .CD(n9456), 
            .Q(wb_smpl_data[27]));   // d:/documents/git_local/fm_modulator/rtl/top.v(214[9] 222[10])
    defparam wb_smpl_data_i27.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i26 (.D(n2114), .CK(i_ref_clk_c), .CD(n9456), 
            .Q(wb_smpl_data[26]));   // d:/documents/git_local/fm_modulator/rtl/top.v(214[9] 222[10])
    defparam wb_smpl_data_i26.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i25 (.D(n2115), .CK(i_ref_clk_c), .CD(n9456), 
            .Q(wb_smpl_data[25]));   // d:/documents/git_local/fm_modulator/rtl/top.v(214[9] 222[10])
    defparam wb_smpl_data_i25.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i24 (.D(n2116), .CK(i_ref_clk_c), .CD(n9456), 
            .Q(wb_smpl_data[24]));   // d:/documents/git_local/fm_modulator/rtl/top.v(214[9] 222[10])
    defparam wb_smpl_data_i24.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i23 (.D(n2117), .CK(i_ref_clk_c), .CD(n9456), 
            .Q(wb_smpl_data[23]));   // d:/documents/git_local/fm_modulator/rtl/top.v(214[9] 222[10])
    defparam wb_smpl_data_i23.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i22 (.D(n2118), .CK(i_ref_clk_c), .CD(n9456), 
            .Q(wb_smpl_data[22]));   // d:/documents/git_local/fm_modulator/rtl/top.v(214[9] 222[10])
    defparam wb_smpl_data_i22.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i29 (.D(wb_addr[29]), .SP(wb_err), .CK(i_ref_clk_c), 
            .Q(bus_err_address[29])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(257[9] 259[31])
    defparam bus_err_address_i0_i29.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i28 (.D(wb_addr[28]), .SP(wb_err), .CK(i_ref_clk_c), 
            .Q(bus_err_address[28])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(257[9] 259[31])
    defparam bus_err_address_i0_i28.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i27 (.D(wb_addr[27]), .SP(wb_err), .CK(i_ref_clk_c), 
            .Q(bus_err_address[27])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(257[9] 259[31])
    defparam bus_err_address_i0_i27.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i26 (.D(wb_addr[26]), .SP(wb_err), .CK(i_ref_clk_c), 
            .Q(bus_err_address[26])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(257[9] 259[31])
    defparam bus_err_address_i0_i26.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i25 (.D(wb_addr[25]), .SP(wb_err), .CK(i_ref_clk_c), 
            .Q(bus_err_address[25])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(257[9] 259[31])
    defparam bus_err_address_i0_i25.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i24 (.D(wb_addr[24]), .SP(wb_err), .CK(i_ref_clk_c), 
            .Q(bus_err_address[24])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(257[9] 259[31])
    defparam bus_err_address_i0_i24.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i23 (.D(wb_addr[23]), .SP(wb_err), .CK(i_ref_clk_c), 
            .Q(bus_err_address[23])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(257[9] 259[31])
    defparam bus_err_address_i0_i23.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i22 (.D(wb_addr[22]), .SP(wb_err), .CK(i_ref_clk_c), 
            .Q(bus_err_address[22])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(257[9] 259[31])
    defparam bus_err_address_i0_i22.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i21 (.D(wb_addr[21]), .SP(wb_err), .CK(i_ref_clk_c), 
            .Q(bus_err_address[21])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(257[9] 259[31])
    defparam bus_err_address_i0_i21.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i20 (.D(wb_addr[20]), .SP(wb_err), .CK(i_ref_clk_c), 
            .Q(bus_err_address[20])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(257[9] 259[31])
    defparam bus_err_address_i0_i20.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i19 (.D(wb_addr[19]), .SP(wb_err), .CK(i_ref_clk_c), 
            .Q(bus_err_address[19])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(257[9] 259[31])
    defparam bus_err_address_i0_i19.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i18 (.D(wb_addr[18]), .SP(wb_err), .CK(i_ref_clk_c), 
            .Q(bus_err_address[18])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(257[9] 259[31])
    defparam bus_err_address_i0_i18.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i17 (.D(wb_addr[17]), .SP(wb_err), .CK(i_ref_clk_c), 
            .Q(bus_err_address[17])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(257[9] 259[31])
    defparam bus_err_address_i0_i17.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i16 (.D(wb_addr[16]), .SP(wb_err), .CK(i_ref_clk_c), 
            .Q(bus_err_address[16])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(257[9] 259[31])
    defparam bus_err_address_i0_i16.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i15 (.D(wb_addr[15]), .SP(wb_err), .CK(i_ref_clk_c), 
            .Q(bus_err_address[15])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(257[9] 259[31])
    defparam bus_err_address_i0_i15.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i14 (.D(wb_addr[14]), .SP(wb_err), .CK(i_ref_clk_c), 
            .Q(bus_err_address[14])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(257[9] 259[31])
    defparam bus_err_address_i0_i14.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i13 (.D(wb_addr[13]), .SP(wb_err), .CK(i_ref_clk_c), 
            .Q(bus_err_address[13])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(257[9] 259[31])
    defparam bus_err_address_i0_i13.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i12 (.D(wb_addr[12]), .SP(wb_err), .CK(i_ref_clk_c), 
            .Q(bus_err_address[12])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(257[9] 259[31])
    defparam bus_err_address_i0_i12.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i11 (.D(wb_addr[11]), .SP(wb_err), .CK(i_ref_clk_c), 
            .Q(bus_err_address[11])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(257[9] 259[31])
    defparam bus_err_address_i0_i11.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i10 (.D(wb_addr[10]), .SP(wb_err), .CK(i_ref_clk_c), 
            .Q(bus_err_address[10])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(257[9] 259[31])
    defparam bus_err_address_i0_i10.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i9 (.D(wb_addr[9]), .SP(wb_err), .CK(i_ref_clk_c), 
            .Q(bus_err_address[9])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(257[9] 259[31])
    defparam bus_err_address_i0_i9.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i8 (.D(wb_addr[8]), .SP(wb_err), .CK(i_ref_clk_c), 
            .Q(bus_err_address[8])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(257[9] 259[31])
    defparam bus_err_address_i0_i8.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i7 (.D(wb_addr[7]), .SP(wb_err), .CK(i_ref_clk_c), 
            .Q(bus_err_address[7])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(257[9] 259[31])
    defparam bus_err_address_i0_i7.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i6 (.D(wb_addr[6]), .SP(wb_err), .CK(i_ref_clk_c), 
            .Q(bus_err_address[6])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(257[9] 259[31])
    defparam bus_err_address_i0_i6.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i5 (.D(wb_addr[5]), .SP(wb_err), .CK(i_ref_clk_c), 
            .Q(bus_err_address[5])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(257[9] 259[31])
    defparam bus_err_address_i0_i5.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i4 (.D(wb_addr[4]), .SP(wb_err), .CK(i_ref_clk_c), 
            .Q(bus_err_address[4])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(257[9] 259[31])
    defparam bus_err_address_i0_i4.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i3 (.D(wb_addr[3]), .SP(wb_err), .CK(i_ref_clk_c), 
            .Q(bus_err_address[3])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(257[9] 259[31])
    defparam bus_err_address_i0_i3.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i2 (.D(wb_addr[2]), .SP(wb_err), .CK(i_ref_clk_c), 
            .Q(bus_err_address[2])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(257[9] 259[31])
    defparam bus_err_address_i0_i2.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i1 (.D(wb_addr[1]), .SP(wb_err), .CK(i_ref_clk_c), 
            .Q(bus_err_address[1])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(257[9] 259[31])
    defparam bus_err_address_i0_i1.GSR = "DISABLED";
    LUT4 m0_lut (.Z(n27529)) /* synthesis lut_function=0, syn_instantiated=1 */ ;
    defparam m0_lut.init = 16'h0000;
    FD1S3IX wb_smpl_data_i21 (.D(n2119), .CK(i_ref_clk_c), .CD(n9456), 
            .Q(wb_smpl_data[21]));   // d:/documents/git_local/fm_modulator/rtl/top.v(214[9] 222[10])
    defparam wb_smpl_data_i21.GSR = "DISABLED";
    OB o_baseband_i_pad_5 (.I(o_baseband_i_c_12), .O(o_baseband_i[5]));   // d:/documents/git_local/fm_modulator/rtl/top.v(27[38:50])
    OB o_baseband_i_pad_4 (.I(o_baseband_i_c_11), .O(o_baseband_i[4]));   // d:/documents/git_local/fm_modulator/rtl/top.v(27[38:50])
    OB o_baseband_i_pad_3 (.I(o_baseband_i_c_10), .O(o_baseband_i[3]));   // d:/documents/git_local/fm_modulator/rtl/top.v(27[38:50])
    OB o_baseband_i_pad_2 (.I(n3607), .O(o_baseband_i[2]));   // d:/documents/git_local/fm_modulator/rtl/top.v(27[38:50])
    OB o_baseband_i_pad_1 (.I(o_baseband_i_c_8), .O(o_baseband_i[1]));   // d:/documents/git_local/fm_modulator/rtl/top.v(27[38:50])
    OB o_baseband_i_pad_0 (.I(o_baseband_i_c_7), .O(o_baseband_i[0]));   // d:/documents/git_local/fm_modulator/rtl/top.v(27[38:50])
    OB o_baseband_q_pad_9 (.I(o_baseband_q_c_9), .O(o_baseband_q[9]));   // d:/documents/git_local/fm_modulator/rtl/top.v(27[52:64])
    OB o_baseband_q_pad_8 (.I(o_baseband_q_c_15), .O(o_baseband_q[8]));   // d:/documents/git_local/fm_modulator/rtl/top.v(27[52:64])
    OB o_baseband_q_pad_7 (.I(o_baseband_q_c_14), .O(o_baseband_q[7]));   // d:/documents/git_local/fm_modulator/rtl/top.v(27[52:64])
    OB o_baseband_q_pad_6 (.I(o_baseband_q_c_13), .O(o_baseband_q[6]));   // d:/documents/git_local/fm_modulator/rtl/top.v(27[52:64])
    OB o_baseband_q_pad_5 (.I(o_baseband_q_c_12), .O(o_baseband_q[5]));   // d:/documents/git_local/fm_modulator/rtl/top.v(27[52:64])
    OB o_baseband_q_pad_4 (.I(o_baseband_q_c_11), .O(o_baseband_q[4]));   // d:/documents/git_local/fm_modulator/rtl/top.v(27[52:64])
    OB o_baseband_q_pad_3 (.I(o_baseband_q_c_10), .O(o_baseband_q[3]));   // d:/documents/git_local/fm_modulator/rtl/top.v(27[52:64])
    OB o_baseband_q_pad_2 (.I(n3608), .O(o_baseband_q[2]));   // d:/documents/git_local/fm_modulator/rtl/top.v(27[52:64])
    OB o_baseband_q_pad_1 (.I(o_baseband_q_c_8), .O(o_baseband_q[1]));   // d:/documents/git_local/fm_modulator/rtl/top.v(27[52:64])
    OB o_baseband_q_pad_0 (.I(o_baseband_q_c_7), .O(o_baseband_q[0]));   // d:/documents/git_local/fm_modulator/rtl/top.v(27[52:64])
    OB dac_clk_p_pad (.I(GND_net), .O(dac_clk_p));   // d:/documents/git_local/fm_modulator/rtl/top.v(28[49:58])
    OB dac_clk_n_pad (.I(VCC_net), .O(dac_clk_n));   // d:/documents/git_local/fm_modulator/rtl/top.v(28[60:69])
    OB i_clk_p_pad (.I(i_clk_p_c), .O(i_clk_p));   // d:/documents/git_local/fm_modulator/rtl/top.v(28[13:20])
    OB i_clk_n_pad (.I(i_clk_n_c), .O(i_clk_n));   // d:/documents/git_local/fm_modulator/rtl/top.v(28[22:29])
    OB q_clk_p_pad (.I(q_clk_p_c), .O(q_clk_p));   // d:/documents/git_local/fm_modulator/rtl/top.v(28[31:38])
    OB q_clk_n_pad (.I(q_clk_n_c), .O(q_clk_n));   // d:/documents/git_local/fm_modulator/rtl/top.v(28[40:47])
    IB i_ref_clk_pad (.I(i_ref_clk), .O(i_ref_clk_c));   // d:/documents/git_local/fm_modulator/rtl/top.v(22[12:21])
    IB i_resetb_pad (.I(i_resetb), .O(i_resetb_c));   // d:/documents/git_local/fm_modulator/rtl/top.v(22[23:31])
    IB i_wbu_uart_rx_pad (.I(i_wbu_uart_rx), .O(i_wbu_uart_rx_c));   // d:/documents/git_local/fm_modulator/rtl/top.v(24[12:25])
    FD1S3IX wb_smpl_data_i3 (.D(n2137), .CK(i_ref_clk_c), .CD(n9456), 
            .Q(wb_smpl_data[3]));   // d:/documents/git_local/fm_modulator/rtl/top.v(214[9] 222[10])
    defparam wb_smpl_data_i3.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i20 (.D(n24794), .CK(i_ref_clk_c), .CD(n9456), 
            .Q(wb_smpl_data[20]));   // d:/documents/git_local/fm_modulator/rtl/top.v(214[9] 222[10])
    defparam wb_smpl_data_i20.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i2 (.D(n2138), .CK(i_ref_clk_c), .CD(n9456), 
            .Q(wb_smpl_data[2]));   // d:/documents/git_local/fm_modulator/rtl/top.v(214[9] 222[10])
    defparam wb_smpl_data_i2.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i19 (.D(n2121), .CK(i_ref_clk_c), .CD(n9456), 
            .Q(wb_smpl_data[19]));   // d:/documents/git_local/fm_modulator/rtl/top.v(214[9] 222[10])
    defparam wb_smpl_data_i19.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i1 (.D(n2139), .CK(i_ref_clk_c), .CD(n9456), 
            .Q(wb_smpl_data[1]));   // d:/documents/git_local/fm_modulator/rtl/top.v(214[9] 222[10])
    defparam wb_smpl_data_i1.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i18 (.D(n24793), .CK(i_ref_clk_c), .CD(n9456), 
            .Q(wb_smpl_data[18]));   // d:/documents/git_local/fm_modulator/rtl/top.v(214[9] 222[10])
    defparam wb_smpl_data_i18.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i17 (.D(n24792), .CK(i_ref_clk_c), .CD(n9456), 
            .Q(wb_smpl_data[17]));   // d:/documents/git_local/fm_modulator/rtl/top.v(214[9] 222[10])
    defparam wb_smpl_data_i17.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i16 (.D(n24791), .CK(i_ref_clk_c), .CD(n9456), 
            .Q(wb_smpl_data[16]));   // d:/documents/git_local/fm_modulator/rtl/top.v(214[9] 222[10])
    defparam wb_smpl_data_i16.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i15 (.D(n2125), .CK(i_ref_clk_c), .CD(n9456), 
            .Q(wb_smpl_data[15]));   // d:/documents/git_local/fm_modulator/rtl/top.v(214[9] 222[10])
    defparam wb_smpl_data_i15.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i14 (.D(n2126), .CK(i_ref_clk_c), .CD(n9456), 
            .Q(wb_smpl_data[14]));   // d:/documents/git_local/fm_modulator/rtl/top.v(214[9] 222[10])
    defparam wb_smpl_data_i14.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i13 (.D(n2127), .CK(i_ref_clk_c), .CD(n9456), 
            .Q(wb_smpl_data[13]));   // d:/documents/git_local/fm_modulator/rtl/top.v(214[9] 222[10])
    defparam wb_smpl_data_i13.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i12 (.D(n2128), .CK(i_ref_clk_c), .CD(n9456), 
            .Q(wb_smpl_data[12]));   // d:/documents/git_local/fm_modulator/rtl/top.v(214[9] 222[10])
    defparam wb_smpl_data_i12.GSR = "DISABLED";
    dynamic_pll lo_gen (.i_clk_2f_N_2249(i_clk_2f_N_2249), .lo_pll_out(lo_pll_out), 
            .i_ref_clk_c(i_ref_clk_c), .pll_clk(pll_clk), .pll_rst(pll_rst), 
            .pll_stb(pll_stb), .pll_we(pll_we), .pll_data_i({pll_data_i}), 
            .pll_addr({pll_addr}), .pll_data_o({pll_data_o}), .pll_ack(pll_ack), 
            .GND_net(GND_net)) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(166[13] 177[5])
    FD1S3IX wb_smpl_data_i11 (.D(n2129), .CK(i_ref_clk_c), .CD(n9456), 
            .Q(wb_smpl_data[11]));   // d:/documents/git_local/fm_modulator/rtl/top.v(214[9] 222[10])
    defparam wb_smpl_data_i11.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i10 (.D(n24790), .CK(i_ref_clk_c), .CD(n9456), 
            .Q(wb_smpl_data[10]));   // d:/documents/git_local/fm_modulator/rtl/top.v(214[9] 222[10])
    defparam wb_smpl_data_i10.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i9 (.D(n24789), .CK(i_ref_clk_c), .CD(n9456), 
            .Q(wb_smpl_data[9]));   // d:/documents/git_local/fm_modulator/rtl/top.v(214[9] 222[10])
    defparam wb_smpl_data_i9.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i8 (.D(n2132), .CK(i_ref_clk_c), .CD(n9456), 
            .Q(wb_smpl_data[8]));   // d:/documents/git_local/fm_modulator/rtl/top.v(214[9] 222[10])
    defparam wb_smpl_data_i8.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i7 (.D(n2133), .CK(i_ref_clk_c), .CD(n9456), 
            .Q(wb_smpl_data[7]));   // d:/documents/git_local/fm_modulator/rtl/top.v(214[9] 222[10])
    defparam wb_smpl_data_i7.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i6 (.D(n2134), .CK(i_ref_clk_c), .CD(n9456), 
            .Q(wb_smpl_data[6]));   // d:/documents/git_local/fm_modulator/rtl/top.v(214[9] 222[10])
    defparam wb_smpl_data_i6.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i5 (.D(n24788), .CK(i_ref_clk_c), .CD(n9456), 
            .Q(wb_smpl_data[5]));   // d:/documents/git_local/fm_modulator/rtl/top.v(214[9] 222[10])
    defparam wb_smpl_data_i5.GSR = "DISABLED";
    \txuartlite(TIMING_BITS=24,CLOCKS_PER_BAUD=20)  txtransport (.i_ref_clk_c(i_ref_clk_c), 
            .i_ref_clk_c_enable_329(i_ref_clk_c_enable_329), .\lcl_data_7__N_511[0] (lcl_data_7__N_511[0]), 
            .zero_baud_counter_N_526(zero_baud_counter_N_526), .zero_baud_counter(zero_baud_counter), 
            .zero_baud_counter_N_525(zero_baud_counter_N_525), .o_wbu_uart_tx_c(o_wbu_uart_tx_c), 
            .n24992(n24992), .GND_net(GND_net), .\lcl_data[7] (lcl_data[7]), 
            .n27530(n27530), .\lcl_data[6] (lcl_data[6]), .\lcl_data_7__N_511[6] (lcl_data_7__N_511[6]), 
            .\lcl_data[5] (lcl_data[5]), .\lcl_data_7__N_511[5] (lcl_data_7__N_511[5]), 
            .\lcl_data[4] (lcl_data[4]), .\lcl_data_7__N_511[4] (lcl_data_7__N_511[4]), 
            .\lcl_data[3] (lcl_data[3]), .\lcl_data_7__N_511[3] (lcl_data_7__N_511[3]), 
            .\lcl_data[2] (lcl_data[2]), .\lcl_data_7__N_511[2] (lcl_data_7__N_511[2]), 
            .\lcl_data[1] (lcl_data[1]), .\lcl_data_7__N_511[1] (lcl_data_7__N_511[1]), 
            .n24890(n24890), .\state[0] (state_adj_3110[0]), .o_busy_N_536(o_busy_N_536), 
            .tx_busy(tx_busy), .n17568(n17568)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(63[55:112])
    FD1S3IX wb_smpl_data_i4 (.D(n2136), .CK(i_ref_clk_c), .CD(n9456), 
            .Q(wb_smpl_data[4]));   // d:/documents/git_local/fm_modulator/rtl/top.v(214[9] 222[10])
    defparam wb_smpl_data_i4.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module hbbus
//

module hbbus (i_ref_clk_c, wb_odata, n27585, wb_addr, wb_we, wb_stb, 
            n27530, GND_net, wb_err, wb_ack, \wb_idata[0] , \wb_idata[2] , 
            \wb_idata[3] , \wb_idata[4] , \wb_idata[5] , \wb_idata[6] , 
            \wb_idata[7] , \wb_idata[8] , \wb_idata[9] , \wb_idata[10] , 
            \wb_idata[11] , \wb_idata[12] , \wb_idata[13] , \wb_idata[14] , 
            \wb_idata[15] , \wb_idata[16] , \wb_idata[17] , \wb_idata[18] , 
            \wb_idata[19] , \wb_idata[20] , \wb_idata[21] , \wb_idata[22] , 
            \wb_idata[23] , \wb_idata[24] , \wb_idata[25] , \wb_idata[26] , 
            \wb_idata[27] , \wb_idata[28] , \wb_idata[29] , \wb_idata[30] , 
            \wb_idata[31] , n2, n12729, VCC_net, \rx_data[6] , \rx_data[0] , 
            \rx_data[5] , \rx_data[1] , \rx_data[2] , rx_stb, \rx_data[3] , 
            \rx_data[4] , tx_busy, n24992, \lcl_data[1] , \lcl_data_7__N_511[0] , 
            \lcl_data[2] , \lcl_data_7__N_511[1] , \lcl_data[3] , \lcl_data_7__N_511[2] , 
            \lcl_data[4] , \lcl_data_7__N_511[3] , \lcl_data[5] , \lcl_data_7__N_511[4] , 
            \lcl_data[6] , \lcl_data_7__N_511[5] , \lcl_data[7] , \lcl_data_7__N_511[6] , 
            n24890, zero_baud_counter_N_526, zero_baud_counter_N_525, 
            zero_baud_counter, i_ref_clk_c_enable_329, o_busy_N_536, \state[0] , 
            n17568) /* synthesis syn_module_defined=1 */ ;
    input i_ref_clk_c;
    output [31:0]wb_odata;
    output n27585;
    output [29:0]wb_addr;
    output wb_we;
    output wb_stb;
    input n27530;
    input GND_net;
    input wb_err;
    input wb_ack;
    input \wb_idata[0] ;
    input \wb_idata[2] ;
    input \wb_idata[3] ;
    input \wb_idata[4] ;
    input \wb_idata[5] ;
    input \wb_idata[6] ;
    input \wb_idata[7] ;
    input \wb_idata[8] ;
    input \wb_idata[9] ;
    input \wb_idata[10] ;
    input \wb_idata[11] ;
    input \wb_idata[12] ;
    input \wb_idata[13] ;
    input \wb_idata[14] ;
    input \wb_idata[15] ;
    input \wb_idata[16] ;
    input \wb_idata[17] ;
    input \wb_idata[18] ;
    input \wb_idata[19] ;
    input \wb_idata[20] ;
    input \wb_idata[21] ;
    input \wb_idata[22] ;
    input \wb_idata[23] ;
    input \wb_idata[24] ;
    input \wb_idata[25] ;
    input \wb_idata[26] ;
    input \wb_idata[27] ;
    input \wb_idata[28] ;
    input \wb_idata[29] ;
    input \wb_idata[30] ;
    input \wb_idata[31] ;
    output n2;
    input n12729;
    input VCC_net;
    input \rx_data[6] ;
    input \rx_data[0] ;
    input \rx_data[5] ;
    input \rx_data[1] ;
    input \rx_data[2] ;
    input rx_stb;
    input \rx_data[3] ;
    input \rx_data[4] ;
    input tx_busy;
    output n24992;
    input \lcl_data[1] ;
    output \lcl_data_7__N_511[0] ;
    input \lcl_data[2] ;
    output \lcl_data_7__N_511[1] ;
    input \lcl_data[3] ;
    output \lcl_data_7__N_511[2] ;
    input \lcl_data[4] ;
    output \lcl_data_7__N_511[3] ;
    input \lcl_data[5] ;
    output \lcl_data_7__N_511[4] ;
    input \lcl_data[6] ;
    output \lcl_data_7__N_511[5] ;
    input \lcl_data[7] ;
    output \lcl_data_7__N_511[6] ;
    input n24890;
    input zero_baud_counter_N_526;
    output zero_baud_counter_N_525;
    input zero_baud_counter;
    output i_ref_clk_c_enable_329;
    input o_busy_N_536;
    input \state[0] ;
    output n17568;
    
    wire i_ref_clk_c /* synthesis SET_AS_NETWORK=i_ref_clk_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(22[12:21])
    
    wire newaddr_N_990;
    wire [33:0]iw_word;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(71[14:21])
    
    wire ow_stb;
    wire [33:0]ow_word;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(73[14:21])
    
    wire n27587, n25103, i_cmd_wr, iw_stb, n27586, n25115, i_ref_clk_c_enable_315, 
        i_ref_clk_c_enable_194;
    wire [4:0]hb_bits;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(79[13:20])
    wire [33:0]idl_word;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(77[14:22])
    
    wire hb_busy, w_reset, n24991, idl_stb, nl_busy, hx_stb, i_ref_clk_c_enable_388;
    wire [4:0]dec_bits;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(69[13:21])
    
    wire o_pck_stb_N_765, cmd_loaded, i_ref_clk_c_enable_192, cmd_loaded_N_768, 
        i_ref_clk_c_enable_357;
    wire [33:0]n14;
    wire [7:0]w_gx_char;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbgenhex.v(80[12:21])
    
    wire n11767;
    wire [33:0]int_word;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(75[14:22])
    
    wire n25186, int_stb;
    
    hbexec wbexec (.i_ref_clk_c(i_ref_clk_c), .newaddr_N_990(newaddr_N_990), 
           .wb_odata({wb_odata}), .iw_word({iw_word}), .ow_stb(ow_stb), 
           .ow_word({ow_word}), .n27587(n27587), .n27585(n27585), .wb_addr({wb_addr}), 
           .n25103(n25103), .wb_we(wb_we), .i_cmd_wr(i_cmd_wr), .wb_stb(wb_stb), 
           .n27530(n27530), .iw_stb(iw_stb), .GND_net(GND_net), .wb_err(wb_err), 
           .n27586(n27586), .wb_ack(wb_ack), .\wb_idata[0] (\wb_idata[0] ), 
           .\wb_idata[2] (\wb_idata[2] ), .\wb_idata[3] (\wb_idata[3] ), 
           .\wb_idata[4] (\wb_idata[4] ), .\wb_idata[5] (\wb_idata[5] ), 
           .\wb_idata[6] (\wb_idata[6] ), .\wb_idata[7] (\wb_idata[7] ), 
           .\wb_idata[8] (\wb_idata[8] ), .\wb_idata[9] (\wb_idata[9] ), 
           .\wb_idata[10] (\wb_idata[10] ), .\wb_idata[11] (\wb_idata[11] ), 
           .\wb_idata[12] (\wb_idata[12] ), .\wb_idata[13] (\wb_idata[13] ), 
           .\wb_idata[14] (\wb_idata[14] ), .\wb_idata[15] (\wb_idata[15] ), 
           .\wb_idata[16] (\wb_idata[16] ), .\wb_idata[17] (\wb_idata[17] ), 
           .\wb_idata[18] (\wb_idata[18] ), .\wb_idata[19] (\wb_idata[19] ), 
           .\wb_idata[20] (\wb_idata[20] ), .\wb_idata[21] (\wb_idata[21] ), 
           .\wb_idata[22] (\wb_idata[22] ), .\wb_idata[23] (\wb_idata[23] ), 
           .\wb_idata[24] (\wb_idata[24] ), .\wb_idata[25] (\wb_idata[25] ), 
           .\wb_idata[26] (\wb_idata[26] ), .\wb_idata[27] (\wb_idata[27] ), 
           .\wb_idata[28] (\wb_idata[28] ), .\wb_idata[29] (\wb_idata[29] ), 
           .\wb_idata[30] (\wb_idata[30] ), .\wb_idata[31] (\wb_idata[31] ), 
           .n2(n2), .n25115(n25115), .n12729(n12729)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(105[15] 109[15])
    hbdeword unpackx (.i_ref_clk_c(i_ref_clk_c), .i_ref_clk_c_enable_315(i_ref_clk_c_enable_315), 
            .i_ref_clk_c_enable_194(i_ref_clk_c_enable_194), .n27587(n27587), 
            .hb_bits({hb_bits}), .idl_word({idl_word}), .n27530(n27530), 
            .hb_busy(hb_busy), .w_reset(w_reset), .n24991(n24991), .idl_stb(idl_stb), 
            .n27586(n27586), .nl_busy(nl_busy), .hx_stb(hx_stb)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(127[11] 129[29])
    hbpack packxi (.i_ref_clk_c(i_ref_clk_c), .i_ref_clk_c_enable_388(i_ref_clk_c_enable_388), 
           .n27587(n27587), .iw_word({iw_word}), .\dec_bits[4] (dec_bits[4]), 
           .iw_stb(iw_stb), .w_reset(w_reset), .o_pck_stb_N_765(o_pck_stb_N_765), 
           .cmd_loaded(cmd_loaded), .i_ref_clk_c_enable_192(i_ref_clk_c_enable_192), 
           .cmd_loaded_N_768(cmd_loaded_N_768), .\dec_bits[0] (dec_bits[0]), 
           .\dec_bits[1] (dec_bits[1]), .i_ref_clk_c_enable_357(i_ref_clk_c_enable_357), 
           .n45(n14[3]), .n46(n14[2]), .n25103(n25103), .n27586(n27586), 
           .newaddr_N_990(newaddr_N_990), .n25115(n25115), .i_cmd_wr(i_cmd_wr)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(99[9] 100[38])
    hbgenhex genhex (.hb_bits({hb_bits}), .\w_gx_char[0] (w_gx_char[0]), 
            .\w_gx_char[1] (w_gx_char[1]), .\w_gx_char[2] (w_gx_char[2]), 
            .\w_gx_char[3] (w_gx_char[3]), .\w_gx_char[4] (w_gx_char[4]), 
            .\w_gx_char[5] (w_gx_char[5]), .\w_gx_char[6] (w_gx_char[6]), 
            .i_ref_clk_c(i_ref_clk_c), .i_ref_clk_c_enable_315(i_ref_clk_c_enable_315), 
            .GND_net(GND_net), .VCC_net(VCC_net), .hx_stb(hx_stb), .w_reset(w_reset), 
            .hb_busy(hb_busy), .n11767(n11767), .nl_busy(nl_busy), .n27586(n27586), 
            .n24991(n24991), .i_ref_clk_c_enable_194(i_ref_clk_c_enable_194)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(132[11] 133[29])
    hbdechex dechxi (.\rx_data[6] (\rx_data[6] ), .i_ref_clk_c(i_ref_clk_c), 
            .dec_bits({dec_bits[4], Open_0, Open_1, Open_2, dec_bits[0]}), 
            .w_reset(w_reset), .n27586(n27586), .\rx_data[0] (\rx_data[0] ), 
            .\rx_data[5] (\rx_data[5] ), .\rx_data[1] (\rx_data[1] ), .\rx_data[2] (\rx_data[2] ), 
            .rx_stb(rx_stb), .\rx_data[3] (\rx_data[3] ), .\rx_data[4] (\rx_data[4] ), 
            .\dec_bits[1] (dec_bits[1]), .n45(n14[3]), .n46(n14[2]), .n27587(n27587), 
            .i_ref_clk_c_enable_388(i_ref_clk_c_enable_388), .i_ref_clk_c_enable_357(i_ref_clk_c_enable_357), 
            .cmd_loaded(cmd_loaded), .o_pck_stb_N_765(o_pck_stb_N_765), 
            .i_ref_clk_c_enable_192(i_ref_clk_c_enable_192), .cmd_loaded_N_768(cmd_loaded_N_768)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(93[11] 95[30])
    hbnewline addnl (.i_ref_clk_c(i_ref_clk_c), .n27587(n27587), .hx_stb(hx_stb), 
            .nl_busy(nl_busy), .\w_gx_char[1] (w_gx_char[1]), .w_reset(w_reset), 
            .n27586(n27586), .\w_gx_char[3] (w_gx_char[3]), .\w_gx_char[6] (w_gx_char[6]), 
            .\w_gx_char[5] (w_gx_char[5]), .n11767(n11767), .tx_busy(tx_busy), 
            .\w_gx_char[4] (w_gx_char[4]), .\w_gx_char[2] (w_gx_char[2]), 
            .\w_gx_char[0] (w_gx_char[0]), .n24992(n24992), .\lcl_data[1] (\lcl_data[1] ), 
            .\lcl_data_7__N_511[0] (\lcl_data_7__N_511[0] ), .\lcl_data[2] (\lcl_data[2] ), 
            .\lcl_data_7__N_511[1] (\lcl_data_7__N_511[1] ), .\lcl_data[3] (\lcl_data[3] ), 
            .\lcl_data_7__N_511[2] (\lcl_data_7__N_511[2] ), .\lcl_data[4] (\lcl_data[4] ), 
            .\lcl_data_7__N_511[3] (\lcl_data_7__N_511[3] ), .\lcl_data[5] (\lcl_data[5] ), 
            .\lcl_data_7__N_511[4] (\lcl_data_7__N_511[4] ), .\lcl_data[6] (\lcl_data[6] ), 
            .\lcl_data_7__N_511[5] (\lcl_data_7__N_511[5] ), .\lcl_data[7] (\lcl_data[7] ), 
            .\lcl_data_7__N_511[6] (\lcl_data_7__N_511[6] ), .n24890(n24890), 
            .zero_baud_counter_N_526(zero_baud_counter_N_526), .zero_baud_counter_N_525(zero_baud_counter_N_525), 
            .zero_baud_counter(zero_baud_counter), .i_ref_clk_c_enable_329(i_ref_clk_c_enable_329), 
            .o_busy_N_536(o_busy_N_536), .\state[0] (\state[0] ), .n17568(n17568)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(138[12] 139[40])
    hbints addints (.int_word({int_word}), .i_ref_clk_c(i_ref_clk_c), .ow_word({ow_word}), 
           .n27586(n27586), .n25186(n25186), .int_stb(int_stb), .n27587(n27587), 
           .ow_stb(ow_stb)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(114[9] 116[32])
    hbidle addidles (.idl_word({idl_word}), .i_ref_clk_c(i_ref_clk_c), .int_word({int_word}), 
           .hb_busy(hb_busy), .int_stb(int_stb), .idl_stb(idl_stb), .n25186(n25186), 
           .n27586(n27586), .n27587(n27587)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(121[9] 123[31])
    
endmodule
//
// Verilog Description of module hbexec
//

module hbexec (i_ref_clk_c, newaddr_N_990, wb_odata, iw_word, ow_stb, 
            ow_word, n27587, n27585, wb_addr, n25103, wb_we, i_cmd_wr, 
            wb_stb, n27530, iw_stb, GND_net, wb_err, n27586, wb_ack, 
            \wb_idata[0] , \wb_idata[2] , \wb_idata[3] , \wb_idata[4] , 
            \wb_idata[5] , \wb_idata[6] , \wb_idata[7] , \wb_idata[8] , 
            \wb_idata[9] , \wb_idata[10] , \wb_idata[11] , \wb_idata[12] , 
            \wb_idata[13] , \wb_idata[14] , \wb_idata[15] , \wb_idata[16] , 
            \wb_idata[17] , \wb_idata[18] , \wb_idata[19] , \wb_idata[20] , 
            \wb_idata[21] , \wb_idata[22] , \wb_idata[23] , \wb_idata[24] , 
            \wb_idata[25] , \wb_idata[26] , \wb_idata[27] , \wb_idata[28] , 
            \wb_idata[29] , \wb_idata[30] , \wb_idata[31] , n2, n25115, 
            n12729) /* synthesis syn_module_defined=1 */ ;
    input i_ref_clk_c;
    input newaddr_N_990;
    output [31:0]wb_odata;
    input [33:0]iw_word;
    output ow_stb;
    output [33:0]ow_word;
    input n27587;
    output n27585;
    output [29:0]wb_addr;
    input n25103;
    output wb_we;
    input i_cmd_wr;
    output wb_stb;
    input n27530;
    input iw_stb;
    input GND_net;
    input wb_err;
    input n27586;
    input wb_ack;
    input \wb_idata[0] ;
    input \wb_idata[2] ;
    input \wb_idata[3] ;
    input \wb_idata[4] ;
    input \wb_idata[5] ;
    input \wb_idata[6] ;
    input \wb_idata[7] ;
    input \wb_idata[8] ;
    input \wb_idata[9] ;
    input \wb_idata[10] ;
    input \wb_idata[11] ;
    input \wb_idata[12] ;
    input \wb_idata[13] ;
    input \wb_idata[14] ;
    input \wb_idata[15] ;
    input \wb_idata[16] ;
    input \wb_idata[17] ;
    input \wb_idata[18] ;
    input \wb_idata[19] ;
    input \wb_idata[20] ;
    input \wb_idata[21] ;
    input \wb_idata[22] ;
    input \wb_idata[23] ;
    input \wb_idata[24] ;
    input \wb_idata[25] ;
    input \wb_idata[26] ;
    input \wb_idata[27] ;
    input \wb_idata[28] ;
    input \wb_idata[29] ;
    input \wb_idata[30] ;
    input \wb_idata[31] ;
    output n2;
    input n25115;
    input n12729;
    
    wire i_ref_clk_c /* synthesis SET_AS_NETWORK=i_ref_clk_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(22[12:21])
    
    wire newaddr, wb_cyc, n8953, o_rsp_stb_N_987;
    wire [33:0]n338;
    wire [33:0]o_rsp_word_33__N_951;
    
    wire i_ref_clk_c_enable_146, n17131, inc, i_ref_clk_c_enable_145, 
        i_cmd_word_0__N_995, i_ref_clk_c_enable_150, n19489, n17127, 
        i_ref_clk_c_enable_449, n17182, n17436, n17125;
    wire [29:0]n125;
    
    wire n17435, n17129, n17434, n17135, n17133, n17433, n17139, 
        n17137, n17432, n17143, n17141, n17431, n17147, n17145, 
        n17430, n17151, n17149, n17429, n17155, n17153, n17428, 
        n17159, n17157, n17427, n17163, n17161, n17426, n17167, 
        n17165, n17425, n17171, n17169, n17424, n17175, n17173, 
        n17423, n17179, n17177, n17422, n17181, i_ref_clk_c_enable_417, 
        o_cmd_busy_N_941, o_cmd_busy_N_933;
    wire [32:0]n2227;
    
    wire n17813;
    
    FD1S3IX newaddr_72 (.D(newaddr_N_990), .CK(i_ref_clk_c), .CD(wb_cyc), 
            .Q(newaddr)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(192[9] 236[5])
    defparam newaddr_72.GSR = "DISABLED";
    FD1S3AX o_wb_data_i0 (.D(iw_word[0]), .CK(i_ref_clk_c), .Q(wb_odata[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i0.GSR = "DISABLED";
    FD1S3JX o_rsp_stb_74 (.D(o_rsp_stb_N_987), .CK(i_ref_clk_c), .PD(n8953), 
            .Q(ow_stb)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_stb_74.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i0 (.D(n338[0]), .CK(i_ref_clk_c), .CD(n8953), 
            .Q(ow_word[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i0.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i2 (.D(n338[2]), .CK(i_ref_clk_c), .CD(n8953), 
            .Q(ow_word[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i2.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i3 (.D(n338[3]), .CK(i_ref_clk_c), .CD(n8953), 
            .Q(ow_word[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i3.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i4 (.D(n338[4]), .CK(i_ref_clk_c), .CD(n8953), 
            .Q(ow_word[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i4.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i5 (.D(n338[5]), .CK(i_ref_clk_c), .CD(n8953), 
            .Q(ow_word[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i5.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i6 (.D(n338[6]), .CK(i_ref_clk_c), .CD(n8953), 
            .Q(ow_word[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i6.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i7 (.D(n338[7]), .CK(i_ref_clk_c), .CD(n8953), 
            .Q(ow_word[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i7.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i8 (.D(n338[8]), .CK(i_ref_clk_c), .CD(n8953), 
            .Q(ow_word[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i8.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i9 (.D(n338[9]), .CK(i_ref_clk_c), .CD(n8953), 
            .Q(ow_word[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i9.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i10 (.D(n338[10]), .CK(i_ref_clk_c), .CD(n8953), 
            .Q(ow_word[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i10.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i11 (.D(n338[11]), .CK(i_ref_clk_c), .CD(n8953), 
            .Q(ow_word[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i11.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i12 (.D(n338[12]), .CK(i_ref_clk_c), .CD(n8953), 
            .Q(ow_word[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i12.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i13 (.D(n338[13]), .CK(i_ref_clk_c), .CD(n8953), 
            .Q(ow_word[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i13.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i14 (.D(n338[14]), .CK(i_ref_clk_c), .CD(n8953), 
            .Q(ow_word[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i14.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i15 (.D(n338[15]), .CK(i_ref_clk_c), .CD(n8953), 
            .Q(ow_word[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i15.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i16 (.D(n338[16]), .CK(i_ref_clk_c), .CD(n8953), 
            .Q(ow_word[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i16.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i17 (.D(n338[17]), .CK(i_ref_clk_c), .CD(n8953), 
            .Q(ow_word[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i17.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i18 (.D(n338[18]), .CK(i_ref_clk_c), .CD(n8953), 
            .Q(ow_word[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i18.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i19 (.D(n338[19]), .CK(i_ref_clk_c), .CD(n8953), 
            .Q(ow_word[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i19.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i20 (.D(n338[20]), .CK(i_ref_clk_c), .CD(n8953), 
            .Q(ow_word[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i20.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i21 (.D(n338[21]), .CK(i_ref_clk_c), .CD(n8953), 
            .Q(ow_word[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i21.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i22 (.D(n338[22]), .CK(i_ref_clk_c), .CD(n8953), 
            .Q(ow_word[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i22.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i23 (.D(n338[23]), .CK(i_ref_clk_c), .CD(n8953), 
            .Q(ow_word[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i23.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i24 (.D(n338[24]), .CK(i_ref_clk_c), .CD(n8953), 
            .Q(ow_word[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i24.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i25 (.D(n338[25]), .CK(i_ref_clk_c), .CD(n8953), 
            .Q(ow_word[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i25.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i26 (.D(n338[26]), .CK(i_ref_clk_c), .CD(n8953), 
            .Q(ow_word[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i26.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i27 (.D(n338[27]), .CK(i_ref_clk_c), .CD(n8953), 
            .Q(ow_word[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i27.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i28 (.D(n338[28]), .CK(i_ref_clk_c), .CD(n8953), 
            .Q(ow_word[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i28.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i29 (.D(o_rsp_word_33__N_951[29]), .CK(i_ref_clk_c), 
            .CD(n27587), .Q(ow_word[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i29.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i30 (.D(n338[30]), .CK(i_ref_clk_c), .CD(n8953), 
            .Q(ow_word[30])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i30.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i31 (.D(n338[31]), .CK(i_ref_clk_c), .CD(n8953), 
            .Q(ow_word[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i31.GSR = "DISABLED";
    FD1S3JX o_rsp_word_i32 (.D(n338[32]), .CK(i_ref_clk_c), .PD(n8953), 
            .Q(ow_word[32])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i32.GSR = "DISABLED";
    FD1S3JX o_rsp_word_i33 (.D(i_ref_clk_c_enable_146), .CK(i_ref_clk_c), 
            .PD(n8953), .Q(ow_word[33])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i33.GSR = "DISABLED";
    LUT4 o_cmd_busy_I_0_1_lut_rep_595 (.A(n27585), .Z(i_ref_clk_c_enable_146)) /* synthesis lut_function=(!(A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(194[21:34])
    defparam o_cmd_busy_I_0_1_lut_rep_595.init = 16'h5555;
    LUT4 i15304_2_lut_3_lut_4_lut_4_lut (.A(n27585), .B(iw_word[1]), .C(wb_addr[26]), 
         .D(n25103), .Z(n17131)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(194[21:34])
    defparam i15304_2_lut_3_lut_4_lut_4_lut.init = 16'he0f0;
    FD1P3AX inc_71 (.D(i_cmd_word_0__N_995), .SP(i_ref_clk_c_enable_145), 
            .CK(i_ref_clk_c), .Q(inc)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(192[9] 236[5])
    defparam inc_71.GSR = "DISABLED";
    FD1P3AX o_wb_we_69 (.D(i_cmd_wr), .SP(i_ref_clk_c_enable_146), .CK(i_ref_clk_c), 
            .Q(wb_we)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(184[9] 186[26])
    defparam o_wb_we_69.GSR = "DISABLED";
    FD1P3IX o_wb_stb_68 (.D(n27530), .SP(i_ref_clk_c_enable_150), .CD(n19489), 
            .CK(i_ref_clk_c), .Q(wb_stb)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(121[9] 168[5])
    defparam o_wb_stb_68.GSR = "DISABLED";
    LUT4 i15309_2_lut_3_lut_4_lut_4_lut (.A(n27585), .B(iw_word[1]), .C(wb_addr[28]), 
         .D(n25103), .Z(n17127)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(194[21:34])
    defparam i15309_2_lut_3_lut_4_lut_4_lut.init = 16'he0f0;
    LUT4 i1_2_lut_3_lut_3_lut (.A(n27585), .B(iw_word[33]), .C(iw_stb), 
         .Z(i_ref_clk_c_enable_150)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(194[21:34])
    defparam i1_2_lut_3_lut_3_lut.init = 16'h1010;
    LUT4 i10924_2_lut_3_lut_3_lut (.A(n27585), .B(wb_stb), .C(n25103), 
         .Z(i_ref_clk_c_enable_449)) /* synthesis lut_function=(A (B)+!A (B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(194[21:34])
    defparam i10924_2_lut_3_lut_3_lut.init = 16'hdcdc;
    LUT4 i15256_3_lut_4_lut_4_lut (.A(n27585), .B(inc), .C(iw_word[2]), 
         .D(n25103), .Z(n17182)) /* synthesis lut_function=(A (B)+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(194[21:34])
    defparam i15256_3_lut_4_lut_4_lut.init = 16'hd8cc;
    CCU2D o_wb_addr_506_add_4_31 (.A0(n17127), .B0(iw_word[1]), .C0(i_ref_clk_c_enable_145), 
          .D0(iw_word[30]), .A1(n17125), .B1(iw_word[1]), .C1(i_ref_clk_c_enable_145), 
          .D1(iw_word[31]), .CIN(n17436), .S0(n125[28]), .S1(n125[29]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_506_add_4_31.INIT0 = 16'h5aaa;
    defparam o_wb_addr_506_add_4_31.INIT1 = 16'h5aaa;
    defparam o_wb_addr_506_add_4_31.INJECT1_0 = "NO";
    defparam o_wb_addr_506_add_4_31.INJECT1_1 = "NO";
    CCU2D o_wb_addr_506_add_4_29 (.A0(n17131), .B0(iw_word[1]), .C0(i_ref_clk_c_enable_145), 
          .D0(iw_word[28]), .A1(n17129), .B1(iw_word[1]), .C1(i_ref_clk_c_enable_145), 
          .D1(iw_word[29]), .CIN(n17435), .COUT(n17436), .S0(n125[26]), 
          .S1(n125[27]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_506_add_4_29.INIT0 = 16'h5aaa;
    defparam o_wb_addr_506_add_4_29.INIT1 = 16'h5aaa;
    defparam o_wb_addr_506_add_4_29.INJECT1_0 = "NO";
    defparam o_wb_addr_506_add_4_29.INJECT1_1 = "NO";
    CCU2D o_wb_addr_506_add_4_27 (.A0(n17135), .B0(iw_word[1]), .C0(i_ref_clk_c_enable_145), 
          .D0(iw_word[26]), .A1(n17133), .B1(iw_word[1]), .C1(i_ref_clk_c_enable_145), 
          .D1(iw_word[27]), .CIN(n17434), .COUT(n17435), .S0(n125[24]), 
          .S1(n125[25]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_506_add_4_27.INIT0 = 16'h5aaa;
    defparam o_wb_addr_506_add_4_27.INIT1 = 16'h5aaa;
    defparam o_wb_addr_506_add_4_27.INJECT1_0 = "NO";
    defparam o_wb_addr_506_add_4_27.INJECT1_1 = "NO";
    CCU2D o_wb_addr_506_add_4_25 (.A0(n17139), .B0(iw_word[1]), .C0(i_ref_clk_c_enable_145), 
          .D0(iw_word[24]), .A1(n17137), .B1(iw_word[1]), .C1(i_ref_clk_c_enable_145), 
          .D1(iw_word[25]), .CIN(n17433), .COUT(n17434), .S0(n125[22]), 
          .S1(n125[23]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_506_add_4_25.INIT0 = 16'h5aaa;
    defparam o_wb_addr_506_add_4_25.INIT1 = 16'h5aaa;
    defparam o_wb_addr_506_add_4_25.INJECT1_0 = "NO";
    defparam o_wb_addr_506_add_4_25.INJECT1_1 = "NO";
    CCU2D o_wb_addr_506_add_4_23 (.A0(n17143), .B0(iw_word[1]), .C0(i_ref_clk_c_enable_145), 
          .D0(iw_word[22]), .A1(n17141), .B1(iw_word[1]), .C1(i_ref_clk_c_enable_145), 
          .D1(iw_word[23]), .CIN(n17432), .COUT(n17433), .S0(n125[20]), 
          .S1(n125[21]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_506_add_4_23.INIT0 = 16'h5aaa;
    defparam o_wb_addr_506_add_4_23.INIT1 = 16'h5aaa;
    defparam o_wb_addr_506_add_4_23.INJECT1_0 = "NO";
    defparam o_wb_addr_506_add_4_23.INJECT1_1 = "NO";
    CCU2D o_wb_addr_506_add_4_21 (.A0(n17147), .B0(iw_word[1]), .C0(i_ref_clk_c_enable_145), 
          .D0(iw_word[20]), .A1(n17145), .B1(iw_word[1]), .C1(i_ref_clk_c_enable_145), 
          .D1(iw_word[21]), .CIN(n17431), .COUT(n17432), .S0(n125[18]), 
          .S1(n125[19]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_506_add_4_21.INIT0 = 16'h5aaa;
    defparam o_wb_addr_506_add_4_21.INIT1 = 16'h5aaa;
    defparam o_wb_addr_506_add_4_21.INJECT1_0 = "NO";
    defparam o_wb_addr_506_add_4_21.INJECT1_1 = "NO";
    CCU2D o_wb_addr_506_add_4_19 (.A0(n17151), .B0(iw_word[1]), .C0(i_ref_clk_c_enable_145), 
          .D0(iw_word[18]), .A1(n17149), .B1(iw_word[1]), .C1(i_ref_clk_c_enable_145), 
          .D1(iw_word[19]), .CIN(n17430), .COUT(n17431), .S0(n125[16]), 
          .S1(n125[17]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_506_add_4_19.INIT0 = 16'h5aaa;
    defparam o_wb_addr_506_add_4_19.INIT1 = 16'h5aaa;
    defparam o_wb_addr_506_add_4_19.INJECT1_0 = "NO";
    defparam o_wb_addr_506_add_4_19.INJECT1_1 = "NO";
    CCU2D o_wb_addr_506_add_4_17 (.A0(n17155), .B0(iw_word[1]), .C0(i_ref_clk_c_enable_145), 
          .D0(iw_word[16]), .A1(n17153), .B1(iw_word[1]), .C1(i_ref_clk_c_enable_145), 
          .D1(iw_word[17]), .CIN(n17429), .COUT(n17430), .S0(n125[14]), 
          .S1(n125[15]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_506_add_4_17.INIT0 = 16'h5aaa;
    defparam o_wb_addr_506_add_4_17.INIT1 = 16'h5aaa;
    defparam o_wb_addr_506_add_4_17.INJECT1_0 = "NO";
    defparam o_wb_addr_506_add_4_17.INJECT1_1 = "NO";
    CCU2D o_wb_addr_506_add_4_15 (.A0(n17159), .B0(iw_word[1]), .C0(i_ref_clk_c_enable_145), 
          .D0(iw_word[14]), .A1(n17157), .B1(iw_word[1]), .C1(i_ref_clk_c_enable_145), 
          .D1(iw_word[15]), .CIN(n17428), .COUT(n17429), .S0(n125[12]), 
          .S1(n125[13]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_506_add_4_15.INIT0 = 16'h5aaa;
    defparam o_wb_addr_506_add_4_15.INIT1 = 16'h5aaa;
    defparam o_wb_addr_506_add_4_15.INJECT1_0 = "NO";
    defparam o_wb_addr_506_add_4_15.INJECT1_1 = "NO";
    CCU2D o_wb_addr_506_add_4_13 (.A0(n17163), .B0(iw_word[1]), .C0(i_ref_clk_c_enable_145), 
          .D0(iw_word[12]), .A1(n17161), .B1(iw_word[1]), .C1(i_ref_clk_c_enable_145), 
          .D1(iw_word[13]), .CIN(n17427), .COUT(n17428), .S0(n125[10]), 
          .S1(n125[11]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_506_add_4_13.INIT0 = 16'h5aaa;
    defparam o_wb_addr_506_add_4_13.INIT1 = 16'h5aaa;
    defparam o_wb_addr_506_add_4_13.INJECT1_0 = "NO";
    defparam o_wb_addr_506_add_4_13.INJECT1_1 = "NO";
    LUT4 i15308_2_lut_3_lut_4_lut_4_lut (.A(n27585), .B(iw_word[1]), .C(wb_addr[27]), 
         .D(n25103), .Z(n17129)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(194[21:34])
    defparam i15308_2_lut_3_lut_4_lut_4_lut.init = 16'he0f0;
    CCU2D o_wb_addr_506_add_4_11 (.A0(n17167), .B0(iw_word[1]), .C0(i_ref_clk_c_enable_145), 
          .D0(iw_word[10]), .A1(n17165), .B1(iw_word[1]), .C1(i_ref_clk_c_enable_145), 
          .D1(iw_word[11]), .CIN(n17426), .COUT(n17427), .S0(n125[8]), 
          .S1(n125[9]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_506_add_4_11.INIT0 = 16'h5aaa;
    defparam o_wb_addr_506_add_4_11.INIT1 = 16'h5aaa;
    defparam o_wb_addr_506_add_4_11.INJECT1_0 = "NO";
    defparam o_wb_addr_506_add_4_11.INJECT1_1 = "NO";
    CCU2D o_wb_addr_506_add_4_9 (.A0(n17171), .B0(iw_word[1]), .C0(i_ref_clk_c_enable_145), 
          .D0(iw_word[8]), .A1(n17169), .B1(iw_word[1]), .C1(i_ref_clk_c_enable_145), 
          .D1(iw_word[9]), .CIN(n17425), .COUT(n17426), .S0(n125[6]), 
          .S1(n125[7]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_506_add_4_9.INIT0 = 16'h5aaa;
    defparam o_wb_addr_506_add_4_9.INIT1 = 16'h5aaa;
    defparam o_wb_addr_506_add_4_9.INJECT1_0 = "NO";
    defparam o_wb_addr_506_add_4_9.INJECT1_1 = "NO";
    LUT4 i15310_2_lut_3_lut_4_lut_4_lut (.A(n27585), .B(iw_word[1]), .C(wb_addr[29]), 
         .D(n25103), .Z(n17125)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(194[21:34])
    defparam i15310_2_lut_3_lut_4_lut_4_lut.init = 16'he0f0;
    CCU2D o_wb_addr_506_add_4_7 (.A0(n17175), .B0(iw_word[1]), .C0(i_ref_clk_c_enable_145), 
          .D0(iw_word[6]), .A1(n17173), .B1(iw_word[1]), .C1(i_ref_clk_c_enable_145), 
          .D1(iw_word[7]), .CIN(n17424), .COUT(n17425), .S0(n125[4]), 
          .S1(n125[5]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_506_add_4_7.INIT0 = 16'h5aaa;
    defparam o_wb_addr_506_add_4_7.INIT1 = 16'h5aaa;
    defparam o_wb_addr_506_add_4_7.INJECT1_0 = "NO";
    defparam o_wb_addr_506_add_4_7.INJECT1_1 = "NO";
    CCU2D o_wb_addr_506_add_4_5 (.A0(n17179), .B0(iw_word[1]), .C0(i_ref_clk_c_enable_145), 
          .D0(iw_word[4]), .A1(n17177), .B1(iw_word[1]), .C1(i_ref_clk_c_enable_145), 
          .D1(iw_word[5]), .CIN(n17423), .COUT(n17424), .S0(n125[2]), 
          .S1(n125[3]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_506_add_4_5.INIT0 = 16'h5aaa;
    defparam o_wb_addr_506_add_4_5.INIT1 = 16'h5aaa;
    defparam o_wb_addr_506_add_4_5.INJECT1_0 = "NO";
    defparam o_wb_addr_506_add_4_5.INJECT1_1 = "NO";
    CCU2D o_wb_addr_506_add_4_3 (.A0(n17182), .B0(i_ref_clk_c_enable_145), 
          .C0(iw_word[1]), .D0(wb_addr[0]), .A1(n17181), .B1(iw_word[1]), 
          .C1(i_ref_clk_c_enable_145), .D1(iw_word[3]), .CIN(n17422), 
          .COUT(n17423), .S0(n125[0]), .S1(n125[1]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_506_add_4_3.INIT0 = 16'h59aa;
    defparam o_wb_addr_506_add_4_3.INIT1 = 16'h5aaa;
    defparam o_wb_addr_506_add_4_3.INJECT1_0 = "NO";
    defparam o_wb_addr_506_add_4_3.INJECT1_1 = "NO";
    CCU2D o_wb_addr_506_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(iw_word[1]), .B1(i_ref_clk_c_enable_145), 
          .C1(GND_net), .D1(GND_net), .COUT(n17422));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_506_add_4_1.INIT0 = 16'hF000;
    defparam o_wb_addr_506_add_4_1.INIT1 = 16'hffff;
    defparam o_wb_addr_506_add_4_1.INJECT1_0 = "NO";
    defparam o_wb_addr_506_add_4_1.INJECT1_1 = "NO";
    LUT4 i15302_2_lut_3_lut_4_lut_4_lut (.A(n27585), .B(iw_word[1]), .C(wb_addr[24]), 
         .D(n25103), .Z(n17135)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(194[21:34])
    defparam i15302_2_lut_3_lut_4_lut_4_lut.init = 16'he0f0;
    LUT4 i15303_2_lut_3_lut_4_lut_4_lut (.A(n27585), .B(iw_word[1]), .C(wb_addr[25]), 
         .D(n25103), .Z(n17133)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(194[21:34])
    defparam i15303_2_lut_3_lut_4_lut_4_lut.init = 16'he0f0;
    LUT4 i15246_2_lut_3_lut_4_lut_4_lut (.A(n27585), .B(iw_word[1]), .C(wb_addr[22]), 
         .D(n25103), .Z(n17139)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(194[21:34])
    defparam i15246_2_lut_3_lut_4_lut_4_lut.init = 16'he0f0;
    FD1S3AX o_wb_data_i31 (.D(iw_word[31]), .CK(i_ref_clk_c), .Q(wb_odata[31])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i31.GSR = "DISABLED";
    LUT4 i15295_2_lut_3_lut_4_lut_4_lut (.A(n27585), .B(iw_word[1]), .C(wb_addr[23]), 
         .D(n25103), .Z(n17137)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(194[21:34])
    defparam i15295_2_lut_3_lut_4_lut_4_lut.init = 16'he0f0;
    FD1P3IX o_wb_cyc_67_rep_687 (.D(o_cmd_busy_N_933), .SP(i_ref_clk_c_enable_417), 
            .CD(o_cmd_busy_N_941), .CK(i_ref_clk_c), .Q(n27585)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(121[9] 168[5])
    defparam o_wb_cyc_67_rep_687.GSR = "DISABLED";
    LUT4 i15260_2_lut_3_lut_4_lut_4_lut (.A(n27585), .B(iw_word[1]), .C(wb_addr[20]), 
         .D(n25103), .Z(n17143)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(194[21:34])
    defparam i15260_2_lut_3_lut_4_lut_4_lut.init = 16'he0f0;
    FD1S3AX o_wb_data_i30 (.D(iw_word[30]), .CK(i_ref_clk_c), .Q(wb_odata[30])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i30.GSR = "DISABLED";
    FD1S3AX o_wb_data_i29 (.D(iw_word[29]), .CK(i_ref_clk_c), .Q(wb_odata[29])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i29.GSR = "DISABLED";
    FD1S3AX o_wb_data_i28 (.D(iw_word[28]), .CK(i_ref_clk_c), .Q(wb_odata[28])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i28.GSR = "DISABLED";
    FD1S3AX o_wb_data_i27 (.D(iw_word[27]), .CK(i_ref_clk_c), .Q(wb_odata[27])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i27.GSR = "DISABLED";
    FD1S3AX o_wb_data_i26 (.D(iw_word[26]), .CK(i_ref_clk_c), .Q(wb_odata[26])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i26.GSR = "DISABLED";
    FD1S3AX o_wb_data_i25 (.D(iw_word[25]), .CK(i_ref_clk_c), .Q(wb_odata[25])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i25.GSR = "DISABLED";
    FD1S3AX o_wb_data_i24 (.D(iw_word[24]), .CK(i_ref_clk_c), .Q(wb_odata[24])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i24.GSR = "DISABLED";
    FD1S3AX o_wb_data_i23 (.D(iw_word[23]), .CK(i_ref_clk_c), .Q(wb_odata[23])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i23.GSR = "DISABLED";
    FD1S3AX o_wb_data_i22 (.D(iw_word[22]), .CK(i_ref_clk_c), .Q(wb_odata[22])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i22.GSR = "DISABLED";
    FD1S3AX o_wb_data_i21 (.D(iw_word[21]), .CK(i_ref_clk_c), .Q(wb_odata[21])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i21.GSR = "DISABLED";
    FD1S3AX o_wb_data_i20 (.D(iw_word[20]), .CK(i_ref_clk_c), .Q(wb_odata[20])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i20.GSR = "DISABLED";
    FD1S3AX o_wb_data_i19 (.D(iw_word[19]), .CK(i_ref_clk_c), .Q(wb_odata[19])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i19.GSR = "DISABLED";
    FD1S3AX o_wb_data_i18 (.D(iw_word[18]), .CK(i_ref_clk_c), .Q(wb_odata[18])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i18.GSR = "DISABLED";
    LUT4 i15307_2_lut_3_lut_4_lut_4_lut (.A(n27585), .B(iw_word[1]), .C(wb_addr[21]), 
         .D(n25103), .Z(n17141)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(194[21:34])
    defparam i15307_2_lut_3_lut_4_lut_4_lut.init = 16'he0f0;
    FD1S3AX o_wb_data_i17 (.D(iw_word[17]), .CK(i_ref_clk_c), .Q(wb_odata[17])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i17.GSR = "DISABLED";
    LUT4 i15248_2_lut_3_lut_4_lut_4_lut (.A(n27585), .B(iw_word[1]), .C(wb_addr[18]), 
         .D(n25103), .Z(n17147)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(194[21:34])
    defparam i15248_2_lut_3_lut_4_lut_4_lut.init = 16'he0f0;
    FD1S3AX o_wb_data_i16 (.D(iw_word[16]), .CK(i_ref_clk_c), .Q(wb_odata[16])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i16.GSR = "DISABLED";
    FD1S3AX o_wb_data_i15 (.D(iw_word[15]), .CK(i_ref_clk_c), .Q(wb_odata[15])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i15.GSR = "DISABLED";
    FD1S3AX o_wb_data_i14 (.D(iw_word[14]), .CK(i_ref_clk_c), .Q(wb_odata[14])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i14.GSR = "DISABLED";
    FD1S3AX o_wb_data_i13 (.D(iw_word[13]), .CK(i_ref_clk_c), .Q(wb_odata[13])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i13.GSR = "DISABLED";
    FD1S3AX o_wb_data_i12 (.D(iw_word[12]), .CK(i_ref_clk_c), .Q(wb_odata[12])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i12.GSR = "DISABLED";
    FD1S3AX o_wb_data_i11 (.D(iw_word[11]), .CK(i_ref_clk_c), .Q(wb_odata[11])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i11.GSR = "DISABLED";
    FD1S3AX o_wb_data_i10 (.D(iw_word[10]), .CK(i_ref_clk_c), .Q(wb_odata[10])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i10.GSR = "DISABLED";
    FD1S3AX o_wb_data_i9 (.D(iw_word[9]), .CK(i_ref_clk_c), .Q(wb_odata[9])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i9.GSR = "DISABLED";
    FD1S3AX o_wb_data_i8 (.D(iw_word[8]), .CK(i_ref_clk_c), .Q(wb_odata[8])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i8.GSR = "DISABLED";
    FD1S3AX o_wb_data_i7 (.D(iw_word[7]), .CK(i_ref_clk_c), .Q(wb_odata[7])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i7.GSR = "DISABLED";
    FD1S3AX o_wb_data_i6 (.D(iw_word[6]), .CK(i_ref_clk_c), .Q(wb_odata[6])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i6.GSR = "DISABLED";
    FD1S3AX o_wb_data_i5 (.D(iw_word[5]), .CK(i_ref_clk_c), .Q(wb_odata[5])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i5.GSR = "DISABLED";
    FD1S3AX o_wb_data_i4 (.D(iw_word[4]), .CK(i_ref_clk_c), .Q(wb_odata[4])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i4.GSR = "DISABLED";
    FD1S3AX o_wb_data_i3 (.D(iw_word[3]), .CK(i_ref_clk_c), .Q(wb_odata[3])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i3.GSR = "DISABLED";
    FD1S3AX o_wb_data_i2 (.D(iw_word[2]), .CK(i_ref_clk_c), .Q(wb_odata[2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i2.GSR = "DISABLED";
    FD1S3AX o_wb_data_i1 (.D(iw_word[1]), .CK(i_ref_clk_c), .Q(wb_odata[1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i1.GSR = "DISABLED";
    LUT4 i6450_2_lut (.A(wb_err), .B(n27586), .Z(n8953)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(283[11] 309[5])
    defparam i6450_2_lut.init = 16'heeee;
    LUT4 newaddr_I_0_3_lut (.A(newaddr), .B(wb_ack), .C(n27585), .Z(o_rsp_stb_N_987)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam newaddr_I_0_3_lut.init = 16'hcaca;
    LUT4 mux_59_i1_4_lut (.A(inc), .B(\wb_idata[0] ), .C(n27585), .D(wb_we), 
         .Z(n338[0])) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A (B (C (D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i1_4_lut.init = 16'h05c5;
    LUT4 mux_59_i3_4_lut (.A(wb_addr[0]), .B(\wb_idata[2] ), .C(n27585), 
         .D(wb_we), .Z(n338[2])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i3_4_lut.init = 16'h0aca;
    LUT4 mux_59_i4_4_lut (.A(wb_addr[1]), .B(\wb_idata[3] ), .C(n27585), 
         .D(wb_we), .Z(n338[3])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i4_4_lut.init = 16'h0aca;
    LUT4 mux_59_i5_4_lut (.A(wb_addr[2]), .B(\wb_idata[4] ), .C(n27585), 
         .D(wb_we), .Z(n338[4])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i5_4_lut.init = 16'h0aca;
    LUT4 mux_59_i6_4_lut (.A(wb_addr[3]), .B(\wb_idata[5] ), .C(n27585), 
         .D(wb_we), .Z(n338[5])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i6_4_lut.init = 16'h0aca;
    LUT4 mux_59_i7_4_lut (.A(wb_addr[4]), .B(\wb_idata[6] ), .C(n27585), 
         .D(wb_we), .Z(n338[6])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i7_4_lut.init = 16'h0aca;
    LUT4 mux_59_i8_4_lut (.A(wb_addr[5]), .B(\wb_idata[7] ), .C(n27585), 
         .D(wb_we), .Z(n338[7])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i8_4_lut.init = 16'h0aca;
    LUT4 mux_59_i9_4_lut (.A(wb_addr[6]), .B(\wb_idata[8] ), .C(n27585), 
         .D(wb_we), .Z(n338[8])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i9_4_lut.init = 16'h0aca;
    LUT4 mux_59_i10_4_lut (.A(wb_addr[7]), .B(\wb_idata[9] ), .C(n27585), 
         .D(wb_we), .Z(n338[9])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i10_4_lut.init = 16'h0aca;
    LUT4 mux_59_i11_4_lut (.A(wb_addr[8]), .B(\wb_idata[10] ), .C(n27585), 
         .D(wb_we), .Z(n338[10])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i11_4_lut.init = 16'h0aca;
    LUT4 mux_59_i12_4_lut (.A(wb_addr[9]), .B(\wb_idata[11] ), .C(n27585), 
         .D(wb_we), .Z(n338[11])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i12_4_lut.init = 16'h0aca;
    LUT4 mux_59_i13_4_lut (.A(wb_addr[10]), .B(\wb_idata[12] ), .C(n27585), 
         .D(wb_we), .Z(n338[12])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i13_4_lut.init = 16'h0aca;
    LUT4 mux_59_i14_4_lut (.A(wb_addr[11]), .B(\wb_idata[13] ), .C(n27585), 
         .D(wb_we), .Z(n338[13])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i14_4_lut.init = 16'h0aca;
    LUT4 mux_59_i15_4_lut (.A(wb_addr[12]), .B(\wb_idata[14] ), .C(n27585), 
         .D(wb_we), .Z(n338[14])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i15_4_lut.init = 16'h0aca;
    LUT4 mux_59_i16_4_lut (.A(wb_addr[13]), .B(\wb_idata[15] ), .C(n27585), 
         .D(wb_we), .Z(n338[15])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i16_4_lut.init = 16'h0aca;
    LUT4 mux_59_i17_4_lut (.A(wb_addr[14]), .B(\wb_idata[16] ), .C(n27585), 
         .D(wb_we), .Z(n338[16])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i17_4_lut.init = 16'h0aca;
    LUT4 mux_59_i18_4_lut (.A(wb_addr[15]), .B(\wb_idata[17] ), .C(n27585), 
         .D(wb_we), .Z(n338[17])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i18_4_lut.init = 16'h0aca;
    LUT4 mux_59_i19_4_lut (.A(wb_addr[16]), .B(\wb_idata[18] ), .C(n27585), 
         .D(wb_we), .Z(n338[18])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i19_4_lut.init = 16'h0aca;
    LUT4 mux_59_i20_4_lut (.A(wb_addr[17]), .B(\wb_idata[19] ), .C(n27585), 
         .D(wb_we), .Z(n338[19])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i20_4_lut.init = 16'h0aca;
    LUT4 mux_59_i21_4_lut (.A(wb_addr[18]), .B(\wb_idata[20] ), .C(n27585), 
         .D(wb_we), .Z(n338[20])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i21_4_lut.init = 16'h0aca;
    LUT4 mux_59_i22_4_lut (.A(wb_addr[19]), .B(\wb_idata[21] ), .C(n27585), 
         .D(wb_we), .Z(n338[21])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i22_4_lut.init = 16'h0aca;
    LUT4 mux_59_i23_4_lut (.A(wb_addr[20]), .B(\wb_idata[22] ), .C(n27585), 
         .D(wb_we), .Z(n338[22])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i23_4_lut.init = 16'h0aca;
    LUT4 mux_59_i24_4_lut (.A(wb_addr[21]), .B(\wb_idata[23] ), .C(n27585), 
         .D(wb_we), .Z(n338[23])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i24_4_lut.init = 16'h0aca;
    LUT4 mux_59_i25_4_lut (.A(wb_addr[22]), .B(\wb_idata[24] ), .C(n27585), 
         .D(wb_we), .Z(n338[24])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i25_4_lut.init = 16'h0aca;
    LUT4 mux_59_i26_4_lut (.A(wb_addr[23]), .B(\wb_idata[25] ), .C(n27585), 
         .D(wb_we), .Z(n338[25])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i26_4_lut.init = 16'h0aca;
    LUT4 mux_59_i27_4_lut (.A(wb_addr[24]), .B(\wb_idata[26] ), .C(n27585), 
         .D(wb_we), .Z(n338[26])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i27_4_lut.init = 16'h0aca;
    LUT4 mux_59_i28_4_lut (.A(wb_addr[25]), .B(\wb_idata[27] ), .C(n27585), 
         .D(wb_we), .Z(n338[27])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i28_4_lut.init = 16'h0aca;
    LUT4 mux_59_i29_4_lut (.A(wb_addr[26]), .B(\wb_idata[28] ), .C(n27585), 
         .D(wb_we), .Z(n338[28])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i29_4_lut.init = 16'h0aca;
    LUT4 i11277_4_lut (.A(wb_addr[27]), .B(wb_err), .C(n2227[29]), .D(n27585), 
         .Z(o_rsp_word_33__N_951[29])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(287[11] 309[5])
    defparam i11277_4_lut.init = 16'hfcee;
    LUT4 i11344_2_lut (.A(\wb_idata[29] ), .B(wb_we), .Z(n2227[29])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(299[4:47])
    defparam i11344_2_lut.init = 16'h2222;
    LUT4 mux_59_i31_4_lut (.A(wb_addr[28]), .B(\wb_idata[30] ), .C(n27585), 
         .D(wb_we), .Z(n338[30])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i31_4_lut.init = 16'h0aca;
    LUT4 mux_59_i32_4_lut (.A(wb_addr[29]), .B(\wb_idata[31] ), .C(n27585), 
         .D(wb_we), .Z(n338[31])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i32_4_lut.init = 16'h0aca;
    LUT4 i11278_2_lut (.A(wb_we), .B(n27585), .Z(n338[32])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam i11278_2_lut.init = 16'h8888;
    FD1P3AX o_wb_addr_506__i0 (.D(n125[0]), .SP(i_ref_clk_c_enable_449), 
            .CK(i_ref_clk_c), .Q(wb_addr[0])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_506__i0.GSR = "DISABLED";
    LUT4 i2_1_lut (.A(wb_stb), .Z(n2)) /* synthesis lut_function=(!(A)) */ ;
    defparam i2_1_lut.init = 16'h5555;
    LUT4 i_cmd_word_0__I_0_1_lut (.A(iw_word[0]), .Z(i_cmd_word_0__N_995)) /* synthesis lut_function=(!(A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(214[11:25])
    defparam i_cmd_word_0__I_0_1_lut.init = 16'h5555;
    LUT4 i15252_2_lut_3_lut_4_lut_4_lut (.A(n27585), .B(iw_word[1]), .C(wb_addr[19]), 
         .D(n25103), .Z(n17145)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(194[21:34])
    defparam i15252_2_lut_3_lut_4_lut_4_lut.init = 16'he0f0;
    LUT4 i15263_2_lut_3_lut_4_lut_4_lut (.A(n27585), .B(iw_word[1]), .C(wb_addr[16]), 
         .D(n25103), .Z(n17151)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(194[21:34])
    defparam i15263_2_lut_3_lut_4_lut_4_lut.init = 16'he0f0;
    LUT4 i15271_2_lut_3_lut_4_lut_4_lut (.A(n27585), .B(iw_word[1]), .C(wb_addr[17]), 
         .D(n25103), .Z(n17149)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(194[21:34])
    defparam i15271_2_lut_3_lut_4_lut_4_lut.init = 16'he0f0;
    LUT4 i15254_2_lut_3_lut_4_lut_4_lut (.A(n27585), .B(iw_word[1]), .C(wb_addr[14]), 
         .D(n25103), .Z(n17155)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(194[21:34])
    defparam i15254_2_lut_3_lut_4_lut_4_lut.init = 16'he0f0;
    LUT4 i15262_2_lut_3_lut_4_lut_4_lut (.A(n27585), .B(iw_word[1]), .C(wb_addr[15]), 
         .D(n25103), .Z(n17153)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(194[21:34])
    defparam i15262_2_lut_3_lut_4_lut_4_lut.init = 16'he0f0;
    LUT4 i15251_2_lut_3_lut_4_lut_4_lut (.A(n27585), .B(iw_word[1]), .C(wb_addr[12]), 
         .D(n25103), .Z(n17159)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(194[21:34])
    defparam i15251_2_lut_3_lut_4_lut_4_lut.init = 16'he0f0;
    LUT4 i15253_2_lut_3_lut_4_lut_4_lut (.A(n27585), .B(iw_word[1]), .C(wb_addr[13]), 
         .D(n25103), .Z(n17157)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(194[21:34])
    defparam i15253_2_lut_3_lut_4_lut_4_lut.init = 16'he0f0;
    LUT4 i15249_2_lut_3_lut_4_lut_4_lut (.A(n27585), .B(iw_word[1]), .C(wb_addr[10]), 
         .D(n25103), .Z(n17163)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(194[21:34])
    defparam i15249_2_lut_3_lut_4_lut_4_lut.init = 16'he0f0;
    LUT4 i15250_2_lut_3_lut_4_lut_4_lut (.A(n27585), .B(iw_word[1]), .C(wb_addr[11]), 
         .D(n25103), .Z(n17161)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(194[21:34])
    defparam i15250_2_lut_3_lut_4_lut_4_lut.init = 16'he0f0;
    LUT4 i3_4_lut (.A(wb_we), .B(n27585), .C(n27586), .D(wb_err), .Z(n17813)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i3_4_lut.init = 16'h0004;
    LUT4 i1_4_lut (.A(n25115), .B(o_cmd_busy_N_941), .C(wb_ack), .D(o_cmd_busy_N_933), 
         .Z(i_ref_clk_c_enable_417)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+!((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(122[6:41])
    defparam i1_4_lut.init = 16'heefc;
    LUT4 i21059_2_lut (.A(n27585), .B(wb_stb), .Z(o_cmd_busy_N_933)) /* synthesis lut_function=(!(A+(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(149[11] 168[5])
    defparam i21059_2_lut.init = 16'h1111;
    LUT4 i15306_2_lut_3_lut_4_lut_4_lut (.A(n27585), .B(iw_word[1]), .C(wb_addr[8]), 
         .D(n25103), .Z(n17167)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(194[21:34])
    defparam i15306_2_lut_3_lut_4_lut_4_lut.init = 16'he0f0;
    LUT4 i15247_2_lut_3_lut_4_lut_4_lut (.A(n27585), .B(iw_word[1]), .C(wb_addr[9]), 
         .D(n25103), .Z(n17165)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(194[21:34])
    defparam i15247_2_lut_3_lut_4_lut_4_lut.init = 16'he0f0;
    LUT4 i15278_2_lut_3_lut_4_lut_4_lut (.A(n27585), .B(iw_word[1]), .C(wb_addr[6]), 
         .D(n25103), .Z(n17171)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(194[21:34])
    defparam i15278_2_lut_3_lut_4_lut_4_lut.init = 16'he0f0;
    LUT4 i15294_2_lut_3_lut_4_lut_4_lut (.A(n27585), .B(iw_word[1]), .C(wb_addr[7]), 
         .D(n25103), .Z(n17169)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(194[21:34])
    defparam i15294_2_lut_3_lut_4_lut_4_lut.init = 16'he0f0;
    LUT4 i15261_2_lut_3_lut_4_lut_4_lut (.A(n27585), .B(iw_word[1]), .C(wb_addr[4]), 
         .D(n25103), .Z(n17175)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(194[21:34])
    defparam i15261_2_lut_3_lut_4_lut_4_lut.init = 16'he0f0;
    LUT4 i15264_2_lut_3_lut_4_lut_4_lut (.A(n27585), .B(iw_word[1]), .C(wb_addr[5]), 
         .D(n25103), .Z(n17173)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(194[21:34])
    defparam i15264_2_lut_3_lut_4_lut_4_lut.init = 16'he0f0;
    LUT4 i15258_2_lut_3_lut_4_lut_4_lut (.A(n27585), .B(iw_word[1]), .C(wb_addr[2]), 
         .D(n25103), .Z(n17179)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(194[21:34])
    defparam i15258_2_lut_3_lut_4_lut_4_lut.init = 16'he0f0;
    LUT4 i15259_2_lut_3_lut_4_lut_4_lut (.A(n27585), .B(iw_word[1]), .C(wb_addr[3]), 
         .D(n25103), .Z(n17177)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(194[21:34])
    defparam i15259_2_lut_3_lut_4_lut_4_lut.init = 16'he0f0;
    LUT4 i15257_2_lut_3_lut_4_lut_4_lut (.A(n27585), .B(iw_word[1]), .C(wb_addr[1]), 
         .D(n25103), .Z(n17181)) /* synthesis lut_function=(A (C)+!A (B (C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(194[21:34])
    defparam i15257_2_lut_3_lut_4_lut_4_lut.init = 16'he0f0;
    LUT4 i1_2_lut_rep_406_4_lut_4_lut (.A(n27585), .B(iw_stb), .C(iw_word[33]), 
         .D(iw_word[32]), .Z(i_ref_clk_c_enable_145)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(194[21:34])
    defparam i1_2_lut_rep_406_4_lut_4_lut.init = 16'h0040;
    FD1S3IX o_rsp_word_i1 (.D(n17813), .CK(i_ref_clk_c), .CD(n12729), 
            .Q(ow_word[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i1.GSR = "DISABLED";
    LUT4 i1_2_lut_3_lut_4_lut (.A(wb_err), .B(n27585), .C(wb_stb), .D(n27586), 
         .Z(n19489)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(122[17:41])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfff8;
    LUT4 i1_2_lut_rep_404_3_lut (.A(wb_err), .B(n27585), .C(n27586), .Z(o_cmd_busy_N_941)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(122[17:41])
    defparam i1_2_lut_rep_404_3_lut.init = 16'hf8f8;
    FD1P3IX o_wb_cyc_67 (.D(o_cmd_busy_N_933), .SP(i_ref_clk_c_enable_417), 
            .CD(o_cmd_busy_N_941), .CK(i_ref_clk_c), .Q(wb_cyc)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(121[9] 168[5])
    defparam o_wb_cyc_67.GSR = "DISABLED";
    FD1P3AX o_wb_addr_506__i29 (.D(n125[29]), .SP(i_ref_clk_c_enable_449), 
            .CK(i_ref_clk_c), .Q(wb_addr[29])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_506__i29.GSR = "DISABLED";
    FD1P3AX o_wb_addr_506__i28 (.D(n125[28]), .SP(i_ref_clk_c_enable_449), 
            .CK(i_ref_clk_c), .Q(wb_addr[28])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_506__i28.GSR = "DISABLED";
    FD1P3AX o_wb_addr_506__i27 (.D(n125[27]), .SP(i_ref_clk_c_enable_449), 
            .CK(i_ref_clk_c), .Q(wb_addr[27])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_506__i27.GSR = "DISABLED";
    FD1P3AX o_wb_addr_506__i26 (.D(n125[26]), .SP(i_ref_clk_c_enable_449), 
            .CK(i_ref_clk_c), .Q(wb_addr[26])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_506__i26.GSR = "DISABLED";
    FD1P3AX o_wb_addr_506__i25 (.D(n125[25]), .SP(i_ref_clk_c_enable_449), 
            .CK(i_ref_clk_c), .Q(wb_addr[25])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_506__i25.GSR = "DISABLED";
    FD1P3AX o_wb_addr_506__i24 (.D(n125[24]), .SP(i_ref_clk_c_enable_449), 
            .CK(i_ref_clk_c), .Q(wb_addr[24])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_506__i24.GSR = "DISABLED";
    FD1P3AX o_wb_addr_506__i23 (.D(n125[23]), .SP(i_ref_clk_c_enable_449), 
            .CK(i_ref_clk_c), .Q(wb_addr[23])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_506__i23.GSR = "DISABLED";
    FD1P3AX o_wb_addr_506__i22 (.D(n125[22]), .SP(i_ref_clk_c_enable_449), 
            .CK(i_ref_clk_c), .Q(wb_addr[22])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_506__i22.GSR = "DISABLED";
    FD1P3AX o_wb_addr_506__i21 (.D(n125[21]), .SP(i_ref_clk_c_enable_449), 
            .CK(i_ref_clk_c), .Q(wb_addr[21])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_506__i21.GSR = "DISABLED";
    FD1P3AX o_wb_addr_506__i20 (.D(n125[20]), .SP(i_ref_clk_c_enable_449), 
            .CK(i_ref_clk_c), .Q(wb_addr[20])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_506__i20.GSR = "DISABLED";
    FD1P3AX o_wb_addr_506__i19 (.D(n125[19]), .SP(i_ref_clk_c_enable_449), 
            .CK(i_ref_clk_c), .Q(wb_addr[19])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_506__i19.GSR = "DISABLED";
    FD1P3AX o_wb_addr_506__i18 (.D(n125[18]), .SP(i_ref_clk_c_enable_449), 
            .CK(i_ref_clk_c), .Q(wb_addr[18])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_506__i18.GSR = "DISABLED";
    FD1P3AX o_wb_addr_506__i17 (.D(n125[17]), .SP(i_ref_clk_c_enable_449), 
            .CK(i_ref_clk_c), .Q(wb_addr[17])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_506__i17.GSR = "DISABLED";
    FD1P3AX o_wb_addr_506__i16 (.D(n125[16]), .SP(i_ref_clk_c_enable_449), 
            .CK(i_ref_clk_c), .Q(wb_addr[16])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_506__i16.GSR = "DISABLED";
    FD1P3AX o_wb_addr_506__i15 (.D(n125[15]), .SP(i_ref_clk_c_enable_449), 
            .CK(i_ref_clk_c), .Q(wb_addr[15])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_506__i15.GSR = "DISABLED";
    FD1P3AX o_wb_addr_506__i14 (.D(n125[14]), .SP(i_ref_clk_c_enable_449), 
            .CK(i_ref_clk_c), .Q(wb_addr[14])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_506__i14.GSR = "DISABLED";
    FD1P3AX o_wb_addr_506__i13 (.D(n125[13]), .SP(i_ref_clk_c_enable_449), 
            .CK(i_ref_clk_c), .Q(wb_addr[13])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_506__i13.GSR = "DISABLED";
    FD1P3AX o_wb_addr_506__i12 (.D(n125[12]), .SP(i_ref_clk_c_enable_449), 
            .CK(i_ref_clk_c), .Q(wb_addr[12])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_506__i12.GSR = "DISABLED";
    FD1P3AX o_wb_addr_506__i11 (.D(n125[11]), .SP(i_ref_clk_c_enable_449), 
            .CK(i_ref_clk_c), .Q(wb_addr[11])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_506__i11.GSR = "DISABLED";
    FD1P3AX o_wb_addr_506__i10 (.D(n125[10]), .SP(i_ref_clk_c_enable_449), 
            .CK(i_ref_clk_c), .Q(wb_addr[10])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_506__i10.GSR = "DISABLED";
    FD1P3AX o_wb_addr_506__i9 (.D(n125[9]), .SP(i_ref_clk_c_enable_449), 
            .CK(i_ref_clk_c), .Q(wb_addr[9])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_506__i9.GSR = "DISABLED";
    FD1P3AX o_wb_addr_506__i8 (.D(n125[8]), .SP(i_ref_clk_c_enable_449), 
            .CK(i_ref_clk_c), .Q(wb_addr[8])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_506__i8.GSR = "DISABLED";
    FD1P3AX o_wb_addr_506__i7 (.D(n125[7]), .SP(i_ref_clk_c_enable_449), 
            .CK(i_ref_clk_c), .Q(wb_addr[7])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_506__i7.GSR = "DISABLED";
    FD1P3AX o_wb_addr_506__i6 (.D(n125[6]), .SP(i_ref_clk_c_enable_449), 
            .CK(i_ref_clk_c), .Q(wb_addr[6])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_506__i6.GSR = "DISABLED";
    FD1P3AX o_wb_addr_506__i5 (.D(n125[5]), .SP(i_ref_clk_c_enable_449), 
            .CK(i_ref_clk_c), .Q(wb_addr[5])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_506__i5.GSR = "DISABLED";
    FD1P3AX o_wb_addr_506__i4 (.D(n125[4]), .SP(i_ref_clk_c_enable_449), 
            .CK(i_ref_clk_c), .Q(wb_addr[4])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_506__i4.GSR = "DISABLED";
    FD1P3AX o_wb_addr_506__i3 (.D(n125[3]), .SP(i_ref_clk_c_enable_449), 
            .CK(i_ref_clk_c), .Q(wb_addr[3])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_506__i3.GSR = "DISABLED";
    FD1P3AX o_wb_addr_506__i2 (.D(n125[2]), .SP(i_ref_clk_c_enable_449), 
            .CK(i_ref_clk_c), .Q(wb_addr[2])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_506__i2.GSR = "DISABLED";
    FD1P3AX o_wb_addr_506__i1 (.D(n125[1]), .SP(i_ref_clk_c_enable_449), 
            .CK(i_ref_clk_c), .Q(wb_addr[1])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_506__i1.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module hbdeword
//

module hbdeword (i_ref_clk_c, i_ref_clk_c_enable_315, i_ref_clk_c_enable_194, 
            n27587, hb_bits, idl_word, n27530, hb_busy, w_reset, 
            n24991, idl_stb, n27586, nl_busy, hx_stb) /* synthesis syn_module_defined=1 */ ;
    input i_ref_clk_c;
    input i_ref_clk_c_enable_315;
    input i_ref_clk_c_enable_194;
    input n27587;
    output [4:0]hb_bits;
    input [33:0]idl_word;
    input n27530;
    output hb_busy;
    input w_reset;
    output n24991;
    input idl_stb;
    input n27586;
    input nl_busy;
    input hx_stb;
    
    wire i_ref_clk_c /* synthesis SET_AS_NETWORK=i_ref_clk_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(22[12:21])
    wire [3:0]r_len;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(58[12:17])
    
    wire n10137;
    wire [3:0]n13;
    wire [3:0]r_len_3__N_1229;
    
    wire i_ref_clk_c_enable_242;
    wire [4:0]o_dw_bits_4__N_1188;
    wire [31:0]r_word;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(59[13:19])
    
    wire n12801;
    wire [31:0]r_word_31__N_1197;
    
    wire o_dw_busy_N_1269;
    wire [4:0]o_dw_bits_4__N_1279;
    
    wire n6, n11575, n11577, n24180, n24674, n24993;
    
    FD1P3IX r_len__i0 (.D(n13[0]), .SP(i_ref_clk_c_enable_315), .CD(n10137), 
            .CK(i_ref_clk_c), .Q(r_len[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(64[9] 81[6])
    defparam r_len__i0.GSR = "DISABLED";
    FD1P3IX r_len__i3 (.D(r_len_3__N_1229[3]), .SP(i_ref_clk_c_enable_194), 
            .CD(n27587), .CK(i_ref_clk_c), .Q(r_len[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(64[9] 81[6])
    defparam r_len__i3.GSR = "DISABLED";
    FD1P3AX o_dw_bits_i0 (.D(o_dw_bits_4__N_1188[0]), .SP(i_ref_clk_c_enable_242), 
            .CK(i_ref_clk_c), .Q(hb_bits[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(95[9] 103[41])
    defparam o_dw_bits_i0.GSR = "DISABLED";
    FD1P3IX r_word_i1 (.D(idl_word[1]), .SP(i_ref_clk_c_enable_242), .CD(n12801), 
            .CK(i_ref_clk_c), .Q(r_word[1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i1.GSR = "DISABLED";
    FD1P3IX r_word_i2 (.D(idl_word[2]), .SP(i_ref_clk_c_enable_242), .CD(n12801), 
            .CK(i_ref_clk_c), .Q(r_word[2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i2.GSR = "DISABLED";
    FD1P3IX r_word_i3 (.D(idl_word[3]), .SP(i_ref_clk_c_enable_242), .CD(n12801), 
            .CK(i_ref_clk_c), .Q(r_word[3])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i3.GSR = "DISABLED";
    FD1P3IX o_dw_bits_i4 (.D(n27530), .SP(i_ref_clk_c_enable_242), .CD(n12801), 
            .CK(i_ref_clk_c), .Q(hb_bits[4])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(95[9] 103[41])
    defparam o_dw_bits_i4.GSR = "DISABLED";
    FD1P3AX o_dw_bits_i3 (.D(o_dw_bits_4__N_1188[3]), .SP(i_ref_clk_c_enable_242), 
            .CK(i_ref_clk_c), .Q(hb_bits[3])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(95[9] 103[41])
    defparam o_dw_bits_i3.GSR = "DISABLED";
    FD1P3AX o_dw_bits_i2 (.D(o_dw_bits_4__N_1188[2]), .SP(i_ref_clk_c_enable_242), 
            .CK(i_ref_clk_c), .Q(hb_bits[2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(95[9] 103[41])
    defparam o_dw_bits_i2.GSR = "DISABLED";
    FD1P3AX o_dw_bits_i1 (.D(o_dw_bits_4__N_1188[1]), .SP(i_ref_clk_c_enable_242), 
            .CK(i_ref_clk_c), .Q(hb_bits[1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(95[9] 103[41])
    defparam o_dw_bits_i1.GSR = "DISABLED";
    FD1P3AX r_word_i31 (.D(r_word_31__N_1197[31]), .SP(i_ref_clk_c_enable_242), 
            .CK(i_ref_clk_c), .Q(r_word[31])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i31.GSR = "DISABLED";
    FD1P3IX o_dw_stb_36 (.D(o_dw_busy_N_1269), .SP(i_ref_clk_c_enable_194), 
            .CD(w_reset), .CK(i_ref_clk_c), .Q(hb_busy)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(64[9] 81[6])
    defparam o_dw_stb_36.GSR = "DISABLED";
    FD1P3IX r_word_i0 (.D(idl_word[0]), .SP(i_ref_clk_c_enable_242), .CD(n12801), 
            .CK(i_ref_clk_c), .Q(r_word[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i0.GSR = "DISABLED";
    FD1P3AX r_word_i30 (.D(r_word_31__N_1197[30]), .SP(i_ref_clk_c_enable_242), 
            .CK(i_ref_clk_c), .Q(r_word[30])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i30.GSR = "DISABLED";
    FD1P3AX r_word_i29 (.D(r_word_31__N_1197[29]), .SP(i_ref_clk_c_enable_242), 
            .CK(i_ref_clk_c), .Q(r_word[29])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i29.GSR = "DISABLED";
    FD1P3AX r_word_i28 (.D(r_word_31__N_1197[28]), .SP(i_ref_clk_c_enable_242), 
            .CK(i_ref_clk_c), .Q(r_word[28])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i28.GSR = "DISABLED";
    FD1P3AX r_word_i27 (.D(r_word_31__N_1197[27]), .SP(i_ref_clk_c_enable_242), 
            .CK(i_ref_clk_c), .Q(r_word[27])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i27.GSR = "DISABLED";
    FD1P3AX r_word_i26 (.D(r_word_31__N_1197[26]), .SP(i_ref_clk_c_enable_242), 
            .CK(i_ref_clk_c), .Q(r_word[26])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i26.GSR = "DISABLED";
    FD1P3AX r_word_i25 (.D(r_word_31__N_1197[25]), .SP(i_ref_clk_c_enable_242), 
            .CK(i_ref_clk_c), .Q(r_word[25])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i25.GSR = "DISABLED";
    FD1P3AX r_word_i24 (.D(r_word_31__N_1197[24]), .SP(i_ref_clk_c_enable_242), 
            .CK(i_ref_clk_c), .Q(r_word[24])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i24.GSR = "DISABLED";
    FD1P3AX r_word_i23 (.D(r_word_31__N_1197[23]), .SP(i_ref_clk_c_enable_242), 
            .CK(i_ref_clk_c), .Q(r_word[23])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i23.GSR = "DISABLED";
    FD1P3AX r_word_i22 (.D(r_word_31__N_1197[22]), .SP(i_ref_clk_c_enable_242), 
            .CK(i_ref_clk_c), .Q(r_word[22])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i22.GSR = "DISABLED";
    FD1P3AX r_word_i21 (.D(r_word_31__N_1197[21]), .SP(i_ref_clk_c_enable_242), 
            .CK(i_ref_clk_c), .Q(r_word[21])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i21.GSR = "DISABLED";
    FD1P3AX r_word_i20 (.D(r_word_31__N_1197[20]), .SP(i_ref_clk_c_enable_242), 
            .CK(i_ref_clk_c), .Q(r_word[20])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i20.GSR = "DISABLED";
    FD1P3AX r_word_i19 (.D(r_word_31__N_1197[19]), .SP(i_ref_clk_c_enable_242), 
            .CK(i_ref_clk_c), .Q(r_word[19])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i19.GSR = "DISABLED";
    FD1P3AX r_word_i18 (.D(r_word_31__N_1197[18]), .SP(i_ref_clk_c_enable_242), 
            .CK(i_ref_clk_c), .Q(r_word[18])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i18.GSR = "DISABLED";
    FD1P3AX r_word_i17 (.D(r_word_31__N_1197[17]), .SP(i_ref_clk_c_enable_242), 
            .CK(i_ref_clk_c), .Q(r_word[17])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i17.GSR = "DISABLED";
    FD1P3AX r_word_i16 (.D(r_word_31__N_1197[16]), .SP(i_ref_clk_c_enable_242), 
            .CK(i_ref_clk_c), .Q(r_word[16])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i16.GSR = "DISABLED";
    FD1P3AX r_word_i15 (.D(r_word_31__N_1197[15]), .SP(i_ref_clk_c_enable_242), 
            .CK(i_ref_clk_c), .Q(r_word[15])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i15.GSR = "DISABLED";
    FD1P3AX r_word_i14 (.D(r_word_31__N_1197[14]), .SP(i_ref_clk_c_enable_242), 
            .CK(i_ref_clk_c), .Q(r_word[14])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i14.GSR = "DISABLED";
    FD1P3AX r_word_i13 (.D(r_word_31__N_1197[13]), .SP(i_ref_clk_c_enable_242), 
            .CK(i_ref_clk_c), .Q(r_word[13])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i13.GSR = "DISABLED";
    FD1P3AX r_word_i12 (.D(r_word_31__N_1197[12]), .SP(i_ref_clk_c_enable_242), 
            .CK(i_ref_clk_c), .Q(r_word[12])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i12.GSR = "DISABLED";
    FD1P3AX r_word_i11 (.D(r_word_31__N_1197[11]), .SP(i_ref_clk_c_enable_242), 
            .CK(i_ref_clk_c), .Q(r_word[11])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i11.GSR = "DISABLED";
    FD1P3AX r_word_i10 (.D(r_word_31__N_1197[10]), .SP(i_ref_clk_c_enable_242), 
            .CK(i_ref_clk_c), .Q(r_word[10])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i10.GSR = "DISABLED";
    FD1P3AX r_word_i9 (.D(r_word_31__N_1197[9]), .SP(i_ref_clk_c_enable_242), 
            .CK(i_ref_clk_c), .Q(r_word[9])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i9.GSR = "DISABLED";
    FD1P3AX r_word_i8 (.D(r_word_31__N_1197[8]), .SP(i_ref_clk_c_enable_242), 
            .CK(i_ref_clk_c), .Q(r_word[8])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i8.GSR = "DISABLED";
    FD1P3AX r_word_i7 (.D(r_word_31__N_1197[7]), .SP(i_ref_clk_c_enable_242), 
            .CK(i_ref_clk_c), .Q(r_word[7])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i7.GSR = "DISABLED";
    FD1P3AX r_word_i6 (.D(r_word_31__N_1197[6]), .SP(i_ref_clk_c_enable_242), 
            .CK(i_ref_clk_c), .Q(r_word[6])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i6.GSR = "DISABLED";
    FD1P3AX r_word_i5 (.D(r_word_31__N_1197[5]), .SP(i_ref_clk_c_enable_242), 
            .CK(i_ref_clk_c), .Q(r_word[5])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i5.GSR = "DISABLED";
    FD1P3AX r_word_i4 (.D(r_word_31__N_1197[4]), .SP(i_ref_clk_c_enable_242), 
            .CK(i_ref_clk_c), .Q(r_word[4])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i4.GSR = "DISABLED";
    LUT4 mux_15_i4_4_lut (.A(r_len[3]), .B(o_dw_bits_4__N_1279[3]), .C(n24991), 
         .D(n6), .Z(r_len_3__N_1229[3])) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(76[12] 81[6])
    defparam mux_15_i4_4_lut.init = 16'h3a35;
    LUT4 i10936_2_lut (.A(idl_word[32]), .B(idl_word[33]), .Z(o_dw_bits_4__N_1279[3])) /* synthesis lut_function=(A (B)) */ ;
    defparam i10936_2_lut.init = 16'h8888;
    FD1P3IX r_len__i2 (.D(n11575), .SP(i_ref_clk_c_enable_315), .CD(n10137), 
            .CK(i_ref_clk_c), .Q(r_len[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(64[9] 81[6])
    defparam r_len__i2.GSR = "DISABLED";
    FD1P3IX r_len__i1 (.D(n11577), .SP(i_ref_clk_c_enable_315), .CD(n10137), 
            .CK(i_ref_clk_c), .Q(r_len[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(64[9] 81[6])
    defparam r_len__i1.GSR = "DISABLED";
    LUT4 o_dw_bits_4__I_0_i3_4_lut (.A(r_word[30]), .B(idl_word[31]), .C(n24991), 
         .D(o_dw_bits_4__N_1279[3]), .Z(o_dw_bits_4__N_1188[2])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(102[12] 103[41])
    defparam o_dw_bits_4__I_0_i3_4_lut.init = 16'hca0a;
    LUT4 r_word_29__bdd_3_lut_22544 (.A(idl_word[30]), .B(idl_word[33]), 
         .C(idl_word[32]), .Z(n24180)) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam r_word_29__bdd_3_lut_22544.init = 16'h8c8c;
    LUT4 r_word_28__bdd_3_lut_22914 (.A(idl_word[29]), .B(idl_word[32]), 
         .C(idl_word[33]), .Z(n24674)) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam r_word_28__bdd_3_lut_22914.init = 16'h8c8c;
    LUT4 i_stb_I_0_2_lut_rep_431 (.A(idl_stb), .B(hb_busy), .Z(n24991)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam i_stb_I_0_2_lut_rep_431.init = 16'h2222;
    LUT4 o_dw_bits_4__I_0_i4_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(o_dw_bits_4__N_1279[3]), 
         .D(r_word[31]), .Z(o_dw_bits_4__N_1188[3])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam o_dw_bits_4__I_0_i4_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_29__bdd_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(n24180), 
         .D(r_word[29]), .Z(o_dw_bits_4__N_1188[1])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_29__bdd_3_lut_4_lut.init = 16'hfd20;
    LUT4 i7634_2_lut_3_lut (.A(idl_stb), .B(hb_busy), .C(n27586), .Z(n10137)) /* synthesis lut_function=(A ((C)+!B)+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam i7634_2_lut_3_lut.init = 16'hf2f2;
    LUT4 i1_2_lut_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(nl_busy), 
         .D(hx_stb), .Z(i_ref_clk_c_enable_242)) /* synthesis lut_function=(!(A (B (C (D)))+!A (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h2fff;
    LUT4 i21072_2_lut_3_lut_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(hx_stb), 
         .D(nl_busy), .Z(n12801)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam i21072_2_lut_3_lut_3_lut_4_lut.init = 16'h0ddd;
    LUT4 r_word_31__I_0_i32_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[31]), 
         .D(r_word[27]), .Z(r_word_31__N_1197[31])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i32_3_lut_4_lut.init = 16'hfd20;
    LUT4 i10944_2_lut_3_lut (.A(idl_stb), .B(hb_busy), .C(n24993), .Z(o_dw_busy_N_1269)) /* synthesis lut_function=(A ((C)+!B)+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam i10944_2_lut_3_lut.init = 16'hf2f2;
    LUT4 r_word_31__I_0_i31_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[30]), 
         .D(r_word[26]), .Z(r_word_31__N_1197[30])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i31_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i30_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[29]), 
         .D(r_word[25]), .Z(r_word_31__N_1197[29])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i30_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i29_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[28]), 
         .D(r_word[24]), .Z(r_word_31__N_1197[28])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i29_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i28_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[27]), 
         .D(r_word[23]), .Z(r_word_31__N_1197[27])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i28_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i27_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[26]), 
         .D(r_word[22]), .Z(r_word_31__N_1197[26])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i27_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i26_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[25]), 
         .D(r_word[21]), .Z(r_word_31__N_1197[25])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i26_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i25_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[24]), 
         .D(r_word[20]), .Z(r_word_31__N_1197[24])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i25_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i24_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[23]), 
         .D(r_word[19]), .Z(r_word_31__N_1197[23])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i24_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i23_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[22]), 
         .D(r_word[18]), .Z(r_word_31__N_1197[22])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i23_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i22_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[21]), 
         .D(r_word[17]), .Z(r_word_31__N_1197[21])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i22_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i21_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[20]), 
         .D(r_word[16]), .Z(r_word_31__N_1197[20])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i21_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i20_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[19]), 
         .D(r_word[15]), .Z(r_word_31__N_1197[19])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i20_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i19_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[18]), 
         .D(r_word[14]), .Z(r_word_31__N_1197[18])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i19_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i18_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[17]), 
         .D(r_word[13]), .Z(r_word_31__N_1197[17])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i18_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i17_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[16]), 
         .D(r_word[12]), .Z(r_word_31__N_1197[16])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i17_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i16_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[15]), 
         .D(r_word[11]), .Z(r_word_31__N_1197[15])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i16_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i15_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[14]), 
         .D(r_word[10]), .Z(r_word_31__N_1197[14])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i15_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i14_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[13]), 
         .D(r_word[9]), .Z(r_word_31__N_1197[13])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i14_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i13_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[12]), 
         .D(r_word[8]), .Z(r_word_31__N_1197[12])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i13_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i12_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[11]), 
         .D(r_word[7]), .Z(r_word_31__N_1197[11])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i12_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i11_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[10]), 
         .D(r_word[6]), .Z(r_word_31__N_1197[10])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i11_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i10_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[9]), 
         .D(r_word[5]), .Z(r_word_31__N_1197[9])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i10_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i9_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[8]), 
         .D(r_word[4]), .Z(r_word_31__N_1197[8])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i9_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i8_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[7]), 
         .D(r_word[3]), .Z(r_word_31__N_1197[7])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i8_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i7_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[6]), 
         .D(r_word[2]), .Z(r_word_31__N_1197[6])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i7_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i6_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[5]), 
         .D(r_word[1]), .Z(r_word_31__N_1197[5])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i6_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i5_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[4]), 
         .D(r_word[0]), .Z(r_word_31__N_1197[4])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i5_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_28__bdd_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(n24674), 
         .D(r_word[28]), .Z(o_dw_bits_4__N_1188[0])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_28__bdd_3_lut_4_lut.init = 16'hfd20;
    LUT4 i3_4_lut_rep_433 (.A(r_len[0]), .B(r_len[2]), .C(r_len[1]), .D(r_len[3]), 
         .Z(n24993)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(78[16:31])
    defparam i3_4_lut_rep_433.init = 16'hfffe;
    LUT4 i1_2_lut_4_lut (.A(r_len[0]), .B(r_len[2]), .C(r_len[1]), .D(r_len[3]), 
         .Z(n13[0])) /* synthesis lut_function=(!(A+!(B+(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(78[16:31])
    defparam i1_2_lut_4_lut.init = 16'h5554;
    LUT4 i1_2_lut_3_lut_4_lut_adj_105 (.A(r_len[0]), .B(r_len[2]), .C(r_len[1]), 
         .D(r_len[3]), .Z(n11577)) /* synthesis lut_function=(A (C)+!A !(B (C)+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(78[16:31])
    defparam i1_2_lut_3_lut_4_lut_adj_105.init = 16'ha5a4;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut (.A(r_len[0]), .B(r_len[2]), .C(r_len[1]), 
         .D(r_len[3]), .Z(n11575)) /* synthesis lut_function=(A (B)+!A (B (C)+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(78[16:31])
    defparam i1_2_lut_3_lut_4_lut_4_lut.init = 16'hc9c8;
    LUT4 i794_2_lut_3_lut_4_lut_4_lut (.A(r_len[0]), .B(r_len[2]), .C(r_len[1]), 
         .D(r_len[3]), .Z(n6)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(78[16:31])
    defparam i794_2_lut_3_lut_4_lut_4_lut.init = 16'hfeff;
    
endmodule
//
// Verilog Description of module hbpack
//

module hbpack (i_ref_clk_c, i_ref_clk_c_enable_388, n27587, iw_word, 
            \dec_bits[4] , iw_stb, w_reset, o_pck_stb_N_765, cmd_loaded, 
            i_ref_clk_c_enable_192, cmd_loaded_N_768, \dec_bits[0] , \dec_bits[1] , 
            i_ref_clk_c_enable_357, n45, n46, n25103, n27586, newaddr_N_990, 
            n25115, i_cmd_wr) /* synthesis syn_module_defined=1 */ ;
    input i_ref_clk_c;
    input i_ref_clk_c_enable_388;
    input n27587;
    output [33:0]iw_word;
    input \dec_bits[4] ;
    output iw_stb;
    input w_reset;
    input o_pck_stb_N_765;
    output cmd_loaded;
    input i_ref_clk_c_enable_192;
    input cmd_loaded_N_768;
    input \dec_bits[0] ;
    input \dec_bits[1] ;
    input i_ref_clk_c_enable_357;
    input n45;
    input n46;
    output n25103;
    input n27586;
    output newaddr_N_990;
    output n25115;
    output i_cmd_wr;
    
    wire i_ref_clk_c /* synthesis SET_AS_NETWORK=i_ref_clk_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(22[12:21])
    wire [33:0]r_word;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(71[13:19])
    wire [33:0]n14;
    
    FD1P3IX r_word__i0 (.D(n14[0]), .SP(i_ref_clk_c_enable_388), .CD(n27587), 
            .CK(i_ref_clk_c), .Q(r_word[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i0.GSR = "DISABLED";
    FD1P3IX o_pck_word__i0 (.D(r_word[0]), .SP(i_ref_clk_c_enable_388), 
            .CD(n27587), .CK(i_ref_clk_c), .Q(iw_word[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i0.GSR = "DISABLED";
    LUT4 i11306_2_lut (.A(r_word[20]), .B(\dec_bits[4] ), .Z(n14[24])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11306_2_lut.init = 16'h2222;
    LUT4 i11307_2_lut (.A(r_word[19]), .B(\dec_bits[4] ), .Z(n14[23])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11307_2_lut.init = 16'h2222;
    LUT4 i11308_2_lut (.A(r_word[18]), .B(\dec_bits[4] ), .Z(n14[22])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11308_2_lut.init = 16'h2222;
    LUT4 i11309_2_lut (.A(r_word[17]), .B(\dec_bits[4] ), .Z(n14[21])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11309_2_lut.init = 16'h2222;
    LUT4 i11310_2_lut (.A(r_word[16]), .B(\dec_bits[4] ), .Z(n14[20])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11310_2_lut.init = 16'h2222;
    FD1S3IX o_pck_stb_24 (.D(o_pck_stb_N_765), .CK(i_ref_clk_c), .CD(w_reset), 
            .Q(iw_stb)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(83[9] 84[65])
    defparam o_pck_stb_24.GSR = "DISABLED";
    LUT4 i11311_2_lut (.A(r_word[15]), .B(\dec_bits[4] ), .Z(n14[19])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11311_2_lut.init = 16'h2222;
    LUT4 i11312_2_lut (.A(r_word[14]), .B(\dec_bits[4] ), .Z(n14[18])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11312_2_lut.init = 16'h2222;
    LUT4 i11313_2_lut (.A(r_word[13]), .B(\dec_bits[4] ), .Z(n14[17])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11313_2_lut.init = 16'h2222;
    LUT4 i11314_2_lut (.A(r_word[12]), .B(\dec_bits[4] ), .Z(n14[16])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11314_2_lut.init = 16'h2222;
    LUT4 i11320_2_lut (.A(r_word[11]), .B(\dec_bits[4] ), .Z(n14[15])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11320_2_lut.init = 16'h2222;
    LUT4 i11321_2_lut (.A(r_word[10]), .B(\dec_bits[4] ), .Z(n14[14])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11321_2_lut.init = 16'h2222;
    LUT4 i11322_2_lut (.A(r_word[9]), .B(\dec_bits[4] ), .Z(n14[13])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11322_2_lut.init = 16'h2222;
    LUT4 i11323_2_lut (.A(r_word[8]), .B(\dec_bits[4] ), .Z(n14[12])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11323_2_lut.init = 16'h2222;
    FD1P3IX cmd_loaded_23 (.D(cmd_loaded_N_768), .SP(i_ref_clk_c_enable_192), 
            .CD(w_reset), .CK(i_ref_clk_c), .Q(cmd_loaded)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(74[9] 80[23])
    defparam cmd_loaded_23.GSR = "DISABLED";
    LUT4 i11328_2_lut (.A(r_word[7]), .B(\dec_bits[4] ), .Z(n14[11])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11328_2_lut.init = 16'h2222;
    LUT4 i11329_2_lut (.A(r_word[6]), .B(\dec_bits[4] ), .Z(n14[10])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11329_2_lut.init = 16'h2222;
    LUT4 i11330_2_lut (.A(r_word[5]), .B(\dec_bits[4] ), .Z(n14[9])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11330_2_lut.init = 16'h2222;
    LUT4 i11331_2_lut (.A(r_word[4]), .B(\dec_bits[4] ), .Z(n14[8])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11331_2_lut.init = 16'h2222;
    LUT4 i11332_2_lut (.A(r_word[3]), .B(\dec_bits[4] ), .Z(n14[7])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11332_2_lut.init = 16'h2222;
    LUT4 i11333_2_lut (.A(r_word[2]), .B(\dec_bits[4] ), .Z(n14[6])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11333_2_lut.init = 16'h2222;
    LUT4 i11334_2_lut (.A(r_word[1]), .B(\dec_bits[4] ), .Z(n14[5])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11334_2_lut.init = 16'h2222;
    LUT4 i11335_2_lut (.A(r_word[0]), .B(\dec_bits[4] ), .Z(n14[4])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11335_2_lut.init = 16'h2222;
    FD1P3IX o_pck_word__i33 (.D(r_word[33]), .SP(i_ref_clk_c_enable_388), 
            .CD(w_reset), .CK(i_ref_clk_c), .Q(iw_word[33])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i33.GSR = "DISABLED";
    FD1P3IX o_pck_word__i32 (.D(r_word[32]), .SP(i_ref_clk_c_enable_388), 
            .CD(w_reset), .CK(i_ref_clk_c), .Q(iw_word[32])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i32.GSR = "DISABLED";
    FD1P3IX o_pck_word__i31 (.D(r_word[31]), .SP(i_ref_clk_c_enable_388), 
            .CD(w_reset), .CK(i_ref_clk_c), .Q(iw_word[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i31.GSR = "DISABLED";
    FD1P3IX o_pck_word__i30 (.D(r_word[30]), .SP(i_ref_clk_c_enable_388), 
            .CD(w_reset), .CK(i_ref_clk_c), .Q(iw_word[30])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i30.GSR = "DISABLED";
    FD1P3IX o_pck_word__i29 (.D(r_word[29]), .SP(i_ref_clk_c_enable_388), 
            .CD(w_reset), .CK(i_ref_clk_c), .Q(iw_word[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i29.GSR = "DISABLED";
    FD1P3IX o_pck_word__i28 (.D(r_word[28]), .SP(i_ref_clk_c_enable_388), 
            .CD(w_reset), .CK(i_ref_clk_c), .Q(iw_word[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i28.GSR = "DISABLED";
    FD1P3IX o_pck_word__i27 (.D(r_word[27]), .SP(i_ref_clk_c_enable_388), 
            .CD(w_reset), .CK(i_ref_clk_c), .Q(iw_word[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i27.GSR = "DISABLED";
    FD1P3IX o_pck_word__i26 (.D(r_word[26]), .SP(i_ref_clk_c_enable_388), 
            .CD(w_reset), .CK(i_ref_clk_c), .Q(iw_word[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i26.GSR = "DISABLED";
    FD1P3IX o_pck_word__i25 (.D(r_word[25]), .SP(i_ref_clk_c_enable_388), 
            .CD(w_reset), .CK(i_ref_clk_c), .Q(iw_word[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i25.GSR = "DISABLED";
    FD1P3IX o_pck_word__i24 (.D(r_word[24]), .SP(i_ref_clk_c_enable_388), 
            .CD(w_reset), .CK(i_ref_clk_c), .Q(iw_word[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i24.GSR = "DISABLED";
    LUT4 i10930_2_lut (.A(\dec_bits[0] ), .B(\dec_bits[4] ), .Z(n14[0])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i10930_2_lut.init = 16'h2222;
    FD1P3IX o_pck_word__i23 (.D(r_word[23]), .SP(i_ref_clk_c_enable_388), 
            .CD(n27587), .CK(i_ref_clk_c), .Q(iw_word[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i23.GSR = "DISABLED";
    FD1P3IX o_pck_word__i22 (.D(r_word[22]), .SP(i_ref_clk_c_enable_388), 
            .CD(n27587), .CK(i_ref_clk_c), .Q(iw_word[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i22.GSR = "DISABLED";
    FD1P3IX o_pck_word__i21 (.D(r_word[21]), .SP(i_ref_clk_c_enable_388), 
            .CD(w_reset), .CK(i_ref_clk_c), .Q(iw_word[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i21.GSR = "DISABLED";
    FD1P3IX o_pck_word__i20 (.D(r_word[20]), .SP(i_ref_clk_c_enable_388), 
            .CD(n27587), .CK(i_ref_clk_c), .Q(iw_word[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i20.GSR = "DISABLED";
    FD1P3IX o_pck_word__i19 (.D(r_word[19]), .SP(i_ref_clk_c_enable_388), 
            .CD(n27587), .CK(i_ref_clk_c), .Q(iw_word[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i19.GSR = "DISABLED";
    FD1P3IX o_pck_word__i18 (.D(r_word[18]), .SP(i_ref_clk_c_enable_388), 
            .CD(n27587), .CK(i_ref_clk_c), .Q(iw_word[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i18.GSR = "DISABLED";
    FD1P3IX o_pck_word__i17 (.D(r_word[17]), .SP(i_ref_clk_c_enable_388), 
            .CD(n27587), .CK(i_ref_clk_c), .Q(iw_word[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i17.GSR = "DISABLED";
    FD1P3IX o_pck_word__i16 (.D(r_word[16]), .SP(i_ref_clk_c_enable_388), 
            .CD(n27587), .CK(i_ref_clk_c), .Q(iw_word[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i16.GSR = "DISABLED";
    FD1P3IX o_pck_word__i15 (.D(r_word[15]), .SP(i_ref_clk_c_enable_388), 
            .CD(n27587), .CK(i_ref_clk_c), .Q(iw_word[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i15.GSR = "DISABLED";
    FD1P3IX o_pck_word__i14 (.D(r_word[14]), .SP(i_ref_clk_c_enable_388), 
            .CD(n27587), .CK(i_ref_clk_c), .Q(iw_word[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i14.GSR = "DISABLED";
    FD1P3IX o_pck_word__i13 (.D(r_word[13]), .SP(i_ref_clk_c_enable_388), 
            .CD(n27587), .CK(i_ref_clk_c), .Q(iw_word[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i13.GSR = "DISABLED";
    FD1P3IX o_pck_word__i12 (.D(r_word[12]), .SP(i_ref_clk_c_enable_388), 
            .CD(n27587), .CK(i_ref_clk_c), .Q(iw_word[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i12.GSR = "DISABLED";
    FD1P3IX o_pck_word__i11 (.D(r_word[11]), .SP(i_ref_clk_c_enable_388), 
            .CD(n27587), .CK(i_ref_clk_c), .Q(iw_word[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i11.GSR = "DISABLED";
    FD1P3IX o_pck_word__i10 (.D(r_word[10]), .SP(i_ref_clk_c_enable_388), 
            .CD(n27587), .CK(i_ref_clk_c), .Q(iw_word[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i10.GSR = "DISABLED";
    FD1P3IX o_pck_word__i9 (.D(r_word[9]), .SP(i_ref_clk_c_enable_388), 
            .CD(n27587), .CK(i_ref_clk_c), .Q(iw_word[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i9.GSR = "DISABLED";
    FD1P3IX o_pck_word__i8 (.D(r_word[8]), .SP(i_ref_clk_c_enable_388), 
            .CD(n27587), .CK(i_ref_clk_c), .Q(iw_word[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i8.GSR = "DISABLED";
    FD1P3IX o_pck_word__i7 (.D(r_word[7]), .SP(i_ref_clk_c_enable_388), 
            .CD(n27587), .CK(i_ref_clk_c), .Q(iw_word[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i7.GSR = "DISABLED";
    FD1P3IX o_pck_word__i6 (.D(r_word[6]), .SP(i_ref_clk_c_enable_388), 
            .CD(n27587), .CK(i_ref_clk_c), .Q(iw_word[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i6.GSR = "DISABLED";
    FD1P3IX o_pck_word__i5 (.D(r_word[5]), .SP(i_ref_clk_c_enable_388), 
            .CD(n27587), .CK(i_ref_clk_c), .Q(iw_word[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i5.GSR = "DISABLED";
    FD1P3IX o_pck_word__i4 (.D(r_word[4]), .SP(i_ref_clk_c_enable_388), 
            .CD(n27587), .CK(i_ref_clk_c), .Q(iw_word[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i4.GSR = "DISABLED";
    FD1P3IX o_pck_word__i3 (.D(r_word[3]), .SP(i_ref_clk_c_enable_388), 
            .CD(n27587), .CK(i_ref_clk_c), .Q(iw_word[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i3.GSR = "DISABLED";
    FD1P3IX o_pck_word__i2 (.D(r_word[2]), .SP(i_ref_clk_c_enable_388), 
            .CD(n27587), .CK(i_ref_clk_c), .Q(iw_word[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i2.GSR = "DISABLED";
    FD1P3IX o_pck_word__i1 (.D(r_word[1]), .SP(i_ref_clk_c_enable_388), 
            .CD(n27587), .CK(i_ref_clk_c), .Q(iw_word[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i1.GSR = "DISABLED";
    LUT4 i11336_2_lut (.A(\dec_bits[1] ), .B(\dec_bits[4] ), .Z(n14[1])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11336_2_lut.init = 16'h2222;
    FD1P3IX r_word__i33 (.D(\dec_bits[1] ), .SP(i_ref_clk_c_enable_357), 
            .CD(n27587), .CK(i_ref_clk_c), .Q(r_word[33])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i33.GSR = "DISABLED";
    FD1P3IX r_word__i32 (.D(\dec_bits[0] ), .SP(i_ref_clk_c_enable_357), 
            .CD(n27587), .CK(i_ref_clk_c), .Q(r_word[32])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i32.GSR = "DISABLED";
    FD1P3IX r_word__i31 (.D(n14[31]), .SP(i_ref_clk_c_enable_388), .CD(n27587), 
            .CK(i_ref_clk_c), .Q(r_word[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i31.GSR = "DISABLED";
    FD1P3IX r_word__i30 (.D(n14[30]), .SP(i_ref_clk_c_enable_388), .CD(n27587), 
            .CK(i_ref_clk_c), .Q(r_word[30])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i30.GSR = "DISABLED";
    FD1P3IX r_word__i29 (.D(n14[29]), .SP(i_ref_clk_c_enable_388), .CD(n27587), 
            .CK(i_ref_clk_c), .Q(r_word[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i29.GSR = "DISABLED";
    FD1P3IX r_word__i28 (.D(n14[28]), .SP(i_ref_clk_c_enable_388), .CD(n27587), 
            .CK(i_ref_clk_c), .Q(r_word[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i28.GSR = "DISABLED";
    FD1P3IX r_word__i27 (.D(n14[27]), .SP(i_ref_clk_c_enable_388), .CD(n27587), 
            .CK(i_ref_clk_c), .Q(r_word[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i27.GSR = "DISABLED";
    FD1P3IX r_word__i26 (.D(n14[26]), .SP(i_ref_clk_c_enable_388), .CD(n27587), 
            .CK(i_ref_clk_c), .Q(r_word[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i26.GSR = "DISABLED";
    FD1P3IX r_word__i25 (.D(n14[25]), .SP(i_ref_clk_c_enable_388), .CD(n27587), 
            .CK(i_ref_clk_c), .Q(r_word[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i25.GSR = "DISABLED";
    FD1P3IX r_word__i24 (.D(n14[24]), .SP(i_ref_clk_c_enable_388), .CD(n27587), 
            .CK(i_ref_clk_c), .Q(r_word[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i24.GSR = "DISABLED";
    FD1P3IX r_word__i23 (.D(n14[23]), .SP(i_ref_clk_c_enable_388), .CD(n27587), 
            .CK(i_ref_clk_c), .Q(r_word[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i23.GSR = "DISABLED";
    FD1P3IX r_word__i22 (.D(n14[22]), .SP(i_ref_clk_c_enable_388), .CD(n27587), 
            .CK(i_ref_clk_c), .Q(r_word[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i22.GSR = "DISABLED";
    FD1P3IX r_word__i21 (.D(n14[21]), .SP(i_ref_clk_c_enable_388), .CD(n27587), 
            .CK(i_ref_clk_c), .Q(r_word[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i21.GSR = "DISABLED";
    FD1P3IX r_word__i20 (.D(n14[20]), .SP(i_ref_clk_c_enable_388), .CD(n27587), 
            .CK(i_ref_clk_c), .Q(r_word[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i20.GSR = "DISABLED";
    FD1P3IX r_word__i19 (.D(n14[19]), .SP(i_ref_clk_c_enable_388), .CD(n27587), 
            .CK(i_ref_clk_c), .Q(r_word[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i19.GSR = "DISABLED";
    FD1P3IX r_word__i18 (.D(n14[18]), .SP(i_ref_clk_c_enable_388), .CD(n27587), 
            .CK(i_ref_clk_c), .Q(r_word[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i18.GSR = "DISABLED";
    FD1P3IX r_word__i17 (.D(n14[17]), .SP(i_ref_clk_c_enable_388), .CD(n27587), 
            .CK(i_ref_clk_c), .Q(r_word[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i17.GSR = "DISABLED";
    FD1P3IX r_word__i16 (.D(n14[16]), .SP(i_ref_clk_c_enable_388), .CD(w_reset), 
            .CK(i_ref_clk_c), .Q(r_word[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i16.GSR = "DISABLED";
    FD1P3IX r_word__i15 (.D(n14[15]), .SP(i_ref_clk_c_enable_388), .CD(w_reset), 
            .CK(i_ref_clk_c), .Q(r_word[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i15.GSR = "DISABLED";
    FD1P3IX r_word__i14 (.D(n14[14]), .SP(i_ref_clk_c_enable_388), .CD(w_reset), 
            .CK(i_ref_clk_c), .Q(r_word[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i14.GSR = "DISABLED";
    FD1P3IX r_word__i13 (.D(n14[13]), .SP(i_ref_clk_c_enable_388), .CD(w_reset), 
            .CK(i_ref_clk_c), .Q(r_word[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i13.GSR = "DISABLED";
    FD1P3IX r_word__i12 (.D(n14[12]), .SP(i_ref_clk_c_enable_388), .CD(w_reset), 
            .CK(i_ref_clk_c), .Q(r_word[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i12.GSR = "DISABLED";
    FD1P3IX r_word__i11 (.D(n14[11]), .SP(i_ref_clk_c_enable_388), .CD(w_reset), 
            .CK(i_ref_clk_c), .Q(r_word[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i11.GSR = "DISABLED";
    FD1P3IX r_word__i10 (.D(n14[10]), .SP(i_ref_clk_c_enable_388), .CD(w_reset), 
            .CK(i_ref_clk_c), .Q(r_word[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i10.GSR = "DISABLED";
    FD1P3IX r_word__i9 (.D(n14[9]), .SP(i_ref_clk_c_enable_388), .CD(w_reset), 
            .CK(i_ref_clk_c), .Q(r_word[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i9.GSR = "DISABLED";
    FD1P3IX r_word__i8 (.D(n14[8]), .SP(i_ref_clk_c_enable_388), .CD(w_reset), 
            .CK(i_ref_clk_c), .Q(r_word[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i8.GSR = "DISABLED";
    FD1P3IX r_word__i7 (.D(n14[7]), .SP(i_ref_clk_c_enable_388), .CD(w_reset), 
            .CK(i_ref_clk_c), .Q(r_word[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i7.GSR = "DISABLED";
    FD1P3IX r_word__i6 (.D(n14[6]), .SP(i_ref_clk_c_enable_388), .CD(w_reset), 
            .CK(i_ref_clk_c), .Q(r_word[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i6.GSR = "DISABLED";
    FD1P3IX r_word__i5 (.D(n14[5]), .SP(i_ref_clk_c_enable_388), .CD(w_reset), 
            .CK(i_ref_clk_c), .Q(r_word[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i5.GSR = "DISABLED";
    FD1P3IX r_word__i4 (.D(n14[4]), .SP(i_ref_clk_c_enable_388), .CD(w_reset), 
            .CK(i_ref_clk_c), .Q(r_word[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i4.GSR = "DISABLED";
    FD1P3IX r_word__i3 (.D(n45), .SP(i_ref_clk_c_enable_388), .CD(w_reset), 
            .CK(i_ref_clk_c), .Q(r_word[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i3.GSR = "DISABLED";
    FD1P3IX r_word__i2 (.D(n46), .SP(i_ref_clk_c_enable_388), .CD(w_reset), 
            .CK(i_ref_clk_c), .Q(r_word[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i2.GSR = "DISABLED";
    FD1P3IX r_word__i1 (.D(n14[1]), .SP(i_ref_clk_c_enable_388), .CD(w_reset), 
            .CK(i_ref_clk_c), .Q(r_word[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i1.GSR = "DISABLED";
    LUT4 i11299_2_lut (.A(r_word[27]), .B(\dec_bits[4] ), .Z(n14[31])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11299_2_lut.init = 16'h2222;
    LUT4 i11300_2_lut (.A(r_word[26]), .B(\dec_bits[4] ), .Z(n14[30])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11300_2_lut.init = 16'h2222;
    LUT4 i11301_2_lut (.A(r_word[25]), .B(\dec_bits[4] ), .Z(n14[29])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11301_2_lut.init = 16'h2222;
    LUT4 i11305_2_lut (.A(r_word[21]), .B(\dec_bits[4] ), .Z(n14[25])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11305_2_lut.init = 16'h2222;
    LUT4 i11304_2_lut (.A(r_word[22]), .B(\dec_bits[4] ), .Z(n14[26])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11304_2_lut.init = 16'h2222;
    LUT4 i11302_2_lut (.A(r_word[24]), .B(\dec_bits[4] ), .Z(n14[28])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11302_2_lut.init = 16'h2222;
    LUT4 i11303_2_lut (.A(r_word[23]), .B(\dec_bits[4] ), .Z(n14[27])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11303_2_lut.init = 16'h2222;
    LUT4 i2_3_lut_rep_543 (.A(iw_word[32]), .B(iw_word[33]), .C(iw_stb), 
         .Z(n25103)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(83[9] 84[65])
    defparam i2_3_lut_rep_543.init = 16'h4040;
    LUT4 i1_2_lut_4_lut (.A(iw_word[32]), .B(iw_word[33]), .C(iw_stb), 
         .D(n27586), .Z(newaddr_N_990)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(83[9] 84[65])
    defparam i1_2_lut_4_lut.init = 16'h0040;
    LUT4 i1_2_lut_rep_555 (.A(iw_stb), .B(iw_word[33]), .Z(n25115)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(83[9] 84[65])
    defparam i1_2_lut_rep_555.init = 16'h2222;
    LUT4 i1_2_lut_3_lut (.A(iw_stb), .B(iw_word[33]), .C(iw_word[32]), 
         .Z(i_cmd_wr)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(83[9] 84[65])
    defparam i1_2_lut_3_lut.init = 16'h2020;
    
endmodule
//
// Verilog Description of module hbgenhex
//

module hbgenhex (hb_bits, \w_gx_char[0] , \w_gx_char[1] , \w_gx_char[2] , 
            \w_gx_char[3] , \w_gx_char[4] , \w_gx_char[5] , \w_gx_char[6] , 
            i_ref_clk_c, i_ref_clk_c_enable_315, GND_net, VCC_net, hx_stb, 
            w_reset, hb_busy, n11767, nl_busy, n27586, n24991, i_ref_clk_c_enable_194) /* synthesis syn_module_defined=1 */ ;
    input [4:0]hb_bits;
    output \w_gx_char[0] ;
    output \w_gx_char[1] ;
    output \w_gx_char[2] ;
    output \w_gx_char[3] ;
    output \w_gx_char[4] ;
    output \w_gx_char[5] ;
    output \w_gx_char[6] ;
    input i_ref_clk_c;
    output i_ref_clk_c_enable_315;
    input GND_net;
    input VCC_net;
    output hx_stb;
    input w_reset;
    input hb_busy;
    output n11767;
    input nl_busy;
    input n27586;
    input n24991;
    output i_ref_clk_c_enable_194;
    
    wire i_ref_clk_c /* synthesis SET_AS_NETWORK=i_ref_clk_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(22[12:21])
    
    wire i_ref_clk_c_enable_148, n19717, n6;
    
    SP8KC mux_105 (.DI0(GND_net), .DI1(GND_net), .DI2(GND_net), .DI3(GND_net), 
          .DI4(GND_net), .DI5(GND_net), .DI6(GND_net), .DI7(GND_net), 
          .DI8(GND_net), .AD0(GND_net), .AD1(GND_net), .AD2(GND_net), 
          .AD3(hb_bits[0]), .AD4(hb_bits[1]), .AD5(hb_bits[2]), .AD6(hb_bits[3]), 
          .AD7(hb_bits[4]), .AD8(GND_net), .AD9(GND_net), .AD10(GND_net), 
          .AD11(GND_net), .AD12(GND_net), .CE(i_ref_clk_c_enable_315), 
          .OCE(VCC_net), .CLK(i_ref_clk_c), .WE(GND_net), .CS0(GND_net), 
          .CS1(GND_net), .CS2(GND_net), .RST(GND_net), .DO0(\w_gx_char[0] ), 
          .DO1(\w_gx_char[1] ), .DO2(\w_gx_char[2] ), .DO3(\w_gx_char[3] ), 
          .DO4(\w_gx_char[4] ), .DO5(\w_gx_char[5] ), .DO6(\w_gx_char[6] ));
    defparam mux_105.DATA_WIDTH = 9;
    defparam mux_105.REGMODE = "NOREG";
    defparam mux_105.CSDECODE = "0b000";
    defparam mux_105.WRITEMODE = "NORMAL";
    defparam mux_105.GSR = "DISABLED";
    defparam mux_105.RESETMODE = "ASYNC";
    defparam mux_105.ASYNC_RESET_RELEASE = "SYNC";
    defparam mux_105.INIT_DATA = "STATIC";
    defparam mux_105.INITVAL_00 = "0x01A0D01A0D0B44908A5401A0D01A0D0A641096520CC650C8630C4610723806E3606A340663206230";
    defparam mux_105.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_105.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_105.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_105.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_105.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_105.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_105.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_105.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_105.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_105.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_105.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_105.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_105.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_105.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_105.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_105.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_105.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_105.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_105.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_105.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_105.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_105.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_105.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_105.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_105.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_105.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_105.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_105.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_105.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_105.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_105.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    FD1P3IX o_gx_stb_13 (.D(hb_busy), .SP(i_ref_clk_c_enable_148), .CD(w_reset), 
            .CK(i_ref_clk_c), .Q(hx_stb)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=132, LSE_RLINE=133 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbgenhex.v(74[9] 78[21])
    defparam o_gx_stb_13.GSR = "DISABLED";
    LUT4 i4_4_lut (.A(\w_gx_char[1] ), .B(n19717), .C(\w_gx_char[5] ), 
         .D(n6), .Z(n11767)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;
    defparam i4_4_lut.init = 16'hfffb;
    LUT4 i17405_3_lut (.A(\w_gx_char[2] ), .B(\w_gx_char[0] ), .C(\w_gx_char[3] ), 
         .Z(n19717)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i17405_3_lut.init = 16'h8080;
    LUT4 i1_2_lut (.A(\w_gx_char[4] ), .B(\w_gx_char[6] ), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i21055_2_lut_rep_329 (.A(hx_stb), .B(nl_busy), .Z(i_ref_clk_c_enable_315)) /* synthesis lut_function=(!(A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(76[16:26])
    defparam i21055_2_lut_rep_329.init = 16'h7777;
    LUT4 i1_2_lut_rep_325_3_lut (.A(hx_stb), .B(nl_busy), .C(n27586), 
         .Z(i_ref_clk_c_enable_148)) /* synthesis lut_function=(((C)+!B)+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(76[16:26])
    defparam i1_2_lut_rep_325_3_lut.init = 16'hf7f7;
    LUT4 i2_2_lut_3_lut_4_lut (.A(hx_stb), .B(nl_busy), .C(n24991), .D(n27586), 
         .Z(i_ref_clk_c_enable_194)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(76[16:26])
    defparam i2_2_lut_3_lut_4_lut.init = 16'hfff7;
    
endmodule
//
// Verilog Description of module hbdechex
//

module hbdechex (\rx_data[6] , i_ref_clk_c, dec_bits, w_reset, n27586, 
            \rx_data[0] , \rx_data[5] , \rx_data[1] , \rx_data[2] , 
            rx_stb, \rx_data[3] , \rx_data[4] , \dec_bits[1] , n45, 
            n46, n27587, i_ref_clk_c_enable_388, i_ref_clk_c_enable_357, 
            cmd_loaded, o_pck_stb_N_765, i_ref_clk_c_enable_192, cmd_loaded_N_768) /* synthesis syn_module_defined=1 */ ;
    input \rx_data[6] ;
    input i_ref_clk_c;
    output [4:0]dec_bits;
    output w_reset;
    output n27586;
    input \rx_data[0] ;
    input \rx_data[5] ;
    input \rx_data[1] ;
    input \rx_data[2] ;
    input rx_stb;
    input \rx_data[3] ;
    input \rx_data[4] ;
    output \dec_bits[1] ;
    output n45;
    output n46;
    output n27587;
    output i_ref_clk_c_enable_388;
    output i_ref_clk_c_enable_357;
    input cmd_loaded;
    output o_pck_stb_N_765;
    output i_ref_clk_c_enable_192;
    output cmd_loaded_N_768;
    
    wire i_ref_clk_c /* synthesis SET_AS_NETWORK=i_ref_clk_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(22[12:21])
    
    wire n22102, n22103;
    wire [4:0]o_dh_bits_4__N_596;
    
    wire dec_stb, o_dh_stb_N_623, o_reset_N_625, n64, n19461, n14506, 
        n19434, n72, n9, n44, n53, n19485, n19617, n47, n12, 
        n11809, n24796, n22929, n22928;
    wire [4:0]dec_bits_c;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(69[13:21])
    
    wire n25002, n25003, n48, n19464, n24837, n24086, n24084, 
        n24983, n6, n56, n24984, n32, n24801, n24, n41, n52, 
        n24127, n25007, n69;
    
    PFUMX i109 (.BLUT(n22102), .ALUT(n22103), .C0(\rx_data[6] ), .Z(o_dh_bits_4__N_596[3]));
    FD1S3AX o_dh_stb_35 (.D(o_dh_stb_N_623), .CK(i_ref_clk_c), .Q(dec_stb)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=30, LSE_LLINE=93, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(57[9] 58[47])
    defparam o_dh_stb_35.GSR = "DISABLED";
    FD1S3AX o_dh_bits_i0 (.D(o_dh_bits_4__N_596[0]), .CK(i_ref_clk_c), .Q(dec_bits[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=30, LSE_LLINE=93, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(60[9] 100[5])
    defparam o_dh_bits_i0.GSR = "DISABLED";
    FD1S3AY o_reset_34 (.D(o_reset_N_625), .CK(i_ref_clk_c), .Q(w_reset)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=30, LSE_LLINE=93, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(53[9] 54[46])
    defparam o_reset_34.GSR = "DISABLED";
    FD1S3AY o_reset_34_rep_688 (.D(o_reset_N_625), .CK(i_ref_clk_c), .Q(n27586)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=30, LSE_LLINE=93, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(53[9] 54[46])
    defparam o_reset_34_rep_688.GSR = "DISABLED";
    LUT4 i1_4_lut_4_lut (.A(\rx_data[0] ), .B(\rx_data[5] ), .C(\rx_data[1] ), 
         .D(\rx_data[2] ), .Z(n64)) /* synthesis lut_function=(!(A (B (C (D))+!B (C+(D)))+!A !(B (C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(65[3] 99[10])
    defparam i1_4_lut_4_lut.init = 16'h4cca;
    LUT4 i_stb_I_0_58_4_lut (.A(rx_stb), .B(\rx_data[6] ), .C(n19461), 
         .D(n14506), .Z(o_dh_stb_N_623)) /* synthesis lut_function=(!((B (C (D)))+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(58[15:46])
    defparam i_stb_I_0_58_4_lut.init = 16'h2aaa;
    LUT4 i1_4_lut (.A(n19434), .B(n72), .C(n9), .D(n44), .Z(o_dh_bits_4__N_596[0])) /* synthesis lut_function=(A+(B+!(C+!(D)))) */ ;
    defparam i1_4_lut.init = 16'hefee;
    LUT4 i2_4_lut (.A(\rx_data[6] ), .B(n53), .C(n19485), .D(n19617), 
         .Z(n19434)) /* synthesis lut_function=(A (B+!(D))+!A (C+!(D))) */ ;
    defparam i2_4_lut.init = 16'hd8ff;
    LUT4 i1_3_lut (.A(\rx_data[3] ), .B(n47), .C(\rx_data[4] ), .Z(n53)) /* synthesis lut_function=(A+!(B+!(C))) */ ;
    defparam i1_3_lut.init = 16'hbaba;
    LUT4 i17316_2_lut (.A(n64), .B(\rx_data[4] ), .Z(n19617)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i17316_2_lut.init = 16'heeee;
    LUT4 i_stb_I_0_4_lut (.A(rx_stb), .B(\rx_data[0] ), .C(n12), .D(n11809), 
         .Z(o_reset_N_625)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(54[14:45])
    defparam i_stb_I_0_4_lut.init = 16'h0002;
    LUT4 i1_2_lut (.A(\rx_data[1] ), .B(\rx_data[2] ), .Z(n11809)) /* synthesis lut_function=(A+!(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(72[3:8])
    defparam i1_2_lut.init = 16'hbbbb;
    LUT4 n61_bdd_4_lut_4_lut (.A(\rx_data[1] ), .B(\rx_data[2] ), .C(\rx_data[0] ), 
         .D(\rx_data[4] ), .Z(n24796)) /* synthesis lut_function=(A (B (C (D))+!B (D))+!A !(B (C+!(D))+!B ((D)+!C))) */ ;
    defparam n61_bdd_4_lut_4_lut.init = 16'ha610;
    FD1S3AX o_dh_bits_i4 (.D(o_dh_bits_4__N_596[4]), .CK(i_ref_clk_c), .Q(dec_bits[4])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=30, LSE_LLINE=93, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(60[9] 100[5])
    defparam o_dh_bits_i4.GSR = "DISABLED";
    LUT4 n19512_bdd_4_lut (.A(\rx_data[0] ), .B(\rx_data[2] ), .C(\rx_data[1] ), 
         .D(\rx_data[5] ), .Z(n22929)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A !(C (D)))) */ ;
    defparam n19512_bdd_4_lut.init = 16'h5800;
    LUT4 n19512_bdd_4_lut_21402 (.A(\rx_data[0] ), .B(\rx_data[2] ), .C(\rx_data[1] ), 
         .D(\rx_data[5] ), .Z(n22928)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A ((C+(D))+!B))) */ ;
    defparam n19512_bdd_4_lut_21402.init = 16'h0024;
    FD1S3AX o_dh_bits_i3 (.D(o_dh_bits_4__N_596[3]), .CK(i_ref_clk_c), .Q(dec_bits_c[3])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=30, LSE_LLINE=93, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(60[9] 100[5])
    defparam o_dh_bits_i3.GSR = "DISABLED";
    FD1S3AX o_dh_bits_i2 (.D(o_dh_bits_4__N_596[2]), .CK(i_ref_clk_c), .Q(dec_bits_c[2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=30, LSE_LLINE=93, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(60[9] 100[5])
    defparam o_dh_bits_i2.GSR = "DISABLED";
    FD1S3AX o_dh_bits_i1 (.D(o_dh_bits_4__N_596[1]), .CK(i_ref_clk_c), .Q(\dec_bits[1] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=30, LSE_LLINE=93, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(60[9] 100[5])
    defparam o_dh_bits_i1.GSR = "DISABLED";
    LUT4 i1_2_lut_adj_93 (.A(dec_bits[4]), .B(dec_bits_c[3]), .Z(n45)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(60[9] 100[5])
    defparam i1_2_lut_adj_93.init = 16'h4444;
    LUT4 i1_2_lut_2_lut_3_lut_4_lut (.A(\rx_data[4] ), .B(n25002), .C(n25003), 
         .D(\rx_data[5] ), .Z(n48)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(87[3:8])
    defparam i1_2_lut_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 i1_2_lut_adj_94 (.A(\rx_data[4] ), .B(\rx_data[5] ), .Z(n19464)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i1_2_lut_adj_94.init = 16'h2222;
    LUT4 i1_2_lut_adj_95 (.A(dec_bits[4]), .B(dec_bits_c[2]), .Z(n46)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(60[9] 100[5])
    defparam i1_2_lut_adj_95.init = 16'h4444;
    LUT4 rx_data_1__bdd_4_lut_24085 (.A(\rx_data[1] ), .B(\rx_data[0] ), 
         .C(\rx_data[2] ), .D(n24837), .Z(n24086)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A (B+((D)+!C)))) */ ;
    defparam rx_data_1__bdd_4_lut_24085.init = 16'h0038;
    LUT4 n9_bdd_4_lut (.A(n9), .B(n25002), .C(\rx_data[4] ), .D(\rx_data[5] ), 
         .Z(n24084)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam n9_bdd_4_lut.init = 16'hfefa;
    LUT4 i1_4_lut_adj_96 (.A(n19617), .B(n24983), .C(n6), .D(n24086), 
         .Z(o_dh_bits_4__N_596[2])) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i1_4_lut_adj_96.init = 16'hfffd;
    LUT4 i2_4_lut_adj_97 (.A(\rx_data[2] ), .B(n56), .C(n24984), .D(n32), 
         .Z(n6)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B)) */ ;
    defparam i2_4_lut_adj_97.init = 16'heeec;
    LUT4 i1_4_lut_adj_98 (.A(n19434), .B(n24801), .C(n24), .D(n24084), 
         .Z(o_dh_bits_4__N_596[1])) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;
    defparam i1_4_lut_adj_98.init = 16'hfeff;
    FD1S3AY o_reset_34_rep_689 (.D(o_reset_N_625), .CK(i_ref_clk_c), .Q(n27587)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=30, LSE_LLINE=93, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(53[9] 54[46])
    defparam o_reset_34_rep_689.GSR = "DISABLED";
    PFUMX i73 (.BLUT(n48), .ALUT(n41), .C0(\rx_data[0] ), .Z(n72));
    LUT4 n22929_bdd_4_lut (.A(n22929), .B(n25002), .C(n22928), .D(\rx_data[4] ), 
         .Z(n24801)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C (D))) */ ;
    defparam n22929_bdd_4_lut.init = 16'hf022;
    LUT4 i1_4_lut_4_lut_adj_99 (.A(n24837), .B(n19464), .C(\rx_data[0] ), 
         .D(\rx_data[1] ), .Z(n32)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A (D))) */ ;
    defparam i1_4_lut_4_lut_adj_99.init = 16'h005d;
    LUT4 dac_clk_n_c_bdd_2_lut_22907_3_lut_4_lut (.A(n24796), .B(\rx_data[5] ), 
         .C(n52), .D(\rx_data[3] ), .Z(n24127)) /* synthesis lut_function=(A (((D)+!C)+!B)+!A ((D)+!C)) */ ;
    defparam dac_clk_n_c_bdd_2_lut_22907_3_lut_4_lut.init = 16'hff2f;
    PFUMX i22491 (.BLUT(n19485), .ALUT(n24127), .C0(\rx_data[6] ), .Z(o_dh_bits_4__N_596[4]));
    LUT4 i1_2_lut_4_lut (.A(n25007), .B(\rx_data[6] ), .C(\rx_data[3] ), 
         .D(\rx_data[1] ), .Z(n24)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_2_lut_4_lut.init = 16'h0200;
    LUT4 i20880_1_lut_3_lut (.A(\rx_data[4] ), .B(\rx_data[3] ), .C(\rx_data[5] ), 
         .Z(n22102)) /* synthesis lut_function=((B+!(C))+!A) */ ;
    defparam i20880_1_lut_3_lut.init = 16'hdfdf;
    LUT4 i11831_2_lut_3_lut (.A(\rx_data[1] ), .B(\rx_data[2] ), .C(\rx_data[0] ), 
         .Z(n14506)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i11831_2_lut_3_lut.init = 16'h8080;
    LUT4 i20881_1_lut_4_lut_4_lut (.A(\rx_data[3] ), .B(n69), .C(n52), 
         .D(n24837), .Z(n22103)) /* synthesis lut_function=(A+!(B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(58[24:46])
    defparam i20881_1_lut_4_lut_4_lut.init = 16'hafbf;
    LUT4 i1_2_lut_rep_442 (.A(\rx_data[3] ), .B(\rx_data[6] ), .Z(n25002)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut_rep_442.init = 16'hbbbb;
    LUT4 i2_3_lut_4_lut (.A(\rx_data[3] ), .B(\rx_data[6] ), .C(\rx_data[5] ), 
         .D(\rx_data[4] ), .Z(n12)) /* synthesis lut_function=(A+((C+!(D))+!B)) */ ;
    defparam i2_3_lut_4_lut.init = 16'hfbff;
    LUT4 i1_2_lut_rep_277_3_lut_4_lut (.A(\rx_data[3] ), .B(\rx_data[6] ), 
         .C(\rx_data[5] ), .D(\rx_data[4] ), .Z(n24837)) /* synthesis lut_function=(A+(((D)+!C)+!B)) */ ;
    defparam i1_2_lut_rep_277_3_lut_4_lut.init = 16'hffbf;
    LUT4 i1_2_lut_rep_443 (.A(\rx_data[1] ), .B(\rx_data[2] ), .Z(n25003)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_443.init = 16'heeee;
    LUT4 i1_4_lut_4_lut_adj_100 (.A(\rx_data[1] ), .B(\rx_data[2] ), .C(n19464), 
         .D(n24984), .Z(n41)) /* synthesis lut_function=(A (C+(D))+!A (B (D))) */ ;
    defparam i1_4_lut_4_lut_adj_100.init = 16'heea0;
    LUT4 i1_2_lut_3_lut_4_lut (.A(\rx_data[1] ), .B(\rx_data[2] ), .C(n25007), 
         .D(\rx_data[3] ), .Z(n19485)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B !(C))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'hef0f;
    LUT4 i1_4_lut_4_lut_3_lut (.A(\rx_data[1] ), .B(\rx_data[2] ), .C(\rx_data[0] ), 
         .Z(n69)) /* synthesis lut_function=(A (B (C))+!A !(B+(C))) */ ;
    defparam i1_4_lut_4_lut_3_lut.init = 16'h8181;
    LUT4 i10965_2_lut_rep_423_3_lut (.A(\rx_data[1] ), .B(\rx_data[2] ), 
         .C(\rx_data[3] ), .Z(n24983)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i10965_2_lut_rep_423_3_lut.init = 16'he0e0;
    LUT4 i_byte_6__I_0_38_i9_2_lut_3_lut (.A(\rx_data[1] ), .B(\rx_data[2] ), 
         .C(\rx_data[0] ), .Z(n9)) /* synthesis lut_function=(A+(B+!(C))) */ ;
    defparam i_byte_6__I_0_38_i9_2_lut_3_lut.init = 16'hefef;
    LUT4 i17300_2_lut_rep_447 (.A(\rx_data[5] ), .B(\rx_data[4] ), .Z(n25007)) /* synthesis lut_function=(A (B)) */ ;
    defparam i17300_2_lut_rep_447.init = 16'h8888;
    LUT4 i1_2_lut_3_lut (.A(\rx_data[5] ), .B(\rx_data[4] ), .C(\rx_data[3] ), 
         .Z(n19461)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_4_lut_adj_101 (.A(\rx_data[5] ), .B(\rx_data[4] ), 
         .C(\rx_data[3] ), .D(\rx_data[6] ), .Z(n44)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A (C)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_101.init = 16'hf0f8;
    LUT4 i21115_3_lut_rep_424_4_lut (.A(\rx_data[5] ), .B(\rx_data[4] ), 
         .C(\rx_data[3] ), .D(\rx_data[6] ), .Z(n24984)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i21115_3_lut_rep_424_4_lut.init = 16'h0008;
    LUT4 i59_3_lut_4_lut (.A(\rx_data[5] ), .B(\rx_data[4] ), .C(\rx_data[6] ), 
         .D(n53), .Z(n56)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C)) */ ;
    defparam i59_3_lut_4_lut.init = 16'hf707;
    LUT4 i82_3_lut (.A(n64), .B(n47), .C(\rx_data[4] ), .Z(n52)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(65[3] 99[10])
    defparam i82_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_489 (.A(n27586), .B(dec_stb), .Z(i_ref_clk_c_enable_388)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(53[9] 54[46])
    defparam i1_2_lut_rep_489.init = 16'heeee;
    LUT4 i8563_2_lut_3_lut (.A(n27586), .B(dec_stb), .C(dec_bits[4]), 
         .Z(i_ref_clk_c_enable_357)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(53[9] 54[46])
    defparam i8563_2_lut_3_lut.init = 16'he0e0;
    LUT4 i1_2_lut_3_lut_adj_102 (.A(dec_stb), .B(dec_bits[4]), .C(cmd_loaded), 
         .Z(o_pck_stb_N_765)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(60[9] 100[5])
    defparam i1_2_lut_3_lut_adj_102.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_103 (.A(dec_stb), .B(dec_bits[4]), .C(n27586), 
         .Z(i_ref_clk_c_enable_192)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(60[9] 100[5])
    defparam i1_2_lut_3_lut_adj_103.init = 16'hf8f8;
    LUT4 i1_3_lut_4_lut (.A(dec_stb), .B(dec_bits[4]), .C(dec_bits_c[3]), 
         .D(dec_bits_c[2]), .Z(cmd_loaded_N_768)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(60[9] 100[5])
    defparam i1_3_lut_4_lut.init = 16'h0008;
    LUT4 i1_4_lut_adj_104 (.A(\rx_data[5] ), .B(\rx_data[2] ), .C(\rx_data[1] ), 
         .D(\rx_data[0] ), .Z(n47)) /* synthesis lut_function=(!(A+!(B (C (D)+!C !(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(65[3] 99[10])
    defparam i1_4_lut_adj_104.init = 16'h5014;
    
endmodule
//
// Verilog Description of module hbnewline
//

module hbnewline (i_ref_clk_c, n27587, hx_stb, nl_busy, \w_gx_char[1] , 
            w_reset, n27586, \w_gx_char[3] , \w_gx_char[6] , \w_gx_char[5] , 
            n11767, tx_busy, \w_gx_char[4] , \w_gx_char[2] , \w_gx_char[0] , 
            n24992, \lcl_data[1] , \lcl_data_7__N_511[0] , \lcl_data[2] , 
            \lcl_data_7__N_511[1] , \lcl_data[3] , \lcl_data_7__N_511[2] , 
            \lcl_data[4] , \lcl_data_7__N_511[3] , \lcl_data[5] , \lcl_data_7__N_511[4] , 
            \lcl_data[6] , \lcl_data_7__N_511[5] , \lcl_data[7] , \lcl_data_7__N_511[6] , 
            n24890, zero_baud_counter_N_526, zero_baud_counter_N_525, 
            zero_baud_counter, i_ref_clk_c_enable_329, o_busy_N_536, \state[0] , 
            n17568) /* synthesis syn_module_defined=1 */ ;
    input i_ref_clk_c;
    input n27587;
    input hx_stb;
    output nl_busy;
    input \w_gx_char[1] ;
    input w_reset;
    input n27586;
    input \w_gx_char[3] ;
    input \w_gx_char[6] ;
    input \w_gx_char[5] ;
    input n11767;
    input tx_busy;
    input \w_gx_char[4] ;
    input \w_gx_char[2] ;
    input \w_gx_char[0] ;
    output n24992;
    input \lcl_data[1] ;
    output \lcl_data_7__N_511[0] ;
    input \lcl_data[2] ;
    output \lcl_data_7__N_511[1] ;
    input \lcl_data[3] ;
    output \lcl_data_7__N_511[2] ;
    input \lcl_data[4] ;
    output \lcl_data_7__N_511[3] ;
    input \lcl_data[5] ;
    output \lcl_data_7__N_511[4] ;
    input \lcl_data[6] ;
    output \lcl_data_7__N_511[5] ;
    input \lcl_data[7] ;
    output \lcl_data_7__N_511[6] ;
    input n24890;
    input zero_baud_counter_N_526;
    output zero_baud_counter_N_525;
    input zero_baud_counter;
    output i_ref_clk_c_enable_329;
    input o_busy_N_536;
    input \state[0] ;
    output n17568;
    
    wire i_ref_clk_c /* synthesis SET_AS_NETWORK=i_ref_clk_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(22[12:21])
    
    wire tx_stb, o_nl_stb_N_1315, last_cr, last_cr_N_1323;
    wire [6:0]o_nl_byte_6__N_1302;
    wire [7:0]tx_data;   // d:/documents/git_local/fm_modulator/rtl/top.v(58[12:19])
    
    wire i_ref_clk_c_enable_197;
    wire [6:0]o_nl_byte_6__N_1295;
    
    wire loaded, n24865, cr_state, cr_state_N_1331;
    wire [6:0]n32;
    
    wire n24975, n25287, n25288, n23954, n23955;
    
    FD1S3IX o_nl_stb_46 (.D(o_nl_stb_N_1315), .CK(i_ref_clk_c), .CD(n27587), 
            .Q(tx_stb)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=12, LSE_RCOL=40, LSE_LLINE=138, LSE_RLINE=139 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam o_nl_stb_46.GSR = "DISABLED";
    FD1S3JX last_cr_45 (.D(last_cr_N_1323), .CK(i_ref_clk_c), .PD(n27587), 
            .Q(last_cr)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=12, LSE_RCOL=40, LSE_LLINE=138, LSE_RLINE=139 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam last_cr_45.GSR = "DISABLED";
    LUT4 i10710_3_lut_4_lut (.A(hx_stb), .B(nl_busy), .C(\w_gx_char[1] ), 
         .D(last_cr), .Z(o_nl_byte_6__N_1302[1])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(90[16:37])
    defparam i10710_3_lut_4_lut.init = 16'hfd20;
    FD1P3JX o_nl_byte_i2 (.D(o_nl_byte_6__N_1302[1]), .SP(i_ref_clk_c_enable_197), 
            .PD(w_reset), .CK(i_ref_clk_c), .Q(tx_data[1])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=12, LSE_RCOL=40, LSE_LLINE=138, LSE_RLINE=139 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam o_nl_byte_i2.GSR = "DISABLED";
    FD1P3JX o_nl_byte_i3 (.D(o_nl_byte_6__N_1302[2]), .SP(i_ref_clk_c_enable_197), 
            .PD(w_reset), .CK(i_ref_clk_c), .Q(tx_data[2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=12, LSE_RCOL=40, LSE_LLINE=138, LSE_RLINE=139 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam o_nl_byte_i3.GSR = "DISABLED";
    FD1P3AY o_nl_byte_i4 (.D(o_nl_byte_6__N_1295[3]), .SP(i_ref_clk_c_enable_197), 
            .CK(i_ref_clk_c), .Q(tx_data[3])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=12, LSE_RCOL=40, LSE_LLINE=138, LSE_RLINE=139 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam o_nl_byte_i4.GSR = "DISABLED";
    FD1P3JX o_nl_byte_i5 (.D(o_nl_byte_6__N_1302[4]), .SP(i_ref_clk_c_enable_197), 
            .PD(w_reset), .CK(i_ref_clk_c), .Q(tx_data[4])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=12, LSE_RCOL=40, LSE_LLINE=138, LSE_RLINE=139 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam o_nl_byte_i5.GSR = "DISABLED";
    FD1P3JX o_nl_byte_i6 (.D(o_nl_byte_6__N_1302[5]), .SP(i_ref_clk_c_enable_197), 
            .PD(w_reset), .CK(i_ref_clk_c), .Q(tx_data[5])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=12, LSE_RCOL=40, LSE_LLINE=138, LSE_RLINE=139 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam o_nl_byte_i6.GSR = "DISABLED";
    FD1P3JX o_nl_byte_i7 (.D(o_nl_byte_6__N_1302[6]), .SP(i_ref_clk_c_enable_197), 
            .PD(w_reset), .CK(i_ref_clk_c), .Q(tx_data[6])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=12, LSE_RCOL=40, LSE_LLINE=138, LSE_RLINE=139 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam o_nl_byte_i7.GSR = "DISABLED";
    LUT4 i2_3_lut_4_lut (.A(hx_stb), .B(nl_busy), .C(n27586), .D(\w_gx_char[3] ), 
         .Z(o_nl_byte_6__N_1295[3])) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(90[16:37])
    defparam i2_3_lut_4_lut.init = 16'hfffd;
    FD1P3IX loaded_47 (.D(n24865), .SP(i_ref_clk_c_enable_197), .CD(w_reset), 
            .CK(i_ref_clk_c), .Q(loaded)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=12, LSE_RCOL=40, LSE_LLINE=138, LSE_RLINE=139 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam loaded_47.GSR = "DISABLED";
    FD1P3IX cr_state_44 (.D(cr_state_N_1331), .SP(i_ref_clk_c_enable_197), 
            .CD(n27587), .CK(i_ref_clk_c), .Q(cr_state)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=12, LSE_RCOL=40, LSE_LLINE=138, LSE_RLINE=139 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam cr_state_44.GSR = "DISABLED";
    FD1P3JX o_nl_byte_i1 (.D(o_nl_byte_6__N_1302[0]), .SP(i_ref_clk_c_enable_197), 
            .PD(n27587), .CK(i_ref_clk_c), .Q(tx_data[0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=12, LSE_RCOL=40, LSE_LLINE=138, LSE_RLINE=139 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam o_nl_byte_i1.GSR = "DISABLED";
    LUT4 mux_24_i7_3_lut_4_lut (.A(hx_stb), .B(nl_busy), .C(\w_gx_char[6] ), 
         .D(n32[4]), .Z(o_nl_byte_6__N_1302[6])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(90[16:37])
    defparam mux_24_i7_3_lut_4_lut.init = 16'hfd20;
    LUT4 i10707_3_lut_4_lut (.A(hx_stb), .B(nl_busy), .C(\w_gx_char[5] ), 
         .D(n32[4]), .Z(o_nl_byte_6__N_1302[5])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(90[16:37])
    defparam i10707_3_lut_4_lut.init = 16'hfd20;
    LUT4 cr_state_I_41_3_lut_4_lut (.A(hx_stb), .B(nl_busy), .C(n11767), 
         .D(last_cr), .Z(cr_state_N_1331)) /* synthesis lut_function=(!(A (B (D)+!B (C))+!A (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(90[16:37])
    defparam cr_state_I_41_3_lut_4_lut.init = 16'h02df;
    LUT4 i_stb_I_0_2_lut_rep_415 (.A(hx_stb), .B(nl_busy), .Z(n24975)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(90[16:37])
    defparam i_stb_I_0_2_lut_rep_415.init = 16'h2222;
    PFUMX i23052 (.BLUT(n25287), .ALUT(n25288), .C0(last_cr), .Z(last_cr_N_1323));
    LUT4 i2_3_lut_4_lut_adj_91 (.A(hx_stb), .B(nl_busy), .C(n27586), .D(tx_busy), 
         .Z(i_ref_clk_c_enable_197)) /* synthesis lut_function=(A ((C+!(D))+!B)+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(90[16:37])
    defparam i2_3_lut_4_lut_adj_91.init = 16'hf2ff;
    LUT4 tx_stb_bdd_2_lut_23394 (.A(tx_stb), .B(hx_stb), .Z(n23954)) /* synthesis lut_function=(A+(B)) */ ;
    defparam tx_stb_bdd_2_lut_23394.init = 16'heeee;
    LUT4 tx_stb_bdd_3_lut (.A(hx_stb), .B(last_cr), .C(cr_state), .Z(n23955)) /* synthesis lut_function=(A (B+!(C))+!A ((C)+!B)) */ ;
    defparam tx_stb_bdd_3_lut.init = 16'hdbdb;
    LUT4 i1_2_lut (.A(last_cr), .B(cr_state), .Z(n32[4])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam i1_2_lut.init = 16'h2222;
    LUT4 mux_24_i5_3_lut_4_lut (.A(hx_stb), .B(nl_busy), .C(\w_gx_char[4] ), 
         .D(n32[4]), .Z(o_nl_byte_6__N_1302[4])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(90[16:37])
    defparam mux_24_i5_3_lut_4_lut.init = 16'hfd20;
    LUT4 i10945_3_lut_rep_305_4_lut (.A(hx_stb), .B(nl_busy), .C(cr_state), 
         .D(last_cr), .Z(n24865)) /* synthesis lut_function=(A ((C (D))+!B)+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(90[16:37])
    defparam i10945_3_lut_rep_305_4_lut.init = 16'hf222;
    LUT4 last_cr_I_39_4_lut_then_3_lut (.A(n11767), .B(hx_stb), .C(nl_busy), 
         .Z(n25288)) /* synthesis lut_function=(((C)+!B)+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(97[12] 120[6])
    defparam last_cr_I_39_4_lut_then_3_lut.init = 16'hf7f7;
    LUT4 last_cr_I_39_4_lut_else_3_lut (.A(n11767), .B(tx_busy), .C(hx_stb), 
         .D(nl_busy), .Z(n25287)) /* synthesis lut_function=(!(A (B+(C))+!A (B ((D)+!C)+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(97[12] 120[6])
    defparam last_cr_I_39_4_lut_else_3_lut.init = 16'h0353;
    LUT4 i1_3_lut_4_lut (.A(last_cr), .B(n24975), .C(cr_state), .D(\w_gx_char[2] ), 
         .Z(o_nl_byte_6__N_1302[2])) /* synthesis lut_function=(A (B (D)+!B !(C))+!A ((D)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(97[12] 120[6])
    defparam i1_3_lut_4_lut.init = 16'hdf13;
    LUT4 i1_3_lut_4_lut_adj_92 (.A(last_cr), .B(n24975), .C(cr_state), 
         .D(\w_gx_char[0] ), .Z(o_nl_byte_6__N_1302[0])) /* synthesis lut_function=(A (B (D)+!B !(C))+!A ((D)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(97[12] 120[6])
    defparam i1_3_lut_4_lut_adj_92.init = 16'hdf13;
    LUT4 i1_2_lut_rep_432 (.A(tx_stb), .B(tx_busy), .Z(n24992)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam i1_2_lut_rep_432.init = 16'h2222;
    LUT4 lcl_data_7__I_0_i1_3_lut_4_lut (.A(tx_stb), .B(tx_busy), .C(tx_data[0]), 
         .D(\lcl_data[1] ), .Z(\lcl_data_7__N_511[0] )) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam lcl_data_7__I_0_i1_3_lut_4_lut.init = 16'hfd20;
    LUT4 lcl_data_7__I_0_i2_3_lut_4_lut (.A(tx_stb), .B(tx_busy), .C(tx_data[1]), 
         .D(\lcl_data[2] ), .Z(\lcl_data_7__N_511[1] )) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam lcl_data_7__I_0_i2_3_lut_4_lut.init = 16'hfd20;
    LUT4 lcl_data_7__I_0_i3_3_lut_4_lut (.A(tx_stb), .B(tx_busy), .C(tx_data[2]), 
         .D(\lcl_data[3] ), .Z(\lcl_data_7__N_511[2] )) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam lcl_data_7__I_0_i3_3_lut_4_lut.init = 16'hfd20;
    LUT4 lcl_data_7__I_0_i4_3_lut_4_lut (.A(tx_stb), .B(tx_busy), .C(tx_data[3]), 
         .D(\lcl_data[4] ), .Z(\lcl_data_7__N_511[3] )) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam lcl_data_7__I_0_i4_3_lut_4_lut.init = 16'hfd20;
    LUT4 lcl_data_7__I_0_i5_3_lut_4_lut (.A(tx_stb), .B(tx_busy), .C(tx_data[4]), 
         .D(\lcl_data[5] ), .Z(\lcl_data_7__N_511[4] )) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam lcl_data_7__I_0_i5_3_lut_4_lut.init = 16'hfd20;
    LUT4 lcl_data_7__I_0_i6_3_lut_4_lut (.A(tx_stb), .B(tx_busy), .C(tx_data[5]), 
         .D(\lcl_data[6] ), .Z(\lcl_data_7__N_511[5] )) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam lcl_data_7__I_0_i6_3_lut_4_lut.init = 16'hfd20;
    LUT4 lcl_data_7__I_0_i7_3_lut_4_lut (.A(tx_stb), .B(tx_busy), .C(tx_data[6]), 
         .D(\lcl_data[7] ), .Z(\lcl_data_7__N_511[6] )) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam lcl_data_7__I_0_i7_3_lut_4_lut.init = 16'hfd20;
    LUT4 zero_baud_counter_I_0_51_3_lut_4_lut (.A(tx_stb), .B(tx_busy), 
         .C(n24890), .D(zero_baud_counter_N_526), .Z(zero_baud_counter_N_525)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam zero_baud_counter_I_0_51_3_lut_4_lut.init = 16'hdfd0;
    LUT4 i519_2_lut_3_lut (.A(tx_stb), .B(tx_busy), .C(zero_baud_counter), 
         .Z(i_ref_clk_c_enable_329)) /* synthesis lut_function=(A ((C)+!B)+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam i519_2_lut_3_lut.init = 16'hf2f2;
    LUT4 state_504_mux_6_i1_3_lut_4_lut (.A(tx_stb), .B(tx_busy), .C(o_busy_N_536), 
         .D(\state[0] ), .Z(n17568)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam state_504_mux_6_i1_3_lut_4_lut.init = 16'hd0df;
    PFUMX i22335 (.BLUT(n23955), .ALUT(n23954), .C0(tx_busy), .Z(o_nl_stb_N_1315));
    LUT4 o_nl_busy_I_0_57_4_lut (.A(tx_stb), .B(cr_state), .C(loaded), 
         .D(tx_busy), .Z(nl_busy)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A !((D)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(123[21] 124[30])
    defparam o_nl_busy_I_0_57_4_lut.init = 16'ha0cc;
    
endmodule
//
// Verilog Description of module hbints
//

module hbints (int_word, i_ref_clk_c, ow_word, n27586, n25186, int_stb, 
            n27587, ow_stb) /* synthesis syn_module_defined=1 */ ;
    output [33:0]int_word;
    input i_ref_clk_c;
    input [33:0]ow_word;
    input n27586;
    input n25186;
    output int_stb;
    input n27587;
    input ow_stb;
    
    wire i_ref_clk_c /* synthesis SET_AS_NETWORK=i_ref_clk_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(22[12:21])
    
    wire i_ref_clk_c_enable_420, n12732, n25028, loaded, i_ref_clk_c_enable_412, 
        i_ref_clk_c_enable_413;
    
    FD1P3IX o_int_word_i8 (.D(ow_word[8]), .SP(i_ref_clk_c_enable_420), 
            .CD(n12732), .CK(i_ref_clk_c), .Q(int_word[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i8.GSR = "DISABLED";
    FD1P3JX o_int_word_i33 (.D(ow_word[33]), .SP(i_ref_clk_c_enable_420), 
            .PD(n12732), .CK(i_ref_clk_c), .Q(int_word[33])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i33.GSR = "DISABLED";
    FD1P3JX o_int_word_i32 (.D(ow_word[32]), .SP(i_ref_clk_c_enable_420), 
            .PD(n12732), .CK(i_ref_clk_c), .Q(int_word[32])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i32.GSR = "DISABLED";
    FD1P3IX o_int_word_i31 (.D(ow_word[31]), .SP(i_ref_clk_c_enable_420), 
            .CD(n12732), .CK(i_ref_clk_c), .Q(int_word[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i31.GSR = "DISABLED";
    FD1P3JX o_int_word_i30 (.D(ow_word[30]), .SP(i_ref_clk_c_enable_420), 
            .PD(n12732), .CK(i_ref_clk_c), .Q(int_word[30])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i30.GSR = "DISABLED";
    FD1P3IX o_int_word_i29 (.D(ow_word[29]), .SP(i_ref_clk_c_enable_420), 
            .CD(n12732), .CK(i_ref_clk_c), .Q(int_word[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i29.GSR = "DISABLED";
    LUT4 i2_3_lut_4_lut (.A(n27586), .B(n25028), .C(n25186), .D(loaded), 
         .Z(i_ref_clk_c_enable_412)) /* synthesis lut_function=(A+(B+!(C (D)))) */ ;
    defparam i2_3_lut_4_lut.init = 16'hefff;
    FD1P3IX o_int_word_i28 (.D(ow_word[28]), .SP(i_ref_clk_c_enable_420), 
            .CD(n12732), .CK(i_ref_clk_c), .Q(int_word[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i28.GSR = "DISABLED";
    LUT4 i1_2_lut_3_lut_4_lut (.A(int_stb), .B(n25186), .C(n25028), .D(n27586), 
         .Z(i_ref_clk_c_enable_413)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(77[12:34])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfff2;
    FD1P3IX o_int_word_i7 (.D(ow_word[7]), .SP(i_ref_clk_c_enable_420), 
            .CD(n12732), .CK(i_ref_clk_c), .Q(int_word[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i7.GSR = "DISABLED";
    FD1P3IX o_int_word_i27 (.D(ow_word[27]), .SP(i_ref_clk_c_enable_420), 
            .CD(n12732), .CK(i_ref_clk_c), .Q(int_word[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i27.GSR = "DISABLED";
    FD1P3IX o_int_word_i26 (.D(ow_word[26]), .SP(i_ref_clk_c_enable_420), 
            .CD(n12732), .CK(i_ref_clk_c), .Q(int_word[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i26.GSR = "DISABLED";
    FD1P3IX o_int_word_i6 (.D(ow_word[6]), .SP(i_ref_clk_c_enable_420), 
            .CD(n12732), .CK(i_ref_clk_c), .Q(int_word[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i6.GSR = "DISABLED";
    FD1P3IX o_int_word_i25 (.D(ow_word[25]), .SP(i_ref_clk_c_enable_420), 
            .CD(n12732), .CK(i_ref_clk_c), .Q(int_word[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i25.GSR = "DISABLED";
    FD1P3IX o_int_word_i5 (.D(ow_word[5]), .SP(i_ref_clk_c_enable_420), 
            .CD(n12732), .CK(i_ref_clk_c), .Q(int_word[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i5.GSR = "DISABLED";
    FD1P3IX o_int_word_i24 (.D(ow_word[24]), .SP(i_ref_clk_c_enable_420), 
            .CD(n12732), .CK(i_ref_clk_c), .Q(int_word[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i24.GSR = "DISABLED";
    FD1P3IX o_int_word_i4 (.D(ow_word[4]), .SP(i_ref_clk_c_enable_420), 
            .CD(n12732), .CK(i_ref_clk_c), .Q(int_word[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i4.GSR = "DISABLED";
    FD1P3IX o_int_word_i3 (.D(ow_word[3]), .SP(i_ref_clk_c_enable_420), 
            .CD(n12732), .CK(i_ref_clk_c), .Q(int_word[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i3.GSR = "DISABLED";
    FD1P3IX o_int_word_i23 (.D(ow_word[23]), .SP(i_ref_clk_c_enable_420), 
            .CD(n12732), .CK(i_ref_clk_c), .Q(int_word[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i23.GSR = "DISABLED";
    FD1P3IX o_int_word_i22 (.D(ow_word[22]), .SP(i_ref_clk_c_enable_420), 
            .CD(n12732), .CK(i_ref_clk_c), .Q(int_word[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i22.GSR = "DISABLED";
    FD1P3IX o_int_word_i2 (.D(ow_word[2]), .SP(i_ref_clk_c_enable_420), 
            .CD(n12732), .CK(i_ref_clk_c), .Q(int_word[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i2.GSR = "DISABLED";
    FD1P3IX o_int_word_i1 (.D(ow_word[1]), .SP(i_ref_clk_c_enable_420), 
            .CD(n12732), .CK(i_ref_clk_c), .Q(int_word[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i1.GSR = "DISABLED";
    FD1P3IX o_int_word_i21 (.D(ow_word[21]), .SP(i_ref_clk_c_enable_420), 
            .CD(n12732), .CK(i_ref_clk_c), .Q(int_word[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i21.GSR = "DISABLED";
    FD1P3IX o_int_word_i0 (.D(ow_word[0]), .SP(i_ref_clk_c_enable_420), 
            .CD(n12732), .CK(i_ref_clk_c), .Q(int_word[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i0.GSR = "DISABLED";
    FD1P3IX o_int_word_i20 (.D(ow_word[20]), .SP(i_ref_clk_c_enable_420), 
            .CD(n12732), .CK(i_ref_clk_c), .Q(int_word[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i20.GSR = "DISABLED";
    FD1P3IX o_int_word_i19 (.D(ow_word[19]), .SP(i_ref_clk_c_enable_420), 
            .CD(n12732), .CK(i_ref_clk_c), .Q(int_word[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i19.GSR = "DISABLED";
    FD1P3IX o_int_word_i18 (.D(ow_word[18]), .SP(i_ref_clk_c_enable_420), 
            .CD(n12732), .CK(i_ref_clk_c), .Q(int_word[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i18.GSR = "DISABLED";
    FD1P3IX o_int_word_i17 (.D(ow_word[17]), .SP(i_ref_clk_c_enable_420), 
            .CD(n12732), .CK(i_ref_clk_c), .Q(int_word[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i17.GSR = "DISABLED";
    FD1P3IX o_int_word_i16 (.D(ow_word[16]), .SP(i_ref_clk_c_enable_420), 
            .CD(n12732), .CK(i_ref_clk_c), .Q(int_word[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i16.GSR = "DISABLED";
    FD1P3IX o_int_word_i15 (.D(ow_word[15]), .SP(i_ref_clk_c_enable_420), 
            .CD(n12732), .CK(i_ref_clk_c), .Q(int_word[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i15.GSR = "DISABLED";
    FD1P3IX o_int_word_i14 (.D(ow_word[14]), .SP(i_ref_clk_c_enable_420), 
            .CD(n12732), .CK(i_ref_clk_c), .Q(int_word[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i14.GSR = "DISABLED";
    FD1P3IX o_int_stb_58 (.D(n25028), .SP(i_ref_clk_c_enable_412), .CD(n27587), 
            .CK(i_ref_clk_c), .Q(int_stb)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(90[9] 98[22])
    defparam o_int_stb_58.GSR = "DISABLED";
    FD1P3IX loaded_57 (.D(n25028), .SP(i_ref_clk_c_enable_413), .CD(n27587), 
            .CK(i_ref_clk_c), .Q(loaded)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(81[9] 87[19])
    defparam loaded_57.GSR = "DISABLED";
    FD1P3IX o_int_word_i13 (.D(ow_word[13]), .SP(i_ref_clk_c_enable_420), 
            .CD(n12732), .CK(i_ref_clk_c), .Q(int_word[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i13.GSR = "DISABLED";
    FD1P3IX o_int_word_i12 (.D(ow_word[12]), .SP(i_ref_clk_c_enable_420), 
            .CD(n12732), .CK(i_ref_clk_c), .Q(int_word[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i12.GSR = "DISABLED";
    FD1P3IX o_int_word_i11 (.D(ow_word[11]), .SP(i_ref_clk_c_enable_420), 
            .CD(n12732), .CK(i_ref_clk_c), .Q(int_word[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i11.GSR = "DISABLED";
    FD1P3IX o_int_word_i10 (.D(ow_word[10]), .SP(i_ref_clk_c_enable_420), 
            .CD(n12732), .CK(i_ref_clk_c), .Q(int_word[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i10.GSR = "DISABLED";
    FD1P3IX o_int_word_i9 (.D(ow_word[9]), .SP(i_ref_clk_c_enable_420), 
            .CD(n12732), .CK(i_ref_clk_c), .Q(int_word[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i9.GSR = "DISABLED";
    LUT4 i_stb_I_0_3_lut_rep_468 (.A(ow_stb), .B(int_stb), .C(loaded), 
         .Z(n25028)) /* synthesis lut_function=(!((B (C))+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(93[12:34])
    defparam i_stb_I_0_3_lut_rep_468.init = 16'h2a2a;
    LUT4 i21051_2_lut_3_lut_3_lut_4_lut (.A(ow_stb), .B(int_stb), .C(loaded), 
         .D(n25186), .Z(n12732)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A (B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(93[12:34])
    defparam i21051_2_lut_3_lut_3_lut_4_lut.init = 16'h11d5;
    LUT4 i1_2_lut_3_lut_4_lut_adj_90 (.A(ow_stb), .B(int_stb), .C(loaded), 
         .D(n25186), .Z(i_ref_clk_c_enable_420)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(93[12:34])
    defparam i1_2_lut_3_lut_4_lut_adj_90.init = 16'h3bff;
    
endmodule
//
// Verilog Description of module hbidle
//

module hbidle (idl_word, i_ref_clk_c, int_word, hb_busy, int_stb, 
            idl_stb, n25186, n27586, n27587) /* synthesis syn_module_defined=1 */ ;
    output [33:0]idl_word;
    input i_ref_clk_c;
    input [33:0]int_word;
    input hb_busy;
    input int_stb;
    output idl_stb;
    output n25186;
    input n27586;
    input n27587;
    
    wire i_ref_clk_c /* synthesis SET_AS_NETWORK=i_ref_clk_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(22[12:21])
    
    wire i_ref_clk_c_enable_353, n12774, n24987, i_ref_clk_c_enable_409;
    
    FD1P3IX o_idl_word_i8 (.D(int_word[8]), .SP(i_ref_clk_c_enable_353), 
            .CD(n12774), .CK(i_ref_clk_c), .Q(idl_word[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i8.GSR = "DISABLED";
    FD1P3IX o_idl_word_i7 (.D(int_word[7]), .SP(i_ref_clk_c_enable_353), 
            .CD(n12774), .CK(i_ref_clk_c), .Q(idl_word[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i7.GSR = "DISABLED";
    FD1P3IX o_idl_word_i6 (.D(int_word[6]), .SP(i_ref_clk_c_enable_353), 
            .CD(n12774), .CK(i_ref_clk_c), .Q(idl_word[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i6.GSR = "DISABLED";
    FD1P3IX o_idl_word_i5 (.D(int_word[5]), .SP(i_ref_clk_c_enable_353), 
            .CD(n12774), .CK(i_ref_clk_c), .Q(idl_word[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i5.GSR = "DISABLED";
    FD1P3IX o_idl_word_i4 (.D(int_word[4]), .SP(i_ref_clk_c_enable_353), 
            .CD(n12774), .CK(i_ref_clk_c), .Q(idl_word[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i4.GSR = "DISABLED";
    FD1P3IX o_idl_word_i3 (.D(int_word[3]), .SP(i_ref_clk_c_enable_353), 
            .CD(n12774), .CK(i_ref_clk_c), .Q(idl_word[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i3.GSR = "DISABLED";
    FD1P3IX o_idl_word_i2 (.D(int_word[2]), .SP(i_ref_clk_c_enable_353), 
            .CD(n12774), .CK(i_ref_clk_c), .Q(idl_word[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i2.GSR = "DISABLED";
    FD1P3IX o_idl_word_i1 (.D(int_word[1]), .SP(i_ref_clk_c_enable_353), 
            .CD(n12774), .CK(i_ref_clk_c), .Q(idl_word[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i1.GSR = "DISABLED";
    FD1P3JX o_idl_word_i33 (.D(int_word[33]), .SP(i_ref_clk_c_enable_353), 
            .PD(n12774), .CK(i_ref_clk_c), .Q(idl_word[33])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i33.GSR = "DISABLED";
    FD1P3JX o_idl_word_i32 (.D(int_word[32]), .SP(i_ref_clk_c_enable_353), 
            .PD(n12774), .CK(i_ref_clk_c), .Q(idl_word[32])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i32.GSR = "DISABLED";
    FD1P3IX o_idl_word_i31 (.D(int_word[31]), .SP(i_ref_clk_c_enable_353), 
            .CD(n12774), .CK(i_ref_clk_c), .Q(idl_word[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i31.GSR = "DISABLED";
    FD1P3JX o_idl_word_i30 (.D(int_word[30]), .SP(i_ref_clk_c_enable_353), 
            .PD(n12774), .CK(i_ref_clk_c), .Q(idl_word[30])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i30.GSR = "DISABLED";
    FD1P3JX o_idl_word_i29 (.D(int_word[29]), .SP(i_ref_clk_c_enable_353), 
            .PD(n12774), .CK(i_ref_clk_c), .Q(idl_word[29])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i29.GSR = "DISABLED";
    FD1P3IX o_idl_word_i28 (.D(int_word[28]), .SP(i_ref_clk_c_enable_353), 
            .CD(n12774), .CK(i_ref_clk_c), .Q(idl_word[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i28.GSR = "DISABLED";
    FD1P3IX o_idl_word_i27 (.D(int_word[27]), .SP(i_ref_clk_c_enable_353), 
            .CD(n12774), .CK(i_ref_clk_c), .Q(idl_word[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i27.GSR = "DISABLED";
    FD1P3IX o_idl_word_i26 (.D(int_word[26]), .SP(i_ref_clk_c_enable_353), 
            .CD(n12774), .CK(i_ref_clk_c), .Q(idl_word[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i26.GSR = "DISABLED";
    FD1P3IX o_idl_word_i25 (.D(int_word[25]), .SP(i_ref_clk_c_enable_353), 
            .CD(n12774), .CK(i_ref_clk_c), .Q(idl_word[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i25.GSR = "DISABLED";
    FD1P3IX o_idl_word_i24 (.D(int_word[24]), .SP(i_ref_clk_c_enable_353), 
            .CD(n12774), .CK(i_ref_clk_c), .Q(idl_word[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i24.GSR = "DISABLED";
    FD1P3IX o_idl_word_i23 (.D(int_word[23]), .SP(i_ref_clk_c_enable_353), 
            .CD(n12774), .CK(i_ref_clk_c), .Q(idl_word[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i23.GSR = "DISABLED";
    FD1P3IX o_idl_word_i22 (.D(int_word[22]), .SP(i_ref_clk_c_enable_353), 
            .CD(n12774), .CK(i_ref_clk_c), .Q(idl_word[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i22.GSR = "DISABLED";
    FD1P3IX o_idl_word_i21 (.D(int_word[21]), .SP(i_ref_clk_c_enable_353), 
            .CD(n12774), .CK(i_ref_clk_c), .Q(idl_word[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i21.GSR = "DISABLED";
    FD1P3IX o_idl_word_i20 (.D(int_word[20]), .SP(i_ref_clk_c_enable_353), 
            .CD(n12774), .CK(i_ref_clk_c), .Q(idl_word[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i20.GSR = "DISABLED";
    FD1P3IX o_idl_word_i19 (.D(int_word[19]), .SP(i_ref_clk_c_enable_353), 
            .CD(n12774), .CK(i_ref_clk_c), .Q(idl_word[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i19.GSR = "DISABLED";
    FD1P3IX o_idl_word_i18 (.D(int_word[18]), .SP(i_ref_clk_c_enable_353), 
            .CD(n12774), .CK(i_ref_clk_c), .Q(idl_word[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i18.GSR = "DISABLED";
    FD1P3IX o_idl_word_i0 (.D(int_word[0]), .SP(i_ref_clk_c_enable_353), 
            .CD(n12774), .CK(i_ref_clk_c), .Q(idl_word[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i0.GSR = "DISABLED";
    LUT4 i21083_2_lut (.A(hb_busy), .B(int_stb), .Z(n12774)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i21083_2_lut.init = 16'h1111;
    LUT4 o_idl_stb_I_0_30_2_lut_rep_626 (.A(idl_stb), .B(hb_busy), .Z(n25186)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(97[22:43])
    defparam o_idl_stb_I_0_30_2_lut_rep_626.init = 16'h8888;
    LUT4 o_int_stb_I_0_66_2_lut_rep_427_3_lut (.A(idl_stb), .B(hb_busy), 
         .C(int_stb), .Z(n24987)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(97[22:43])
    defparam o_int_stb_I_0_66_2_lut_rep_427_3_lut.init = 16'h7070;
    LUT4 i2_3_lut_4_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(n27586), .D(int_stb), 
         .Z(i_ref_clk_c_enable_409)) /* synthesis lut_function=(A ((C)+!B)+!A ((C+(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(97[22:43])
    defparam i2_3_lut_4_lut_4_lut.init = 16'hf7f3;
    LUT4 i1_2_lut_3_lut_3_lut (.A(idl_stb), .B(hb_busy), .C(int_stb), 
         .Z(i_ref_clk_c_enable_353)) /* synthesis lut_function=(!(A (B)+!A !((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(97[22:43])
    defparam i1_2_lut_3_lut_3_lut.init = 16'h7373;
    FD1P3IX o_idl_word_i12 (.D(int_word[12]), .SP(i_ref_clk_c_enable_353), 
            .CD(n12774), .CK(i_ref_clk_c), .Q(idl_word[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i12.GSR = "DISABLED";
    FD1P3IX o_idl_word_i17 (.D(int_word[17]), .SP(i_ref_clk_c_enable_353), 
            .CD(n12774), .CK(i_ref_clk_c), .Q(idl_word[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i17.GSR = "DISABLED";
    FD1P3IX o_idl_word_i16 (.D(int_word[16]), .SP(i_ref_clk_c_enable_353), 
            .CD(n12774), .CK(i_ref_clk_c), .Q(idl_word[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i16.GSR = "DISABLED";
    FD1P3IX o_idl_word_i15 (.D(int_word[15]), .SP(i_ref_clk_c_enable_353), 
            .CD(n12774), .CK(i_ref_clk_c), .Q(idl_word[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i15.GSR = "DISABLED";
    FD1P3IX o_idl_word_i14 (.D(int_word[14]), .SP(i_ref_clk_c_enable_353), 
            .CD(n12774), .CK(i_ref_clk_c), .Q(idl_word[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i14.GSR = "DISABLED";
    FD1P3IX o_idl_word_i13 (.D(int_word[13]), .SP(i_ref_clk_c_enable_353), 
            .CD(n12774), .CK(i_ref_clk_c), .Q(idl_word[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i13.GSR = "DISABLED";
    FD1P3IX o_idl_word_i11 (.D(int_word[11]), .SP(i_ref_clk_c_enable_353), 
            .CD(n12774), .CK(i_ref_clk_c), .Q(idl_word[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i11.GSR = "DISABLED";
    FD1P3IX o_idl_word_i10 (.D(int_word[10]), .SP(i_ref_clk_c_enable_353), 
            .CD(n12774), .CK(i_ref_clk_c), .Q(idl_word[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i10.GSR = "DISABLED";
    FD1P3IX o_idl_word_i9 (.D(int_word[9]), .SP(i_ref_clk_c_enable_353), 
            .CD(n12774), .CK(i_ref_clk_c), .Q(idl_word[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i9.GSR = "DISABLED";
    FD1P3IX o_idl_stb_28 (.D(n24987), .SP(i_ref_clk_c_enable_409), .CD(n27587), 
            .CK(i_ref_clk_c), .Q(idl_stb)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(80[9] 88[22])
    defparam o_idl_stb_28.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module fm_generator_wb_slave
//

module fm_generator_wb_slave (i_ref_clk_c, i_ref_clk_c_enable_106, i_resetb_N_301, 
            wb_odata, i_ref_clk_c_enable_66, i_ref_clk_c_enable_98, wb_fm_data, 
            wb_fm_ack, wb_fm_data_31__N_63, GND_net, \wb_addr[1] , \wb_addr[0] , 
            \power_counter[1] , \smpl_register[1] , n2139, i_resetb_c, 
            n24803, n2, \smpl_register[5] , n24788, n2_adj_1, \smpl_register[29] , 
            n24795, n2_adj_2, \smpl_register[20] , n24794, n2_adj_3, 
            \smpl_register[18] , n24793, n2_adj_4, \smpl_register[17] , 
            n24792, n2_adj_5, \smpl_register[16] , n24791, n2_adj_6, 
            \smpl_register[10] , n24790, n2_adj_7, \smpl_register[9] , 
            n24789, o_baseband_i_c_15, o_baseband_i_c_14, o_baseband_i_c_13, 
            o_baseband_i_c_12, o_baseband_i_c_11, o_baseband_i_c_10, n3607, 
            o_baseband_q_c_7, o_baseband_i_c_7, o_baseband_i_c_8, n27529, 
            o_baseband_q_c_15, o_baseband_q_c_14, o_baseband_q_c_13, o_baseband_q_c_12, 
            o_baseband_q_c_11, o_baseband_q_c_10, n3608, o_baseband_q_c_8) /* synthesis syn_module_defined=1 */ ;
    input i_ref_clk_c;
    input i_ref_clk_c_enable_106;
    input i_resetb_N_301;
    input [31:0]wb_odata;
    input i_ref_clk_c_enable_66;
    input i_ref_clk_c_enable_98;
    output [31:0]wb_fm_data;
    output wb_fm_ack;
    input wb_fm_data_31__N_63;
    input GND_net;
    input \wb_addr[1] ;
    input \wb_addr[0] ;
    input \power_counter[1] ;
    input \smpl_register[1] ;
    output n2139;
    input i_resetb_c;
    input n24803;
    input n2;
    input \smpl_register[5] ;
    output n24788;
    input n2_adj_1;
    input \smpl_register[29] ;
    output n24795;
    input n2_adj_2;
    input \smpl_register[20] ;
    output n24794;
    input n2_adj_3;
    input \smpl_register[18] ;
    output n24793;
    input n2_adj_4;
    input \smpl_register[17] ;
    output n24792;
    input n2_adj_5;
    input \smpl_register[16] ;
    output n24791;
    input n2_adj_6;
    input \smpl_register[10] ;
    output n24790;
    input n2_adj_7;
    input \smpl_register[9] ;
    output n24789;
    output o_baseband_i_c_15;
    output o_baseband_i_c_14;
    output o_baseband_i_c_13;
    output o_baseband_i_c_12;
    output o_baseband_i_c_11;
    output o_baseband_i_c_10;
    output n3607;
    output o_baseband_q_c_7;
    output o_baseband_i_c_7;
    output o_baseband_i_c_8;
    input n27529;
    output o_baseband_q_c_15;
    output o_baseband_q_c_14;
    output o_baseband_q_c_13;
    output o_baseband_q_c_12;
    output o_baseband_q_c_11;
    output o_baseband_q_c_10;
    output n3608;
    output o_baseband_q_c_8;
    
    wire i_ref_clk_c /* synthesis SET_AS_NETWORK=i_ref_clk_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(22[12:21])
    wire [15:0]modulation_output /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(62[39:56])
    wire o_baseband_i_c_15 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[37:47])
    wire o_baseband_i_c_14 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[37:47])
    wire o_baseband_i_c_13 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[37:47])
    wire o_baseband_i_c_12 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[37:47])
    wire o_baseband_i_c_11 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[37:47])
    wire o_baseband_i_c_10 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[37:47])
    wire n3607 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[37:47])
    wire o_baseband_q_c_7 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[49:59])
    wire o_baseband_i_c_7 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[37:47])
    wire o_baseband_i_c_8 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[37:47])
    wire o_baseband_q_c_15 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[49:59])
    wire o_baseband_q_c_14 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[49:59])
    wire o_baseband_q_c_13 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[49:59])
    wire o_baseband_q_c_12 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[49:59])
    wire o_baseband_q_c_11 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[49:59])
    wire o_baseband_q_c_10 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[49:59])
    wire n3608 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[49:59])
    wire o_baseband_q_c_8 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[49:59])
    wire [31:0]\addr_space[0] ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(25[12:22])
    wire [31:0]\addr_space[1] ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(25[12:22])
    wire [31:0]\addr_space[2] ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(25[12:22])
    wire [31:0]\addr_space[3] ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(25[12:22])
    
    wire i_ref_clk_c_enable_149;
    wire [30:0]carrier_center_increment_offset_ls;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(52[31:65])
    wire [30:0]n64;
    wire [31:0]o_wb_data_31__N_1337;
    wire [30:0]carrier_center_increment_offset_rs;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(52[67:101])
    wire [30:0]carrier_center_increment_offset_rs_30__N_1560;
    wire [30:0]carrier_increment;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(53[31:48])
    wire [30:0]carrier_increment_30__N_1591;
    wire [16:0]sine_lookup_width_minus_modulation_deviation_amount;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(74[27:78])
    wire [31:0]sine_lookup_width_minus_modulation_deviation_amount_16__N_1622;
    wire [16:0]modulation_deviation_amount_minus_sine_lookup_width;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(74[80:131])
    
    wire n178, n24526, n22763, n13476, n6, n24516, n24539, n24549, 
        n17361, n14286, n17360, n17359, n17358, n17357, n17356, 
        n17355, n17354, n17353, n17352, n17351, n17350, n17349, 
        n17348, n17347, n17345, n20020, n20021, n17344, n17343, 
        n17342, n17341, n43, n24515, n17340, n17339, n20023, n20024, 
        n17338, n20026, n20027, n20029, n20030, n20032, n20033, 
        n20035, n20036, n17400;
    wire [17:0]modulation_deviation_amount_minus_sine_lookup_width_16__N_1639;
    
    wire n17399, n17398, n17397, n17396, n17395, n24823, n44, 
        n22, n18, n178_adj_3009, n20, n14, n20038, n20039, n20041, 
        n20042, n20066, n22761, n36, n22762, n20065, n20063, n20062, 
        n40, n71, n9, n11, n22760, n13, n15, n20060, n20059, 
        n13468, n13470, n7, n22_adj_3010, n18_adj_3011, n20_adj_3012, 
        n14_adj_3013, n20057, n41, n45, n72, n14_adj_3014, n10, 
        n12, n8, n37, n38, n42, n46, n73, n20056, n73_adj_3015, 
        n104, n19807, n135, n72_adj_3016, n103, n134, n20044, 
        n20045, n22765, n22766, n22767, n24988, n85, n24819, n24517, 
        n24518, n22770, n24548, n24547, n22771, n22772, n17801, 
        n24, n20_adj_3027, n22_adj_3028, n16, n24538, n24537, n24525, 
        n24524, n39_adj_3029, n20054, n78, n101, n79, n102, n25008, 
        n60_adj_3030, n59_adj_3031, n82, n105, n47_adj_3032, n74, 
        n83, n106, n48_adj_3033, n75, n20053, n55_adj_3034, n24846, 
        n56_adj_3035, n24850, n20051, n25012, n24888, n24834, n81, 
        n89, n24820, n80, n88, n24821, n24822, n25187, n29, 
        n20015, n20014, n20012, n20011, n20009, n20008, n20006, 
        n20005, n20047, n20048, n21575, n21574, n20003, n20002, 
        n20000, n19999, n19997, n19996, n21566, n21565, n21563, 
        n21562, n19991, n19990, n20050, n19988, n19987, n19985, 
        n19984, n19982, n19981, n17, n19979, n50_adj_3036, n54_adj_3037, 
        n19978, n27, n58_adj_3038, n19, n21, n23, n25, n49_adj_3039, 
        n53_adj_3040, n57_adj_3041, n30, n26, n28, n18_adj_3042, 
        n20_adj_3043, n22_adj_3044, n24_adj_3045, n9012, n9010, n70, 
        n52_adj_3046, n95, n24901, n96, n25015, n97, n113, n16_adj_3047, 
        n51_adj_3048, n98, n114, n99, n115, n76, n45_adj_3049, 
        n84, n25009, n100, n77, n46_adj_3050, n132, n133, n136, 
        n137, n107, n4, n108, n24835, n22768, n25133, n20018, 
        n118, n117, n20017;
    wire [15:0]quarter_wave_sample_register_q;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(22[56:86])
    
    FD1P3DX \addr_space_0[[30__162  (.D(wb_odata[30]), .SP(i_ref_clk_c_enable_106), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[0] [30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[30__162 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[29__163  (.D(wb_odata[29]), .SP(i_ref_clk_c_enable_106), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[0] [29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[29__163 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[28__164  (.D(wb_odata[28]), .SP(i_ref_clk_c_enable_106), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[0] [28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[28__164 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[27__165  (.D(wb_odata[27]), .SP(i_ref_clk_c_enable_106), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[0] [27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[27__165 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[26__166  (.D(wb_odata[26]), .SP(i_ref_clk_c_enable_106), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[0] [26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[26__166 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[25__167  (.D(wb_odata[25]), .SP(i_ref_clk_c_enable_106), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[0] [25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[25__167 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[24__168  (.D(wb_odata[24]), .SP(i_ref_clk_c_enable_106), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[0] [24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[24__168 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[23__169  (.D(wb_odata[23]), .SP(i_ref_clk_c_enable_106), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[0] [23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[23__169 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[21__172  (.D(wb_odata[21]), .SP(i_ref_clk_c_enable_106), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[0] [21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[21__172 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[20__173  (.D(wb_odata[20]), .SP(i_ref_clk_c_enable_106), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[0] [20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[20__173 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[19__174  (.D(wb_odata[19]), .SP(i_ref_clk_c_enable_106), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[0] [19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[19__174 .GSR = "DISABLED";
    FD1P3BX \addr_space_0[[18__175  (.D(wb_odata[18]), .SP(i_ref_clk_c_enable_106), 
            .CK(i_ref_clk_c), .PD(i_resetb_N_301), .Q(\addr_space[0] [18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[18__175 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[17__176  (.D(wb_odata[17]), .SP(i_ref_clk_c_enable_106), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[0] [17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[17__176 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[16__177  (.D(wb_odata[16]), .SP(i_ref_clk_c_enable_106), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[0] [16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[16__177 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[15__178  (.D(wb_odata[15]), .SP(i_ref_clk_c_enable_106), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[0] [15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[15__178 .GSR = "DISABLED";
    FD1P3BX \addr_space_0[[14__179  (.D(wb_odata[14]), .SP(i_ref_clk_c_enable_106), 
            .CK(i_ref_clk_c), .PD(i_resetb_N_301), .Q(\addr_space[0] [14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[14__179 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[13__180  (.D(wb_odata[13]), .SP(i_ref_clk_c_enable_106), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[0] [13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[13__180 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[12__181  (.D(wb_odata[12]), .SP(i_ref_clk_c_enable_106), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[0] [12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[12__181 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[11__182  (.D(wb_odata[11]), .SP(i_ref_clk_c_enable_106), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[0] [11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[11__182 .GSR = "DISABLED";
    FD1P3BX \addr_space_0[[10__183  (.D(wb_odata[10]), .SP(i_ref_clk_c_enable_106), 
            .CK(i_ref_clk_c), .PD(i_resetb_N_301), .Q(\addr_space[0] [10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[10__183 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[9__184  (.D(wb_odata[9]), .SP(i_ref_clk_c_enable_106), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[0] [9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[9__184 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[8__185  (.D(wb_odata[8]), .SP(i_ref_clk_c_enable_106), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[0] [8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[8__185 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[7__186  (.D(wb_odata[7]), .SP(i_ref_clk_c_enable_106), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[0] [7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[7__186 .GSR = "DISABLED";
    FD1P3BX \addr_space_0[[6__187  (.D(wb_odata[6]), .SP(i_ref_clk_c_enable_106), 
            .CK(i_ref_clk_c), .PD(i_resetb_N_301), .Q(\addr_space[0] [6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[6__187 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[5__188  (.D(wb_odata[5]), .SP(i_ref_clk_c_enable_106), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[0] [5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[5__188 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[4__189  (.D(wb_odata[4]), .SP(i_ref_clk_c_enable_106), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[0] [4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[4__189 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[3__190  (.D(wb_odata[3]), .SP(i_ref_clk_c_enable_106), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[0] [3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[3__190 .GSR = "DISABLED";
    FD1P3BX \addr_space_0[[2__191  (.D(wb_odata[2]), .SP(i_ref_clk_c_enable_106), 
            .CK(i_ref_clk_c), .PD(i_resetb_N_301), .Q(\addr_space[0] [2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[2__191 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[1__192  (.D(wb_odata[1]), .SP(i_ref_clk_c_enable_106), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[0] [1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[1__192 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[0__193  (.D(wb_odata[0]), .SP(i_ref_clk_c_enable_106), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[0] [0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[0__193 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[31__194  (.D(wb_odata[31]), .SP(i_ref_clk_c_enable_66), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[1] [31])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[31__194 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[30__195  (.D(wb_odata[30]), .SP(i_ref_clk_c_enable_66), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[1] [30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[30__195 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[29__196  (.D(wb_odata[29]), .SP(i_ref_clk_c_enable_66), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[1] [29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[29__196 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[28__197  (.D(wb_odata[28]), .SP(i_ref_clk_c_enable_66), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[1] [28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[28__197 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[27__198  (.D(wb_odata[27]), .SP(i_ref_clk_c_enable_66), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[1] [27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[27__198 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[26__199  (.D(wb_odata[26]), .SP(i_ref_clk_c_enable_66), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[1] [26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[26__199 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[25__200  (.D(wb_odata[25]), .SP(i_ref_clk_c_enable_66), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[1] [25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[25__200 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[24__201  (.D(wb_odata[24]), .SP(i_ref_clk_c_enable_66), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[1] [24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[24__201 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[23__202  (.D(wb_odata[23]), .SP(i_ref_clk_c_enable_66), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[1] [23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[23__202 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[22__203  (.D(wb_odata[22]), .SP(i_ref_clk_c_enable_66), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[1] [22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[22__203 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[21__204  (.D(wb_odata[21]), .SP(i_ref_clk_c_enable_66), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[1] [21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[21__204 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[20__205  (.D(wb_odata[20]), .SP(i_ref_clk_c_enable_66), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[1] [20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[20__205 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[19__206  (.D(wb_odata[19]), .SP(i_ref_clk_c_enable_66), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[1] [19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[19__206 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[18__207  (.D(wb_odata[18]), .SP(i_ref_clk_c_enable_66), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[1] [18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[18__207 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[17__208  (.D(wb_odata[17]), .SP(i_ref_clk_c_enable_66), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[1] [17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[17__208 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[16__209  (.D(wb_odata[16]), .SP(i_ref_clk_c_enable_66), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[1] [16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[16__209 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[15__210  (.D(wb_odata[15]), .SP(i_ref_clk_c_enable_66), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[1] [15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[15__210 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[14__211  (.D(wb_odata[14]), .SP(i_ref_clk_c_enable_66), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[1] [14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[14__211 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[13__212  (.D(wb_odata[13]), .SP(i_ref_clk_c_enable_66), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[1] [13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[13__212 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[12__213  (.D(wb_odata[12]), .SP(i_ref_clk_c_enable_66), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[1] [12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[12__213 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[11__214  (.D(wb_odata[11]), .SP(i_ref_clk_c_enable_66), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[1] [11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[11__214 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[10__215  (.D(wb_odata[10]), .SP(i_ref_clk_c_enable_66), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[1] [10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[10__215 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[9__216  (.D(wb_odata[9]), .SP(i_ref_clk_c_enable_66), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[1] [9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[9__216 .GSR = "DISABLED";
    FD1P3BX \addr_space_1[[8__217  (.D(wb_odata[8]), .SP(i_ref_clk_c_enable_66), 
            .CK(i_ref_clk_c), .PD(i_resetb_N_301), .Q(\addr_space[1] [8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[8__217 .GSR = "DISABLED";
    FD1P3BX \addr_space_1[[7__218  (.D(wb_odata[7]), .SP(i_ref_clk_c_enable_66), 
            .CK(i_ref_clk_c), .PD(i_resetb_N_301), .Q(\addr_space[1] [7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[7__218 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[6__219  (.D(wb_odata[6]), .SP(i_ref_clk_c_enable_66), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[1] [6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[6__219 .GSR = "DISABLED";
    FD1P3BX \addr_space_1[[5__220  (.D(wb_odata[5]), .SP(i_ref_clk_c_enable_66), 
            .CK(i_ref_clk_c), .PD(i_resetb_N_301), .Q(\addr_space[1] [5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[5__220 .GSR = "DISABLED";
    FD1P3BX \addr_space_1[[4__221  (.D(wb_odata[4]), .SP(i_ref_clk_c_enable_66), 
            .CK(i_ref_clk_c), .PD(i_resetb_N_301), .Q(\addr_space[1] [4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[4__221 .GSR = "DISABLED";
    FD1P3BX \addr_space_1[[3__222  (.D(wb_odata[3]), .SP(i_ref_clk_c_enable_66), 
            .CK(i_ref_clk_c), .PD(i_resetb_N_301), .Q(\addr_space[1] [3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[3__222 .GSR = "DISABLED";
    FD1P3BX \addr_space_1[[2__223  (.D(wb_odata[2]), .SP(i_ref_clk_c_enable_66), 
            .CK(i_ref_clk_c), .PD(i_resetb_N_301), .Q(\addr_space[1] [2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[2__223 .GSR = "DISABLED";
    FD1P3BX \addr_space_1[[1__224  (.D(wb_odata[1]), .SP(i_ref_clk_c_enable_66), 
            .CK(i_ref_clk_c), .PD(i_resetb_N_301), .Q(\addr_space[1] [1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[1__224 .GSR = "DISABLED";
    FD1P3BX \addr_space_1[[0__225  (.D(wb_odata[0]), .SP(i_ref_clk_c_enable_66), 
            .CK(i_ref_clk_c), .PD(i_resetb_N_301), .Q(\addr_space[1] [0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[0__225 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[31__226  (.D(wb_odata[31]), .SP(i_ref_clk_c_enable_98), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [31])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[31__226 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[30__227  (.D(wb_odata[30]), .SP(i_ref_clk_c_enable_98), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[30__227 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[29__228  (.D(wb_odata[29]), .SP(i_ref_clk_c_enable_98), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[29__228 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[28__229  (.D(wb_odata[28]), .SP(i_ref_clk_c_enable_98), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[28__229 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[27__230  (.D(wb_odata[27]), .SP(i_ref_clk_c_enable_98), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[27__230 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[26__231  (.D(wb_odata[26]), .SP(i_ref_clk_c_enable_98), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[26__231 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[25__232  (.D(wb_odata[25]), .SP(i_ref_clk_c_enable_98), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[25__232 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[24__233  (.D(wb_odata[24]), .SP(i_ref_clk_c_enable_98), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[24__233 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[23__234  (.D(wb_odata[23]), .SP(i_ref_clk_c_enable_98), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[23__234 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[22__235  (.D(wb_odata[22]), .SP(i_ref_clk_c_enable_98), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[22__235 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[21__236  (.D(wb_odata[21]), .SP(i_ref_clk_c_enable_98), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[21__236 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[20__237  (.D(wb_odata[20]), .SP(i_ref_clk_c_enable_98), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[20__237 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[19__238  (.D(wb_odata[19]), .SP(i_ref_clk_c_enable_98), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[19__238 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[18__239  (.D(wb_odata[18]), .SP(i_ref_clk_c_enable_98), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[18__239 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[17__240  (.D(wb_odata[17]), .SP(i_ref_clk_c_enable_98), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[17__240 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[16__241  (.D(wb_odata[16]), .SP(i_ref_clk_c_enable_98), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[16__241 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[15__242  (.D(wb_odata[15]), .SP(i_ref_clk_c_enable_98), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[15__242 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[14__243  (.D(wb_odata[14]), .SP(i_ref_clk_c_enable_98), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[14__243 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[13__244  (.D(wb_odata[13]), .SP(i_ref_clk_c_enable_98), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[13__244 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[12__245  (.D(wb_odata[12]), .SP(i_ref_clk_c_enable_98), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[12__245 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[11__246  (.D(wb_odata[11]), .SP(i_ref_clk_c_enable_98), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[11__246 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[10__247  (.D(wb_odata[10]), .SP(i_ref_clk_c_enable_98), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[10__247 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[9__248  (.D(wb_odata[9]), .SP(i_ref_clk_c_enable_98), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[9__248 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[8__249  (.D(wb_odata[8]), .SP(i_ref_clk_c_enable_98), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[8__249 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[7__250  (.D(wb_odata[7]), .SP(i_ref_clk_c_enable_98), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[7__250 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[6__251  (.D(wb_odata[6]), .SP(i_ref_clk_c_enable_98), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[6__251 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[5__252  (.D(wb_odata[5]), .SP(i_ref_clk_c_enable_98), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[5__252 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[4__253  (.D(wb_odata[4]), .SP(i_ref_clk_c_enable_98), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[4__253 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[3__254  (.D(wb_odata[3]), .SP(i_ref_clk_c_enable_98), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[3__254 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[2__255  (.D(wb_odata[2]), .SP(i_ref_clk_c_enable_98), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[2__255 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[1__256  (.D(wb_odata[1]), .SP(i_ref_clk_c_enable_98), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[1__256 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[0__257  (.D(wb_odata[0]), .SP(i_ref_clk_c_enable_98), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[0__257 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[30__261  (.D(wb_odata[30]), .SP(i_ref_clk_c_enable_149), 
            .CK(i_ref_clk_c), .Q(\addr_space[3] [30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[30__261 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[29__263  (.D(wb_odata[29]), .SP(i_ref_clk_c_enable_149), 
            .CK(i_ref_clk_c), .Q(\addr_space[3] [29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[29__263 .GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i0 (.D(n64[0]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_ls[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_ls__i0.GSR = "DISABLED";
    FD1S3AX o_wb_data_i0 (.D(o_wb_data_31__N_1337[0]), .CK(i_ref_clk_c), 
            .Q(wb_fm_data[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i0.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_rs_i1 (.D(carrier_center_increment_offset_rs_30__N_1560[0]), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_rs[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_rs_i1.GSR = "DISABLED";
    FD1S3DX carrier_increment_i0 (.D(carrier_increment_30__N_1591[0]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(carrier_increment[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_increment_i0.GSR = "DISABLED";
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i0 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[0]), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(sine_lookup_width_minus_modulation_deviation_amount[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i0.GSR = "DISABLED";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i0 (.D(\addr_space[2] [0]), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(modulation_deviation_amount_minus_sine_lookup_width[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i0.GSR = "DISABLED";
    FD1P3DX \addr_space_0[[31__161  (.D(wb_odata[31]), .SP(i_ref_clk_c_enable_106), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(\addr_space[0] [31])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[31__161 .GSR = "DISABLED";
    FD1P3BX \addr_space_0[[22__171  (.D(wb_odata[22]), .SP(i_ref_clk_c_enable_106), 
            .CK(i_ref_clk_c), .PD(i_resetb_N_301), .Q(\addr_space[0] [22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[22__171 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[28__265  (.D(wb_odata[28]), .SP(i_ref_clk_c_enable_149), 
            .CK(i_ref_clk_c), .Q(\addr_space[3] [28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[28__265 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[27__267  (.D(wb_odata[27]), .SP(i_ref_clk_c_enable_149), 
            .CK(i_ref_clk_c), .Q(\addr_space[3] [27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[27__267 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[26__269  (.D(wb_odata[26]), .SP(i_ref_clk_c_enable_149), 
            .CK(i_ref_clk_c), .Q(\addr_space[3] [26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[26__269 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[25__271  (.D(wb_odata[25]), .SP(i_ref_clk_c_enable_149), 
            .CK(i_ref_clk_c), .Q(\addr_space[3] [25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[25__271 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[24__273  (.D(wb_odata[24]), .SP(i_ref_clk_c_enable_149), 
            .CK(i_ref_clk_c), .Q(\addr_space[3] [24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[24__273 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[23__275  (.D(wb_odata[23]), .SP(i_ref_clk_c_enable_149), 
            .CK(i_ref_clk_c), .Q(\addr_space[3] [23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[23__275 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[22__277  (.D(wb_odata[22]), .SP(i_ref_clk_c_enable_149), 
            .CK(i_ref_clk_c), .Q(\addr_space[3] [22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[22__277 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[21__279  (.D(wb_odata[21]), .SP(i_ref_clk_c_enable_149), 
            .CK(i_ref_clk_c), .Q(\addr_space[3] [21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[21__279 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[20__281  (.D(wb_odata[20]), .SP(i_ref_clk_c_enable_149), 
            .CK(i_ref_clk_c), .Q(\addr_space[3] [20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[20__281 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[19__283  (.D(wb_odata[19]), .SP(i_ref_clk_c_enable_149), 
            .CK(i_ref_clk_c), .Q(\addr_space[3] [19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[19__283 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[18__285  (.D(wb_odata[18]), .SP(i_ref_clk_c_enable_149), 
            .CK(i_ref_clk_c), .Q(\addr_space[3] [18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[18__285 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[17__287  (.D(wb_odata[17]), .SP(i_ref_clk_c_enable_149), 
            .CK(i_ref_clk_c), .Q(\addr_space[3] [17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[17__287 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[16__289  (.D(wb_odata[16]), .SP(i_ref_clk_c_enable_149), 
            .CK(i_ref_clk_c), .Q(\addr_space[3] [16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[16__289 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[15__291  (.D(wb_odata[15]), .SP(i_ref_clk_c_enable_149), 
            .CK(i_ref_clk_c), .Q(\addr_space[3] [15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[15__291 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[14__293  (.D(wb_odata[14]), .SP(i_ref_clk_c_enable_149), 
            .CK(i_ref_clk_c), .Q(\addr_space[3] [14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[14__293 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[13__295  (.D(wb_odata[13]), .SP(i_ref_clk_c_enable_149), 
            .CK(i_ref_clk_c), .Q(\addr_space[3] [13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[13__295 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[12__297  (.D(wb_odata[12]), .SP(i_ref_clk_c_enable_149), 
            .CK(i_ref_clk_c), .Q(\addr_space[3] [12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[12__297 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[11__299  (.D(wb_odata[11]), .SP(i_ref_clk_c_enable_149), 
            .CK(i_ref_clk_c), .Q(\addr_space[3] [11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[11__299 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[10__301  (.D(wb_odata[10]), .SP(i_ref_clk_c_enable_149), 
            .CK(i_ref_clk_c), .Q(\addr_space[3] [10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[10__301 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[9__303  (.D(wb_odata[9]), .SP(i_ref_clk_c_enable_149), 
            .CK(i_ref_clk_c), .Q(\addr_space[3] [9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[9__303 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[8__305  (.D(wb_odata[8]), .SP(i_ref_clk_c_enable_149), 
            .CK(i_ref_clk_c), .Q(\addr_space[3] [8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[8__305 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[7__307  (.D(wb_odata[7]), .SP(i_ref_clk_c_enable_149), 
            .CK(i_ref_clk_c), .Q(\addr_space[3] [7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[7__307 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[6__309  (.D(wb_odata[6]), .SP(i_ref_clk_c_enable_149), 
            .CK(i_ref_clk_c), .Q(\addr_space[3] [6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[6__309 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[5__311  (.D(wb_odata[5]), .SP(i_ref_clk_c_enable_149), 
            .CK(i_ref_clk_c), .Q(\addr_space[3] [5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[5__311 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[4__313  (.D(wb_odata[4]), .SP(i_ref_clk_c_enable_149), 
            .CK(i_ref_clk_c), .Q(\addr_space[3] [4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[4__313 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[3__315  (.D(wb_odata[3]), .SP(i_ref_clk_c_enable_149), 
            .CK(i_ref_clk_c), .Q(\addr_space[3] [3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[3__315 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[2__317  (.D(wb_odata[2]), .SP(i_ref_clk_c_enable_149), 
            .CK(i_ref_clk_c), .Q(\addr_space[3] [2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[2__317 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[1__319  (.D(wb_odata[1]), .SP(i_ref_clk_c_enable_149), 
            .CK(i_ref_clk_c), .Q(\addr_space[3] [1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[1__319 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[0__321  (.D(wb_odata[0]), .SP(i_ref_clk_c_enable_149), 
            .CK(i_ref_clk_c), .Q(\addr_space[3] [0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[0__321 .GSR = "DISABLED";
    LUT4 n24526_bdd_3_lut_4_lut (.A(sine_lookup_width_minus_modulation_deviation_amount[4]), 
         .B(n178), .C(modulation_output[15]), .D(n24526), .Z(carrier_center_increment_offset_rs_30__N_1560[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam n24526_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n22763_bdd_3_lut_4_lut (.A(sine_lookup_width_minus_modulation_deviation_amount[4]), 
         .B(n178), .C(modulation_output[15]), .D(n22763), .Z(carrier_center_increment_offset_rs_30__N_1560[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam n22763_bdd_3_lut_4_lut.init = 16'hf1e0;
    FD1S3IX o_wb_ack_323 (.D(wb_fm_data_31__N_63), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(wb_fm_ack)) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[8] 48[4])
    defparam o_wb_ack_323.GSR = "DISABLED";
    FD1P3AX \addr_space_3[[31__259  (.D(wb_odata[31]), .SP(i_ref_clk_c_enable_149), 
            .CK(i_ref_clk_c), .Q(\addr_space[3] [31])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[31__259 .GSR = "DISABLED";
    LUT4 n39_bdd_3_lut_23815 (.A(n13476), .B(n6), .C(sine_lookup_width_minus_modulation_deviation_amount[1]), 
         .Z(n24516)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n39_bdd_3_lut_23815.init = 16'hcaca;
    LUT4 n24539_bdd_3_lut_4_lut (.A(sine_lookup_width_minus_modulation_deviation_amount[4]), 
         .B(n178), .C(modulation_output[15]), .D(n24539), .Z(carrier_center_increment_offset_rs_30__N_1560[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam n24539_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n24549_bdd_3_lut_4_lut (.A(sine_lookup_width_minus_modulation_deviation_amount[4]), 
         .B(n178), .C(modulation_output[15]), .D(n24549), .Z(carrier_center_increment_offset_rs_30__N_1560[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam n24549_bdd_3_lut_4_lut.init = 16'hf1e0;
    CCU2D add_365_31 (.A0(\addr_space[0] [29]), .B0(n14286), .C0(carrier_center_increment_offset_rs[30]), 
          .D0(carrier_center_increment_offset_ls[29]), .A1(\addr_space[0] [30]), 
          .B1(n14286), .C1(carrier_center_increment_offset_rs[30]), .D1(carrier_center_increment_offset_ls[30]), 
          .CIN(n17361), .S0(carrier_increment_30__N_1591[29]), .S1(carrier_increment_30__N_1591[30]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(92[4:87])
    defparam add_365_31.INIT0 = 16'h569a;
    defparam add_365_31.INIT1 = 16'h569a;
    defparam add_365_31.INJECT1_0 = "NO";
    defparam add_365_31.INJECT1_1 = "NO";
    CCU2D add_365_29 (.A0(\addr_space[0] [27]), .B0(n14286), .C0(carrier_center_increment_offset_rs[30]), 
          .D0(carrier_center_increment_offset_ls[27]), .A1(\addr_space[0] [28]), 
          .B1(n14286), .C1(carrier_center_increment_offset_rs[30]), .D1(carrier_center_increment_offset_ls[28]), 
          .CIN(n17360), .COUT(n17361), .S0(carrier_increment_30__N_1591[27]), 
          .S1(carrier_increment_30__N_1591[28]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(92[4:87])
    defparam add_365_29.INIT0 = 16'h569a;
    defparam add_365_29.INIT1 = 16'h569a;
    defparam add_365_29.INJECT1_0 = "NO";
    defparam add_365_29.INJECT1_1 = "NO";
    CCU2D add_365_27 (.A0(\addr_space[0] [25]), .B0(n14286), .C0(carrier_center_increment_offset_rs[30]), 
          .D0(carrier_center_increment_offset_ls[25]), .A1(\addr_space[0] [26]), 
          .B1(n14286), .C1(carrier_center_increment_offset_rs[30]), .D1(carrier_center_increment_offset_ls[26]), 
          .CIN(n17359), .COUT(n17360), .S0(carrier_increment_30__N_1591[25]), 
          .S1(carrier_increment_30__N_1591[26]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(92[4:87])
    defparam add_365_27.INIT0 = 16'h569a;
    defparam add_365_27.INIT1 = 16'h569a;
    defparam add_365_27.INJECT1_0 = "NO";
    defparam add_365_27.INJECT1_1 = "NO";
    CCU2D add_365_25 (.A0(\addr_space[0] [23]), .B0(n14286), .C0(carrier_center_increment_offset_rs[30]), 
          .D0(carrier_center_increment_offset_ls[23]), .A1(\addr_space[0] [24]), 
          .B1(n14286), .C1(carrier_center_increment_offset_rs[30]), .D1(carrier_center_increment_offset_ls[24]), 
          .CIN(n17358), .COUT(n17359), .S0(carrier_increment_30__N_1591[23]), 
          .S1(carrier_increment_30__N_1591[24]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(92[4:87])
    defparam add_365_25.INIT0 = 16'h569a;
    defparam add_365_25.INIT1 = 16'h569a;
    defparam add_365_25.INJECT1_0 = "NO";
    defparam add_365_25.INJECT1_1 = "NO";
    CCU2D add_365_23 (.A0(\addr_space[0] [21]), .B0(n14286), .C0(carrier_center_increment_offset_rs[30]), 
          .D0(carrier_center_increment_offset_ls[21]), .A1(\addr_space[0] [22]), 
          .B1(n14286), .C1(carrier_center_increment_offset_rs[30]), .D1(carrier_center_increment_offset_ls[22]), 
          .CIN(n17357), .COUT(n17358), .S0(carrier_increment_30__N_1591[21]), 
          .S1(carrier_increment_30__N_1591[22]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(92[4:87])
    defparam add_365_23.INIT0 = 16'h569a;
    defparam add_365_23.INIT1 = 16'h569a;
    defparam add_365_23.INJECT1_0 = "NO";
    defparam add_365_23.INJECT1_1 = "NO";
    CCU2D add_365_21 (.A0(\addr_space[0] [19]), .B0(n14286), .C0(carrier_center_increment_offset_rs[30]), 
          .D0(carrier_center_increment_offset_ls[19]), .A1(\addr_space[0] [20]), 
          .B1(n14286), .C1(carrier_center_increment_offset_rs[30]), .D1(carrier_center_increment_offset_ls[20]), 
          .CIN(n17356), .COUT(n17357), .S0(carrier_increment_30__N_1591[19]), 
          .S1(carrier_increment_30__N_1591[20]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(92[4:87])
    defparam add_365_21.INIT0 = 16'h569a;
    defparam add_365_21.INIT1 = 16'h569a;
    defparam add_365_21.INJECT1_0 = "NO";
    defparam add_365_21.INJECT1_1 = "NO";
    CCU2D add_365_19 (.A0(\addr_space[0] [17]), .B0(n14286), .C0(carrier_center_increment_offset_rs[30]), 
          .D0(carrier_center_increment_offset_ls[17]), .A1(\addr_space[0] [18]), 
          .B1(n14286), .C1(carrier_center_increment_offset_rs[30]), .D1(carrier_center_increment_offset_ls[18]), 
          .CIN(n17355), .COUT(n17356), .S0(carrier_increment_30__N_1591[17]), 
          .S1(carrier_increment_30__N_1591[18]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(92[4:87])
    defparam add_365_19.INIT0 = 16'h569a;
    defparam add_365_19.INIT1 = 16'h569a;
    defparam add_365_19.INJECT1_0 = "NO";
    defparam add_365_19.INJECT1_1 = "NO";
    CCU2D add_365_17 (.A0(\addr_space[0] [15]), .B0(n14286), .C0(carrier_center_increment_offset_rs[30]), 
          .D0(carrier_center_increment_offset_ls[15]), .A1(\addr_space[0] [16]), 
          .B1(n14286), .C1(carrier_center_increment_offset_rs[30]), .D1(carrier_center_increment_offset_ls[16]), 
          .CIN(n17354), .COUT(n17355), .S0(carrier_increment_30__N_1591[15]), 
          .S1(carrier_increment_30__N_1591[16]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(92[4:87])
    defparam add_365_17.INIT0 = 16'h569a;
    defparam add_365_17.INIT1 = 16'h569a;
    defparam add_365_17.INJECT1_0 = "NO";
    defparam add_365_17.INJECT1_1 = "NO";
    CCU2D add_365_15 (.A0(\addr_space[0] [13]), .B0(n14286), .C0(carrier_center_increment_offset_rs[13]), 
          .D0(carrier_center_increment_offset_ls[13]), .A1(\addr_space[0] [14]), 
          .B1(n14286), .C1(carrier_center_increment_offset_rs[14]), .D1(carrier_center_increment_offset_ls[14]), 
          .CIN(n17353), .COUT(n17354), .S0(carrier_increment_30__N_1591[13]), 
          .S1(carrier_increment_30__N_1591[14]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(92[4:87])
    defparam add_365_15.INIT0 = 16'h569a;
    defparam add_365_15.INIT1 = 16'h569a;
    defparam add_365_15.INJECT1_0 = "NO";
    defparam add_365_15.INJECT1_1 = "NO";
    CCU2D add_365_13 (.A0(\addr_space[0] [11]), .B0(n14286), .C0(carrier_center_increment_offset_rs[11]), 
          .D0(carrier_center_increment_offset_ls[11]), .A1(\addr_space[0] [12]), 
          .B1(n14286), .C1(carrier_center_increment_offset_rs[12]), .D1(carrier_center_increment_offset_ls[12]), 
          .CIN(n17352), .COUT(n17353), .S0(carrier_increment_30__N_1591[11]), 
          .S1(carrier_increment_30__N_1591[12]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(92[4:87])
    defparam add_365_13.INIT0 = 16'h569a;
    defparam add_365_13.INIT1 = 16'h569a;
    defparam add_365_13.INJECT1_0 = "NO";
    defparam add_365_13.INJECT1_1 = "NO";
    CCU2D add_365_11 (.A0(\addr_space[0] [9]), .B0(n14286), .C0(carrier_center_increment_offset_rs[9]), 
          .D0(carrier_center_increment_offset_ls[9]), .A1(\addr_space[0] [10]), 
          .B1(n14286), .C1(carrier_center_increment_offset_rs[10]), .D1(carrier_center_increment_offset_ls[10]), 
          .CIN(n17351), .COUT(n17352), .S0(carrier_increment_30__N_1591[9]), 
          .S1(carrier_increment_30__N_1591[10]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(92[4:87])
    defparam add_365_11.INIT0 = 16'h569a;
    defparam add_365_11.INIT1 = 16'h569a;
    defparam add_365_11.INJECT1_0 = "NO";
    defparam add_365_11.INJECT1_1 = "NO";
    CCU2D add_365_9 (.A0(\addr_space[0] [7]), .B0(n14286), .C0(carrier_center_increment_offset_rs[7]), 
          .D0(carrier_center_increment_offset_ls[7]), .A1(\addr_space[0] [8]), 
          .B1(n14286), .C1(carrier_center_increment_offset_rs[8]), .D1(carrier_center_increment_offset_ls[8]), 
          .CIN(n17350), .COUT(n17351), .S0(carrier_increment_30__N_1591[7]), 
          .S1(carrier_increment_30__N_1591[8]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(92[4:87])
    defparam add_365_9.INIT0 = 16'h569a;
    defparam add_365_9.INIT1 = 16'h569a;
    defparam add_365_9.INJECT1_0 = "NO";
    defparam add_365_9.INJECT1_1 = "NO";
    CCU2D add_365_7 (.A0(\addr_space[0] [5]), .B0(n14286), .C0(carrier_center_increment_offset_rs[5]), 
          .D0(carrier_center_increment_offset_ls[5]), .A1(\addr_space[0] [6]), 
          .B1(n14286), .C1(carrier_center_increment_offset_rs[6]), .D1(carrier_center_increment_offset_ls[6]), 
          .CIN(n17349), .COUT(n17350), .S0(carrier_increment_30__N_1591[5]), 
          .S1(carrier_increment_30__N_1591[6]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(92[4:87])
    defparam add_365_7.INIT0 = 16'h569a;
    defparam add_365_7.INIT1 = 16'h569a;
    defparam add_365_7.INJECT1_0 = "NO";
    defparam add_365_7.INJECT1_1 = "NO";
    CCU2D add_365_5 (.A0(\addr_space[0] [3]), .B0(n14286), .C0(carrier_center_increment_offset_rs[3]), 
          .D0(carrier_center_increment_offset_ls[3]), .A1(\addr_space[0] [4]), 
          .B1(n14286), .C1(carrier_center_increment_offset_rs[4]), .D1(carrier_center_increment_offset_ls[4]), 
          .CIN(n17348), .COUT(n17349), .S0(carrier_increment_30__N_1591[3]), 
          .S1(carrier_increment_30__N_1591[4]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(92[4:87])
    defparam add_365_5.INIT0 = 16'h569a;
    defparam add_365_5.INIT1 = 16'h569a;
    defparam add_365_5.INJECT1_0 = "NO";
    defparam add_365_5.INJECT1_1 = "NO";
    CCU2D add_365_3 (.A0(\addr_space[0] [1]), .B0(n14286), .C0(carrier_center_increment_offset_rs[1]), 
          .D0(carrier_center_increment_offset_ls[1]), .A1(\addr_space[0] [2]), 
          .B1(n14286), .C1(carrier_center_increment_offset_rs[2]), .D1(carrier_center_increment_offset_ls[2]), 
          .CIN(n17347), .COUT(n17348), .S0(carrier_increment_30__N_1591[1]), 
          .S1(carrier_increment_30__N_1591[2]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(92[4:87])
    defparam add_365_3.INIT0 = 16'h569a;
    defparam add_365_3.INIT1 = 16'h569a;
    defparam add_365_3.INJECT1_0 = "NO";
    defparam add_365_3.INJECT1_1 = "NO";
    CCU2D add_365_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\addr_space[0] [0]), .B1(n14286), .C1(carrier_center_increment_offset_rs[0]), 
          .D1(carrier_center_increment_offset_ls[0]), .COUT(n17347), .S1(carrier_increment_30__N_1591[0]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(92[4:87])
    defparam add_365_1.INIT0 = 16'hF000;
    defparam add_365_1.INIT1 = 16'h569a;
    defparam add_365_1.INJECT1_0 = "NO";
    defparam add_365_1.INJECT1_1 = "NO";
    CCU2D sub_377_add_2_17 (.A0(\addr_space[2] [15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\addr_space[2] [16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17345), .S0(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[15]), 
          .S1(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[16]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(85[58:109])
    defparam sub_377_add_2_17.INIT0 = 16'hf555;
    defparam sub_377_add_2_17.INIT1 = 16'hf555;
    defparam sub_377_add_2_17.INJECT1_0 = "NO";
    defparam sub_377_add_2_17.INJECT1_1 = "NO";
    PFUMX i17692 (.BLUT(n20020), .ALUT(n20021), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[16]));
    CCU2D sub_377_add_2_15 (.A0(\addr_space[2] [13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\addr_space[2] [14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17344), .COUT(n17345), .S0(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[13]), 
          .S1(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[14]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(85[58:109])
    defparam sub_377_add_2_15.INIT0 = 16'hf555;
    defparam sub_377_add_2_15.INIT1 = 16'hf555;
    defparam sub_377_add_2_15.INJECT1_0 = "NO";
    defparam sub_377_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_377_add_2_13 (.A0(\addr_space[2] [11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\addr_space[2] [12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17343), .COUT(n17344), .S0(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[11]), 
          .S1(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[12]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(85[58:109])
    defparam sub_377_add_2_13.INIT0 = 16'hf555;
    defparam sub_377_add_2_13.INIT1 = 16'hf555;
    defparam sub_377_add_2_13.INJECT1_0 = "NO";
    defparam sub_377_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_377_add_2_11 (.A0(\addr_space[2] [9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\addr_space[2] [10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17342), .COUT(n17343), .S0(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[9]), 
          .S1(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[10]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(85[58:109])
    defparam sub_377_add_2_11.INIT0 = 16'hf555;
    defparam sub_377_add_2_11.INIT1 = 16'hf555;
    defparam sub_377_add_2_11.INJECT1_0 = "NO";
    defparam sub_377_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_377_add_2_9 (.A0(\addr_space[2] [7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\addr_space[2] [8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17341), .COUT(n17342), .S0(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[7]), 
          .S1(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[8]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(85[58:109])
    defparam sub_377_add_2_9.INIT0 = 16'hf555;
    defparam sub_377_add_2_9.INIT1 = 16'hf555;
    defparam sub_377_add_2_9.INJECT1_0 = "NO";
    defparam sub_377_add_2_9.INJECT1_1 = "NO";
    LUT4 n39_bdd_3_lut_22812 (.A(n43), .B(modulation_output[15]), .C(sine_lookup_width_minus_modulation_deviation_amount[2]), 
         .Z(n24515)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n39_bdd_3_lut_22812.init = 16'hcaca;
    CCU2D sub_377_add_2_7 (.A0(\addr_space[2] [5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\addr_space[2] [6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17340), .COUT(n17341), .S0(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[5]), 
          .S1(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[6]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(85[58:109])
    defparam sub_377_add_2_7.INIT0 = 16'hf555;
    defparam sub_377_add_2_7.INIT1 = 16'hf555;
    defparam sub_377_add_2_7.INJECT1_0 = "NO";
    defparam sub_377_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_377_add_2_5 (.A0(\addr_space[2] [3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\addr_space[2] [4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17339), .COUT(n17340), .S0(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[3]), 
          .S1(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[4]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(85[58:109])
    defparam sub_377_add_2_5.INIT0 = 16'hf555;
    defparam sub_377_add_2_5.INIT1 = 16'h0aaa;
    defparam sub_377_add_2_5.INJECT1_0 = "NO";
    defparam sub_377_add_2_5.INJECT1_1 = "NO";
    PFUMX i17695 (.BLUT(n20023), .ALUT(n20024), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[15]));
    CCU2D sub_377_add_2_3 (.A0(\addr_space[2] [1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\addr_space[2] [2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17338), .COUT(n17339), .S0(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[1]), 
          .S1(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[2]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(85[58:109])
    defparam sub_377_add_2_3.INIT0 = 16'hf555;
    defparam sub_377_add_2_3.INIT1 = 16'hf555;
    defparam sub_377_add_2_3.INJECT1_0 = "NO";
    defparam sub_377_add_2_3.INJECT1_1 = "NO";
    PFUMX i17698 (.BLUT(n20026), .ALUT(n20027), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[14]));
    CCU2D sub_377_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\addr_space[2] [0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n17338));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(85[58:109])
    defparam sub_377_add_2_1.INIT0 = 16'h0000;
    defparam sub_377_add_2_1.INIT1 = 16'h0aaa;
    defparam sub_377_add_2_1.INJECT1_0 = "NO";
    defparam sub_377_add_2_1.INJECT1_1 = "NO";
    PFUMX i17701 (.BLUT(n20029), .ALUT(n20030), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[13]));
    PFUMX i17704 (.BLUT(n20032), .ALUT(n20033), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[12]));
    PFUMX i17707 (.BLUT(n20035), .ALUT(n20036), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[11]));
    CCU2D sub_113_add_2_13 (.A0(\addr_space[2] [15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\addr_space[2] [16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17400), .S0(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[15]), 
          .S1(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[16]));
    defparam sub_113_add_2_13.INIT0 = 16'h5555;
    defparam sub_113_add_2_13.INIT1 = 16'h5555;
    defparam sub_113_add_2_13.INJECT1_0 = "NO";
    defparam sub_113_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_113_add_2_11 (.A0(\addr_space[2] [13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\addr_space[2] [14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17399), .COUT(n17400), .S0(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[13]), 
          .S1(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[14]));
    defparam sub_113_add_2_11.INIT0 = 16'h5555;
    defparam sub_113_add_2_11.INIT1 = 16'h5555;
    defparam sub_113_add_2_11.INJECT1_0 = "NO";
    defparam sub_113_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_113_add_2_9 (.A0(\addr_space[2] [11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\addr_space[2] [12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17398), .COUT(n17399), .S0(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[11]), 
          .S1(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[12]));
    defparam sub_113_add_2_9.INIT0 = 16'h5555;
    defparam sub_113_add_2_9.INIT1 = 16'h5555;
    defparam sub_113_add_2_9.INJECT1_0 = "NO";
    defparam sub_113_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_113_add_2_7 (.A0(\addr_space[2] [9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\addr_space[2] [10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17397), .COUT(n17398), .S0(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[9]), 
          .S1(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[10]));
    defparam sub_113_add_2_7.INIT0 = 16'h5555;
    defparam sub_113_add_2_7.INIT1 = 16'h5555;
    defparam sub_113_add_2_7.INJECT1_0 = "NO";
    defparam sub_113_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_113_add_2_5 (.A0(\addr_space[2] [7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\addr_space[2] [8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17396), .COUT(n17397), .S0(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[7]), 
          .S1(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[8]));
    defparam sub_113_add_2_5.INIT0 = 16'h5555;
    defparam sub_113_add_2_5.INIT1 = 16'h5555;
    defparam sub_113_add_2_5.INJECT1_0 = "NO";
    defparam sub_113_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_113_add_2_3 (.A0(\addr_space[2] [5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\addr_space[2] [6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17395), .COUT(n17396), .S0(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[5]), 
          .S1(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[6]));
    defparam sub_113_add_2_3.INIT0 = 16'h5555;
    defparam sub_113_add_2_3.INIT1 = 16'h5555;
    defparam sub_113_add_2_3.INJECT1_0 = "NO";
    defparam sub_113_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_113_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\addr_space[2] [4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n17395), .S1(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[4]));
    defparam sub_113_add_2_1.INIT0 = 16'hF000;
    defparam sub_113_add_2_1.INIT1 = 16'h5555;
    defparam sub_113_add_2_1.INJECT1_0 = "NO";
    defparam sub_113_add_2_1.INJECT1_1 = "NO";
    LUT4 mux_374_Mux_1_i3_4_lut_4_lut_4_lut (.A(\wb_addr[0] ), .B(\wb_addr[1] ), 
         .C(\power_counter[1] ), .D(\smpl_register[1] ), .Z(n2139)) /* synthesis lut_function=(A (B (C)+!B (D))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(34[4:25])
    defparam mux_374_Mux_1_i3_4_lut_4_lut_4_lut.init = 16'hb391;
    LUT4 i6563_3_lut_4_lut (.A(sine_lookup_width_minus_modulation_deviation_amount[2]), 
         .B(n24823), .C(modulation_output[15]), .D(n44), .Z(carrier_center_increment_offset_rs_30__N_1560[12])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam i6563_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i3_4_lut (.A(i_resetb_c), .B(n24803), .C(\wb_addr[0] ), .D(\wb_addr[1] ), 
         .Z(i_ref_clk_c_enable_149)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i3_4_lut.init = 16'h8000;
    LUT4 i11_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[9]), 
         .B(n22), .C(n18), .D(modulation_deviation_amount_minus_sine_lookup_width[12]), 
         .Z(n178_adj_3009)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam i11_4_lut.init = 16'hfffe;
    LUT4 i10_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[15]), 
         .B(n20), .C(n14), .D(modulation_deviation_amount_minus_sine_lookup_width[5]), 
         .Z(n22)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam i10_4_lut.init = 16'hfffe;
    LUT4 i6_2_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[6]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[7]), .Z(n18)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam i6_2_lut.init = 16'heeee;
    LUT4 i8_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[14]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[11]), .C(modulation_deviation_amount_minus_sine_lookup_width[8]), 
         .D(modulation_deviation_amount_minus_sine_lookup_width[16]), .Z(n20)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam i8_4_lut.init = 16'hfffe;
    LUT4 i2_2_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[10]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[13]), .Z(n14)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam i2_2_lut.init = 16'heeee;
    LUT4 sub_377_inv_0_i1_1_lut (.A(\addr_space[2] [0]), .Z(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[0])) /* synthesis lut_function=(!(A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(85[58:109])
    defparam sub_377_inv_0_i1_1_lut.init = 16'h5555;
    PFUMX i17710 (.BLUT(n20038), .ALUT(n20039), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[10]));
    PFUMX i17713 (.BLUT(n20041), .ALUT(n20042), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[9]));
    LUT4 i17736_3_lut (.A(\addr_space[2] [1]), .B(\addr_space[3] [1]), .C(\wb_addr[0] ), 
         .Z(n20066)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17736_3_lut.init = 16'hcaca;
    LUT4 n22761_bdd_3_lut (.A(n22761), .B(n36), .C(sine_lookup_width_minus_modulation_deviation_amount[2]), 
         .Z(n22762)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n22761_bdd_3_lut.init = 16'hcaca;
    LUT4 i17735_3_lut (.A(\addr_space[0] [1]), .B(\addr_space[1] [1]), .C(\wb_addr[0] ), 
         .Z(n20065)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17735_3_lut.init = 16'hcaca;
    LUT4 i17733_3_lut (.A(\addr_space[2] [2]), .B(\addr_space[3] [2]), .C(\wb_addr[0] ), 
         .Z(n20063)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17733_3_lut.init = 16'hcaca;
    LUT4 i17732_3_lut (.A(\addr_space[0] [2]), .B(\addr_space[1] [2]), .C(\wb_addr[0] ), 
         .Z(n20062)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17732_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i71_3_lut (.A(n40), .B(n44), .C(sine_lookup_width_minus_modulation_deviation_amount[2]), 
         .Z(n71)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam modulation_output_15__I_0_i71_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i40_3_lut (.A(n9), .B(n11), .C(sine_lookup_width_minus_modulation_deviation_amount[1]), 
         .Z(n40)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam modulation_output_15__I_0_i40_3_lut.init = 16'hcaca;
    LUT4 n13468_bdd_3_lut_22879 (.A(modulation_output[1]), .B(modulation_output[0]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[0]), .Z(n22760)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n13468_bdd_3_lut_22879.init = 16'hacac;
    LUT4 modulation_output_15__I_0_i44_3_lut (.A(n13), .B(n15), .C(sine_lookup_width_minus_modulation_deviation_amount[1]), 
         .Z(n44)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam modulation_output_15__I_0_i44_3_lut.init = 16'hcaca;
    LUT4 i17730_3_lut (.A(\addr_space[2] [3]), .B(\addr_space[3] [3]), .C(\wb_addr[0] ), 
         .Z(n20060)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17730_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i15_3_lut (.A(modulation_output[14]), .B(modulation_output[15]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[0]), .Z(n15)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam modulation_output_15__I_0_i15_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i13_3_lut (.A(modulation_output[12]), .B(modulation_output[13]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[0]), .Z(n13)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam modulation_output_15__I_0_i13_3_lut.init = 16'hcaca;
    LUT4 i17729_3_lut (.A(\addr_space[0] [3]), .B(\addr_space[1] [3]), .C(\wb_addr[0] ), 
         .Z(n20059)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17729_3_lut.init = 16'hcaca;
    LUT4 i10811_3_lut (.A(modulation_output[2]), .B(modulation_output[3]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[0]), .Z(n13468)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(74[27:78])
    defparam i10811_3_lut.init = 16'hcaca;
    LUT4 i10815_3_lut (.A(n13470), .B(n7), .C(sine_lookup_width_minus_modulation_deviation_amount[1]), 
         .Z(n36)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(74[27:78])
    defparam i10815_3_lut.init = 16'hcaca;
    LUT4 i10813_3_lut (.A(modulation_output[4]), .B(modulation_output[5]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[0]), .Z(n13470)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(74[27:78])
    defparam i10813_3_lut.init = 16'hcaca;
    LUT4 i10814_3_lut (.A(modulation_output[6]), .B(modulation_output[7]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[0]), .Z(n7)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(74[27:78])
    defparam i10814_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i9_3_lut (.A(modulation_output[8]), .B(modulation_output[9]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[0]), .Z(n9)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam modulation_output_15__I_0_i9_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i11_3_lut (.A(modulation_output[10]), .B(modulation_output[11]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[0]), .Z(n11)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam modulation_output_15__I_0_i11_3_lut.init = 16'hcaca;
    LUT4 i11_4_lut_adj_84 (.A(sine_lookup_width_minus_modulation_deviation_amount[9]), 
         .B(n22_adj_3010), .C(n18_adj_3011), .D(sine_lookup_width_minus_modulation_deviation_amount[12]), 
         .Z(n178)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam i11_4_lut_adj_84.init = 16'hfffe;
    LUT4 i10_4_lut_adj_85 (.A(sine_lookup_width_minus_modulation_deviation_amount[15]), 
         .B(n20_adj_3012), .C(n14_adj_3013), .D(sine_lookup_width_minus_modulation_deviation_amount[5]), 
         .Z(n22_adj_3010)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam i10_4_lut_adj_85.init = 16'hfffe;
    LUT4 i6_2_lut_adj_86 (.A(sine_lookup_width_minus_modulation_deviation_amount[6]), 
         .B(sine_lookup_width_minus_modulation_deviation_amount[7]), .Z(n18_adj_3011)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam i6_2_lut_adj_86.init = 16'heeee;
    LUT4 i8_4_lut_adj_87 (.A(sine_lookup_width_minus_modulation_deviation_amount[14]), 
         .B(sine_lookup_width_minus_modulation_deviation_amount[11]), .C(sine_lookup_width_minus_modulation_deviation_amount[8]), 
         .D(sine_lookup_width_minus_modulation_deviation_amount[16]), .Z(n20_adj_3012)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam i8_4_lut_adj_87.init = 16'hfffe;
    LUT4 i2_2_lut_adj_88 (.A(sine_lookup_width_minus_modulation_deviation_amount[10]), 
         .B(sine_lookup_width_minus_modulation_deviation_amount[13]), .Z(n14_adj_3013)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam i2_2_lut_adj_88.init = 16'heeee;
    LUT4 i17727_3_lut (.A(\addr_space[2] [4]), .B(\addr_space[3] [4]), .C(\wb_addr[0] ), 
         .Z(n20057)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17727_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i72_3_lut (.A(n41), .B(n45), .C(sine_lookup_width_minus_modulation_deviation_amount[2]), 
         .Z(n72)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam modulation_output_15__I_0_i72_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i45_3_lut (.A(n14_adj_3014), .B(modulation_output[15]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[1]), .Z(n45)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam modulation_output_15__I_0_i45_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i14_3_lut (.A(modulation_output[13]), .B(modulation_output[14]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[0]), .Z(n14_adj_3014)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam modulation_output_15__I_0_i14_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i41_3_lut (.A(n10), .B(n12), .C(sine_lookup_width_minus_modulation_deviation_amount[1]), 
         .Z(n41)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam modulation_output_15__I_0_i41_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i10_3_lut (.A(modulation_output[9]), .B(modulation_output[10]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[0]), .Z(n10)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam modulation_output_15__I_0_i10_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i12_3_lut (.A(modulation_output[11]), .B(modulation_output[12]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[0]), .Z(n12)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam modulation_output_15__I_0_i12_3_lut.init = 16'hcaca;
    LUT4 i10819_3_lut (.A(modulation_output[3]), .B(modulation_output[4]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[0]), .Z(n13476)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(74[27:78])
    defparam i10819_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i37_3_lut (.A(n6), .B(n8), .C(sine_lookup_width_minus_modulation_deviation_amount[1]), 
         .Z(n37)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam modulation_output_15__I_0_i37_3_lut.init = 16'hcaca;
    LUT4 i10821_3_lut (.A(modulation_output[5]), .B(modulation_output[6]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[0]), .Z(n6)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(74[27:78])
    defparam i10821_3_lut.init = 16'hcaca;
    LUT4 i10827_3_lut (.A(modulation_output[7]), .B(modulation_output[8]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[0]), .Z(n8)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(74[27:78])
    defparam i10827_3_lut.init = 16'hcaca;
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i16 (.D(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[16]), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(modulation_deviation_amount_minus_sine_lookup_width[16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i16.GSR = "DISABLED";
    LUT4 modulation_output_15__I_0_i38_3_lut (.A(n7), .B(n9), .C(sine_lookup_width_minus_modulation_deviation_amount[1]), 
         .Z(n38)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam modulation_output_15__I_0_i38_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i73_3_lut (.A(n42), .B(n46), .C(sine_lookup_width_minus_modulation_deviation_amount[2]), 
         .Z(n73)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam modulation_output_15__I_0_i73_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i42_3_lut (.A(n11), .B(n13), .C(sine_lookup_width_minus_modulation_deviation_amount[1]), 
         .Z(n42)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam modulation_output_15__I_0_i42_3_lut.init = 16'hcaca;
    LUT4 i17726_3_lut (.A(\addr_space[0] [4]), .B(\addr_space[1] [4]), .C(\wb_addr[0] ), 
         .Z(n20056)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17726_3_lut.init = 16'hcaca;
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i15 (.D(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[15]), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(modulation_deviation_amount_minus_sine_lookup_width[15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i15.GSR = "DISABLED";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i14 (.D(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[14]), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(modulation_deviation_amount_minus_sine_lookup_width[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i14.GSR = "DISABLED";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i13 (.D(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[13]), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(modulation_deviation_amount_minus_sine_lookup_width[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i13.GSR = "DISABLED";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i12 (.D(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[12]), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(modulation_deviation_amount_minus_sine_lookup_width[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i12.GSR = "DISABLED";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i11 (.D(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[11]), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(modulation_deviation_amount_minus_sine_lookup_width[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i11.GSR = "DISABLED";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i10 (.D(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[10]), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(modulation_deviation_amount_minus_sine_lookup_width[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i10.GSR = "DISABLED";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i9 (.D(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[9]), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(modulation_deviation_amount_minus_sine_lookup_width[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i9.GSR = "DISABLED";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i8 (.D(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[8]), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(modulation_deviation_amount_minus_sine_lookup_width[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i8.GSR = "DISABLED";
    PFUMX modulation_output_15__I_0_332_i135 (.BLUT(n73_adj_3015), .ALUT(n104), 
          .C0(n19807), .Z(n135)) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i7 (.D(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[7]), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(modulation_deviation_amount_minus_sine_lookup_width[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i7.GSR = "DISABLED";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i6 (.D(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[6]), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(modulation_deviation_amount_minus_sine_lookup_width[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i6.GSR = "DISABLED";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i5 (.D(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[5]), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(modulation_deviation_amount_minus_sine_lookup_width[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i5.GSR = "DISABLED";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i4 (.D(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[4]), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(modulation_deviation_amount_minus_sine_lookup_width[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i4.GSR = "DISABLED";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i3 (.D(\addr_space[2] [3]), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(modulation_deviation_amount_minus_sine_lookup_width[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i3.GSR = "DISABLED";
    PFUMX modulation_output_15__I_0_332_i134 (.BLUT(n72_adj_3016), .ALUT(n103), 
          .C0(n19807), .Z(n134)) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i2 (.D(\addr_space[2] [2]), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(modulation_deviation_amount_minus_sine_lookup_width[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i2.GSR = "DISABLED";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i1 (.D(\addr_space[2] [1]), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(modulation_deviation_amount_minus_sine_lookup_width[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i1.GSR = "DISABLED";
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i16 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[16]), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(sine_lookup_width_minus_modulation_deviation_amount[16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i16.GSR = "DISABLED";
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i15 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[15]), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(sine_lookup_width_minus_modulation_deviation_amount[15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i15.GSR = "DISABLED";
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i14 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[14]), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(sine_lookup_width_minus_modulation_deviation_amount[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i14.GSR = "DISABLED";
    PFUMX i17716 (.BLUT(n20044), .ALUT(n20045), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[8]));
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i13 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[13]), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(sine_lookup_width_minus_modulation_deviation_amount[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i13.GSR = "DISABLED";
    LUT4 n13476_bdd_3_lut_22815 (.A(modulation_output[2]), .B(modulation_output[1]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[0]), .Z(n22765)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n13476_bdd_3_lut_22815.init = 16'hacac;
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i12 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[12]), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(sine_lookup_width_minus_modulation_deviation_amount[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i12.GSR = "DISABLED";
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i11 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[11]), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(sine_lookup_width_minus_modulation_deviation_amount[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i11.GSR = "DISABLED";
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i10 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[10]), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(sine_lookup_width_minus_modulation_deviation_amount[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i10.GSR = "DISABLED";
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i9 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[9]), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(sine_lookup_width_minus_modulation_deviation_amount[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i9.GSR = "DISABLED";
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i8 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[8]), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(sine_lookup_width_minus_modulation_deviation_amount[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i8.GSR = "DISABLED";
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i7 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[7]), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(sine_lookup_width_minus_modulation_deviation_amount[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i7.GSR = "DISABLED";
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i6 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[6]), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(sine_lookup_width_minus_modulation_deviation_amount[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i6.GSR = "DISABLED";
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i5 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[5]), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(sine_lookup_width_minus_modulation_deviation_amount[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i5.GSR = "DISABLED";
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i4 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[4]), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(sine_lookup_width_minus_modulation_deviation_amount[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i4.GSR = "DISABLED";
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i3 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[3]), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(sine_lookup_width_minus_modulation_deviation_amount[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i3.GSR = "DISABLED";
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i2 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[2]), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(sine_lookup_width_minus_modulation_deviation_amount[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i2.GSR = "DISABLED";
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i1 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[1]), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(sine_lookup_width_minus_modulation_deviation_amount[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i1.GSR = "DISABLED";
    FD1S3DX carrier_increment_i30 (.D(carrier_increment_30__N_1591[30]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(carrier_increment[30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_increment_i30.GSR = "DISABLED";
    FD1S3DX carrier_increment_i29 (.D(carrier_increment_30__N_1591[29]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(carrier_increment[29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_increment_i29.GSR = "DISABLED";
    FD1S3DX carrier_increment_i28 (.D(carrier_increment_30__N_1591[28]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(carrier_increment[28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_increment_i28.GSR = "DISABLED";
    FD1S3DX carrier_increment_i27 (.D(carrier_increment_30__N_1591[27]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(carrier_increment[27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_increment_i27.GSR = "DISABLED";
    FD1S3DX carrier_increment_i26 (.D(carrier_increment_30__N_1591[26]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(carrier_increment[26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_increment_i26.GSR = "DISABLED";
    FD1S3DX carrier_increment_i25 (.D(carrier_increment_30__N_1591[25]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(carrier_increment[25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_increment_i25.GSR = "DISABLED";
    FD1S3DX carrier_increment_i24 (.D(carrier_increment_30__N_1591[24]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(carrier_increment[24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_increment_i24.GSR = "DISABLED";
    FD1S3DX carrier_increment_i23 (.D(carrier_increment_30__N_1591[23]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(carrier_increment[23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_increment_i23.GSR = "DISABLED";
    FD1S3DX carrier_increment_i22 (.D(carrier_increment_30__N_1591[22]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(carrier_increment[22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_increment_i22.GSR = "DISABLED";
    FD1S3DX carrier_increment_i21 (.D(carrier_increment_30__N_1591[21]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(carrier_increment[21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_increment_i21.GSR = "DISABLED";
    FD1S3DX carrier_increment_i20 (.D(carrier_increment_30__N_1591[20]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(carrier_increment[20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_increment_i20.GSR = "DISABLED";
    FD1S3DX carrier_increment_i19 (.D(carrier_increment_30__N_1591[19]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(carrier_increment[19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_increment_i19.GSR = "DISABLED";
    FD1S3DX carrier_increment_i18 (.D(carrier_increment_30__N_1591[18]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(carrier_increment[18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_increment_i18.GSR = "DISABLED";
    FD1S3DX carrier_increment_i17 (.D(carrier_increment_30__N_1591[17]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(carrier_increment[17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_increment_i17.GSR = "DISABLED";
    FD1S3DX carrier_increment_i16 (.D(carrier_increment_30__N_1591[16]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(carrier_increment[16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_increment_i16.GSR = "DISABLED";
    FD1S3DX carrier_increment_i15 (.D(carrier_increment_30__N_1591[15]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(carrier_increment[15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_increment_i15.GSR = "DISABLED";
    FD1S3DX carrier_increment_i14 (.D(carrier_increment_30__N_1591[14]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(carrier_increment[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_increment_i14.GSR = "DISABLED";
    LUT4 n22766_bdd_3_lut (.A(n22766), .B(n37), .C(sine_lookup_width_minus_modulation_deviation_amount[2]), 
         .Z(n22767)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n22766_bdd_3_lut.init = 16'hcaca;
    LUT4 i10817_3_lut_rep_259_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[2]), 
         .B(n24988), .C(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .D(n85), .Z(n24819)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i10817_3_lut_rep_259_4_lut.init = 16'h4f40;
    FD1S3DX carrier_increment_i13 (.D(carrier_increment_30__N_1591[13]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(carrier_increment[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_increment_i13.GSR = "DISABLED";
    FD1S3DX carrier_increment_i12 (.D(carrier_increment_30__N_1591[12]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(carrier_increment[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_increment_i12.GSR = "DISABLED";
    FD1S3DX carrier_increment_i11 (.D(carrier_increment_30__N_1591[11]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(carrier_increment[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_increment_i11.GSR = "DISABLED";
    FD1S3DX carrier_increment_i10 (.D(carrier_increment_30__N_1591[10]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(carrier_increment[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_increment_i10.GSR = "DISABLED";
    FD1S3DX carrier_increment_i9 (.D(carrier_increment_30__N_1591[9]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(carrier_increment[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_increment_i9.GSR = "DISABLED";
    LUT4 n24517_bdd_3_lut (.A(n24517), .B(n24515), .C(sine_lookup_width_minus_modulation_deviation_amount[3]), 
         .Z(n24518)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n24517_bdd_3_lut.init = 16'hcaca;
    FD1S3DX carrier_increment_i8 (.D(carrier_increment_30__N_1591[8]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(carrier_increment[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_increment_i8.GSR = "DISABLED";
    FD1S3DX carrier_increment_i7 (.D(carrier_increment_30__N_1591[7]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(carrier_increment[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_increment_i7.GSR = "DISABLED";
    FD1S3DX carrier_increment_i6 (.D(carrier_increment_30__N_1591[6]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(carrier_increment[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_increment_i6.GSR = "DISABLED";
    FD1S3DX carrier_increment_i5 (.D(carrier_increment_30__N_1591[5]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(carrier_increment[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_increment_i5.GSR = "DISABLED";
    FD1S3DX carrier_increment_i4 (.D(carrier_increment_30__N_1591[4]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(carrier_increment[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_increment_i4.GSR = "DISABLED";
    FD1S3DX carrier_increment_i3 (.D(carrier_increment_30__N_1591[3]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(carrier_increment[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_increment_i3.GSR = "DISABLED";
    FD1S3DX carrier_increment_i2 (.D(carrier_increment_30__N_1591[2]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(carrier_increment[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_increment_i2.GSR = "DISABLED";
    FD1S3DX carrier_increment_i1 (.D(carrier_increment_30__N_1591[1]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(carrier_increment[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_increment_i1.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_rs_i16 (.D(modulation_output[15]), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_rs[30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_rs_i16.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_rs_i15 (.D(carrier_center_increment_offset_rs_30__N_1560[14]), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_rs[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_rs_i15.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_rs_i14 (.D(carrier_center_increment_offset_rs_30__N_1560[13]), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_rs[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_rs_i14.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_rs_i13 (.D(carrier_center_increment_offset_rs_30__N_1560[12]), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_rs[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_rs_i13.GSR = "DISABLED";
    LUT4 n38_bdd_3_lut_22704 (.A(n13468), .B(n13470), .C(sine_lookup_width_minus_modulation_deviation_amount[1]), 
         .Z(n22770)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n38_bdd_3_lut_22704.init = 16'hcaca;
    FD1S3DX carrier_center_increment_offset_rs_i12 (.D(carrier_center_increment_offset_rs_30__N_1560[11]), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_rs[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_rs_i12.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_rs_i11 (.D(carrier_center_increment_offset_rs_30__N_1560[10]), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_rs[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_rs_i11.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_rs_i10 (.D(carrier_center_increment_offset_rs_30__N_1560[9]), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_rs[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_rs_i10.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_rs_i9 (.D(carrier_center_increment_offset_rs_30__N_1560[8]), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_rs[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_rs_i9.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_rs_i8 (.D(carrier_center_increment_offset_rs_30__N_1560[7]), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_rs[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_rs_i8.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_rs_i7 (.D(carrier_center_increment_offset_rs_30__N_1560[6]), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_rs[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_rs_i7.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_rs_i6 (.D(carrier_center_increment_offset_rs_30__N_1560[5]), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_rs[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_rs_i6.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_rs_i5 (.D(carrier_center_increment_offset_rs_30__N_1560[4]), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_rs[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_rs_i5.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_rs_i4 (.D(carrier_center_increment_offset_rs_30__N_1560[3]), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_rs[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_rs_i4.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_rs_i3 (.D(carrier_center_increment_offset_rs_30__N_1560[2]), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_rs[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_rs_i3.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_rs_i2 (.D(carrier_center_increment_offset_rs_30__N_1560[1]), 
            .CK(i_ref_clk_c), .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_rs[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_rs_i2.GSR = "DISABLED";
    FD1S3AX o_wb_data_i31 (.D(o_wb_data_31__N_1337[31]), .CK(i_ref_clk_c), 
            .Q(wb_fm_data[31])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i31.GSR = "DISABLED";
    FD1S3AX o_wb_data_i30 (.D(o_wb_data_31__N_1337[30]), .CK(i_ref_clk_c), 
            .Q(wb_fm_data[30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i30.GSR = "DISABLED";
    FD1S3AX o_wb_data_i29 (.D(o_wb_data_31__N_1337[29]), .CK(i_ref_clk_c), 
            .Q(wb_fm_data[29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i29.GSR = "DISABLED";
    FD1S3AX o_wb_data_i28 (.D(o_wb_data_31__N_1337[28]), .CK(i_ref_clk_c), 
            .Q(wb_fm_data[28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i28.GSR = "DISABLED";
    FD1S3AX o_wb_data_i27 (.D(o_wb_data_31__N_1337[27]), .CK(i_ref_clk_c), 
            .Q(wb_fm_data[27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i27.GSR = "DISABLED";
    FD1S3AX o_wb_data_i26 (.D(o_wb_data_31__N_1337[26]), .CK(i_ref_clk_c), 
            .Q(wb_fm_data[26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i26.GSR = "DISABLED";
    FD1S3AX o_wb_data_i25 (.D(o_wb_data_31__N_1337[25]), .CK(i_ref_clk_c), 
            .Q(wb_fm_data[25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i25.GSR = "DISABLED";
    FD1S3AX o_wb_data_i24 (.D(o_wb_data_31__N_1337[24]), .CK(i_ref_clk_c), 
            .Q(wb_fm_data[24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i24.GSR = "DISABLED";
    FD1S3AX o_wb_data_i23 (.D(o_wb_data_31__N_1337[23]), .CK(i_ref_clk_c), 
            .Q(wb_fm_data[23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i23.GSR = "DISABLED";
    FD1S3AX o_wb_data_i22 (.D(o_wb_data_31__N_1337[22]), .CK(i_ref_clk_c), 
            .Q(wb_fm_data[22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i22.GSR = "DISABLED";
    FD1S3AX o_wb_data_i21 (.D(o_wb_data_31__N_1337[21]), .CK(i_ref_clk_c), 
            .Q(wb_fm_data[21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i21.GSR = "DISABLED";
    FD1S3AX o_wb_data_i20 (.D(o_wb_data_31__N_1337[20]), .CK(i_ref_clk_c), 
            .Q(wb_fm_data[20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i20.GSR = "DISABLED";
    FD1S3AX o_wb_data_i19 (.D(o_wb_data_31__N_1337[19]), .CK(i_ref_clk_c), 
            .Q(wb_fm_data[19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i19.GSR = "DISABLED";
    FD1S3AX o_wb_data_i18 (.D(o_wb_data_31__N_1337[18]), .CK(i_ref_clk_c), 
            .Q(wb_fm_data[18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i18.GSR = "DISABLED";
    FD1S3AX o_wb_data_i17 (.D(o_wb_data_31__N_1337[17]), .CK(i_ref_clk_c), 
            .Q(wb_fm_data[17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i17.GSR = "DISABLED";
    FD1S3AX o_wb_data_i16 (.D(o_wb_data_31__N_1337[16]), .CK(i_ref_clk_c), 
            .Q(wb_fm_data[16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i16.GSR = "DISABLED";
    FD1S3AX o_wb_data_i15 (.D(o_wb_data_31__N_1337[15]), .CK(i_ref_clk_c), 
            .Q(wb_fm_data[15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i15.GSR = "DISABLED";
    FD1S3AX o_wb_data_i14 (.D(o_wb_data_31__N_1337[14]), .CK(i_ref_clk_c), 
            .Q(wb_fm_data[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i14.GSR = "DISABLED";
    FD1S3AX o_wb_data_i13 (.D(o_wb_data_31__N_1337[13]), .CK(i_ref_clk_c), 
            .Q(wb_fm_data[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i13.GSR = "DISABLED";
    FD1S3AX o_wb_data_i12 (.D(o_wb_data_31__N_1337[12]), .CK(i_ref_clk_c), 
            .Q(wb_fm_data[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i12.GSR = "DISABLED";
    FD1S3AX o_wb_data_i11 (.D(o_wb_data_31__N_1337[11]), .CK(i_ref_clk_c), 
            .Q(wb_fm_data[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i11.GSR = "DISABLED";
    FD1S3AX o_wb_data_i10 (.D(o_wb_data_31__N_1337[10]), .CK(i_ref_clk_c), 
            .Q(wb_fm_data[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i10.GSR = "DISABLED";
    FD1S3AX o_wb_data_i9 (.D(o_wb_data_31__N_1337[9]), .CK(i_ref_clk_c), 
            .Q(wb_fm_data[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i9.GSR = "DISABLED";
    FD1S3AX o_wb_data_i8 (.D(o_wb_data_31__N_1337[8]), .CK(i_ref_clk_c), 
            .Q(wb_fm_data[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i8.GSR = "DISABLED";
    FD1S3AX o_wb_data_i7 (.D(o_wb_data_31__N_1337[7]), .CK(i_ref_clk_c), 
            .Q(wb_fm_data[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i7.GSR = "DISABLED";
    FD1S3AX o_wb_data_i6 (.D(o_wb_data_31__N_1337[6]), .CK(i_ref_clk_c), 
            .Q(wb_fm_data[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i6.GSR = "DISABLED";
    FD1S3AX o_wb_data_i5 (.D(o_wb_data_31__N_1337[5]), .CK(i_ref_clk_c), 
            .Q(wb_fm_data[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i5.GSR = "DISABLED";
    FD1S3AX o_wb_data_i4 (.D(o_wb_data_31__N_1337[4]), .CK(i_ref_clk_c), 
            .Q(wb_fm_data[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i4.GSR = "DISABLED";
    FD1S3AX o_wb_data_i3 (.D(o_wb_data_31__N_1337[3]), .CK(i_ref_clk_c), 
            .Q(wb_fm_data[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i3.GSR = "DISABLED";
    FD1S3AX o_wb_data_i2 (.D(o_wb_data_31__N_1337[2]), .CK(i_ref_clk_c), 
            .Q(wb_fm_data[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i2.GSR = "DISABLED";
    FD1S3AX o_wb_data_i1 (.D(o_wb_data_31__N_1337[1]), .CK(i_ref_clk_c), 
            .Q(wb_fm_data[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i1.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i30 (.D(n64[30]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_ls[30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_ls__i30.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i29 (.D(n64[29]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_ls[29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_ls__i29.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i28 (.D(n64[28]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_ls[28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_ls__i28.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i27 (.D(n64[27]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_ls[27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_ls__i27.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i26 (.D(n64[26]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_ls[26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_ls__i26.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i25 (.D(n64[25]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_ls[25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_ls__i25.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i24 (.D(n64[24]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_ls[24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_ls__i24.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i23 (.D(n64[23]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_ls[23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_ls__i23.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i22 (.D(n64[22]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_ls[22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_ls__i22.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i21 (.D(n64[21]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_ls[21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_ls__i21.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i20 (.D(n64[20]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_ls[20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_ls__i20.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i19 (.D(n64[19]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_ls[19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_ls__i19.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i18 (.D(n64[18]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_ls[18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_ls__i18.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i17 (.D(n64[17]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_ls[17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_ls__i17.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i16 (.D(n64[16]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_ls[16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_ls__i16.GSR = "DISABLED";
    PFUMX i22838 (.BLUT(n24548), .ALUT(n24547), .C0(sine_lookup_width_minus_modulation_deviation_amount[3]), 
          .Z(n24549));
    FD1S3DX carrier_center_increment_offset_ls__i15 (.D(n64[15]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_ls[15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_ls__i15.GSR = "DISABLED";
    LUT4 n22771_bdd_3_lut (.A(n22771), .B(n73), .C(sine_lookup_width_minus_modulation_deviation_amount[3]), 
         .Z(n22772)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n22771_bdd_3_lut.init = 16'hcaca;
    FD1S3DX carrier_center_increment_offset_ls__i14 (.D(n64[14]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_ls[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_ls__i14.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i13 (.D(n64[13]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_ls[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_ls__i13.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i12 (.D(n64[12]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_ls[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_ls__i12.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i11 (.D(n64[11]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_ls[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_ls__i11.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i10 (.D(n64[10]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_ls[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_ls__i10.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i9 (.D(n64[9]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_ls[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_ls__i9.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i8 (.D(n64[8]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_ls[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_ls__i8.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i7 (.D(n64[7]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_ls[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_ls__i7.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i6 (.D(n64[6]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_ls[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_ls__i6.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i5 (.D(n64[5]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_ls[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_ls__i5.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i4 (.D(n64[4]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_ls[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_ls__i4.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i3 (.D(n64[3]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_ls[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_ls__i3.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i2 (.D(n64[2]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_ls[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_ls__i2.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i1 (.D(n17801), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_ls[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_ls__i1.GSR = "DISABLED";
    LUT4 i12_4_lut (.A(\addr_space[2] [8]), .B(n24), .C(n20_adj_3027), 
         .D(\addr_space[2] [11]), .Z(n14286)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i12_4_lut.init = 16'hfffe;
    LUT4 i11_4_lut_adj_89 (.A(\addr_space[2] [5]), .B(n22_adj_3028), .C(n16), 
         .D(\addr_space[2] [10]), .Z(n24)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i11_4_lut_adj_89.init = 16'hfffe;
    LUT4 i7_3_lut (.A(\addr_space[2] [16]), .B(\addr_space[2] [4]), .C(\addr_space[2] [14]), 
         .Z(n20_adj_3027)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i7_3_lut.init = 16'hfefe;
    LUT4 i9_4_lut (.A(\addr_space[2] [13]), .B(\addr_space[2] [7]), .C(\addr_space[2] [15]), 
         .D(\addr_space[2] [6]), .Z(n22_adj_3028)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i9_4_lut.init = 16'hfffe;
    LUT4 i3_2_lut (.A(\addr_space[2] [12]), .B(\addr_space[2] [9]), .Z(n16)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i3_2_lut.init = 16'heeee;
    PFUMX i22829 (.BLUT(n24538), .ALUT(n24537), .C0(sine_lookup_width_minus_modulation_deviation_amount[3]), 
          .Z(n24539));
    PFUMX i22821 (.BLUT(n24525), .ALUT(n24524), .C0(sine_lookup_width_minus_modulation_deviation_amount[3]), 
          .Z(n24526));
    PFUMX i22813 (.BLUT(n24516), .ALUT(n39_adj_3029), .C0(sine_lookup_width_minus_modulation_deviation_amount[2]), 
          .Z(n24517));
    LUT4 i17724_3_lut (.A(\addr_space[2] [5]), .B(\addr_space[3] [5]), .C(\wb_addr[0] ), 
         .Z(n20054)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17724_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_332_i101_3_lut (.A(modulation_output[15]), 
         .B(n78), .C(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .Z(n101)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i101_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_332_i102_3_lut (.A(modulation_output[15]), 
         .B(n79), .C(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .Z(n102)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i102_3_lut.init = 16'hcaca;
    LUT4 i11512_2_lut_3_lut_4_lut_4_lut (.A(n25008), .B(n60_adj_3030), .C(n178_adj_3009), 
         .D(modulation_deviation_amount_minus_sine_lookup_width[4]), .Z(n64[2])) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam i11512_2_lut_3_lut_4_lut_4_lut.init = 16'h0008;
    LUT4 i11513_2_lut_3_lut_4_lut_4_lut (.A(n25008), .B(n59_adj_3031), .C(n178_adj_3009), 
         .D(modulation_deviation_amount_minus_sine_lookup_width[4]), .Z(n64[3])) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam i11513_2_lut_3_lut_4_lut_4_lut.init = 16'h0008;
    LUT4 modulation_output_15__I_0_332_i105_4_lut (.A(n82), .B(n59_adj_3031), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[4]), .D(n25008), 
         .Z(n105)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i105_4_lut.init = 16'hca0a;
    LUT4 modulation_output_15__I_0_332_i74_3_lut (.A(modulation_output[15]), 
         .B(n47_adj_3032), .C(modulation_deviation_amount_minus_sine_lookup_width[2]), 
         .Z(n74)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i74_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_332_i106_4_lut (.A(n83), .B(n60_adj_3030), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[4]), .D(n25008), 
         .Z(n106)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i106_4_lut.init = 16'hca0a;
    LUT4 modulation_output_15__I_0_332_i75_3_lut (.A(modulation_output[15]), 
         .B(n48_adj_3033), .C(modulation_deviation_amount_minus_sine_lookup_width[2]), 
         .Z(n75)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i75_3_lut.init = 16'hcaca;
    LUT4 i17723_3_lut (.A(\addr_space[0] [5]), .B(\addr_space[1] [5]), .C(\wb_addr[0] ), 
         .Z(n20053)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17723_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_332_i86_3_lut_rep_286 (.A(n55_adj_3034), 
         .B(n59_adj_3031), .C(modulation_deviation_amount_minus_sine_lookup_width[2]), 
         .Z(n24846)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i86_3_lut_rep_286.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_332_i87_3_lut_rep_290 (.A(n56_adj_3035), 
         .B(n60_adj_3030), .C(modulation_deviation_amount_minus_sine_lookup_width[2]), 
         .Z(n24850)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i87_3_lut_rep_290.init = 16'hcaca;
    LUT4 i17721_3_lut (.A(\addr_space[2] [6]), .B(\addr_space[3] [6]), .C(\wb_addr[0] ), 
         .Z(n20051)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17721_3_lut.init = 16'hcaca;
    LUT4 i6466_3_lut_4_lut (.A(n25012), .B(modulation_deviation_amount_minus_sine_lookup_width[2]), 
         .C(modulation_output[14]), .D(modulation_output[15]), .Z(n72_adj_3016)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam i6466_3_lut_4_lut.init = 16'hf780;
    LUT4 i11519_2_lut_4_lut (.A(n85), .B(n24888), .C(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .D(n24834), .Z(n64[8])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(74[80:131])
    defparam i11519_2_lut_4_lut.init = 16'h00ca;
    LUT4 modulation_output_15__I_0_332_i112_3_lut_rep_260 (.A(n81), .B(n89), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[3]), .Z(n24820)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i112_3_lut_rep_260.init = 16'hcaca;
    LUT4 i11523_2_lut_4_lut (.A(n81), .B(n89), .C(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .D(n24834), .Z(n64[12])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam i11523_2_lut_4_lut.init = 16'h00ca;
    LUT4 modulation_output_15__I_0_332_i111_3_lut_rep_261 (.A(n80), .B(n88), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[3]), .Z(n24821)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i111_3_lut_rep_261.init = 16'hcaca;
    LUT4 i11524_2_lut_4_lut (.A(n80), .B(n88), .C(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .D(n24834), .Z(n64[13])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam i11524_2_lut_4_lut.init = 16'h00ca;
    LUT4 modulation_output_15__I_0_332_i110_3_lut_rep_262 (.A(n79), .B(n24850), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[3]), .Z(n24822)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i110_3_lut_rep_262.init = 16'hcaca;
    LUT4 i11525_2_lut_4_lut (.A(n79), .B(n24850), .C(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .D(n24834), .Z(n64[14])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam i11525_2_lut_4_lut.init = 16'h00ca;
    LUT4 i2_3_lut_rep_263 (.A(n178), .B(sine_lookup_width_minus_modulation_deviation_amount[4]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[3]), .Z(n24823)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam i2_3_lut_rep_263.init = 16'hfefe;
    LUT4 i1_2_lut_rep_627 (.A(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .B(modulation_output[0]), .Z(n25187)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i1_2_lut_rep_627.init = 16'h4444;
    LUT4 i1_2_lut_rep_428_3_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .B(modulation_output[0]), .C(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .Z(n24988)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i1_2_lut_rep_428_3_lut.init = 16'h0404;
    LUT4 i1_2_lut_rep_328_3_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .B(modulation_output[0]), .C(modulation_deviation_amount_minus_sine_lookup_width[2]), 
         .D(modulation_deviation_amount_minus_sine_lookup_width[1]), .Z(n24888)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i1_2_lut_rep_328_3_lut_4_lut.init = 16'h0004;
    LUT4 modulation_output_15__I_0_332_i60_3_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .B(modulation_output[0]), .C(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .D(n29), .Z(n60_adj_3030)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam modulation_output_15__I_0_332_i60_3_lut_4_lut.init = 16'h4f40;
    LUT4 i17685_3_lut (.A(\addr_space[2] [18]), .B(\addr_space[3] [18]), 
         .C(\wb_addr[0] ), .Z(n20015)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17685_3_lut.init = 16'hcaca;
    LUT4 i17684_3_lut (.A(\addr_space[0] [18]), .B(\addr_space[1] [18]), 
         .C(\wb_addr[0] ), .Z(n20014)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17684_3_lut.init = 16'hcaca;
    LUT4 i17682_3_lut (.A(\addr_space[2] [19]), .B(\addr_space[3] [19]), 
         .C(\wb_addr[0] ), .Z(n20012)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17682_3_lut.init = 16'hcaca;
    LUT4 i17681_3_lut (.A(\addr_space[0] [19]), .B(\addr_space[1] [19]), 
         .C(\wb_addr[0] ), .Z(n20011)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17681_3_lut.init = 16'hcaca;
    LUT4 i17679_3_lut (.A(\addr_space[2] [20]), .B(\addr_space[3] [20]), 
         .C(\wb_addr[0] ), .Z(n20009)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17679_3_lut.init = 16'hcaca;
    LUT4 i17678_3_lut (.A(\addr_space[0] [20]), .B(\addr_space[1] [20]), 
         .C(\wb_addr[0] ), .Z(n20008)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17678_3_lut.init = 16'hcaca;
    LUT4 i17676_3_lut (.A(\addr_space[2] [21]), .B(\addr_space[3] [21]), 
         .C(\wb_addr[0] ), .Z(n20006)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17676_3_lut.init = 16'hcaca;
    LUT4 i17675_3_lut (.A(\addr_space[0] [21]), .B(\addr_space[1] [21]), 
         .C(\wb_addr[0] ), .Z(n20005)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17675_3_lut.init = 16'hcaca;
    PFUMX i17719 (.BLUT(n20047), .ALUT(n20048), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[7]));
    LUT4 i19245_3_lut (.A(\addr_space[2] [30]), .B(\addr_space[3] [30]), 
         .C(\wb_addr[0] ), .Z(n21575)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19245_3_lut.init = 16'hcaca;
    LUT4 i19244_3_lut (.A(\addr_space[0] [30]), .B(\addr_space[1] [30]), 
         .C(\wb_addr[0] ), .Z(n21574)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19244_3_lut.init = 16'hcaca;
    LUT4 i17673_3_lut (.A(\addr_space[2] [22]), .B(\addr_space[3] [22]), 
         .C(\wb_addr[0] ), .Z(n20003)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17673_3_lut.init = 16'hcaca;
    LUT4 i17672_3_lut (.A(\addr_space[0] [22]), .B(\addr_space[1] [22]), 
         .C(\wb_addr[0] ), .Z(n20002)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17672_3_lut.init = 16'hcaca;
    LUT4 i17670_3_lut (.A(\addr_space[2] [23]), .B(\addr_space[3] [23]), 
         .C(\wb_addr[0] ), .Z(n20000)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17670_3_lut.init = 16'hcaca;
    LUT4 i17669_3_lut (.A(\addr_space[0] [23]), .B(\addr_space[1] [23]), 
         .C(\wb_addr[0] ), .Z(n19999)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17669_3_lut.init = 16'hcaca;
    LUT4 i17667_3_lut (.A(\addr_space[2] [24]), .B(\addr_space[3] [24]), 
         .C(\wb_addr[0] ), .Z(n19997)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17667_3_lut.init = 16'hcaca;
    LUT4 i17666_3_lut (.A(\addr_space[0] [24]), .B(\addr_space[1] [24]), 
         .C(\wb_addr[0] ), .Z(n19996)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17666_3_lut.init = 16'hcaca;
    LUT4 i19236_3_lut (.A(\addr_space[2] [31]), .B(\addr_space[3] [31]), 
         .C(\wb_addr[0] ), .Z(n21566)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19236_3_lut.init = 16'hcaca;
    LUT4 i19235_3_lut (.A(\addr_space[0] [31]), .B(\addr_space[1] [31]), 
         .C(\wb_addr[0] ), .Z(n21565)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19235_3_lut.init = 16'hcaca;
    LUT4 i19233_3_lut (.A(\addr_space[2] [0]), .B(\addr_space[3] [0]), .C(\wb_addr[0] ), 
         .Z(n21563)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19233_3_lut.init = 16'hcaca;
    LUT4 i19232_3_lut (.A(\addr_space[0] [0]), .B(\addr_space[1] [0]), .C(\wb_addr[0] ), 
         .Z(n21562)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19232_3_lut.init = 16'hcaca;
    LUT4 i17661_3_lut (.A(\addr_space[2] [25]), .B(\addr_space[3] [25]), 
         .C(\wb_addr[0] ), .Z(n19991)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17661_3_lut.init = 16'hcaca;
    LUT4 i17660_3_lut (.A(\addr_space[0] [25]), .B(\addr_space[1] [25]), 
         .C(\wb_addr[0] ), .Z(n19990)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17660_3_lut.init = 16'hcaca;
    PFUMX i17722 (.BLUT(n20050), .ALUT(n20051), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[6]));
    LUT4 i17658_3_lut (.A(\addr_space[2] [26]), .B(\addr_space[3] [26]), 
         .C(\wb_addr[0] ), .Z(n19988)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17658_3_lut.init = 16'hcaca;
    LUT4 i17657_3_lut (.A(\addr_space[0] [26]), .B(\addr_space[1] [26]), 
         .C(\wb_addr[0] ), .Z(n19987)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17657_3_lut.init = 16'hcaca;
    LUT4 i17655_3_lut (.A(\addr_space[2] [27]), .B(\addr_space[3] [27]), 
         .C(\wb_addr[0] ), .Z(n19985)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17655_3_lut.init = 16'hcaca;
    LUT4 i17654_3_lut (.A(\addr_space[0] [27]), .B(\addr_space[1] [27]), 
         .C(\wb_addr[0] ), .Z(n19984)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17654_3_lut.init = 16'hcaca;
    LUT4 i17652_3_lut (.A(\addr_space[2] [28]), .B(\addr_space[3] [28]), 
         .C(\wb_addr[0] ), .Z(n19982)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17652_3_lut.init = 16'hcaca;
    LUT4 i17651_3_lut (.A(\addr_space[0] [28]), .B(\addr_space[1] [28]), 
         .C(\wb_addr[0] ), .Z(n19981)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17651_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_332_i17_3_lut (.A(modulation_output[14]), 
         .B(modulation_output[13]), .C(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .Z(n17)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i17_3_lut.init = 16'hcaca;
    LUT4 i17649_3_lut (.A(\addr_space[2] [29]), .B(\addr_space[3] [29]), 
         .C(\wb_addr[0] ), .Z(n19979)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17649_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_332_i81_3_lut (.A(n50_adj_3036), .B(n54_adj_3037), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[2]), .Z(n81)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i81_3_lut.init = 16'hcaca;
    LUT4 i17648_3_lut (.A(\addr_space[0] [29]), .B(\addr_space[1] [29]), 
         .C(\wb_addr[0] ), .Z(n19978)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17648_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_332_i58_3_lut (.A(n27), .B(n29), .C(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .Z(n58_adj_3038)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i58_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_332_i50_3_lut (.A(n19), .B(n21), .C(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .Z(n50_adj_3036)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i50_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_332_i54_3_lut (.A(n23), .B(n25), .C(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .Z(n54_adj_3037)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i54_3_lut.init = 16'hcaca;
    LUT4 i10826_3_lut (.A(modulation_output[8]), .B(modulation_output[7]), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[0]), .Z(n23)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(74[80:131])
    defparam i10826_3_lut.init = 16'hcaca;
    LUT4 i10829_3_lut (.A(modulation_output[6]), .B(modulation_output[5]), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[0]), .Z(n25)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(74[80:131])
    defparam i10829_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_332_i19_3_lut (.A(modulation_output[12]), 
         .B(modulation_output[11]), .C(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .Z(n19)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i19_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_332_i21_3_lut (.A(modulation_output[10]), 
         .B(modulation_output[9]), .C(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .Z(n21)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i21_3_lut.init = 16'hcaca;
    LUT4 i10834_3_lut (.A(modulation_output[4]), .B(modulation_output[3]), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[0]), .Z(n27)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(74[80:131])
    defparam i10834_3_lut.init = 16'hcaca;
    LUT4 i10828_3_lut (.A(modulation_output[2]), .B(modulation_output[1]), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[0]), .Z(n29)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(74[80:131])
    defparam i10828_3_lut.init = 16'hcaca;
    LUT4 i21161_2_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[3]), .Z(n19807)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam i21161_2_lut.init = 16'heeee;
    LUT4 modulation_output_15__I_0_332_i80_3_lut (.A(n49_adj_3039), .B(n53_adj_3040), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[2]), .Z(n80)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i80_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_332_i88_4_lut (.A(n57_adj_3041), .B(n30), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[2]), .D(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .Z(n88)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i88_4_lut.init = 16'h0aca;
    LUT4 modulation_output_15__I_0_332_i57_3_lut (.A(n26), .B(n28), .C(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .Z(n57_adj_3041)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i57_3_lut.init = 16'hcaca;
    LUT4 i10830_3_lut (.A(modulation_output[1]), .B(modulation_output[0]), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[0]), .Z(n30)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(74[80:131])
    defparam i10830_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_332_i49_3_lut (.A(n18_adj_3042), .B(n20_adj_3043), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[1]), .Z(n49_adj_3039)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i49_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_332_i53_3_lut (.A(n22_adj_3044), .B(n24_adj_3045), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[1]), .Z(n53_adj_3040)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i53_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_332_i18_3_lut (.A(modulation_output[13]), 
         .B(modulation_output[12]), .C(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .Z(n18_adj_3042)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i18_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_332_i20_3_lut (.A(modulation_output[11]), 
         .B(modulation_output[10]), .C(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .Z(n20_adj_3043)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i20_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_332_i22_3_lut (.A(modulation_output[9]), 
         .B(modulation_output[8]), .C(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .Z(n22_adj_3044)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i22_3_lut.init = 16'hcaca;
    LUT4 i10831_3_lut (.A(modulation_output[7]), .B(modulation_output[6]), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[0]), .Z(n24_adj_3045)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(74[80:131])
    defparam i10831_3_lut.init = 16'hcaca;
    LUT4 i10832_3_lut (.A(modulation_output[5]), .B(modulation_output[4]), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[0]), .Z(n26)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(74[80:131])
    defparam i10832_3_lut.init = 16'hcaca;
    LUT4 i10833_3_lut (.A(modulation_output[3]), .B(modulation_output[2]), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[0]), .Z(n28)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(74[80:131])
    defparam i10833_3_lut.init = 16'hcaca;
    LUT4 n36_bdd_3_lut (.A(n36), .B(n40), .C(sine_lookup_width_minus_modulation_deviation_amount[2]), 
         .Z(n24525)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n36_bdd_3_lut.init = 16'hcaca;
    LUT4 i6567_4_lut (.A(modulation_output[14]), .B(modulation_output[15]), 
         .C(n9012), .D(n24823), .Z(carrier_center_increment_offset_rs_30__N_1560[14])) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam i6567_4_lut.init = 16'hccca;
    LUT4 i6565_4_lut (.A(n14_adj_3014), .B(modulation_output[15]), .C(n9010), 
         .D(n24823), .Z(carrier_center_increment_offset_rs_30__N_1560[13])) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam i6565_4_lut.init = 16'hccca;
    LUT4 i6507_2_lut (.A(sine_lookup_width_minus_modulation_deviation_amount[1]), 
         .B(sine_lookup_width_minus_modulation_deviation_amount[2]), .Z(n9010)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam i6507_2_lut.init = 16'heeee;
    LUT4 modulation_output_15__I_0_i43_3_lut (.A(n12), .B(n14_adj_3014), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[1]), .Z(n43)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam modulation_output_15__I_0_i43_3_lut.init = 16'hcaca;
    LUT4 i6559_3_lut (.A(n73), .B(modulation_output[15]), .C(n24823), 
         .Z(carrier_center_increment_offset_rs_30__N_1560[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam i6559_3_lut.init = 16'hcaca;
    LUT4 i6557_3_lut (.A(n72), .B(modulation_output[15]), .C(n24823), 
         .Z(carrier_center_increment_offset_rs_30__N_1560[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam i6557_3_lut.init = 16'hcaca;
    LUT4 i6555_3_lut (.A(n71), .B(modulation_output[15]), .C(n24823), 
         .Z(carrier_center_increment_offset_rs_30__N_1560[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam i6555_3_lut.init = 16'hcaca;
    LUT4 i6553_3_lut (.A(n70), .B(modulation_output[15]), .C(n24823), 
         .Z(carrier_center_increment_offset_rs_30__N_1560[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam i6553_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i70_3_lut (.A(n39_adj_3029), .B(n43), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[2]), .Z(n70)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam modulation_output_15__I_0_i70_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i39_3_lut (.A(n8), .B(n10), .C(sine_lookup_width_minus_modulation_deviation_amount[1]), 
         .Z(n39_adj_3029)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam modulation_output_15__I_0_i39_3_lut.init = 16'hcaca;
    LUT4 i11802_4_lut (.A(modulation_output[15]), .B(n178_adj_3009), .C(n24822), 
         .D(modulation_deviation_amount_minus_sine_lookup_width[4]), .Z(n64[30])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i11802_4_lut.init = 16'h3022;
    LUT4 modulation_output_15__I_0_332_i79_3_lut (.A(n48_adj_3033), .B(n52_adj_3046), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[2]), .Z(n79)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i79_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_332_i48_3_lut (.A(n17), .B(n19), .C(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .Z(n48_adj_3033)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i48_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_332_i52_3_lut (.A(n21), .B(n23), .C(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .Z(n52_adj_3046)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i52_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_332_i56_3_lut (.A(n25), .B(n27), .C(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .Z(n56_adj_3035)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i56_3_lut.init = 16'hcaca;
    LUT4 i11803_4_lut (.A(n95), .B(n178_adj_3009), .C(n24821), .D(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .Z(n64[29])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i11803_4_lut.init = 16'h3022;
    LUT4 i6474_4_lut (.A(modulation_output[15]), .B(modulation_output[14]), 
         .C(n24901), .D(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .Z(n95)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C (D)))) */ ;
    defparam i6474_4_lut.init = 16'hcaaa;
    LUT4 i11804_4_lut (.A(n96), .B(n178_adj_3009), .C(n24820), .D(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .Z(n64[28])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i11804_4_lut.init = 16'h3022;
    LUT4 i6476_4_lut (.A(modulation_output[15]), .B(n17), .C(n25015), 
         .D(modulation_deviation_amount_minus_sine_lookup_width[3]), .Z(n96)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C (D)))) */ ;
    defparam i6476_4_lut.init = 16'hcaaa;
    LUT4 i17720_3_lut (.A(\addr_space[0] [6]), .B(\addr_space[1] [6]), .C(\wb_addr[0] ), 
         .Z(n20050)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17720_3_lut.init = 16'hcaca;
    LUT4 i11805_4_lut (.A(n97), .B(n178_adj_3009), .C(n113), .D(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .Z(n64[27])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i11805_4_lut.init = 16'h3022;
    LUT4 modulation_output_15__I_0_332_i47_3_lut (.A(n16_adj_3047), .B(n18_adj_3042), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[1]), .Z(n47_adj_3032)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i47_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_332_i16_3_lut (.A(modulation_output[15]), 
         .B(modulation_output[14]), .C(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .Z(n16_adj_3047)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i16_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_332_i113_4_lut (.A(n82), .B(n59_adj_3031), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[3]), .D(modulation_deviation_amount_minus_sine_lookup_width[2]), 
         .Z(n113)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i113_4_lut.init = 16'h0aca;
    LUT4 modulation_output_15__I_0_332_i82_3_lut (.A(n51_adj_3048), .B(n55_adj_3034), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[2]), .Z(n82)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i82_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_332_i59_3_lut (.A(n28), .B(n30), .C(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .Z(n59_adj_3031)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i59_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_332_i51_3_lut (.A(n20_adj_3043), .B(n22_adj_3044), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[1]), .Z(n51_adj_3048)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i51_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_332_i55_3_lut (.A(n24_adj_3045), .B(n26), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[1]), .Z(n55_adj_3034)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i55_3_lut.init = 16'hcaca;
    LUT4 i11806_4_lut (.A(n98), .B(n178_adj_3009), .C(n114), .D(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .Z(n64[26])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i11806_4_lut.init = 16'h3022;
    LUT4 modulation_output_15__I_0_332_i114_4_lut (.A(n83), .B(n60_adj_3030), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[3]), .D(modulation_deviation_amount_minus_sine_lookup_width[2]), 
         .Z(n114)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i114_4_lut.init = 16'h0aca;
    LUT4 modulation_output_15__I_0_332_i83_3_lut (.A(n52_adj_3046), .B(n56_adj_3035), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[2]), .Z(n83)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i83_3_lut.init = 16'hcaca;
    LUT4 i11807_4_lut (.A(n99), .B(n178_adj_3009), .C(n115), .D(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .Z(n64[25])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i11807_4_lut.init = 16'h3022;
    LUT4 modulation_output_15__I_0_332_i99_3_lut (.A(modulation_output[15]), 
         .B(n76), .C(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .Z(n99)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i99_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_332_i76_3_lut (.A(n45_adj_3049), .B(n49_adj_3039), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[2]), .Z(n76)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i76_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_332_i115_4_lut (.A(n84), .B(n30), .C(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .D(n25009), .Z(n115)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i115_4_lut.init = 16'h0aca;
    LUT4 modulation_output_15__I_0_332_i84_3_lut (.A(n53_adj_3040), .B(n57_adj_3041), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[2]), .Z(n84)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i84_3_lut.init = 16'hcaca;
    LUT4 i11808_4_lut (.A(n100), .B(n178_adj_3009), .C(n24819), .D(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .Z(n64[24])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i11808_4_lut.init = 16'h3022;
    LUT4 modulation_output_15__I_0_332_i100_3_lut (.A(modulation_output[15]), 
         .B(n77), .C(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .Z(n100)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i100_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_332_i77_3_lut (.A(n46_adj_3050), .B(n50_adj_3036), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[2]), .Z(n77)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i77_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_332_i46_3_lut (.A(modulation_output[15]), 
         .B(n17), .C(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .Z(n46_adj_3050)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i46_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_332_i85_3_lut (.A(n54_adj_3037), .B(n58_adj_3038), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[2]), .Z(n85)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i85_3_lut.init = 16'hcaca;
    LUT4 i11809_2_lut (.A(n132), .B(n178_adj_3009), .Z(n64[23])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i11809_2_lut.init = 16'h2222;
    LUT4 i11810_2_lut (.A(n133), .B(n178_adj_3009), .Z(n64[22])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i11810_2_lut.init = 16'h2222;
    LUT4 i11811_2_lut (.A(n134), .B(n178_adj_3009), .Z(n64[21])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i11811_2_lut.init = 16'h2222;
    LUT4 i11812_2_lut (.A(n135), .B(n178_adj_3009), .Z(n64[20])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i11812_2_lut.init = 16'h2222;
    LUT4 i11813_2_lut (.A(n136), .B(n178_adj_3009), .Z(n64[19])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i11813_2_lut.init = 16'h2222;
    LUT4 i11814_2_lut (.A(n137), .B(n178_adj_3009), .Z(n64[18])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i11814_2_lut.init = 16'h2222;
    LUT4 i11815_4_lut (.A(n107), .B(n178_adj_3009), .C(n4), .D(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .Z(n64[17])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i11815_4_lut.init = 16'h3022;
    LUT4 modulation_output_15__I_0_332_i107_3_lut (.A(n76), .B(n84), .C(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .Z(n107)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i107_3_lut.init = 16'hcaca;
    LUT4 i11816_4_lut (.A(n108), .B(n178_adj_3009), .C(n24835), .D(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .Z(n64[16])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i11816_4_lut.init = 16'h3022;
    LUT4 modulation_output_15__I_0_332_i108_3_lut (.A(n77), .B(n85), .C(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .Z(n108)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i108_3_lut.init = 16'hcaca;
    LUT4 i11526_4_lut (.A(n78), .B(n24834), .C(n24846), .D(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .Z(n64[15])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i11526_4_lut.init = 16'h3022;
    LUT4 modulation_output_15__I_0_332_i78_3_lut (.A(n47_adj_3032), .B(n51_adj_3048), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[2]), .Z(n78)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i78_3_lut.init = 16'hcaca;
    LUT4 i6561_3_lut_4_lut (.A(sine_lookup_width_minus_modulation_deviation_amount[2]), 
         .B(n24823), .C(modulation_output[15]), .D(n43), .Z(carrier_center_increment_offset_rs_30__N_1560[11])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam i6561_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i17718_3_lut (.A(\addr_space[2] [7]), .B(\addr_space[3] [7]), .C(\wb_addr[0] ), 
         .Z(n20048)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17718_3_lut.init = 16'hcaca;
    LUT4 i17717_3_lut (.A(\addr_space[0] [7]), .B(\addr_space[1] [7]), .C(\wb_addr[0] ), 
         .Z(n20047)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17717_3_lut.init = 16'hcaca;
    LUT4 n36_bdd_3_lut_22820 (.A(n44), .B(modulation_output[15]), .C(sine_lookup_width_minus_modulation_deviation_amount[2]), 
         .Z(n24524)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n36_bdd_3_lut_22820.init = 16'hcaca;
    LUT4 i8579_2_lut_rep_274 (.A(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .B(n178_adj_3009), .Z(n24834)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i8579_2_lut_rep_274.init = 16'heeee;
    PFUMX i17650 (.BLUT(n19978), .ALUT(n19979), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[29]));
    PFUMX i17653 (.BLUT(n19981), .ALUT(n19982), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[28]));
    PFUMX i17656 (.BLUT(n19984), .ALUT(n19985), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[27]));
    PFUMX i17659 (.BLUT(n19987), .ALUT(n19988), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[26]));
    LUT4 n22768_bdd_3_lut_4_lut (.A(sine_lookup_width_minus_modulation_deviation_amount[4]), 
         .B(n178), .C(modulation_output[15]), .D(n22768), .Z(carrier_center_increment_offset_rs_30__N_1560[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam n22768_bdd_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i17662 (.BLUT(n19990), .ALUT(n19991), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[25]));
    LUT4 n24518_bdd_3_lut_4_lut (.A(sine_lookup_width_minus_modulation_deviation_amount[4]), 
         .B(n178), .C(modulation_output[15]), .D(n24518), .Z(carrier_center_increment_offset_rs_30__N_1560[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam n24518_bdd_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i19234 (.BLUT(n21562), .ALUT(n21563), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[0]));
    LUT4 n22772_bdd_3_lut_4_lut (.A(sine_lookup_width_minus_modulation_deviation_amount[4]), 
         .B(n178), .C(modulation_output[15]), .D(n22772), .Z(carrier_center_increment_offset_rs_30__N_1560[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam n22772_bdd_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i19237 (.BLUT(n21565), .ALUT(n21566), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[31]));
    LUT4 i11515_2_lut_3_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .B(n178_adj_3009), .C(n89), .D(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .Z(n64[4])) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i11515_2_lut_3_lut_4_lut.init = 16'h0010;
    PFUMX i17668 (.BLUT(n19996), .ALUT(n19997), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[24]));
    LUT4 i11518_2_lut_3_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .B(n178_adj_3009), .C(n24846), .D(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .Z(n64[7])) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i11518_2_lut_3_lut_4_lut.init = 16'h0010;
    PFUMX i17671 (.BLUT(n19999), .ALUT(n20000), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[23]));
    PFUMX i17674 (.BLUT(n20002), .ALUT(n20003), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[22]));
    LUT4 i11516_2_lut_3_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .B(n178_adj_3009), .C(n88), .D(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .Z(n64[5])) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i11516_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 i11517_2_lut_3_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .B(n178_adj_3009), .C(n24850), .D(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .Z(n64[6])) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i11517_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 i11522_2_lut_3_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .B(n178_adj_3009), .C(n113), .Z(n64[11])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i11522_2_lut_3_lut.init = 16'h1010;
    PFUMX i19246 (.BLUT(n21574), .ALUT(n21575), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[30]));
    PFUMX i17677 (.BLUT(n20005), .ALUT(n20006), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[21]));
    PFUMX i17680 (.BLUT(n20008), .ALUT(n20009), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[20]));
    LUT4 n37_bdd_3_lut (.A(n37), .B(n41), .C(sine_lookup_width_minus_modulation_deviation_amount[2]), 
         .Z(n24538)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n37_bdd_3_lut.init = 16'hcaca;
    LUT4 n37_bdd_4_lut (.A(n14_adj_3014), .B(modulation_output[15]), .C(sine_lookup_width_minus_modulation_deviation_amount[2]), 
         .D(sine_lookup_width_minus_modulation_deviation_amount[1]), .Z(n24537)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;
    defparam n37_bdd_4_lut.init = 16'hccca;
    PFUMX i17683 (.BLUT(n20011), .ALUT(n20012), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[19]));
    PFUMX i17686 (.BLUT(n20014), .ALUT(n20015), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[18]));
    LUT4 n38_bdd_3_lut_23804 (.A(n38), .B(n42), .C(sine_lookup_width_minus_modulation_deviation_amount[2]), 
         .Z(n24548)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n38_bdd_3_lut_23804.init = 16'hcaca;
    LUT4 n38_bdd_4_lut (.A(modulation_output[14]), .B(modulation_output[15]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[2]), .D(n25133), 
         .Z(n24547)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;
    defparam n38_bdd_4_lut.init = 16'hccca;
    LUT4 i11521_2_lut_3_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .B(n178_adj_3009), .C(n114), .Z(n64[10])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i11521_2_lut_3_lut.init = 16'h1010;
    LUT4 i11520_2_lut_3_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .B(n178_adj_3009), .C(n115), .Z(n64[9])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i11520_2_lut_3_lut.init = 16'h1010;
    LUT4 i2_2_lut_3_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .B(n178_adj_3009), .C(n4), .Z(n17801)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i2_2_lut_3_lut.init = 16'h1010;
    LUT4 i17715_3_lut (.A(\addr_space[2] [8]), .B(\addr_space[3] [8]), .C(\wb_addr[0] ), 
         .Z(n20045)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17715_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .B(n24888), .C(n178_adj_3009), .D(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .Z(n64[0])) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0004;
    LUT4 i17714_3_lut (.A(\addr_space[0] [8]), .B(\addr_space[1] [8]), .C(\wb_addr[0] ), 
         .Z(n20044)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17714_3_lut.init = 16'hcaca;
    LUT4 i17712_3_lut (.A(\addr_space[2] [9]), .B(\addr_space[3] [9]), .C(\wb_addr[0] ), 
         .Z(n20042)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17712_3_lut.init = 16'hcaca;
    PFUMX i17725 (.BLUT(n20053), .ALUT(n20054), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[5]));
    LUT4 i17711_3_lut (.A(\addr_space[0] [9]), .B(\addr_space[1] [9]), .C(\wb_addr[0] ), 
         .Z(n20041)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17711_3_lut.init = 16'hcaca;
    LUT4 i17709_3_lut (.A(\addr_space[2] [10]), .B(\addr_space[3] [10]), 
         .C(\wb_addr[0] ), .Z(n20039)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17709_3_lut.init = 16'hcaca;
    LUT4 i17708_3_lut (.A(\addr_space[0] [10]), .B(\addr_space[1] [10]), 
         .C(\wb_addr[0] ), .Z(n20038)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17708_3_lut.init = 16'hcaca;
    LUT4 i17688_3_lut (.A(\addr_space[2] [17]), .B(\addr_space[3] [17]), 
         .C(\wb_addr[0] ), .Z(n20018)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17688_3_lut.init = 16'hcaca;
    LUT4 i17706_3_lut (.A(\addr_space[2] [11]), .B(\addr_space[3] [11]), 
         .C(\wb_addr[0] ), .Z(n20036)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17706_3_lut.init = 16'hcaca;
    LUT4 i10825_3_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .B(n25187), .C(modulation_deviation_amount_minus_sine_lookup_width[2]), 
         .D(n58_adj_3038), .Z(n89)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i10825_3_lut_4_lut.init = 16'h4f40;
    LUT4 i1_2_lut_rep_275_3_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .B(n25187), .C(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .D(modulation_deviation_amount_minus_sine_lookup_width[2]), .Z(n24835)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i1_2_lut_rep_275_3_lut_4_lut.init = 16'h0004;
    PFUMX modulation_output_15__I_0_332_i137 (.BLUT(n75), .ALUT(n106), .C0(n19807), 
          .Z(n137)) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;
    PFUMX modulation_output_15__I_0_332_i136 (.BLUT(n74), .ALUT(n105), .C0(n19807), 
          .Z(n136)) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;
    PFUMX modulation_output_15__I_0_332_i133 (.BLUT(n102), .ALUT(n118), 
          .C0(modulation_deviation_amount_minus_sine_lookup_width[4]), .Z(n133)) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;
    PFUMX modulation_output_15__I_0_332_i132 (.BLUT(n101), .ALUT(n117), 
          .C0(modulation_deviation_amount_minus_sine_lookup_width[4]), .Z(n132)) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=123, LSE_RLINE=134 */ ;
    LUT4 i17705_3_lut (.A(\addr_space[0] [11]), .B(\addr_space[1] [11]), 
         .C(\wb_addr[0] ), .Z(n20035)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17705_3_lut.init = 16'hcaca;
    LUT4 i6505_2_lut_rep_573 (.A(sine_lookup_width_minus_modulation_deviation_amount[0]), 
         .B(sine_lookup_width_minus_modulation_deviation_amount[1]), .Z(n25133)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam i6505_2_lut_rep_573.init = 16'heeee;
    LUT4 i6506_3_lut_4_lut (.A(sine_lookup_width_minus_modulation_deviation_amount[0]), 
         .B(sine_lookup_width_minus_modulation_deviation_amount[1]), .C(modulation_output[15]), 
         .D(modulation_output[14]), .Z(n46)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam i6506_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i6509_2_lut_3_lut (.A(sine_lookup_width_minus_modulation_deviation_amount[0]), 
         .B(sine_lookup_width_minus_modulation_deviation_amount[1]), .C(sine_lookup_width_minus_modulation_deviation_amount[2]), 
         .Z(n9012)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam i6509_2_lut_3_lut.init = 16'hfefe;
    LUT4 i17703_3_lut (.A(\addr_space[2] [12]), .B(\addr_space[3] [12]), 
         .C(\wb_addr[0] ), .Z(n20033)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17703_3_lut.init = 16'hcaca;
    LUT4 i17702_3_lut (.A(\addr_space[0] [12]), .B(\addr_space[1] [12]), 
         .C(\wb_addr[0] ), .Z(n20032)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17702_3_lut.init = 16'hcaca;
    LUT4 i17700_3_lut (.A(\addr_space[2] [13]), .B(\addr_space[3] [13]), 
         .C(\wb_addr[0] ), .Z(n20030)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17700_3_lut.init = 16'hcaca;
    PFUMX i21285 (.BLUT(n22770), .ALUT(n38), .C0(sine_lookup_width_minus_modulation_deviation_amount[2]), 
          .Z(n22771));
    LUT4 i17699_3_lut (.A(\addr_space[0] [13]), .B(\addr_space[1] [13]), 
         .C(\wb_addr[0] ), .Z(n20029)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17699_3_lut.init = 16'hcaca;
    LUT4 i17697_3_lut (.A(\addr_space[2] [14]), .B(\addr_space[3] [14]), 
         .C(\wb_addr[0] ), .Z(n20027)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17697_3_lut.init = 16'hcaca;
    LUT4 i17696_3_lut (.A(\addr_space[0] [14]), .B(\addr_space[1] [14]), 
         .C(\wb_addr[0] ), .Z(n20026)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17696_3_lut.init = 16'hcaca;
    LUT4 i17694_3_lut (.A(\addr_space[2] [15]), .B(\addr_space[3] [15]), 
         .C(\wb_addr[0] ), .Z(n20024)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17694_3_lut.init = 16'hcaca;
    PFUMX i21283 (.BLUT(n22767), .ALUT(n72), .C0(sine_lookup_width_minus_modulation_deviation_amount[3]), 
          .Z(n22768));
    LUT4 i17693_3_lut (.A(\addr_space[0] [15]), .B(\addr_space[1] [15]), 
         .C(\wb_addr[0] ), .Z(n20023)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17693_3_lut.init = 16'hcaca;
    LUT4 i17691_3_lut (.A(\addr_space[2] [16]), .B(\addr_space[3] [16]), 
         .C(\wb_addr[0] ), .Z(n20021)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17691_3_lut.init = 16'hcaca;
    PFUMX i17728 (.BLUT(n20056), .ALUT(n20057), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[4]));
    PFUMX i21281 (.BLUT(n22765), .ALUT(n13476), .C0(sine_lookup_width_minus_modulation_deviation_amount[1]), 
          .Z(n22766));
    LUT4 smpl_register_5__bdd_4_lut_4_lut (.A(\wb_addr[0] ), .B(\wb_addr[1] ), 
         .C(n2), .D(\smpl_register[5] ), .Z(n24788)) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(34[4:25])
    defparam smpl_register_5__bdd_4_lut_4_lut.init = 16'hf3d1;
    LUT4 smpl_register_29__bdd_4_lut_4_lut (.A(\wb_addr[0] ), .B(\wb_addr[1] ), 
         .C(n2_adj_1), .D(\smpl_register[29] ), .Z(n24795)) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(34[4:25])
    defparam smpl_register_29__bdd_4_lut_4_lut.init = 16'hf3d1;
    LUT4 smpl_register_20__bdd_4_lut_4_lut (.A(\wb_addr[0] ), .B(\wb_addr[1] ), 
         .C(n2_adj_2), .D(\smpl_register[20] ), .Z(n24794)) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(34[4:25])
    defparam smpl_register_20__bdd_4_lut_4_lut.init = 16'hf3d1;
    LUT4 smpl_register_18__bdd_4_lut_4_lut (.A(\wb_addr[0] ), .B(\wb_addr[1] ), 
         .C(n2_adj_3), .D(\smpl_register[18] ), .Z(n24793)) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(34[4:25])
    defparam smpl_register_18__bdd_4_lut_4_lut.init = 16'hf3d1;
    LUT4 smpl_register_17__bdd_4_lut_4_lut (.A(\wb_addr[0] ), .B(\wb_addr[1] ), 
         .C(n2_adj_4), .D(\smpl_register[17] ), .Z(n24792)) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(34[4:25])
    defparam smpl_register_17__bdd_4_lut_4_lut.init = 16'hf3d1;
    LUT4 i17687_3_lut (.A(\addr_space[0] [17]), .B(\addr_space[1] [17]), 
         .C(\wb_addr[0] ), .Z(n20017)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17687_3_lut.init = 16'hcaca;
    LUT4 smpl_register_16__bdd_4_lut_4_lut (.A(\wb_addr[0] ), .B(\wb_addr[1] ), 
         .C(n2_adj_5), .D(\smpl_register[16] ), .Z(n24791)) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(34[4:25])
    defparam smpl_register_16__bdd_4_lut_4_lut.init = 16'hf3d1;
    LUT4 smpl_register_10__bdd_4_lut_4_lut (.A(\wb_addr[0] ), .B(\wb_addr[1] ), 
         .C(n2_adj_6), .D(\smpl_register[10] ), .Z(n24790)) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(34[4:25])
    defparam smpl_register_10__bdd_4_lut_4_lut.init = 16'hf3d1;
    LUT4 smpl_register_9__bdd_4_lut_4_lut (.A(\wb_addr[0] ), .B(\wb_addr[1] ), 
         .C(n2_adj_7), .D(\smpl_register[9] ), .Z(n24789)) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(34[4:25])
    defparam smpl_register_9__bdd_4_lut_4_lut.init = 16'hf3d1;
    LUT4 i21171_2_lut_rep_448 (.A(modulation_deviation_amount_minus_sine_lookup_width[2]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[3]), .Z(n25008)) /* synthesis lut_function=(!(A+(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam i21171_2_lut_rep_448.init = 16'h1111;
    LUT4 i6469_2_lut_rep_449 (.A(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[2]), .Z(n25009)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam i6469_2_lut_rep_449.init = 16'heeee;
    LUT4 i1_3_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[2]), .C(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .D(n30), .Z(n4)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam i1_3_lut_4_lut.init = 16'h0100;
    LUT4 i6478_3_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[2]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[3]), .C(n47_adj_3032), 
         .D(modulation_output[15]), .Z(n97)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam i6478_3_lut_4_lut.init = 16'hf780;
    LUT4 i6480_3_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[2]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[3]), .C(n48_adj_3033), 
         .D(modulation_output[15]), .Z(n98)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam i6480_3_lut_4_lut.init = 16'hf780;
    LUT4 i6461_2_lut_rep_452 (.A(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[1]), .Z(n25012)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam i6461_2_lut_rep_452.init = 16'h8888;
    LUT4 i6465_2_lut_rep_341_3_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[1]), .C(modulation_deviation_amount_minus_sine_lookup_width[2]), 
         .Z(n24901)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam i6465_2_lut_rep_341_3_lut.init = 16'h8080;
    LUT4 i6462_3_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[1]), .C(modulation_output[14]), 
         .D(modulation_output[15]), .Z(n45_adj_3049)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam i6462_3_lut_4_lut.init = 16'hf780;
    LUT4 i17690_3_lut (.A(\addr_space[0] [16]), .B(\addr_space[1] [16]), 
         .C(\wb_addr[0] ), .Z(n20020)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17690_3_lut.init = 16'hcaca;
    LUT4 i10950_2_lut_4_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[2]), .C(n59_adj_3031), 
         .D(n55_adj_3034), .Z(n117)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i10950_2_lut_4_lut_4_lut.init = 16'h5140;
    LUT4 modulation_output_15__I_0_332_i104_4_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[4]), .C(n89), 
         .D(n81), .Z(n104)) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C)+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam modulation_output_15__I_0_332_i104_4_lut_4_lut.init = 16'h7340;
    LUT4 i10951_2_lut_4_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[2]), .C(n60_adj_3030), 
         .D(n56_adj_3035), .Z(n118)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i10951_2_lut_4_lut_4_lut.init = 16'h5140;
    LUT4 modulation_output_15__I_0_332_i103_4_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[4]), .C(n88), 
         .D(n80), .Z(n103)) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C)+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam modulation_output_15__I_0_332_i103_4_lut_4_lut.init = 16'h7340;
    LUT4 i6467_2_lut_rep_455 (.A(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[2]), .Z(n25015)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam i6467_2_lut_rep_455.init = 16'h8888;
    LUT4 i6468_3_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[2]), .C(n17), 
         .D(modulation_output[15]), .Z(n73_adj_3015)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam i6468_3_lut_4_lut.init = 16'hf780;
    PFUMX i21279 (.BLUT(n22762), .ALUT(n71), .C0(sine_lookup_width_minus_modulation_deviation_amount[3]), 
          .Z(n22763));
    PFUMX i17731 (.BLUT(n20059), .ALUT(n20060), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[3]));
    PFUMX i17734 (.BLUT(n20062), .ALUT(n20063), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[2]));
    PFUMX i17737 (.BLUT(n20065), .ALUT(n20066), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[1]));
    PFUMX i21277 (.BLUT(n22760), .ALUT(n13468), .C0(sine_lookup_width_minus_modulation_deviation_amount[1]), 
          .Z(n22761));
    PFUMX i17689 (.BLUT(n20017), .ALUT(n20018), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[17]));
    dds modulation (.i_ref_clk_c(i_ref_clk_c), .i_resetb_N_301(i_resetb_N_301), 
        .\addr_space[1][0] (\addr_space[1] [0]), .\addr_space[1][30] (\addr_space[1] [30]), 
        .\addr_space[1][29] (\addr_space[1] [29]), .\addr_space[1][28] (\addr_space[1] [28]), 
        .\addr_space[1][27] (\addr_space[1] [27]), .\addr_space[1][26] (\addr_space[1] [26]), 
        .\addr_space[1][25] (\addr_space[1] [25]), .\addr_space[1][24] (\addr_space[1] [24]), 
        .\addr_space[1][23] (\addr_space[1] [23]), .\addr_space[1][22] (\addr_space[1] [22]), 
        .\addr_space[1][21] (\addr_space[1] [21]), .\addr_space[1][20] (\addr_space[1] [20]), 
        .\addr_space[1][19] (\addr_space[1] [19]), .\addr_space[1][18] (\addr_space[1] [18]), 
        .\addr_space[1][17] (\addr_space[1] [17]), .\addr_space[1][16] (\addr_space[1] [16]), 
        .\addr_space[1][15] (\addr_space[1] [15]), .\addr_space[1][14] (\addr_space[1] [14]), 
        .\addr_space[1][13] (\addr_space[1] [13]), .\addr_space[1][12] (\addr_space[1] [12]), 
        .\addr_space[1][11] (\addr_space[1] [11]), .\addr_space[1][10] (\addr_space[1] [10]), 
        .\addr_space[1][9] (\addr_space[1] [9]), .\addr_space[1][8] (\addr_space[1] [8]), 
        .\addr_space[1][7] (\addr_space[1] [7]), .\addr_space[1][6] (\addr_space[1] [6]), 
        .\addr_space[1][5] (\addr_space[1] [5]), .\addr_space[1][4] (\addr_space[1] [4]), 
        .\addr_space[1][3] (\addr_space[1] [3]), .\addr_space[1][2] (\addr_space[1] [2]), 
        .\addr_space[1][1] (\addr_space[1] [1]), .modulation_output({modulation_output}), 
        .i_resetb_c(i_resetb_c), .GND_net(GND_net), .\quarter_wave_sample_register_q[15] (quarter_wave_sample_register_q[15])) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(72[4:161])
    dds_U2 carrier (.i_ref_clk_c(i_ref_clk_c), .i_resetb_N_301(i_resetb_N_301), 
           .carrier_increment({carrier_increment}), .o_baseband_i_c_15(o_baseband_i_c_15), 
           .o_baseband_i_c_14(o_baseband_i_c_14), .o_baseband_i_c_13(o_baseband_i_c_13), 
           .o_baseband_i_c_12(o_baseband_i_c_12), .o_baseband_i_c_11(o_baseband_i_c_11), 
           .o_baseband_i_c_10(o_baseband_i_c_10), .n3607(n3607), .i_resetb_c(i_resetb_c), 
           .o_baseband_q_c_7(o_baseband_q_c_7), .o_baseband_i_c_7(o_baseband_i_c_7), 
           .o_baseband_i_c_8(o_baseband_i_c_8), .\quarter_wave_sample_register_q[15] (quarter_wave_sample_register_q[15]), 
           .n27529(n27529), .o_baseband_q_c_15(o_baseband_q_c_15), .o_baseband_q_c_14(o_baseband_q_c_14), 
           .o_baseband_q_c_13(o_baseband_q_c_13), .o_baseband_q_c_12(o_baseband_q_c_12), 
           .o_baseband_q_c_11(o_baseband_q_c_11), .o_baseband_q_c_10(o_baseband_q_c_10), 
           .n3608(n3608), .o_baseband_q_c_8(o_baseband_q_c_8), .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(67[4:158])
    
endmodule
//
// Verilog Description of module dds
//

module dds (i_ref_clk_c, i_resetb_N_301, \addr_space[1][0] , \addr_space[1][30] , 
            \addr_space[1][29] , \addr_space[1][28] , \addr_space[1][27] , 
            \addr_space[1][26] , \addr_space[1][25] , \addr_space[1][24] , 
            \addr_space[1][23] , \addr_space[1][22] , \addr_space[1][21] , 
            \addr_space[1][20] , \addr_space[1][19] , \addr_space[1][18] , 
            \addr_space[1][17] , \addr_space[1][16] , \addr_space[1][15] , 
            \addr_space[1][14] , \addr_space[1][13] , \addr_space[1][12] , 
            \addr_space[1][11] , \addr_space[1][10] , \addr_space[1][9] , 
            \addr_space[1][8] , \addr_space[1][7] , \addr_space[1][6] , 
            \addr_space[1][5] , \addr_space[1][4] , \addr_space[1][3] , 
            \addr_space[1][2] , \addr_space[1][1] , modulation_output, 
            i_resetb_c, GND_net, \quarter_wave_sample_register_q[15] ) /* synthesis syn_module_defined=1 */ ;
    input i_ref_clk_c;
    input i_resetb_N_301;
    input \addr_space[1][0] ;
    input \addr_space[1][30] ;
    input \addr_space[1][29] ;
    input \addr_space[1][28] ;
    input \addr_space[1][27] ;
    input \addr_space[1][26] ;
    input \addr_space[1][25] ;
    input \addr_space[1][24] ;
    input \addr_space[1][23] ;
    input \addr_space[1][22] ;
    input \addr_space[1][21] ;
    input \addr_space[1][20] ;
    input \addr_space[1][19] ;
    input \addr_space[1][18] ;
    input \addr_space[1][17] ;
    input \addr_space[1][16] ;
    input \addr_space[1][15] ;
    input \addr_space[1][14] ;
    input \addr_space[1][13] ;
    input \addr_space[1][12] ;
    input \addr_space[1][11] ;
    input \addr_space[1][10] ;
    input \addr_space[1][9] ;
    input \addr_space[1][8] ;
    input \addr_space[1][7] ;
    input \addr_space[1][6] ;
    input \addr_space[1][5] ;
    input \addr_space[1][4] ;
    input \addr_space[1][3] ;
    input \addr_space[1][2] ;
    input \addr_space[1][1] ;
    output [15:0]modulation_output;
    input i_resetb_c;
    input GND_net;
    input \quarter_wave_sample_register_q[15] ;
    
    wire i_ref_clk_c /* synthesis SET_AS_NETWORK=i_ref_clk_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(22[12:21])
    wire [15:0]modulation_output_c /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(62[39:56])
    wire [30:0]increment;   // d:/documents/git_local/fm_modulator/rtl/dds.v(14[31:40])
    wire [11:0]o_phase;   // d:/documents/git_local/fm_modulator/rtl/dds.v(18[26:33])
    
    FD1S3DX increment_i0 (.D(\addr_space[1][0] ), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(increment[0])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i0.GSR = "DISABLED";
    FD1S3DX increment_i30 (.D(\addr_space[1][30] ), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(increment[30])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i30.GSR = "DISABLED";
    FD1S3DX increment_i29 (.D(\addr_space[1][29] ), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(increment[29])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i29.GSR = "DISABLED";
    FD1S3DX increment_i28 (.D(\addr_space[1][28] ), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(increment[28])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i28.GSR = "DISABLED";
    FD1S3DX increment_i27 (.D(\addr_space[1][27] ), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(increment[27])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i27.GSR = "DISABLED";
    FD1S3DX increment_i26 (.D(\addr_space[1][26] ), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(increment[26])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i26.GSR = "DISABLED";
    FD1S3DX increment_i25 (.D(\addr_space[1][25] ), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(increment[25])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i25.GSR = "DISABLED";
    FD1S3DX increment_i24 (.D(\addr_space[1][24] ), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(increment[24])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i24.GSR = "DISABLED";
    FD1S3DX increment_i23 (.D(\addr_space[1][23] ), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(increment[23])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i23.GSR = "DISABLED";
    FD1S3DX increment_i22 (.D(\addr_space[1][22] ), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(increment[22])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i22.GSR = "DISABLED";
    FD1S3DX increment_i21 (.D(\addr_space[1][21] ), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(increment[21])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i21.GSR = "DISABLED";
    FD1S3DX increment_i20 (.D(\addr_space[1][20] ), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(increment[20])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i20.GSR = "DISABLED";
    FD1S3DX increment_i19 (.D(\addr_space[1][19] ), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(increment[19])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i19.GSR = "DISABLED";
    FD1S3DX increment_i18 (.D(\addr_space[1][18] ), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(increment[18])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i18.GSR = "DISABLED";
    FD1S3DX increment_i17 (.D(\addr_space[1][17] ), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(increment[17])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i17.GSR = "DISABLED";
    FD1S3DX increment_i16 (.D(\addr_space[1][16] ), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(increment[16])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i16.GSR = "DISABLED";
    FD1S3DX increment_i15 (.D(\addr_space[1][15] ), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(increment[15])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i15.GSR = "DISABLED";
    FD1S3DX increment_i14 (.D(\addr_space[1][14] ), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(increment[14])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i14.GSR = "DISABLED";
    FD1S3DX increment_i13 (.D(\addr_space[1][13] ), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(increment[13])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i13.GSR = "DISABLED";
    FD1S3DX increment_i12 (.D(\addr_space[1][12] ), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(increment[12])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i12.GSR = "DISABLED";
    FD1S3DX increment_i11 (.D(\addr_space[1][11] ), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(increment[11])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i11.GSR = "DISABLED";
    FD1S3DX increment_i10 (.D(\addr_space[1][10] ), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(increment[10])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i10.GSR = "DISABLED";
    FD1S3DX increment_i9 (.D(\addr_space[1][9] ), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(increment[9])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i9.GSR = "DISABLED";
    FD1S3DX increment_i8 (.D(\addr_space[1][8] ), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(increment[8])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i8.GSR = "DISABLED";
    FD1S3DX increment_i7 (.D(\addr_space[1][7] ), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(increment[7])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i7.GSR = "DISABLED";
    FD1S3DX increment_i6 (.D(\addr_space[1][6] ), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(increment[6])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i6.GSR = "DISABLED";
    FD1S3DX increment_i5 (.D(\addr_space[1][5] ), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(increment[5])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i5.GSR = "DISABLED";
    FD1S3DX increment_i4 (.D(\addr_space[1][4] ), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(increment[4])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i4.GSR = "DISABLED";
    FD1S3DX increment_i3 (.D(\addr_space[1][3] ), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(increment[3])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i3.GSR = "DISABLED";
    FD1S3DX increment_i2 (.D(\addr_space[1][2] ), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(increment[2])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i2.GSR = "DISABLED";
    FD1S3DX increment_i1 (.D(\addr_space[1][1] ), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(increment[1])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i1.GSR = "DISABLED";
    quarter_wave_sine_lookup qtr_inst (.i_ref_clk_c(i_ref_clk_c), .i_resetb_N_301(i_resetb_N_301), 
            .modulation_output({modulation_output}), .i_resetb_c(i_resetb_c), 
            .o_phase({o_phase}), .GND_net(GND_net), .\quarter_wave_sample_register_q[15] (\quarter_wave_sample_register_q[15] )) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(21[70:134])
    \nco(OW=12)  nco_inst (.i_ref_clk_c(i_ref_clk_c), .i_resetb_N_301(i_resetb_N_301), 
            .increment({increment}), .o_phase({o_phase}), .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(20[49:100])
    
endmodule
//
// Verilog Description of module quarter_wave_sine_lookup
//

module quarter_wave_sine_lookup (i_ref_clk_c, i_resetb_N_301, modulation_output, 
            i_resetb_c, o_phase, GND_net, \quarter_wave_sample_register_q[15] ) /* synthesis syn_module_defined=1 */ ;
    input i_ref_clk_c;
    input i_resetb_N_301;
    output [15:0]modulation_output;
    input i_resetb_c;
    input [11:0]o_phase;
    input GND_net;
    input \quarter_wave_sample_register_q[15] ;
    
    wire i_ref_clk_c /* synthesis SET_AS_NETWORK=i_ref_clk_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(22[12:21])
    wire [15:0]\o_val_pipeline_i[0]  /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(15[24:40])
    wire [15:0]modulation_output_c /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(62[39:56])
    
    wire n20077, n20078;
    wire [9:0]index_i;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(31[17:24])
    
    wire n20079;
    wire [15:0]quarter_wave_sample_register_i;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(22[24:54])
    wire [14:0]quarter_wave_sample_register_i_15__N_2126;
    
    wire n21669, n21656, n20092;
    wire [15:0]n1205;
    
    wire n21713, n21714, n21715, n20080, n20081, n20082, n20083, 
        n20084, n20085, n21707, n21708, n21709, n25098, n24995, 
        n27516, n653, n557, n572, n21717, n25107, n684, n589, 
        n604, n21718, n30, n620, n635, n21719, n20800, n404, 
        n25139, n653_adj_2797, n668, n21720, n24892, n93, n20765;
    wire [11:0]phase_i;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(11[17:24])
    wire [1:0]phase_negation_i;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(23[12:28])
    wire [9:0]index_i_9__N_2106;
    
    wire n684_adj_2798, n699, n21721, n716, n731, n21722, n21603, 
        n21604, n21609, n21620, n21621, n21628, n21624, n21625, 
        n21630, n21626, n21627, n21631, n747, n762, n21723, n382, 
        n509, n20580, n781, n796, n21724, n812, n11935, n21725, 
        n875, n890, n21727, n22968, n908, n923, n21728, n25144, 
        n325, n939, n954, n21729, n21654, n21655, n23000, n971, 
        n986, n21730, n24994, n491, n23116, n20591, n20592, n20593, 
        n20594, n20595, n20596, n24996, n19936, n1002, n1017, 
        n21731, n526, n541, n21716, n21667, n21668, n20613, n20614, 
        n20624, n20615, n20616, n20625, n20621, n20622, n20628, 
        n21750, n21751, n21752, n21753, n21754, n21755, n20133, 
        n20134, n20141, n17363;
    wire [15:0]o_val_pipeline_i_0__15__N_2157;
    
    wire n17364, n20135, n20136, n20142, n20195, n20196, n20203, 
        n20197, n20198, n20204, n24925, n317, n25101, n443, n20201, 
        n20202, n20206, n20228, n20229, n20235, n20230, n20231, 
        n20236, n20232, n20233, n20237, n859, n860, n25126, n25149, 
        n21787, n21788, n21789, n21790, n21791, n21792, n21591, 
        n21592, n21796, n21797, n21798, n21593, n21594, n21595, 
        n21596, n21605, n221, n252, n20120, n11940, n20744, n20757, 
        n20760, n21623, n574, n20763, n20766, n764, n27500, n27505, 
        n21650, n21651, n21652, n21653, n701, n764_adj_2799, n21663, 
        n21664, n21665, n21666, n732, n763, n24868, n21616, n891, 
        n20603, n20604, n20619, n20607, n20608, n20609, n20610, 
        n20748, n20749, n20752, n20617, n20618, n20626, n20750, 
        n20751, n20753, n316, n20653, n316_adj_2800, n412, n924, 
        n20773, n20780, n20102, n21732, n21733, n21740, n158, 
        n189, n20150, n21734, n21735, n21741, n21736, n21737, 
        n21742, n21738, n21739, n21743, n20793, n20796, n20105, 
        n20656, n20657, n382_adj_2801, n20799, n20802, n20106, n20805, 
        n20808, n20107, n20663, n20664, n509_adj_2802, n20738, n20741, 
        n20767, n20768, n20771, n20769, n20770, n20772, n20774, 
        n20775, n20778, n20776, n20777, n20779, n20781, n20782, 
        n20785, n20783, n20784, n20786, n20117, n20118, n20119, 
        n20121, n20122, n20123, n20124, n20125, n20126, n20137, 
        n20129, n20130, n20139, n20148, n20149, n20164, n20151, 
        n20165, n20152, n20153, n20166, n20156, n20157, n20168, 
        n20158, n20159, n20169, n20160, n20161, n20170, n20162, 
        n20163, n20171, n25151, n17552, n21571, n21572, n21573, 
        n17551, n20179, n20180, n20181, n20182, n20183, n20184, 
        n20185, n20186, n20187, n20188, n20199, n20191, n20192, 
        n20193, n20194, n25269, n20212, n20213, n20227, n20214, 
        n20215, n20216, n20217, n20218, n20219, n20220, n20221, 
        n428, n762_adj_2803, n844, n27515, n11976, n890_adj_2804, 
        n11938, n21800, n781_adj_2805, n21039, n21040, n21047, n25138, 
        n21045, n21046, n21050, n17554, n23026, n25110, n25108, 
        n20072, n19916, n635_adj_2806, n30_adj_2807, n506, n46, 
        n19958, n716_adj_2808, n348, n349, n23752, n23749, n781_adj_2809, 
        n747_adj_2810, n23711, n25299, n25300, n62, n491_adj_2811, 
        n443_adj_2812, n251, n20071, n20073, n24844, n251_adj_2813, 
        n21049, n21052, n21614, n21335, n109, n460, n301, n908_adj_2814, 
        n317_adj_2815, n21048, n21051, n25120, n27508, n21748, n699_adj_2816, 
        n412_adj_2817, n684_adj_2818, n24978, n445, n716_adj_2819, 
        n21747, n21749, n20068, n20069, n20070, n19957, n379, 
        n443_adj_2820, n24952, n22865, n25092, n254, n24891, n14964, 
        n252_adj_2821, n24960, n62_adj_2822, n860_adj_2823, n364, 
        n20655, n24810, n25137, n23674, n24843, n24831, n189_adj_2824, 
        n24951, n127, n27502, n23677, n125, n25152, n23693, n27504, 
        n23694, n25143, n23697, n21642, n332, n21641, n20175, 
        n25153, n23705, n25099, n25150, n23714, n25275, n25276, 
        n25277, n25131, n21635, n21636, n21637, n1001, n588, n21617, 
        n22970, n22971, n21618, n21619, n252_adj_2825, n23816, n24800, 
        n413, n574_adj_2826, n637, n157, n828, n20659, n318, n381, 
        n25136, n23737, n25121, n21578, n254_adj_2827, n20579, n23108, 
        n20144, n24961, n20138, n20143, n24869, n924_adj_2828, n956, 
        n20146, n21745, n21744, n17787, n24878, n653_adj_2829, n27501, 
        n142, n157_adj_2830, n21027, n25004, n24893, n766, n20090, 
        n25272, n25273, n25274, n173, n188, n21028, n638, n765, 
        n986_adj_2831, n987, n333, n348_adj_2832, n21033, n85, n23813, 
        n24805, n364_adj_2833, n21034, n25125, n397, n21035, n21036, 
        n475, n21037, n491_adj_2834, n11113, n21038, n23825, n12166, 
        n23827, n27510, n900, n19975, n24997, n124, n11943, n475_adj_2835, 
        n25283, n19973, n19974, n23029, n20761, n12159, n12160, 
        n25029, n24827, n24998, n19966, n19967, n19968, n21333, 
        n21336, n21584, n25270, n25271, n19961, n21643, n17553, 
        n21588, n11952, n21589, n19959, n23104, n19955, n20239, 
        n20234, n20238, n19954, n19956, n19951, n19952, n19953, 
        n20205, n20208, n20207, n20764, n542, n573, n605, n636, 
        n25094, n892, n893, n669, n700, n25093, n19943, n732_adj_2836, 
        n797, n828_adj_2837, n19942, n19944, n860_adj_2838, n891_adj_2839, 
        n20145, n511, n508, n526_adj_2840, n542_adj_2841, n20762, 
        n731_adj_2842, n94, n25148, n19940, n23033, n19977, n19995, 
        n20605, n23036, n23037, n19937, n19938, n22797, n20089, 
        n21633, n21629, n21632, n20076, n19931, n19930, n19932, 
        n21570, n636_adj_2843, n20612, n700_adj_2844, n25141, n19928, 
        n19927, n684_adj_2845, n21579, n21582, n19929, n25027, n24976, 
        n444, n20629, n20630, n20632, n26428, n26429, n20627, 
        n20631, n21726, n20652, n20654, n20660, n20661, n20662, 
        n22784, n157_adj_2846, n22785, n17674, n20109, n251_adj_2847, 
        n27527, n747_adj_2848, n14960, n732_adj_2849, n94_adj_2850, 
        n125_adj_2851, n17544, n14348, n25129, n23675, n890_adj_2852, 
        n21332, n25266, n25267, n25268, n25249, n25436, n25431, 
        n25437, n15, n31, n24999, n61, n62_adj_2853, n15_adj_2854, 
        n24841, n31_adj_2855, n620_adj_2856, n635_adj_2857, n413_adj_2858, 
        n30_adj_2859, n31_adj_2860, n26967, n25434, n25433, n25435, 
        n25248, n476, n507, n17556, n573_adj_2861, n26966, n26968, 
        n26969, n605_adj_2862, n636_adj_2863, n26970, n26971, n26972, 
        n26973, n875_adj_2864, n891_adj_2865, n124_adj_2866, n46_adj_2867, 
        n20737, n27039, n859_adj_2868, n860_adj_2869, n21795, n700_adj_2870, 
        n20127, n732_adj_2871, n20128, n797_adj_2872, n828_adj_2873, 
        n27041, n25263, n25264, n25265, n860_adj_2874, n891_adj_2875, 
        n844_adj_2876, n124_adj_2877, n11998, n25147, n11999, n747_adj_2878, 
        n763_adj_2879, n14932, n22792, n24797, n21331, n21334, n954_adj_2880, 
        n173_adj_2881, n23106, n20736, n20739, n20740, n476_adj_2882, 
        n23117, n20742, n20743, n731_adj_2883, n94_adj_2884, n21801, 
        n20754, n20755, n20756, n221_adj_2885, n252_adj_2886, n20758, 
        n20759, n286, n19899, n15_adj_2887, n890_adj_2888, n349_adj_2889, 
        n19902, n6, n669_adj_2890, n700_adj_2891, n19914, n763_adj_2892, 
        n19917, n828_adj_2893, n860_adj_2894, n19920, n24376, n24373, 
        n24874, n24799, n20787, n20788, n20789, n20790, n20791, 
        n20792, n20794, n20795, n24372, n20797, n20798, n20801, 
        n24375, n24374, n22796, n20803, n20804, n24350, n24347, 
        n20806, n20807, n24349, n24348, n94_adj_2895, n125_adj_2896, 
        n158_adj_2897, n24346, n20098, n221_adj_2898, n286_adj_2899, 
        n349_adj_2900, n413_adj_2901, n444_adj_2902, n444_adj_2903, 
        n23120, n476_adj_2904, n507_adj_2905, n19935, n573_adj_2906, 
        n11986, n669_adj_2907, n700_adj_2908, n20189, n24310, n24307, 
        n24311, n19941, n20190, n797_adj_2909, n24309, n24308, n891_adj_2910, 
        n924_adj_2911, n19947, n1018, n24306, n21602, n158_adj_2912, 
        n189_adj_2913, n24826, n221_adj_2914, n286_adj_2915, n317_adj_2916, 
        n349_adj_2917, n413_adj_2918, n19962, n507_adj_2919, n19965, 
        n573_adj_2920, n605_adj_2921, n669_adj_2922, n700_adj_2923, 
        n732_adj_2924, n763_adj_2925, n20223, n24283, n24281, n24282, 
        n20111, n25261, n25260, n141, n25430, n236, n21030, n15_adj_2926, 
        n21023, n23157, n23158, n11139, n24926, n23159, n23162, 
        n19906, n19907, n19919, n19918, n24280, n24279, n653_adj_2927, 
        n108, n27509, n668_adj_2928, n23163, n93_adj_2929, n25262, 
        n19915, n812_adj_2930, n22869, n19913, n716_adj_2931, n731_adj_2932, 
        n653_adj_2933, n475_adj_2934, n142_adj_2935, n604_adj_2936, 
        n21024, n892_adj_2937, n25281, n19964, n19960, n397_adj_2938, 
        n668_adj_2939, n316_adj_2940, n270, n21025, n21026, n19901, 
        n19900, n142_adj_2941, n13831, n21041, n21029, n21042, n25127, 
        n19898, n23679, n19897, n22786, n21586, n21044, n397_adj_2942, 
        n844_adj_2943, n506_adj_2944, n25429, n24855, n25146, n859_adj_2945, 
        n875_adj_2946, n19945, n25279, n23740, n908_adj_2947, n541_adj_2948, 
        n796_adj_2949, n14719, n19492, n19933, n19934, n460_adj_2950, 
        n285, n25111, n25154, n397_adj_2951, n270_adj_2952, n93_adj_2953, 
        n14729, n348_adj_2954, n684_adj_2955, n25030, n491_adj_2956, 
        n526_adj_2957, n173_adj_2958, n333_adj_2959, n27517, n348_adj_2960, 
        n397_adj_2961, n23004, n23032, n762_adj_2962, n716_adj_2963, 
        n14712, n93_adj_2964, n23121, n11944, n23030, n526_adj_2965, 
        n475_adj_2966, n23002, n364_adj_2967, n379_adj_2968, n348_adj_2969, 
        n1002_adj_2970, n15_adj_2971, n684_adj_2972, n25428, n19912, 
        n17370, n668_adj_2973, n542_adj_2974, n25432, n24927, n17369, 
        n17368, n460_adj_2975, n285_adj_2976, n25142, n17367, n557_adj_2977, 
        n491_adj_2978, n17366, n22999, n573_adj_2979, n236_adj_2980, 
        n205, n301_adj_2981, n24866, n25124, n781_adj_2982, n251_adj_2983, 
        n21793, n21794, n12162, n12163, n157_adj_2984, n24928, n17555, 
        n491_adj_2985, n220, n460_adj_2986, n475_adj_2987, n24880, 
        n24879, n17542, n17543, n109_adj_2988, n635_adj_2989, n17365, 
        n19821, n812_adj_2990, n13817, n24818, n526_adj_2991, n882, 
        n890_adj_2992, n252_adj_2993, n23673, n25250, n23107, n23105, 
        n924_adj_2994, n24867, n19809, n20620, n23710, n20623, n62_adj_2995, 
        n23716, n20104, n25061, n21622, n23754, n20200, n101, 
        n19633, n27043, n27040, n27044, n25233, n27042, n27038, 
        n25112, n21615, n24852, n62_adj_2996, n25135, n23734, n20581, 
        n766_adj_2997, n20093, n23735, n21569, n25062, n286_adj_2998, 
        n27511, n20224, n23829, n985, n23706, n23672, n23035, 
        n23034, n22969, n205_adj_2999, n23751, n19939, n23031, n124_adj_3000, 
        n14349, n620_adj_3001, n25117, n22783, n21799, n21053, n21746, 
        n25140, n506_adj_3002, n11990, n23003, n23001, n13813, n348_adj_3003, 
        n19976, n21581, n572_adj_3004, n19993, n19994, n21612, n21610, 
        n20075, n23828, n23826, n23812, n142_adj_3005, n572_adj_3006, 
        n23824, n21580, n23814, n23818, n19630, n93_adj_3007, n25105, 
        n491_adj_3008, n20074, n21568, n23753, n23750, n25119, n12165, 
        n19862, n11945, n21577, n23739, n23736, n20087, n23712, 
        n23699, n22867, n23715, n23713, n20813, n23709, n23707, 
        n23708, n23698, n23695, n23678, n23676, n746, n22868, 
        n22866;
    
    PFUMX i17749 (.BLUT(n20077), .ALUT(n20078), .C0(index_i[4]), .Z(n20079));
    FD1S3BX quarter_wave_sample_register_i_i9 (.D(quarter_wave_sample_register_i_15__N_2126[9]), 
            .CK(i_ref_clk_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_i[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i9.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i8 (.D(quarter_wave_sample_register_i_15__N_2126[8]), 
            .CK(i_ref_clk_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_i[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i8.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i7 (.D(quarter_wave_sample_register_i_15__N_2126[7]), 
            .CK(i_ref_clk_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_i[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i7.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i6 (.D(quarter_wave_sample_register_i_15__N_2126[6]), 
            .CK(i_ref_clk_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_i[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i6.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i5 (.D(quarter_wave_sample_register_i_15__N_2126[5]), 
            .CK(i_ref_clk_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_i[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i5.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i4 (.D(quarter_wave_sample_register_i_15__N_2126[4]), 
            .CK(i_ref_clk_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_i[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i4.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i3 (.D(quarter_wave_sample_register_i_15__N_2126[3]), 
            .CK(i_ref_clk_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_i[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i3.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i2 (.D(quarter_wave_sample_register_i_15__N_2126[2]), 
            .CK(i_ref_clk_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_i[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i2.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i1 (.D(quarter_wave_sample_register_i_15__N_2126[1]), 
            .CK(i_ref_clk_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_i[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i1.GSR = "DISABLED";
    L6MUX21 i17762 (.D0(n21669), .D1(n21656), .SD(index_i[8]), .Z(n20092));
    FD1S3DX o_val_pipeline_i_1__i32 (.D(n1205[15]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(\o_val_pipeline_i[0] [15])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i32.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i31 (.D(n1205[14]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(\o_val_pipeline_i[0] [14])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i31.GSR = "DISABLED";
    LUT4 i20440_3_lut (.A(n21713), .B(n21714), .C(index_i[4]), .Z(n21715)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20440_3_lut.init = 16'hcaca;
    PFUMX i17752 (.BLUT(n20080), .ALUT(n20081), .C0(index_i[4]), .Z(n20082));
    PFUMX i17755 (.BLUT(n20083), .ALUT(n20084), .C0(index_i[4]), .Z(n20085));
    PFUMX i19379 (.BLUT(n21707), .ALUT(n21708), .C0(index_i[4]), .Z(n21709));
    LUT4 i19384_3_lut_4_lut (.A(n25098), .B(index_i[2]), .C(index_i[3]), 
         .D(n24995), .Z(n21714)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19384_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_194_Mux_7_i653_3_lut_4_lut (.A(n25098), .B(index_i[2]), .C(index_i[3]), 
         .D(n27516), .Z(n653)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_7_i653_3_lut_4_lut.init = 16'hf606;
    PFUMX i19387 (.BLUT(n557), .ALUT(n572), .C0(index_i[4]), .Z(n21717));
    FD1S3DX o_val_pipeline_i_1__i30 (.D(n1205[13]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(\o_val_pipeline_i[0] [13])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i30.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i29 (.D(n1205[12]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(\o_val_pipeline_i[0] [12])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i29.GSR = "DISABLED";
    LUT4 mux_194_Mux_2_i684_3_lut_4_lut (.A(n25098), .B(index_i[2]), .C(index_i[3]), 
         .D(n25107), .Z(n684)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_2_i684_3_lut_4_lut.init = 16'h6f60;
    PFUMX i19388 (.BLUT(n589), .ALUT(n604), .C0(index_i[4]), .Z(n21718));
    LUT4 mux_194_Mux_5_i30_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n30)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A (B+!(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_5_i30_3_lut_4_lut.init = 16'hcc67;
    FD1S3DX o_val_pipeline_i_1__i28 (.D(n1205[11]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(\o_val_pipeline_i[0] [11])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i28.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i27 (.D(n1205[10]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(\o_val_pipeline_i[0] [10])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i27.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i26 (.D(n1205[9]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(\o_val_pipeline_i[0] [9])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i26.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i25 (.D(n1205[8]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(\o_val_pipeline_i[0] [8])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i25.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i24 (.D(n1205[7]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(\o_val_pipeline_i[0] [7])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i24.GSR = "DISABLED";
    PFUMX i19389 (.BLUT(n620), .ALUT(n635), .C0(index_i[4]), .Z(n21719));
    LUT4 i18470_4_lut_4_lut_4_lut (.A(n25098), .B(index_i[2]), .C(index_i[4]), 
         .D(index_i[3]), .Z(n20800)) /* synthesis lut_function=(A (B)+!A !(B (C+(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18470_4_lut_4_lut_4_lut.init = 16'h999c;
    FD1S3DX o_val_pipeline_i_1__i23 (.D(n1205[6]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(\o_val_pipeline_i[0] [6])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i23.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i22 (.D(n1205[5]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(\o_val_pipeline_i[0] [5])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i22.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i21 (.D(n1205[4]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(\o_val_pipeline_i[0] [4])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i21.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i20 (.D(n1205[3]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(\o_val_pipeline_i[0] [3])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i20.GSR = "DISABLED";
    LUT4 i19378_3_lut (.A(n404), .B(n25139), .C(index_i[3]), .Z(n21708)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19378_3_lut.init = 16'hcaca;
    FD1S3DX o_val_pipeline_i_1__i19 (.D(n1205[2]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(\o_val_pipeline_i[0] [2])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i19.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i18 (.D(n1205[1]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(\o_val_pipeline_i[0] [1])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i18.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i17 (.D(n1205[0]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(\o_val_pipeline_i[0] [0])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i17.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i16 (.D(\o_val_pipeline_i[0] [15]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(modulation_output[15])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i16.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i15 (.D(\o_val_pipeline_i[0] [14]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(modulation_output[14])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i15.GSR = "DISABLED";
    PFUMX i19390 (.BLUT(n653_adj_2797), .ALUT(n668), .C0(index_i[4]), 
          .Z(n21720));
    FD1S3DX o_val_pipeline_i_1__i14 (.D(\o_val_pipeline_i[0] [13]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(modulation_output[13])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i14.GSR = "DISABLED";
    LUT4 i18435_3_lut_3_lut_4_lut (.A(n24892), .B(index_i[3]), .C(n93), 
         .D(index_i[4]), .Z(n20765)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18435_3_lut_3_lut_4_lut.init = 16'h11f0;
    FD1S3DX o_val_pipeline_i_1__i13 (.D(\o_val_pipeline_i[0] [12]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(modulation_output[12])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i13.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i0 (.D(o_phase[0]), .SP(i_resetb_c), .CK(i_ref_clk_c), 
            .Q(phase_i[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i0.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i12 (.D(\o_val_pipeline_i[0] [11]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(modulation_output[11])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i12.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i11 (.D(\o_val_pipeline_i[0] [10]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(modulation_output[10])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i11.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i10 (.D(\o_val_pipeline_i[0] [9]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(modulation_output[9])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i10.GSR = "DISABLED";
    FD1S3DX phase_negation_i_i0 (.D(phase_i[11]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(phase_negation_i[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_negation_i_i0.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i9 (.D(\o_val_pipeline_i[0] [8]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(modulation_output[8])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i9.GSR = "DISABLED";
    FD1S3DX index_i_i0 (.D(index_i_9__N_2106[0]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(index_i[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_i_i0.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i1 (.D(\o_val_pipeline_i[0] [0]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(modulation_output[0])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i1.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i0 (.D(quarter_wave_sample_register_i_15__N_2126[0]), 
            .CK(i_ref_clk_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_i[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i0.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i8 (.D(\o_val_pipeline_i[0] [7]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(modulation_output[7])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i8.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i7 (.D(\o_val_pipeline_i[0] [6]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(modulation_output[6])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i7.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i6 (.D(\o_val_pipeline_i[0] [5]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(modulation_output[5])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i6.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i5 (.D(\o_val_pipeline_i[0] [4]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(modulation_output[4])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i5.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i4 (.D(\o_val_pipeline_i[0] [3]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(modulation_output[3])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i4.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i3 (.D(\o_val_pipeline_i[0] [2]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(modulation_output[2])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i3.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i2 (.D(\o_val_pipeline_i[0] [1]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(modulation_output[1])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i2.GSR = "DISABLED";
    PFUMX i19391 (.BLUT(n684_adj_2798), .ALUT(n699), .C0(index_i[4]), 
          .Z(n21721));
    FD1S3DX index_i_i9 (.D(index_i_9__N_2106[9]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(index_i[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_i_i9.GSR = "DISABLED";
    FD1S3DX index_i_i8 (.D(index_i_9__N_2106[8]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(index_i[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_i_i8.GSR = "DISABLED";
    FD1S3DX index_i_i7 (.D(index_i_9__N_2106[7]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(index_i[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_i_i7.GSR = "DISABLED";
    FD1S3DX index_i_i6 (.D(index_i_9__N_2106[6]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(index_i[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_i_i6.GSR = "DISABLED";
    FD1S3DX index_i_i5 (.D(index_i_9__N_2106[5]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(index_i[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_i_i5.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i11 (.D(o_phase[11]), .SP(i_resetb_c), .CK(i_ref_clk_c), 
            .Q(phase_i[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i11.GSR = "DISABLED";
    FD1S3DX index_i_i4 (.D(index_i_9__N_2106[4]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(index_i[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_i_i4.GSR = "DISABLED";
    FD1S3DX index_i_i3 (.D(index_i_9__N_2106[3]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(index_i[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_i_i3.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i10 (.D(o_phase[10]), .SP(i_resetb_c), .CK(i_ref_clk_c), 
            .Q(phase_i[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i10.GSR = "DISABLED";
    FD1S3DX index_i_i2 (.D(index_i_9__N_2106[2]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(index_i[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_i_i2.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i9 (.D(o_phase[9]), .SP(i_resetb_c), .CK(i_ref_clk_c), 
            .Q(phase_i[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i9.GSR = "DISABLED";
    FD1S3DX index_i_i1 (.D(index_i_9__N_2106[1]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(index_i[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_i_i1.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i8 (.D(o_phase[8]), .SP(i_resetb_c), .CK(i_ref_clk_c), 
            .Q(phase_i[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i8.GSR = "DISABLED";
    FD1S3DX phase_negation_i_i1 (.D(phase_negation_i[0]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(phase_negation_i[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_negation_i_i1.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i7 (.D(o_phase[7]), .SP(i_resetb_c), .CK(i_ref_clk_c), 
            .Q(phase_i[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i7.GSR = "DISABLED";
    PFUMX i19392 (.BLUT(n716), .ALUT(n731), .C0(index_i[4]), .Z(n21722));
    L6MUX21 i19279 (.D0(n21603), .D1(n21604), .SD(index_i[7]), .Z(n21609));
    L6MUX21 i19298 (.D0(n21620), .D1(n21621), .SD(index_i[7]), .Z(n21628));
    L6MUX21 i19300 (.D0(n21624), .D1(n21625), .SD(index_i[7]), .Z(n21630));
    PFUMX i19301 (.BLUT(n21626), .ALUT(n21627), .C0(index_i[7]), .Z(n21631));
    FD1P3AX phase_i_i0_i6 (.D(o_phase[6]), .SP(i_resetb_c), .CK(i_ref_clk_c), 
            .Q(phase_i[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i6.GSR = "DISABLED";
    PFUMX i19393 (.BLUT(n747), .ALUT(n762), .C0(index_i[4]), .Z(n21723));
    FD1P3AX phase_i_i0_i5 (.D(o_phase[5]), .SP(i_resetb_c), .CK(i_ref_clk_c), 
            .Q(phase_i[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i5.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i4 (.D(o_phase[4]), .SP(i_resetb_c), .CK(i_ref_clk_c), 
            .Q(phase_i[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i4.GSR = "DISABLED";
    PFUMX i18250 (.BLUT(n382), .ALUT(n509), .C0(index_i[7]), .Z(n20580));
    FD1P3AX phase_i_i0_i3 (.D(o_phase[3]), .SP(i_resetb_c), .CK(i_ref_clk_c), 
            .Q(phase_i[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i3.GSR = "DISABLED";
    PFUMX i19394 (.BLUT(n781), .ALUT(n796), .C0(index_i[4]), .Z(n21724));
    PFUMX i19395 (.BLUT(n812), .ALUT(n11935), .C0(index_i[4]), .Z(n21725));
    PFUMX i19397 (.BLUT(n875), .ALUT(n890), .C0(index_i[4]), .Z(n21727));
    LUT4 n699_bdd_4_lut_21434_4_lut (.A(n24892), .B(index_i[3]), .C(index_i[2]), 
         .D(index_i[6]), .Z(n22968)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C+(D)))+!A (B ((D)+!C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n699_bdd_4_lut_21434_4_lut.init = 16'hee3c;
    FD1P3AX phase_i_i0_i2 (.D(o_phase[2]), .SP(i_resetb_c), .CK(i_ref_clk_c), 
            .Q(phase_i[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i2.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i1 (.D(o_phase[1]), .SP(i_resetb_c), .CK(i_ref_clk_c), 
            .Q(phase_i[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i1.GSR = "DISABLED";
    PFUMX i19398 (.BLUT(n908), .ALUT(n923), .C0(index_i[4]), .Z(n21728));
    LUT4 i19377_3_lut (.A(n25144), .B(n325), .C(index_i[3]), .Z(n21707)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19377_3_lut.init = 16'hcaca;
    PFUMX i19399 (.BLUT(n939), .ALUT(n954), .C0(index_i[4]), .Z(n21729));
    L6MUX21 i19326 (.D0(n21654), .D1(n21655), .SD(index_i[7]), .Z(n21656));
    LUT4 n124_bdd_3_lut_22767_4_lut (.A(n24892), .B(index_i[3]), .C(index_i[4]), 
         .D(n93), .Z(n23000)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n124_bdd_3_lut_22767_4_lut.init = 16'hfe0e;
    PFUMX i19400 (.BLUT(n971), .ALUT(n986), .C0(index_i[4]), .Z(n21730));
    LUT4 n476_bdd_3_lut_21573_3_lut_4_lut (.A(index_i[2]), .B(n24994), .C(n491), 
         .D(index_i[4]), .Z(n23116)) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))+!A !(B ((D)+!C)+!B !(C+(D)))) */ ;
    defparam n476_bdd_3_lut_21573_3_lut_4_lut.init = 16'h99f0;
    L6MUX21 i18263 (.D0(n20591), .D1(n20592), .SD(index_i[7]), .Z(n20593));
    L6MUX21 i18266 (.D0(n20594), .D1(n20595), .SD(index_i[7]), .Z(n20596));
    LUT4 i17606_3_lut_3_lut_4_lut (.A(index_i[2]), .B(n24994), .C(n24996), 
         .D(index_i[3]), .Z(n19936)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (B (C (D))+!B (C+!(D)))) */ ;
    defparam i17606_3_lut_3_lut_4_lut.init = 16'hf099;
    PFUMX i19401 (.BLUT(n1002), .ALUT(n1017), .C0(index_i[4]), .Z(n21731));
    PFUMX i19386 (.BLUT(n526), .ALUT(n541), .C0(index_i[4]), .Z(n21716));
    L6MUX21 i19339 (.D0(n21667), .D1(n21668), .SD(index_i[7]), .Z(n21669));
    L6MUX21 i18294 (.D0(n20613), .D1(n20614), .SD(index_i[6]), .Z(n20624));
    L6MUX21 i18295 (.D0(n20615), .D1(n20616), .SD(index_i[6]), .Z(n20625));
    L6MUX21 i18298 (.D0(n20621), .D1(n20622), .SD(index_i[7]), .Z(n20628));
    PFUMX i19422 (.BLUT(n21750), .ALUT(n21751), .C0(index_i[4]), .Z(n21752));
    PFUMX i19425 (.BLUT(n21753), .ALUT(n21754), .C0(index_i[4]), .Z(n21755));
    L6MUX21 i17811 (.D0(n20133), .D1(n20134), .SD(index_i[7]), .Z(n20141));
    CCU2D unary_minus_10_add_3_3 (.A0(quarter_wave_sample_register_i[1]), 
          .B0(GND_net), .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[2]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17363), .COUT(n17364), 
          .S0(o_val_pipeline_i_0__15__N_2157[1]), .S1(o_val_pipeline_i_0__15__N_2157[2]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam unary_minus_10_add_3_3.INIT0 = 16'hf555;
    defparam unary_minus_10_add_3_3.INIT1 = 16'hf555;
    defparam unary_minus_10_add_3_3.INJECT1_0 = "NO";
    defparam unary_minus_10_add_3_3.INJECT1_1 = "NO";
    CCU2D unary_minus_10_add_3_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(quarter_wave_sample_register_i[0]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .COUT(n17363), .S1(o_val_pipeline_i_0__15__N_2157[0]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam unary_minus_10_add_3_1.INIT0 = 16'hF000;
    defparam unary_minus_10_add_3_1.INIT1 = 16'h0aaa;
    defparam unary_minus_10_add_3_1.INJECT1_0 = "NO";
    defparam unary_minus_10_add_3_1.INJECT1_1 = "NO";
    L6MUX21 i17812 (.D0(n20135), .D1(n20136), .SD(index_i[7]), .Z(n20142));
    L6MUX21 i17873 (.D0(n20195), .D1(n20196), .SD(index_i[7]), .Z(n20203));
    L6MUX21 i17874 (.D0(n20197), .D1(n20198), .SD(index_i[7]), .Z(n20204));
    LUT4 mux_194_Mux_10_i317_3_lut_3_lut_4_lut (.A(n24892), .B(index_i[3]), 
         .C(n24925), .D(index_i[4]), .Z(n317)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_10_i317_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 mux_194_Mux_7_i443_3_lut_4_lut (.A(index_i[2]), .B(n24994), .C(index_i[3]), 
         .D(n25101), .Z(n443)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;
    defparam mux_194_Mux_7_i443_3_lut_4_lut.init = 16'h6f60;
    L6MUX21 i17876 (.D0(n20201), .D1(n20202), .SD(index_i[7]), .Z(n20206));
    L6MUX21 i17905 (.D0(n20228), .D1(n20229), .SD(index_i[7]), .Z(n20235));
    L6MUX21 i17906 (.D0(n20230), .D1(n20231), .SD(index_i[7]), .Z(n20236));
    PFUMX i17907 (.BLUT(n20232), .ALUT(n20233), .C0(index_i[7]), .Z(n20237));
    LUT4 mux_194_Mux_3_i860_3_lut_4_lut (.A(index_i[2]), .B(n24994), .C(index_i[4]), 
         .D(n859), .Z(n860)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam mux_194_Mux_3_i860_3_lut_4_lut.init = 16'hf606;
    LUT4 i17751_3_lut (.A(n25126), .B(n25149), .C(index_i[3]), .Z(n20081)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17751_3_lut.init = 16'hcaca;
    PFUMX i19459 (.BLUT(n21787), .ALUT(n21788), .C0(index_i[4]), .Z(n21789));
    PFUMX i19462 (.BLUT(n21790), .ALUT(n21791), .C0(index_i[4]), .Z(n21792));
    L6MUX21 i19273 (.D0(n21591), .D1(n21592), .SD(index_i[6]), .Z(n21603));
    PFUMX i19468 (.BLUT(n21796), .ALUT(n21797), .C0(index_i[4]), .Z(n21798));
    L6MUX21 i19274 (.D0(n21593), .D1(n21594), .SD(index_i[6]), .Z(n21604));
    L6MUX21 i19275 (.D0(n21595), .D1(n21596), .SD(index_i[6]), .Z(n21605));
    PFUMX i17790 (.BLUT(n221), .ALUT(n252), .C0(index_i[5]), .Z(n20120));
    L6MUX21 i19291 (.D0(n11940), .D1(n20744), .SD(index_i[6]), .Z(n21621));
    L6MUX21 i19293 (.D0(n20757), .D1(n20760), .SD(index_i[6]), .Z(n21623));
    L6MUX21 i19294 (.D0(n574), .D1(n20763), .SD(index_i[6]), .Z(n21624));
    L6MUX21 i19295 (.D0(n20766), .D1(n764), .SD(index_i[6]), .Z(n21625));
    LUT4 i19424_3_lut (.A(n27500), .B(n27505), .C(index_i[3]), .Z(n21754)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19424_3_lut.init = 16'hcaca;
    PFUMX i19324 (.BLUT(n21650), .ALUT(n21651), .C0(index_i[6]), .Z(n21654));
    PFUMX i19325 (.BLUT(n21652), .ALUT(n21653), .C0(index_i[6]), .Z(n21655));
    PFUMX i18265 (.BLUT(n701), .ALUT(n764_adj_2799), .C0(index_i[6]), 
          .Z(n20595));
    PFUMX i19337 (.BLUT(n21663), .ALUT(n21664), .C0(index_i[6]), .Z(n21667));
    PFUMX i19338 (.BLUT(n21665), .ALUT(n21666), .C0(index_i[6]), .Z(n21668));
    PFUMX i18284 (.BLUT(n732), .ALUT(n763), .C0(index_i[5]), .Z(n20614));
    LUT4 i19323_3_lut_4_lut_4_lut (.A(n24925), .B(index_i[4]), .C(index_i[5]), 
         .D(n24868), .Z(n21653)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A (B (C+(D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19323_3_lut_4_lut_4_lut.init = 16'h101c;
    L6MUX21 i18286 (.D0(n21616), .D1(n891), .SD(index_i[5]), .Z(n20616));
    L6MUX21 i18289 (.D0(n20603), .D1(n20604), .SD(index_i[6]), .Z(n20619));
    L6MUX21 i18291 (.D0(n20607), .D1(n20608), .SD(index_i[6]), .Z(n20621));
    L6MUX21 i18292 (.D0(n20609), .D1(n20610), .SD(index_i[6]), .Z(n20622));
    PFUMX i18422 (.BLUT(n20748), .ALUT(n20749), .C0(index_i[4]), .Z(n20752));
    L6MUX21 i18296 (.D0(n20617), .D1(n20618), .SD(index_i[6]), .Z(n20626));
    PFUMX i18423 (.BLUT(n20750), .ALUT(n20751), .C0(index_i[4]), .Z(n20753));
    LUT4 i18323_3_lut_3_lut_4_lut (.A(n24892), .B(index_i[3]), .C(n316), 
         .D(index_i[4]), .Z(n20653)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18323_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 i19383_3_lut_3_lut_4_lut (.A(index_i[2]), .B(n24994), .C(n25101), 
         .D(index_i[3]), .Z(n21713)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (B (C (D))+!B (C+!(D)))) */ ;
    defparam i19383_3_lut_3_lut_4_lut.init = 16'hf099;
    LUT4 mux_194_Mux_1_i924_3_lut (.A(n316_adj_2800), .B(n412), .C(index_i[4]), 
         .Z(n924)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_1_i924_3_lut.init = 16'hcaca;
    L6MUX21 i17772 (.D0(n20773), .D1(n20780), .SD(index_i[6]), .Z(n20102));
    L6MUX21 i19410 (.D0(n21732), .D1(n21733), .SD(index_i[6]), .Z(n21740));
    PFUMX i17820 (.BLUT(n158), .ALUT(n189), .C0(index_i[5]), .Z(n20150));
    L6MUX21 i19411 (.D0(n21734), .D1(n21735), .SD(index_i[6]), .Z(n21741));
    L6MUX21 i19412 (.D0(n21736), .D1(n21737), .SD(index_i[6]), .Z(n21742));
    L6MUX21 i19413 (.D0(n21738), .D1(n21739), .SD(index_i[6]), .Z(n21743));
    L6MUX21 i17775 (.D0(n20793), .D1(n20796), .SD(index_i[6]), .Z(n20105));
    L6MUX21 i18328 (.D0(n20656), .D1(n20657), .SD(index_i[6]), .Z(n382_adj_2801));
    L6MUX21 i17776 (.D0(n20799), .D1(n20802), .SD(index_i[6]), .Z(n20106));
    L6MUX21 i17777 (.D0(n20805), .D1(n20808), .SD(index_i[6]), .Z(n20107));
    L6MUX21 i18335 (.D0(n20663), .D1(n20664), .SD(index_i[6]), .Z(n509_adj_2802));
    L6MUX21 i19290 (.D0(n20738), .D1(n20741), .SD(index_i[6]), .Z(n21620));
    PFUMX i18441 (.BLUT(n20767), .ALUT(n20768), .C0(index_i[4]), .Z(n20771));
    PFUMX i18442 (.BLUT(n20769), .ALUT(n20770), .C0(index_i[4]), .Z(n20772));
    PFUMX i18448 (.BLUT(n20774), .ALUT(n20775), .C0(index_i[4]), .Z(n20778));
    PFUMX i18449 (.BLUT(n20776), .ALUT(n20777), .C0(index_i[4]), .Z(n20779));
    PFUMX i18455 (.BLUT(n20781), .ALUT(n20782), .C0(index_i[4]), .Z(n20785));
    PFUMX i18456 (.BLUT(n20783), .ALUT(n20784), .C0(index_i[4]), .Z(n20786));
    L6MUX21 i17803 (.D0(n20117), .D1(n20118), .SD(index_i[6]), .Z(n20133));
    L6MUX21 i17804 (.D0(n20119), .D1(n20120), .SD(index_i[6]), .Z(n20134));
    L6MUX21 i17805 (.D0(n20121), .D1(n20122), .SD(index_i[6]), .Z(n20135));
    L6MUX21 i17806 (.D0(n20123), .D1(n20124), .SD(index_i[6]), .Z(n20136));
    L6MUX21 i17807 (.D0(n20125), .D1(n20126), .SD(index_i[6]), .Z(n20137));
    L6MUX21 i17809 (.D0(n20129), .D1(n20130), .SD(index_i[6]), .Z(n20139));
    L6MUX21 i17834 (.D0(n20148), .D1(n20149), .SD(index_i[6]), .Z(n20164));
    L6MUX21 i17835 (.D0(n20150), .D1(n20151), .SD(index_i[6]), .Z(n20165));
    L6MUX21 i17836 (.D0(n20152), .D1(n20153), .SD(index_i[6]), .Z(n20166));
    PFUMX i17838 (.BLUT(n20156), .ALUT(n20157), .C0(index_i[6]), .Z(n20168));
    L6MUX21 i17839 (.D0(n20158), .D1(n20159), .SD(index_i[6]), .Z(n20169));
    L6MUX21 i17840 (.D0(n20160), .D1(n20161), .SD(index_i[6]), .Z(n20170));
    PFUMX i17841 (.BLUT(n20162), .ALUT(n20163), .C0(index_i[6]), .Z(n20171));
    LUT4 i15289_3_lut (.A(n25139), .B(n25151), .C(index_i[3]), .Z(n17552)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15289_3_lut.init = 16'hcaca;
    LUT4 i20419_3_lut (.A(n21571), .B(n21572), .C(index_i[4]), .Z(n21573)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20419_3_lut.init = 16'hcaca;
    LUT4 i15288_3_lut (.A(n25151), .B(n25144), .C(index_i[3]), .Z(n17551)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15288_3_lut.init = 16'hcaca;
    L6MUX21 i17865 (.D0(n20179), .D1(n20180), .SD(index_i[6]), .Z(n20195));
    L6MUX21 i17866 (.D0(n20181), .D1(n20182), .SD(index_i[6]), .Z(n20196));
    L6MUX21 i17867 (.D0(n20183), .D1(n20184), .SD(index_i[6]), .Z(n20197));
    L6MUX21 i17868 (.D0(n20185), .D1(n20186), .SD(index_i[6]), .Z(n20198));
    L6MUX21 i17869 (.D0(n20187), .D1(n20188), .SD(index_i[6]), .Z(n20199));
    L6MUX21 i17871 (.D0(n20191), .D1(n20192), .SD(index_i[6]), .Z(n20201));
    L6MUX21 i17872 (.D0(n20193), .D1(n20194), .SD(index_i[6]), .Z(n20202));
    LUT4 i17581_else_4_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[4]), 
         .D(index_i[3]), .Z(n25269)) /* synthesis lut_function=(!(A (B (C)+!B !(C (D)+!C !(D)))+!A (B (C+(D))+!B !(C+!(D))))) */ ;
    defparam i17581_else_4_lut.init = 16'h381f;
    L6MUX21 i17897 (.D0(n20212), .D1(n20213), .SD(index_i[6]), .Z(n20227));
    L6MUX21 i17898 (.D0(n20214), .D1(n20215), .SD(index_i[6]), .Z(n20228));
    L6MUX21 i17899 (.D0(n20216), .D1(n20217), .SD(index_i[6]), .Z(n20229));
    L6MUX21 i17900 (.D0(n20218), .D1(n20219), .SD(index_i[6]), .Z(n20230));
    L6MUX21 i17901 (.D0(n20220), .D1(n20221), .SD(index_i[6]), .Z(n20231));
    LUT4 mux_194_Mux_0_i428_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[2]), .D(index_i[3]), .Z(n428)) /* synthesis lut_function=(A (B (C+(D))+!B !(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_0_i428_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h8fe1;
    LUT4 mux_194_Mux_0_i604_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n604)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)+!C !(D)))+!A (B (C (D))+!B (C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_0_i604_3_lut_4_lut_4_lut.init = 16'h0e65;
    LUT4 i9422_3_lut_3_lut_4_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n762_adj_2803)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9422_3_lut_3_lut_4_lut_3_lut_4_lut.init = 16'h1999;
    LUT4 i9427_3_lut_4_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n844)) /* synthesis lut_function=(A (B)+!A !(B+!(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9427_3_lut_4_lut_3_lut_4_lut.init = 16'h9998;
    LUT4 mux_194_Mux_0_i653_3_lut (.A(n24996), .B(n27515), .C(index_i[3]), 
         .Z(n653_adj_2797)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_0_i653_3_lut.init = 16'hcaca;
    LUT4 i9410_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n11976)) /* synthesis lut_function=(!(A (B (C)+!B ((D)+!C))+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9410_3_lut_4_lut_4_lut.init = 16'h4969;
    LUT4 mux_194_Mux_2_i890_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n890_adj_2804)) /* synthesis lut_function=(A (B (C)+!B !(C+!(D)))+!A !(B (C+(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_2_i890_3_lut_4_lut_4_lut.init = 16'h9394;
    LUT4 i9369_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n11935)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))+!A !(B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9369_3_lut_4_lut_4_lut.init = 16'hb5b3;
    LUT4 i9372_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n11938)) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B ((D)+!C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9372_3_lut_4_lut_4_lut.init = 16'hcdad;
    LUT4 i19470_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[1]), .Z(n21800)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C))+!A (B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19470_3_lut_4_lut_4_lut_4_lut.init = 16'h29a9;
    LUT4 mux_194_Mux_6_i781_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), 
         .B(index_i[2]), .C(index_i[3]), .D(index_i[0]), .Z(n781_adj_2805)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+(D)))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_6_i781_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h9993;
    L6MUX21 i18717 (.D0(n21039), .D1(n21040), .SD(index_i[6]), .Z(n21047));
    LUT4 i19420_3_lut (.A(n25138), .B(n27505), .C(index_i[3]), .Z(n21750)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19420_3_lut.init = 16'hcaca;
    L6MUX21 i18720 (.D0(n21045), .D1(n21046), .SD(index_i[6]), .Z(n21050));
    LUT4 mux_194_Mux_5_i252_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[4]), .Z(n252)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+(D)))+!A (B (C (D))+!B !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_5_i252_3_lut_4_lut.init = 16'hc993;
    LUT4 i15291_3_lut_4_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[1]), .D(index_i[3]), .Z(n17554)) /* synthesis lut_function=(A (B (C (D))+!B !(D))+!A (B+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i15291_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'hd566;
    LUT4 n557_bdd_3_lut_21486_4_lut_4_lut_4_lut (.A(index_i[3]), .B(index_i[2]), 
         .C(index_i[4]), .D(index_i[1]), .Z(n23026)) /* synthesis lut_function=(A (B (C)+!B !(C+(D)))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n557_bdd_3_lut_21486_4_lut_4_lut_4_lut.init = 16'h8587;
    LUT4 mux_194_Mux_4_i93_3_lut_4_lut_3_lut_rep_550_4_lut (.A(index_i[0]), 
         .B(index_i[3]), .C(index_i[1]), .D(index_i[2]), .Z(n25110)) /* synthesis lut_function=(!(A (B+(C (D)))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_4_i93_3_lut_4_lut_3_lut_rep_550_4_lut.init = 16'h4666;
    LUT4 mux_194_Mux_4_i236_3_lut_4_lut_4_lut_3_lut_rep_548_4_lut (.A(index_i[0]), 
         .B(index_i[3]), .C(index_i[1]), .D(index_i[2]), .Z(n25108)) /* synthesis lut_function=(A (B)+!A !(B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_4_i236_3_lut_4_lut_4_lut_3_lut_rep_548_4_lut.init = 16'h999d;
    LUT4 i17742_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n20072)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(D))+!A (B (D)+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i17742_3_lut_4_lut_4_lut_4_lut.init = 16'hd52b;
    LUT4 i17586_3_lut_4_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[3]), 
         .C(index_i[1]), .D(index_i[2]), .Z(n19916)) /* synthesis lut_function=(A (B+(C (D)))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i17586_3_lut_4_lut_3_lut_4_lut.init = 16'hb999;
    LUT4 mux_194_Mux_8_i635_3_lut_4_lut_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[0]), .D(index_i[1]), .Z(n635_adj_2806)) /* synthesis lut_function=(!(A (B)+!A !(B+(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_8_i635_3_lut_4_lut_3_lut_4_lut.init = 16'h7666;
    LUT4 mux_194_Mux_9_i30_3_lut_4_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n30_adj_2807)) /* synthesis lut_function=(A (B (C (D)))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_9_i30_3_lut_4_lut_4_lut_4_lut.init = 16'h9111;
    LUT4 mux_194_Mux_8_i506_3_lut_4_lut_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[0]), .D(index_i[1]), .Z(n506)) /* synthesis lut_function=(!(A (B+!(C+(D)))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_8_i506_3_lut_4_lut_3_lut_4_lut.init = 16'h6664;
    LUT4 mux_194_Mux_0_i46_3_lut_4_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n46)) /* synthesis lut_function=(A (B)+!A ((C+(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_0_i46_3_lut_4_lut_4_lut_4_lut.init = 16'hddd9;
    LUT4 i17628_3_lut_4_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n19958)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i17628_3_lut_4_lut_4_lut_4_lut.init = 16'h6444;
    LUT4 mux_194_Mux_8_i716_3_lut_4_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n716_adj_2808)) /* synthesis lut_function=(!(A (B)+!A !(B+(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_8_i716_3_lut_4_lut_4_lut_4_lut.init = 16'h7776;
    LUT4 mux_194_Mux_0_i890_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n890)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)+!C !(D)))+!A !(B (C)+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_0_i890_3_lut_4_lut_4_lut.init = 16'h70ca;
    LUT4 mux_194_Mux_1_i349_3_lut (.A(n506), .B(n348), .C(index_i[4]), 
         .Z(n349)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_1_i349_3_lut.init = 16'hcaca;
    LUT4 n9595_bdd_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n23752)) /* synthesis lut_function=(A (B (C)+!B ((D)+!C))+!A (B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n9595_bdd_3_lut_4_lut_4_lut_4_lut.init = 16'he7c7;
    LUT4 n301_bdd_3_lut_22890_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n23749)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A !((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n301_bdd_3_lut_22890_4_lut_4_lut_4_lut.init = 16'h7173;
    LUT4 mux_194_Mux_9_i316_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n316)) /* synthesis lut_function=(!(A (B (C)+!B !(C+(D)))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_9_i316_3_lut_4_lut_4_lut_4_lut.init = 16'h7e7c;
    LUT4 mux_194_Mux_7_i781_3_lut_4_lut_4_lut_4_lut_4_lut (.A(index_i[1]), 
         .B(index_i[2]), .C(index_i[0]), .D(index_i[3]), .Z(n781_adj_2809)) /* synthesis lut_function=(!(A (B (D)+!B ((D)+!C))+!A (B (D)+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_7_i781_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'h11ec;
    LUT4 mux_194_Mux_7_i747_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), 
         .B(index_i[2]), .C(index_i[3]), .D(index_i[0]), .Z(n747_adj_2810)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))+!A (B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_7_i747_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'he1e3;
    LUT4 i18418_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[3]), 
         .C(index_i[2]), .D(index_i[0]), .Z(n20748)) /* synthesis lut_function=(A (B (C (D))+!B (C))+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18418_3_lut_4_lut_4_lut_4_lut.init = 16'hb434;
    LUT4 n676_bdd_2_lut_22926_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[3]), 
         .C(index_i[2]), .D(index_i[0]), .Z(n23711)) /* synthesis lut_function=(!(A (B+(C+!(D)))+!A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n676_bdd_2_lut_22926_4_lut_4_lut_4_lut.init = 16'h1210;
    PFUMX i23060 (.BLUT(n25299), .ALUT(n25300), .C0(index_i[3]), .Z(n62));
    LUT4 mux_194_Mux_7_i491_3_lut_4_lut_4_lut_4_lut_4_lut (.A(index_i[1]), 
         .B(index_i[3]), .C(index_i[2]), .D(index_i[0]), .Z(n491_adj_2811)) /* synthesis lut_function=(!(A (B (C+!(D))+!B ((D)+!C))+!A !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_7_i491_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'h5870;
    LUT4 mux_194_Mux_1_i348_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[3]), 
         .C(index_i[2]), .D(index_i[0]), .Z(n348)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_1_i348_3_lut_4_lut_4_lut_4_lut.init = 16'h7870;
    LUT4 mux_194_Mux_0_i443_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .D(index_i[3]), .Z(n443_adj_2812)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C (D))+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_0_i443_3_lut_4_lut_4_lut_4_lut.init = 16'h0ed5;
    LUT4 i17748_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[3]), 
         .C(index_i[2]), .D(index_i[0]), .Z(n20078)) /* synthesis lut_function=(!(A (B+!((D)+!C))+!A !(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i17748_3_lut_4_lut_4_lut_4_lut.init = 16'h6747;
    LUT4 mux_194_Mux_0_i251_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n251)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A !(B ((D)+!C)+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_0_i251_3_lut_4_lut_4_lut_4_lut.init = 16'h543c;
    LUT4 i20426_3_lut (.A(n20071), .B(n20072), .C(index_i[4]), .Z(n20073)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20426_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_8_i61_3_lut_rep_284_4_lut_4_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[2]), .D(index_i[3]), .Z(n24844)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A (B (C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_8_i61_3_lut_rep_284_4_lut_4_lut_4_lut.init = 16'he0f8;
    LUT4 mux_194_Mux_8_i251_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[2]), .D(index_i[3]), .Z(n251_adj_2813)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_8_i251_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h07e0;
    LUT4 i18722_3_lut (.A(n21049), .B(n21050), .C(index_i[7]), .Z(n21052)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18722_3_lut.init = 16'hcaca;
    LUT4 i18419_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n20749)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18419_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hf81f;
    LUT4 i19284_3_lut_4_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n21614)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(D))+!A !(B (D)+!B ((D)+!C)))) */ ;
    defparam i19284_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'h7f01;
    LUT4 i19005_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21335)) /* synthesis lut_function=(A (C)+!A !(B (C)+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19005_3_lut_4_lut_4_lut.init = 16'hb4b5;
    LUT4 mux_194_Mux_8_i109_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n109)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C+!(D)))+!A (B (C (D)+!C !(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_8_i109_3_lut_4_lut_4_lut.init = 16'hf83e;
    LUT4 mux_194_Mux_0_i460_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n460)) /* synthesis lut_function=(A (B+(C (D)+!C !(D)))+!A (B (C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_0_i460_3_lut_4_lut_4_lut.init = 16'hf8cb;
    LUT4 mux_194_Mux_1_i317_3_lut (.A(n301), .B(n908_adj_2814), .C(index_i[4]), 
         .Z(n317_adj_2815)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_1_i317_3_lut.init = 16'hcaca;
    LUT4 i18721_3_lut (.A(n21047), .B(n21048), .C(index_i[7]), .Z(n21051)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18721_3_lut.init = 16'hcaca;
    LUT4 i19418_3_lut (.A(n25120), .B(n27508), .C(index_i[3]), .Z(n21748)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19418_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_7_i699_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n699_adj_2816)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C+!(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_7_i699_3_lut_4_lut_4_lut.init = 16'hf07e;
    LUT4 mux_194_Mux_0_i412_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[1]), .D(index_i[3]), .Z(n412_adj_2817)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C (D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_0_i412_3_lut_4_lut_4_lut.init = 16'hf12a;
    LUT4 mux_194_Mux_1_i684_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n684_adj_2818)) /* synthesis lut_function=(A (B ((D)+!C)+!B !((D)+!C))+!A !(B (C+(D))+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_1_i684_3_lut_4_lut_4_lut.init = 16'h992d;
    LUT4 mux_194_Mux_11_i445_3_lut_4_lut_4_lut_4_lut (.A(index_i[3]), .B(index_i[4]), 
         .C(index_i[5]), .D(n24978), .Z(n445)) /* synthesis lut_function=(!(A (B (C))+!A !(B+(C+(D))))) */ ;
    defparam mux_194_Mux_11_i445_3_lut_4_lut_4_lut_4_lut.init = 16'h7f7e;
    LUT4 mux_194_Mux_1_i716_3_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[1]), .D(index_i[3]), .Z(n716_adj_2819)) /* synthesis lut_function=(!(A (B (D)+!B !(C))+!A !(B (C (D))+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_1_i716_3_lut_4_lut_4_lut.init = 16'h70a9;
    LUT4 i20008_3_lut (.A(n21747), .B(n21748), .C(index_i[4]), .Z(n21749)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20008_3_lut.init = 16'hcaca;
    LUT4 i17747_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n20077)) /* synthesis lut_function=(A (B (C (D)))+!A !(B+(C+(D)))) */ ;
    defparam i17747_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h8001;
    LUT4 i20428_3_lut (.A(n20068), .B(n20069), .C(index_i[4]), .Z(n20070)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20428_3_lut.init = 16'hcaca;
    LUT4 i17627_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n19957)) /* synthesis lut_function=(!(A (B (C (D)))+!A !(B+(C+(D))))) */ ;
    defparam i17627_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h7ffe;
    LUT4 mux_194_Mux_0_i379_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n379)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !((D)+!C))+!A !(B ((D)+!C)+!B (D))) */ ;
    defparam mux_194_Mux_0_i379_3_lut_4_lut_4_lut.init = 16'h8079;
    LUT4 mux_194_Mux_8_i443_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n443_adj_2820)) /* synthesis lut_function=(A (B (C+!(D))+!B !((D)+!C))+!A !(B (D)+!B ((D)+!C))) */ ;
    defparam mux_194_Mux_8_i443_3_lut_4_lut_4_lut.init = 16'h80fc;
    LUT4 n62_bdd_3_lut_21460_4_lut_4_lut (.A(n24952), .B(index_i[3]), .C(n24892), 
         .D(index_i[4]), .Z(n22865)) /* synthesis lut_function=(A (B (C+!(D))+!B !((D)+!C))+!A (B (C+!(D))+!B (C+(D)))) */ ;
    defparam n62_bdd_3_lut_21460_4_lut_4_lut.init = 16'hd1fc;
    LUT4 i11106_2_lut_3_lut_4_lut (.A(n24978), .B(n25092), .C(index_i[6]), 
         .D(index_i[5]), .Z(n254)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i11106_2_lut_3_lut_4_lut.init = 16'hfef0;
    LUT4 mux_194_Mux_3_i252_3_lut_4_lut (.A(n24891), .B(index_i[3]), .C(index_i[4]), 
         .D(n14964), .Z(n252_adj_2821)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_3_i252_3_lut_4_lut.init = 16'h08f8;
    LUT4 mux_194_Mux_10_i62_3_lut_3_lut_4_lut (.A(n24891), .B(index_i[3]), 
         .C(n24960), .D(index_i[4]), .Z(n62_adj_2822)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_10_i62_3_lut_3_lut_4_lut.init = 16'hf077;
    LUT4 mux_194_Mux_8_i860_3_lut_4_lut (.A(n24891), .B(index_i[3]), .C(index_i[4]), 
         .D(n24960), .Z(n860_adj_2823)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_8_i860_3_lut_4_lut.init = 16'h08f8;
    LUT4 i18325_3_lut_4_lut (.A(n24891), .B(index_i[3]), .C(index_i[4]), 
         .D(n364), .Z(n20655)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18325_3_lut_4_lut.init = 16'h8f80;
    LUT4 i11054_2_lut_rep_250_3_lut_4_lut (.A(n24891), .B(index_i[3]), .C(index_i[5]), 
         .D(index_i[4]), .Z(n24810)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11054_2_lut_rep_250_3_lut_4_lut.init = 16'hf080;
    LUT4 n347_bdd_3_lut_22071 (.A(n25149), .B(n25137), .C(index_i[3]), 
         .Z(n23674)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n347_bdd_3_lut_22071.init = 16'hcaca;
    LUT4 index_i_6__bdd_3_lut_21493_rep_271_4_lut (.A(n24891), .B(index_i[3]), 
         .C(index_i[4]), .D(n24843), .Z(n24831)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam index_i_6__bdd_3_lut_21493_rep_271_4_lut.init = 16'h8f80;
    LUT4 mux_194_Mux_3_i189_3_lut_3_lut_4_lut (.A(n24891), .B(index_i[3]), 
         .C(index_i[4]), .D(n24925), .Z(n189_adj_2824)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_3_i189_3_lut_3_lut_4_lut.init = 16'h08f8;
    LUT4 i11037_3_lut_4_lut (.A(n24951), .B(index_i[4]), .C(index_i[5]), 
         .D(index_i[6]), .Z(n127)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11037_3_lut_4_lut.init = 16'hf800;
    LUT4 n396_bdd_3_lut_22953 (.A(n27502), .B(n25137), .C(index_i[3]), 
         .Z(n23677)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n396_bdd_3_lut_22953.init = 16'hcaca;
    LUT4 i19334_3_lut_3_lut_4_lut (.A(n24951), .B(index_i[4]), .C(n125), 
         .D(index_i[5]), .Z(n21664)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19334_3_lut_3_lut_4_lut.init = 16'hf077;
    LUT4 n123_bdd_3_lut_22091 (.A(n25152), .B(n404), .C(index_i[3]), .Z(n23693)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n123_bdd_3_lut_22091.init = 16'hacac;
    LUT4 n123_bdd_3_lut_22939 (.A(n27504), .B(n27505), .C(index_i[3]), 
         .Z(n23694)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n123_bdd_3_lut_22939.init = 16'hcaca;
    LUT4 n452_bdd_3_lut_22285 (.A(n25143), .B(n27500), .C(index_i[3]), 
         .Z(n23697)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n452_bdd_3_lut_22285.init = 16'hcaca;
    LUT4 i19312_3_lut (.A(n25144), .B(n25139), .C(index_i[3]), .Z(n21642)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19312_3_lut.init = 16'hcaca;
    LUT4 i19311_3_lut (.A(n325), .B(n332), .C(index_i[3]), .Z(n21641)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19311_3_lut.init = 16'hcaca;
    LUT4 mux_191_i16_3_lut (.A(\quarter_wave_sample_register_q[15] ), .B(o_val_pipeline_i_0__15__N_2157[15]), 
         .C(phase_negation_i[1]), .Z(n1205[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam mux_191_i16_3_lut.init = 16'hcaca;
    LUT4 mux_191_i15_3_lut (.A(quarter_wave_sample_register_i[14]), .B(o_val_pipeline_i_0__15__N_2157[14]), 
         .C(phase_negation_i[1]), .Z(n1205[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam mux_191_i15_3_lut.init = 16'hcaca;
    LUT4 i17845_3_lut (.A(n20170), .B(n20171), .C(index_i[7]), .Z(n20175)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17845_3_lut.init = 16'hcaca;
    LUT4 n77_bdd_3_lut_22104 (.A(n25153), .B(n27505), .C(index_i[3]), 
         .Z(n23705)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n77_bdd_3_lut_22104.init = 16'hacac;
    LUT4 n20087_bdd_3_lut (.A(n25099), .B(n25150), .C(index_i[3]), .Z(n23714)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n20087_bdd_3_lut.init = 16'hcaca;
    PFUMX i23043 (.BLUT(n25275), .ALUT(n25276), .C0(index_i[1]), .Z(n25277));
    LUT4 i19305_3_lut (.A(n27515), .B(n25131), .C(index_i[3]), .Z(n21635)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19305_3_lut.init = 16'hcaca;
    LUT4 i20414_3_lut (.A(n21635), .B(n21636), .C(index_i[4]), .Z(n21637)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20414_3_lut.init = 16'hcaca;
    LUT4 i19287_3_lut (.A(n1001), .B(n588), .C(index_i[3]), .Z(n21617)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19287_3_lut.init = 16'hcaca;
    LUT4 n22970_bdd_3_lut_4_lut (.A(n24831), .B(index_i[6]), .C(index_i[5]), 
         .D(n22970), .Z(n22971)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam n22970_bdd_3_lut_4_lut.init = 16'hefe0;
    LUT4 i20416_3_lut (.A(n21617), .B(n21618), .C(index_i[4]), .Z(n21619)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20416_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_10_i252_3_lut_4_lut_4_lut (.A(n24978), .B(index_i[3]), 
         .C(index_i[4]), .D(n24952), .Z(n252_adj_2825)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B (C (D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_10_i252_3_lut_4_lut_4_lut.init = 16'h3efe;
    LUT4 n348_bdd_3_lut_4_lut (.A(n24978), .B(index_i[3]), .C(index_i[5]), 
         .D(n23816), .Z(n24800)) /* synthesis lut_function=(!(A (C+!(D))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n348_bdd_3_lut_4_lut.init = 16'h1f10;
    LUT4 mux_194_Mux_10_i413_3_lut_4_lut (.A(n24978), .B(index_i[3]), .C(index_i[4]), 
         .D(n24925), .Z(n413)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_10_i413_3_lut_4_lut.init = 16'hf101;
    PFUMX i18264 (.BLUT(n574_adj_2826), .ALUT(n637), .C0(index_i[6]), 
          .Z(n20594));
    LUT4 mux_194_Mux_3_i828_3_lut_3_lut_4_lut (.A(n24978), .B(index_i[3]), 
         .C(n157), .D(index_i[4]), .Z(n828)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_3_i828_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 i18329_3_lut_3_lut_4_lut (.A(n24978), .B(index_i[3]), .C(n412), 
         .D(index_i[4]), .Z(n20659)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18329_3_lut_3_lut_4_lut.init = 16'hf011;
    PFUMX i18261 (.BLUT(n318), .ALUT(n381), .C0(index_i[6]), .Z(n20591));
    LUT4 n22_bdd_3_lut_22134 (.A(n25136), .B(n25153), .C(index_i[3]), 
         .Z(n23737)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n22_bdd_3_lut_22134.init = 16'hcaca;
    LUT4 i19248_3_lut (.A(n25121), .B(n25152), .C(index_i[3]), .Z(n21578)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19248_3_lut.init = 16'hcaca;
    LUT4 i12251_1_lut_2_lut_3_lut_4_lut (.A(n24978), .B(index_i[3]), .C(index_i[5]), 
         .D(index_i[4]), .Z(n381)) /* synthesis lut_function=(!(A (C+(D))+!A (B (C+(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i12251_1_lut_2_lut_3_lut_4_lut.init = 16'h010f;
    PFUMX i18249 (.BLUT(n127), .ALUT(n254_adj_2827), .C0(index_i[7]), 
          .Z(n20579));
    LUT4 i17814_3_lut (.A(n20139), .B(n23108), .C(index_i[7]), .Z(n20144)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17814_3_lut.init = 16'hcaca;
    LUT4 i19336_3_lut_3_lut_4_lut (.A(n24961), .B(index_i[4]), .C(n252_adj_2825), 
         .D(index_i[5]), .Z(n21666)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19336_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 i17813_3_lut (.A(n20137), .B(n20138), .C(index_i[7]), .Z(n20143)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17813_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_10_i701_4_lut_4_lut (.A(n24961), .B(index_i[4]), .C(index_i[5]), 
         .D(n24869), .Z(n701)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B (C (D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_10_i701_4_lut_4_lut.init = 16'h3efe;
    LUT4 mux_194_Mux_7_i956_3_lut_3_lut_4_lut (.A(n24961), .B(index_i[4]), 
         .C(n924_adj_2828), .D(index_i[5]), .Z(n956)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_7_i956_3_lut_3_lut_4_lut.init = 16'h11f0;
    LUT4 i20947_3_lut (.A(n20143), .B(n20144), .C(index_i[8]), .Z(n20146)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20947_3_lut.init = 16'hcaca;
    LUT4 i19415_3_lut (.A(n21742), .B(n21743), .C(index_i[7]), .Z(n21745)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19415_3_lut.init = 16'hcaca;
    LUT4 i19414_3_lut (.A(n21740), .B(n21741), .C(index_i[7]), .Z(n21744)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19414_3_lut.init = 16'hcaca;
    LUT4 i3_3_lut_4_lut (.A(n24960), .B(index_i[4]), .C(index_i[6]), .D(index_i[5]), 
         .Z(n17787)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i3_3_lut_4_lut.init = 16'hfffe;
    LUT4 mux_194_Mux_0_i526_3_lut (.A(n25144), .B(n25121), .C(index_i[3]), 
         .Z(n526)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_0_i526_3_lut.init = 16'hcaca;
    LUT4 i19321_3_lut_4_lut_4_lut (.A(n24960), .B(index_i[4]), .C(index_i[5]), 
         .D(n24878), .Z(n21651)) /* synthesis lut_function=(A ((C+!(D))+!B)+!A (B (C+!(D))+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19321_3_lut_4_lut_4_lut.init = 16'he3ef;
    LUT4 mux_191_i14_3_lut (.A(quarter_wave_sample_register_i[13]), .B(o_val_pipeline_i_0__15__N_2157[13]), 
         .C(phase_negation_i[1]), .Z(n1205[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam mux_191_i14_3_lut.init = 16'hcaca;
    LUT4 mux_191_i13_3_lut (.A(quarter_wave_sample_register_i[12]), .B(o_val_pipeline_i_0__15__N_2157[12]), 
         .C(phase_negation_i[1]), .Z(n1205[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam mux_191_i13_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_2_i284_3_lut_4_lut_3_lut_rep_660 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27500)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_2_i284_3_lut_4_lut_3_lut_rep_660.init = 16'h4d4d;
    LUT4 mux_194_Mux_3_i653_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n653_adj_2829)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A !(B (D)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_3_i653_3_lut_4_lut_4_lut.init = 16'h4d99;
    LUT4 mux_191_i12_3_lut (.A(quarter_wave_sample_register_i[11]), .B(o_val_pipeline_i_0__15__N_2157[11]), 
         .C(phase_negation_i[1]), .Z(n1205[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam mux_191_i12_3_lut.init = 16'hcaca;
    LUT4 mux_191_i11_3_lut (.A(quarter_wave_sample_register_i[10]), .B(o_val_pipeline_i_0__15__N_2157[10]), 
         .C(phase_negation_i[1]), .Z(n1205[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam mux_191_i11_3_lut.init = 16'hcaca;
    LUT4 mux_191_i10_3_lut (.A(quarter_wave_sample_register_i[9]), .B(o_val_pipeline_i_0__15__N_2157[9]), 
         .C(phase_negation_i[1]), .Z(n1205[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam mux_191_i10_3_lut.init = 16'hcaca;
    LUT4 mux_191_i9_3_lut (.A(quarter_wave_sample_register_i[8]), .B(o_val_pipeline_i_0__15__N_2157[8]), 
         .C(phase_negation_i[1]), .Z(n1205[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam mux_191_i9_3_lut.init = 16'hcaca;
    LUT4 mux_191_i8_3_lut (.A(quarter_wave_sample_register_i[7]), .B(o_val_pipeline_i_0__15__N_2157[7]), 
         .C(phase_negation_i[1]), .Z(n1205[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam mux_191_i8_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_0_i363_3_lut_4_lut_3_lut_rep_661 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27501)) /* synthesis lut_function=(A (B+!(C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_0_i363_3_lut_4_lut_3_lut_rep_661.init = 16'hdbdb;
    PFUMX i18697 (.BLUT(n142), .ALUT(n157_adj_2830), .C0(index_i[4]), 
          .Z(n21027));
    LUT4 i20952_3_lut_4_lut (.A(n25004), .B(n24893), .C(index_i[8]), .D(n766), 
         .Z(n20090)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20952_3_lut_4_lut.init = 16'hefe0;
    LUT4 mux_191_i7_3_lut (.A(quarter_wave_sample_register_i[6]), .B(o_val_pipeline_i_0__15__N_2157[6]), 
         .C(phase_negation_i[1]), .Z(n1205[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam mux_191_i7_3_lut.init = 16'hcaca;
    LUT4 mux_191_i6_3_lut (.A(quarter_wave_sample_register_i[5]), .B(o_val_pipeline_i_0__15__N_2157[5]), 
         .C(phase_negation_i[1]), .Z(n1205[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam mux_191_i6_3_lut.init = 16'hcaca;
    LUT4 mux_191_i5_3_lut (.A(quarter_wave_sample_register_i[4]), .B(o_val_pipeline_i_0__15__N_2157[4]), 
         .C(phase_negation_i[1]), .Z(n1205[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam mux_191_i5_3_lut.init = 16'hcaca;
    LUT4 mux_191_i4_3_lut (.A(quarter_wave_sample_register_i[3]), .B(o_val_pipeline_i_0__15__N_2157[3]), 
         .C(phase_negation_i[1]), .Z(n1205[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam mux_191_i4_3_lut.init = 16'hcaca;
    LUT4 mux_191_i3_3_lut (.A(quarter_wave_sample_register_i[2]), .B(o_val_pipeline_i_0__15__N_2157[2]), 
         .C(phase_negation_i[1]), .Z(n1205[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam mux_191_i3_3_lut.init = 16'hcaca;
    LUT4 mux_191_i2_3_lut (.A(quarter_wave_sample_register_i[1]), .B(o_val_pipeline_i_0__15__N_2157[1]), 
         .C(phase_negation_i[1]), .Z(n1205[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam mux_191_i2_3_lut.init = 16'hcaca;
    LUT4 mux_191_i1_3_lut (.A(quarter_wave_sample_register_i[0]), .B(o_val_pipeline_i_0__15__N_2157[0]), 
         .C(phase_negation_i[1]), .Z(n1205[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam mux_191_i1_3_lut.init = 16'hcaca;
    PFUMX i23041 (.BLUT(n25272), .ALUT(n25273), .C0(index_i[2]), .Z(n25274));
    PFUMX i18698 (.BLUT(n173), .ALUT(n188), .C0(index_i[4]), .Z(n21028));
    LUT4 mux_194_Mux_11_i766_3_lut (.A(n638), .B(n765), .C(index_i[7]), 
         .Z(n766)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_11_i766_3_lut.init = 16'h3a3a;
    LUT4 mux_194_Mux_1_i987_3_lut_4_lut (.A(n24995), .B(index_i[3]), .C(index_i[4]), 
         .D(n986_adj_2831), .Z(n987)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_1_i987_3_lut_4_lut.init = 16'hf202;
    PFUMX i18703 (.BLUT(n333), .ALUT(n348_adj_2832), .C0(index_i[4]), 
          .Z(n21033));
    LUT4 index_i_5__bdd_4_lut_23805 (.A(n85), .B(index_i[2]), .C(index_i[3]), 
         .D(n25098), .Z(n23813)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (B+!(C (D))))) */ ;
    defparam index_i_5__bdd_4_lut_23805.init = 16'h3a0a;
    LUT4 i11104_3_lut_4_lut (.A(n24805), .B(index_i[7]), .C(index_i[8]), 
         .D(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2126[14])) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11104_3_lut_4_lut.init = 16'hffe0;
    LUT4 i6361_2_lut (.A(phase_i[0]), .B(phase_i[10]), .Z(index_i_9__N_2106[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i6361_2_lut.init = 16'h6666;
    PFUMX i18704 (.BLUT(n364_adj_2833), .ALUT(n379), .C0(index_i[4]), 
          .Z(n21034));
    LUT4 n348_bdd_3_lut_22718 (.A(n25125), .B(n27505), .C(index_i[3]), 
         .Z(n23816)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n348_bdd_3_lut_22718.init = 16'hcaca;
    PFUMX i18705 (.BLUT(n397), .ALUT(n412_adj_2817), .C0(index_i[4]), 
          .Z(n21035));
    LUT4 i6362_2_lut (.A(phase_i[9]), .B(phase_i[10]), .Z(index_i_9__N_2106[9])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i6362_2_lut.init = 16'h6666;
    LUT4 i6363_2_lut (.A(phase_i[8]), .B(phase_i[10]), .Z(index_i_9__N_2106[8])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i6363_2_lut.init = 16'h6666;
    LUT4 i6364_2_lut (.A(phase_i[7]), .B(phase_i[10]), .Z(index_i_9__N_2106[7])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i6364_2_lut.init = 16'h6666;
    LUT4 i6365_2_lut (.A(phase_i[6]), .B(phase_i[10]), .Z(index_i_9__N_2106[6])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i6365_2_lut.init = 16'h6666;
    PFUMX i18706 (.BLUT(n428), .ALUT(n443_adj_2812), .C0(index_i[4]), 
          .Z(n21036));
    LUT4 i6366_2_lut (.A(phase_i[5]), .B(phase_i[10]), .Z(index_i_9__N_2106[5])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i6366_2_lut.init = 16'h6666;
    LUT4 i6367_2_lut (.A(phase_i[4]), .B(phase_i[10]), .Z(index_i_9__N_2106[4])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i6367_2_lut.init = 16'h6666;
    PFUMX i18707 (.BLUT(n460), .ALUT(n475), .C0(index_i[4]), .Z(n21037));
    PFUMX i18708 (.BLUT(n491_adj_2834), .ALUT(n11113), .C0(index_i[4]), 
          .Z(n21038));
    LUT4 i6368_2_lut (.A(phase_i[3]), .B(phase_i[10]), .Z(index_i_9__N_2106[3])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i6368_2_lut.init = 16'h6666;
    LUT4 i6369_2_lut (.A(phase_i[2]), .B(phase_i[10]), .Z(index_i_9__N_2106[2])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i6369_2_lut.init = 16'h6666;
    LUT4 i6370_2_lut (.A(phase_i[1]), .B(phase_i[10]), .Z(index_i_9__N_2106[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i6370_2_lut.init = 16'h6666;
    LUT4 n22_bdd_3_lut_23228 (.A(n27508), .B(n25138), .C(index_i[3]), 
         .Z(n23825)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n22_bdd_3_lut_23228.init = 16'hacac;
    LUT4 i9596_3_lut_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n12166)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A !(B (C+(D))+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9596_3_lut_3_lut_4_lut_4_lut.init = 16'h44db;
    LUT4 n572_bdd_3_lut_22842 (.A(n588), .B(n25125), .C(index_i[3]), .Z(n23827)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n572_bdd_3_lut_22842.init = 16'hcaca;
    LUT4 mux_194_Mux_4_i491_3_lut_4_lut (.A(n24994), .B(index_i[2]), .C(index_i[3]), 
         .D(n27510), .Z(n491)) /* synthesis lut_function=(A (C+(D))+!A !(B (C+!(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_4_i491_3_lut_4_lut.init = 16'hbfb0;
    LUT4 i17645_3_lut (.A(n900), .B(n25152), .C(index_i[3]), .Z(n19975)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17645_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_9_i124_3_lut_3_lut_4_lut (.A(index_i[0]), .B(n24997), 
         .C(index_i[3]), .D(n24952), .Z(n124)) /* synthesis lut_function=(!(A (C (D))+!A (B (C (D))+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_9_i124_3_lut_3_lut_4_lut.init = 16'h0efe;
    LUT4 mux_194_Mux_0_i572_3_lut_4_lut (.A(index_i[0]), .B(n24997), .C(index_i[3]), 
         .D(n27505), .Z(n572)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_0_i572_3_lut_4_lut.init = 16'hefe0;
    LUT4 mux_194_Mux_9_i364_3_lut_3_lut_4_lut (.A(index_i[0]), .B(n24997), 
         .C(index_i[3]), .D(n24978), .Z(n364)) /* synthesis lut_function=(!(A (C (D))+!A (B (C (D))+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_9_i364_3_lut_3_lut_4_lut.init = 16'h0efe;
    LUT4 mux_194_Mux_3_i251_3_lut_4_lut (.A(index_i[0]), .B(n24997), .C(index_i[3]), 
         .D(n24978), .Z(n14964)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_3_i251_3_lut_4_lut.init = 16'hfe0e;
    LUT4 i9377_3_lut_4_lut (.A(index_i[0]), .B(n24997), .C(index_i[3]), 
         .D(index_i[4]), .Z(n11943)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9377_3_lut_4_lut.init = 16'h0e1e;
    LUT4 mux_194_Mux_8_i475_3_lut_3_lut_4_lut (.A(index_i[0]), .B(n24997), 
         .C(index_i[3]), .D(n24952), .Z(n475_adj_2835)) /* synthesis lut_function=(A (C+!(D))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_8_i475_3_lut_3_lut_4_lut.init = 16'he0ef;
    LUT4 i20433_3_lut (.A(n25283), .B(n19973), .C(index_i[4]), .Z(n19974)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20433_3_lut.init = 16'hcaca;
    LUT4 n557_bdd_3_lut_21487_3_lut_4_lut (.A(index_i[0]), .B(n24997), .C(index_i[4]), 
         .D(index_i[3]), .Z(n23029)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n557_bdd_3_lut_21487_3_lut_4_lut.init = 16'hf10f;
    LUT4 i18431_4_lut_4_lut_3_lut_4_lut (.A(index_i[0]), .B(n24997), .C(index_i[4]), 
         .D(index_i[3]), .Z(n20761)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18431_4_lut_4_lut_3_lut_4_lut.init = 16'h11ef;
    PFUMX i9374 (.BLUT(n12159), .ALUT(n12160), .C0(n25029), .Z(n11940));
    LUT4 i11053_2_lut_rep_267_3_lut_4_lut (.A(index_i[0]), .B(n24997), .C(index_i[4]), 
         .D(index_i[3]), .Z(n24827)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11053_2_lut_rep_267_3_lut_4_lut.init = 16'hfef0;
    LUT4 mux_194_Mux_8_i653_3_lut_rep_283_4_lut (.A(index_i[0]), .B(n24998), 
         .C(index_i[3]), .D(n24978), .Z(n24843)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(C+(D)))) */ ;
    defparam mux_194_Mux_8_i653_3_lut_rep_283_4_lut.init = 16'h7f70;
    LUT4 i17636_3_lut (.A(n404), .B(n25137), .C(index_i[3]), .Z(n19966)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17636_3_lut.init = 16'hcaca;
    LUT4 i20238_3_lut (.A(n19966), .B(n19967), .C(index_i[4]), .Z(n19968)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20238_3_lut.init = 16'hcaca;
    L6MUX21 i19254 (.D0(n21333), .D1(n21336), .SD(index_i[5]), .Z(n21584));
    PFUMX i23039 (.BLUT(n25269), .ALUT(n25270), .C0(index_i[0]), .Z(n25271));
    LUT4 i17631_3_lut (.A(n404), .B(n27500), .C(index_i[3]), .Z(n19961)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17631_3_lut.init = 16'hcaca;
    L6MUX21 i19258 (.D0(n21643), .D1(n17553), .SD(index_i[5]), .Z(n21588));
    L6MUX21 i19259 (.D0(n21709), .D1(n11952), .SD(index_i[5]), .Z(n21589));
    LUT4 i20244_3_lut (.A(n19957), .B(n19958), .C(index_i[4]), .Z(n19959)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20244_3_lut.init = 16'hcaca;
    LUT4 n1018_bdd_4_lut_4_lut_4_lut (.A(index_i[0]), .B(n24998), .C(index_i[4]), 
         .D(index_i[3]), .Z(n23104)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (D))+!A (B (C (D)+!C !(D))+!B (D)))) */ ;
    defparam n1018_bdd_4_lut_4_lut_4_lut.init = 16'h0c73;
    LUT4 i17625_3_lut (.A(n27500), .B(n25120), .C(index_i[3]), .Z(n19955)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17625_3_lut.init = 16'hcaca;
    LUT4 i17909_3_lut (.A(n20236), .B(n20237), .C(index_i[8]), .Z(n20239)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17909_3_lut.init = 16'hcaca;
    LUT4 i17908_3_lut (.A(n20234), .B(n20235), .C(index_i[8]), .Z(n20238)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17908_3_lut.init = 16'hcaca;
    LUT4 i20246_3_lut (.A(n19954), .B(n19955), .C(index_i[4]), .Z(n19956)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20246_3_lut.init = 16'hcaca;
    LUT4 i20249_3_lut (.A(n19951), .B(n19952), .C(index_i[4]), .Z(n19953)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20249_3_lut.init = 16'hcaca;
    LUT4 i11058_3_lut_4_lut (.A(index_i[0]), .B(n24998), .C(n25092), .D(index_i[5]), 
         .Z(n318)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (C (D))) */ ;
    defparam i11058_3_lut_4_lut.init = 16'hf800;
    LUT4 i17878_3_lut (.A(n20205), .B(n20206), .C(index_i[8]), .Z(n20208)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17878_3_lut.init = 16'hcaca;
    LUT4 i17877_3_lut (.A(n20203), .B(n20204), .C(index_i[8]), .Z(n20207)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17877_3_lut.init = 16'hcaca;
    LUT4 i18434_3_lut_4_lut (.A(n24978), .B(n24892), .C(index_i[3]), .D(index_i[4]), 
         .Z(n20764)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C (D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18434_3_lut_4_lut.init = 16'hf03a;
    PFUMX i19261 (.BLUT(n542), .ALUT(n573), .C0(index_i[5]), .Z(n21591));
    PFUMX i19262 (.BLUT(n605), .ALUT(n636), .C0(index_i[5]), .Z(n21592));
    LUT4 mux_194_Mux_0_i396_3_lut_4_lut_3_lut_rep_662 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27502)) /* synthesis lut_function=(A ((C)+!B)+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_0_i396_3_lut_4_lut_3_lut_rep_662.init = 16'hb6b6;
    LUT4 mux_194_Mux_10_i893_3_lut_4_lut (.A(n25094), .B(index_i[5]), .C(index_i[6]), 
         .D(n892), .Z(n893)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_10_i893_3_lut_4_lut.init = 16'hf101;
    LUT4 mux_194_Mux_1_i301_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n301)) /* synthesis lut_function=(A (B (C+(D))+!B !(D))+!A !(B (C+(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_1_i301_3_lut_4_lut_4_lut.init = 16'h99b6;
    PFUMX i19263 (.BLUT(n669), .ALUT(n700), .C0(index_i[5]), .Z(n21593));
    LUT4 i20732_3_lut_4_lut (.A(n25093), .B(index_i[4]), .C(index_i[5]), 
         .D(n62_adj_2822), .Z(n21663)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20732_3_lut_4_lut.init = 16'hf808;
    LUT4 i17613_3_lut (.A(n325), .B(n25152), .C(index_i[3]), .Z(n19943)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17613_3_lut.init = 16'hcaca;
    PFUMX i19264 (.BLUT(n732_adj_2836), .ALUT(n21715), .C0(index_i[5]), 
          .Z(n21594));
    PFUMX i19265 (.BLUT(n797), .ALUT(n828_adj_2837), .C0(index_i[5]), 
          .Z(n21595));
    LUT4 i20269_3_lut (.A(n19942), .B(n19943), .C(index_i[4]), .Z(n19944)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20269_3_lut.init = 16'hcaca;
    PFUMX i19266 (.BLUT(n860_adj_2838), .ALUT(n891_adj_2839), .C0(index_i[5]), 
          .Z(n21596));
    LUT4 i17815_3_lut (.A(n20141), .B(n20142), .C(index_i[8]), .Z(n20145)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17815_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_13_i511_4_lut_4_lut (.A(n24805), .B(index_i[7]), .C(index_i[8]), 
         .D(n254), .Z(n511)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (B (C+!(D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_13_i511_4_lut_4_lut.init = 16'h1c10;
    PFUMX i18262 (.BLUT(n445), .ALUT(n508), .C0(index_i[6]), .Z(n20592));
    LUT4 mux_194_Mux_8_i542_3_lut_4_lut (.A(n24997), .B(index_i[3]), .C(index_i[4]), 
         .D(n526_adj_2840), .Z(n542_adj_2841)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_8_i542_3_lut_4_lut.init = 16'h6f60;
    LUT4 i18432_3_lut_4_lut (.A(n24997), .B(index_i[3]), .C(index_i[4]), 
         .D(n635_adj_2806), .Z(n20762)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18432_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_194_Mux_6_i732_3_lut_4_lut (.A(n25099), .B(index_i[3]), .C(index_i[4]), 
         .D(n731_adj_2842), .Z(n732_adj_2836)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_6_i732_3_lut_4_lut.init = 16'hf909;
    PFUMX i18274 (.BLUT(n94), .ALUT(n19974), .C0(index_i[5]), .Z(n20604));
    LUT4 i17610_3_lut (.A(n25148), .B(n27502), .C(index_i[3]), .Z(n19940)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17610_3_lut.init = 16'hcaca;
    LUT4 n699_bdd_4_lut_22658 (.A(n24869), .B(index_i[6]), .C(n24960), 
         .D(index_i[5]), .Z(n23033)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C+!(D))+!B (D))) */ ;
    defparam n699_bdd_4_lut_22658.init = 16'hd1cc;
    L6MUX21 i18275 (.D0(n19977), .D1(n19995), .SD(index_i[5]), .Z(n20605));
    LUT4 n23036_bdd_3_lut (.A(n23036), .B(n23033), .C(index_i[4]), .Z(n23037)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n23036_bdd_3_lut.init = 16'hcaca;
    LUT4 i20278_3_lut (.A(n19936), .B(n19937), .C(index_i[4]), .Z(n19938)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20278_3_lut.init = 16'hcaca;
    LUT4 i17759_3_lut (.A(n22797), .B(n20593), .C(index_i[8]), .Z(n20089)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17759_3_lut.init = 16'hcaca;
    PFUMX i18277 (.BLUT(n20070), .ALUT(n317_adj_2815), .C0(index_i[5]), 
          .Z(n20607));
    PFUMX i18278 (.BLUT(n349), .ALUT(n20073), .C0(index_i[5]), .Z(n20608));
    LUT4 i19303_3_lut (.A(n21630), .B(n21631), .C(index_i[8]), .Z(n21633)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19303_3_lut.init = 16'hcaca;
    LUT4 i19302_3_lut (.A(n21628), .B(n21629), .C(index_i[8]), .Z(n21632)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19302_3_lut.init = 16'hcaca;
    L6MUX21 i18279 (.D0(n20076), .D1(n20079), .SD(index_i[5]), .Z(n20609));
    L6MUX21 i18280 (.D0(n20082), .D1(n20085), .SD(index_i[5]), .Z(n20610));
    LUT4 i17601_3_lut (.A(n27501), .B(n27515), .C(index_i[3]), .Z(n19931)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17601_3_lut.init = 16'hcaca;
    LUT4 i17600_3_lut (.A(n27505), .B(n25151), .C(index_i[3]), .Z(n19930)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17600_3_lut.init = 16'hcaca;
    LUT4 i20285_3_lut (.A(n19930), .B(n19931), .C(index_i[4]), .Z(n19932)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20285_3_lut.init = 16'hcaca;
    PFUMX i15290 (.BLUT(n17551), .ALUT(n17552), .C0(index_i[4]), .Z(n17553));
    L6MUX21 i18282 (.D0(n21570), .D1(n636_adj_2843), .SD(index_i[5]), 
            .Z(n20612));
    PFUMX i18283 (.BLUT(n21573), .ALUT(n700_adj_2844), .C0(index_i[5]), 
          .Z(n20613));
    LUT4 i17598_3_lut (.A(n27508), .B(n25141), .C(index_i[3]), .Z(n19928)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17598_3_lut.init = 16'hcaca;
    LUT4 i17597_3_lut (.A(n25099), .B(n85), .C(index_i[3]), .Z(n19927)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17597_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_6_i700_3_lut_4_lut (.A(n25099), .B(index_i[3]), .C(index_i[4]), 
         .D(n684_adj_2845), .Z(n700)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_6_i700_3_lut_4_lut.init = 16'h9f90;
    L6MUX21 i18285 (.D0(n21579), .D1(n21582), .SD(index_i[5]), .Z(n20615));
    LUT4 i20287_3_lut (.A(n19927), .B(n19928), .C(index_i[4]), .Z(n19929)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20287_3_lut.init = 16'hcaca;
    PFUMX i18287 (.BLUT(n924), .ALUT(n21619), .C0(index_i[5]), .Z(n20617));
    PFUMX i18288 (.BLUT(n987), .ALUT(n21637), .C0(index_i[5]), .Z(n20618));
    LUT4 mux_194_Mux_1_i700_3_lut_4_lut (.A(n25027), .B(index_i[3]), .C(index_i[4]), 
         .D(n684_adj_2818), .Z(n700_adj_2844)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_1_i700_3_lut_4_lut.init = 16'hefe0;
    LUT4 i9404_3_lut_4_lut (.A(n24976), .B(index_i[2]), .C(n25094), .D(n25149), 
         .Z(n444)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9404_3_lut_4_lut.init = 16'h6f60;
    LUT4 i18302_3_lut (.A(n20629), .B(n20630), .C(index_i[8]), .Z(n20632)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18302_3_lut.init = 16'hcaca;
    LUT4 n26428_bdd_3_lut (.A(n26428), .B(index_i[1]), .C(index_i[4]), 
         .Z(n26429)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n26428_bdd_3_lut.init = 16'hcaca;
    LUT4 i18301_3_lut (.A(n20627), .B(n20628), .C(index_i[8]), .Z(n20631)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18301_3_lut.init = 16'hcaca;
    LUT4 index_i_1__bdd_4_lut (.A(index_i[1]), .B(index_i[3]), .C(index_i[0]), 
         .D(index_i[2]), .Z(n26428)) /* synthesis lut_function=(A (B (C+(D))+!B (C (D)))+!A !(B (C)+!B !(C+(D)))) */ ;
    defparam index_i_1__bdd_4_lut.init = 16'hbd94;
    L6MUX21 i19402 (.D0(n21716), .D1(n21717), .SD(index_i[5]), .Z(n21732));
    L6MUX21 i19403 (.D0(n21718), .D1(n21719), .SD(index_i[5]), .Z(n21733));
    L6MUX21 i19404 (.D0(n21720), .D1(n21721), .SD(index_i[5]), .Z(n21734));
    L6MUX21 i19405 (.D0(n21722), .D1(n21723), .SD(index_i[5]), .Z(n21735));
    L6MUX21 i19406 (.D0(n21724), .D1(n21725), .SD(index_i[5]), .Z(n21736));
    L6MUX21 i19407 (.D0(n21726), .D1(n21727), .SD(index_i[5]), .Z(n21737));
    L6MUX21 i19408 (.D0(n21728), .D1(n21729), .SD(index_i[5]), .Z(n21738));
    L6MUX21 i19409 (.D0(n21730), .D1(n21731), .SD(index_i[5]), .Z(n21739));
    PFUMX i18326 (.BLUT(n20652), .ALUT(n20653), .C0(index_i[5]), .Z(n20656));
    PFUMX i18327 (.BLUT(n20654), .ALUT(n20655), .C0(index_i[5]), .Z(n20657));
    PFUMX i18333 (.BLUT(n20659), .ALUT(n20660), .C0(index_i[5]), .Z(n20663));
    PFUMX i18334 (.BLUT(n20661), .ALUT(n20662), .C0(index_i[5]), .Z(n20664));
    LUT4 n22784_bdd_3_lut (.A(n22784), .B(n157_adj_2846), .C(index_i[4]), 
         .Z(n22785)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n22784_bdd_3_lut.init = 16'hcaca;
    PFUMX i17779 (.BLUT(n956), .ALUT(n17674), .C0(index_i[6]), .Z(n20109));
    LUT4 mux_194_Mux_6_i251_3_lut_4_lut (.A(n24976), .B(index_i[2]), .C(index_i[3]), 
         .D(n25149), .Z(n251_adj_2847)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_6_i251_3_lut_4_lut.init = 16'hf606;
    LUT4 index_i_2__bdd_4_lut (.A(index_i[2]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[0]), .Z(n27527)) /* synthesis lut_function=(A (B ((D)+!C))+!A !(B+!(C+!(D)))) */ ;
    defparam index_i_2__bdd_4_lut.init = 16'h9819;
    LUT4 mux_194_Mux_4_i747_3_lut_4_lut (.A(n24976), .B(index_i[2]), .C(index_i[3]), 
         .D(n27502), .Z(n747_adj_2848)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_4_i747_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_194_Mux_8_i732_3_lut (.A(index_i[3]), .B(n14960), .C(index_i[5]), 
         .Z(n732_adj_2849)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_8_i732_3_lut.init = 16'h3a3a;
    PFUMX i17788 (.BLUT(n94_adj_2850), .ALUT(n125_adj_2851), .C0(index_i[5]), 
          .Z(n20118));
    LUT4 i19467_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21797)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A (B (C (D)+!C !(D))+!B (D))) */ ;
    defparam i19467_3_lut_4_lut.init = 16'hd926;
    PFUMX i17789 (.BLUT(n17544), .ALUT(n14348), .C0(index_i[5]), .Z(n20119));
    LUT4 n347_bdd_3_lut_22949_4_lut (.A(n25129), .B(index_i[2]), .C(index_i[3]), 
         .D(n25125), .Z(n23675)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n347_bdd_3_lut_22949_4_lut.init = 16'hf606;
    LUT4 mux_194_Mux_3_i890_3_lut_4_lut (.A(n25129), .B(index_i[2]), .C(index_i[3]), 
         .D(n325), .Z(n890_adj_2852)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_3_i890_3_lut_4_lut.init = 16'h6f60;
    LUT4 i19002_3_lut_4_lut (.A(n25129), .B(index_i[2]), .C(index_i[3]), 
         .D(n25153), .Z(n21332)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19002_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_194_Mux_0_i348_3_lut_4_lut (.A(n25129), .B(index_i[2]), .C(index_i[3]), 
         .D(n25107), .Z(n348_adj_2832)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_0_i348_3_lut_4_lut.init = 16'h6f60;
    PFUMX i23037 (.BLUT(n25266), .ALUT(n25267), .C0(index_i[1]), .Z(n25268));
    L6MUX21 i17791 (.D0(n21752), .D1(n21755), .SD(index_i[5]), .Z(n20121));
    LUT4 mux_194_Mux_2_i955_then_4_lut (.A(index_i[4]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n25249)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B (C+!(D))+!B !(C (D)))) */ ;
    defparam mux_194_Mux_2_i955_then_4_lut.init = 16'he95d;
    LUT4 mux_194_Mux_0_i123_3_lut_3_lut_rep_664 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27504)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_0_i123_3_lut_3_lut_rep_664.init = 16'h6c6c;
    PFUMX i23143 (.BLUT(n25436), .ALUT(n25431), .C0(index_i[3]), .Z(n25437));
    LUT4 mux_194_Mux_0_i684_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n684_adj_2798)) /* synthesis lut_function=(!(A ((D)+!B)+!A !(B (D)+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_0_i684_3_lut_4_lut_4_lut.init = 16'h5498;
    LUT4 mux_194_Mux_5_i31_3_lut (.A(n15), .B(n30), .C(index_i[4]), .Z(n31)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_5_i31_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_4_i62_4_lut (.A(n24999), .B(n61), .C(index_i[4]), 
         .D(index_i[3]), .Z(n62_adj_2853)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_4_i62_4_lut.init = 16'hc5ca;
    LUT4 mux_194_Mux_4_i31_4_lut (.A(n15_adj_2854), .B(n24841), .C(index_i[4]), 
         .D(index_i[3]), .Z(n31_adj_2855)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_4_i31_4_lut.init = 16'h3aca;
    L6MUX21 i17792 (.D0(n21789), .D1(n21792), .SD(index_i[5]), .Z(n20122));
    PFUMX mux_194_Mux_1_i636 (.BLUT(n620_adj_2856), .ALUT(n635_adj_2857), 
          .C0(index_i[4]), .Z(n636_adj_2843)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    PFUMX i17793 (.BLUT(n413_adj_2858), .ALUT(n444), .C0(index_i[5]), 
          .Z(n20123));
    LUT4 mux_194_Mux_3_i31_3_lut (.A(n781_adj_2805), .B(n30_adj_2859), .C(index_i[4]), 
         .Z(n31_adj_2860)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_3_i31_3_lut.init = 16'hcaca;
    LUT4 index_i_6__bdd_4_lut_24346 (.A(index_i[6]), .B(index_i[5]), .C(index_i[1]), 
         .D(index_i[0]), .Z(n26967)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C))+!A (B (C)+!B !(C)))) */ ;
    defparam index_i_6__bdd_4_lut_24346.init = 16'h3cbc;
    PFUMX i23141 (.BLUT(n25434), .ALUT(n25433), .C0(index_i[6]), .Z(n25435));
    LUT4 mux_194_Mux_2_i955_else_4_lut (.A(index_i[4]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n25248)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+(D)))+!A !(B (C+!(D))+!B !(C+!(D))))) */ ;
    defparam mux_194_Mux_2_i955_else_4_lut.init = 16'h49c6;
    PFUMX i17794 (.BLUT(n476), .ALUT(n507), .C0(index_i[5]), .Z(n20124));
    PFUMX i17795 (.BLUT(n17556), .ALUT(n573_adj_2861), .C0(index_i[5]), 
          .Z(n20125));
    LUT4 index_i_6__bdd_1_lut (.A(index_i[5]), .Z(n26966)) /* synthesis lut_function=(!(A)) */ ;
    defparam index_i_6__bdd_1_lut.init = 16'h5555;
    LUT4 index_i_5__bdd_3_lut_24565 (.A(index_i[5]), .B(n26968), .C(index_i[3]), 
         .Z(n26969)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam index_i_5__bdd_3_lut_24565.init = 16'hcaca;
    PFUMX i17796 (.BLUT(n605_adj_2862), .ALUT(n636_adj_2863), .C0(index_i[5]), 
          .Z(n20126));
    LUT4 n25098_bdd_4_lut_24277 (.A(n24878), .B(n24892), .C(index_i[6]), 
         .D(index_i[5]), .Z(n26970)) /* synthesis lut_function=(!(A (B (C)+!B (D))+!A !(B (D)+!B (C)))) */ ;
    defparam n25098_bdd_4_lut_24277.init = 16'h5c3a;
    LUT4 n25098_bdd_4_lut (.A(n25098), .B(index_i[6]), .C(index_i[2]), 
         .D(index_i[5]), .Z(n26971)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A !(B (C+(D))+!B (D)))) */ ;
    defparam n25098_bdd_4_lut.init = 16'h5fe0;
    LUT4 n26972_bdd_3_lut (.A(n26972), .B(n26969), .C(index_i[4]), .Z(n26973)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n26972_bdd_3_lut.init = 16'hcaca;
    PFUMX mux_194_Mux_2_i891 (.BLUT(n875_adj_2864), .ALUT(n890_adj_2804), 
          .C0(index_i[4]), .Z(n891_adj_2865)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 mux_194_Mux_5_i124_3_lut (.A(n24996), .B(n25120), .C(index_i[3]), 
         .Z(n124_adj_2866)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_5_i124_3_lut.init = 16'hcaca;
    LUT4 i18407_3_lut_3_lut (.A(n24844), .B(index_i[4]), .C(n46_adj_2867), 
         .Z(n20737)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam i18407_3_lut_3_lut.init = 16'h7474;
    LUT4 n22_bdd_4_lut (.A(index_i[2]), .B(index_i[0]), .C(index_i[1]), 
         .D(index_i[5]), .Z(n27039)) /* synthesis lut_function=(!(A (B (C)+!B (D))+!A !(B (C+!(D))+!B (C+(D))))) */ ;
    defparam n22_bdd_4_lut.init = 16'h597e;
    PFUMX mux_194_Mux_2_i860 (.BLUT(n844), .ALUT(n859_adj_2868), .C0(index_i[4]), 
          .Z(n860_adj_2869)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    PFUMX i17797 (.BLUT(n21795), .ALUT(n700_adj_2870), .C0(index_i[5]), 
          .Z(n20127));
    L6MUX21 i17798 (.D0(n732_adj_2871), .D1(n21798), .SD(index_i[5]), 
            .Z(n20128));
    PFUMX i17799 (.BLUT(n797_adj_2872), .ALUT(n828_adj_2873), .C0(index_i[5]), 
          .Z(n20129));
    LUT4 n262_bdd_4_lut (.A(index_i[2]), .B(index_i[0]), .C(index_i[1]), 
         .D(index_i[3]), .Z(n27041)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(D))+!A (B ((D)+!C)+!B !(C+(D))))) */ ;
    defparam n262_bdd_4_lut.init = 16'h3358;
    PFUMX i23035 (.BLUT(n25263), .ALUT(n25264), .C0(index_i[1]), .Z(n25265));
    PFUMX i17800 (.BLUT(n860_adj_2874), .ALUT(n891_adj_2875), .C0(index_i[5]), 
          .Z(n20130));
    LUT4 i18420_3_lut_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n20750)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C+!(D))+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18420_3_lut_3_lut_4_lut_4_lut.init = 16'h1f81;
    LUT4 mux_194_Mux_6_i860_3_lut_3_lut (.A(n24844), .B(index_i[4]), .C(n844_adj_2876), 
         .Z(n860_adj_2838)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam mux_194_Mux_6_i860_3_lut_3_lut.init = 16'h7474;
    LUT4 mux_194_Mux_0_i124_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n124_adj_2877)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A !(B (D)+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_0_i124_3_lut_4_lut_4_lut.init = 16'h6c99;
    LUT4 i9433_3_lut (.A(n11998), .B(n25147), .C(index_i[3]), .Z(n11999)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9433_3_lut.init = 16'hcaca;
    PFUMX mux_194_Mux_3_i763 (.BLUT(n747_adj_2878), .ALUT(n762_adj_2803), 
          .C0(index_i[4]), .Z(n763_adj_2879)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 index_i_7__bdd_4_lut (.A(index_i[7]), .B(n14932), .C(n22792), 
         .D(index_i[5]), .Z(n24797)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(B (C+(D))+!B !((D)+!C)))) */ ;
    defparam index_i_7__bdd_4_lut.init = 16'h66f0;
    PFUMX i19003 (.BLUT(n21331), .ALUT(n21332), .C0(index_i[4]), .Z(n21333));
    PFUMX i19006 (.BLUT(n21334), .ALUT(n21335), .C0(index_i[4]), .Z(n21336));
    LUT4 n954_bdd_3_lut (.A(n954_adj_2880), .B(n173_adj_2881), .C(index_i[4]), 
         .Z(n23106)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n954_bdd_3_lut.init = 16'hacac;
    PFUMX i18408 (.BLUT(n20736), .ALUT(n20737), .C0(index_i[5]), .Z(n20738));
    PFUMX i18411 (.BLUT(n20739), .ALUT(n20740), .C0(index_i[5]), .Z(n20741));
    LUT4 index_i_4__bdd_4_lut_21646 (.A(index_i[4]), .B(n24961), .C(index_i[7]), 
         .D(n24951), .Z(n22792)) /* synthesis lut_function=(A (C+!(D))+!A (B+!(C))) */ ;
    defparam index_i_4__bdd_4_lut_21646.init = 16'he5ef;
    LUT4 n476_bdd_3_lut_21606 (.A(n476_adj_2882), .B(n23116), .C(index_i[5]), 
         .Z(n23117)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n476_bdd_3_lut_21606.init = 16'hcaca;
    PFUMX i18414 (.BLUT(n20742), .ALUT(n20743), .C0(index_i[5]), .Z(n20744));
    PFUMX mux_194_Mux_5_i732 (.BLUT(n11976), .ALUT(n731_adj_2883), .C0(index_i[4]), 
          .Z(n732_adj_2871)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    PFUMX i17819 (.BLUT(n94_adj_2884), .ALUT(n21801), .C0(index_i[5]), 
          .Z(n20149));
    L6MUX21 i18424 (.D0(n20752), .D1(n20753), .SD(index_i[5]), .Z(n20754));
    PFUMX i18427 (.BLUT(n20755), .ALUT(n20756), .C0(index_i[5]), .Z(n20757));
    PFUMX i17821 (.BLUT(n221_adj_2885), .ALUT(n252_adj_2886), .C0(index_i[5]), 
          .Z(n20151));
    PFUMX i18430 (.BLUT(n20758), .ALUT(n20759), .C0(index_i[5]), .Z(n20760));
    PFUMX i17822 (.BLUT(n286), .ALUT(n19899), .C0(index_i[5]), .Z(n20152));
    PFUMX i18433 (.BLUT(n20761), .ALUT(n20762), .C0(index_i[5]), .Z(n20763));
    LUT4 mux_194_Mux_8_i157_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n15_adj_2887)) /* synthesis lut_function=(A (B (C)+!B !(C (D)+!C !(D)))+!A !(B ((D)+!C)+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_8_i157_3_lut_4_lut_4_lut.init = 16'h83e0;
    LUT4 mux_194_Mux_0_i908_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n908)) /* synthesis lut_function=(!(A (B (C (D))+!B !(D))+!A (B+((D)+!C)))) */ ;
    defparam mux_194_Mux_0_i908_3_lut_4_lut_4_lut.init = 16'h2a98;
    LUT4 mux_194_Mux_6_i890_3_lut_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n890_adj_2888)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !((D)+!C))+!A !(B ((D)+!C)+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_6_i890_3_lut_3_lut_4_lut_4_lut.init = 16'h7e07;
    PFUMX i17823 (.BLUT(n349_adj_2889), .ALUT(n19902), .C0(index_i[5]), 
          .Z(n20153));
    LUT4 i18421_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n20751)) /* synthesis lut_function=(A (B (C+!(D))+!B !((D)+!C))+!A !(B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18421_3_lut_4_lut_4_lut.init = 16'h81f8;
    PFUMX i18436 (.BLUT(n20764), .ALUT(n20765), .C0(index_i[5]), .Z(n20766));
    LUT4 i2_2_lut (.A(index_i[3]), .B(index_i[5]), .Z(n6)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2_2_lut.init = 16'h8888;
    PFUMX i17828 (.BLUT(n669_adj_2890), .ALUT(n700_adj_2891), .C0(index_i[5]), 
          .Z(n20158));
    L6MUX21 i18443 (.D0(n20771), .D1(n20772), .SD(index_i[5]), .Z(n20773));
    PFUMX i17829 (.BLUT(n19914), .ALUT(n763_adj_2892), .C0(index_i[5]), 
          .Z(n20159));
    PFUMX i17830 (.BLUT(n19917), .ALUT(n828_adj_2893), .C0(index_i[5]), 
          .Z(n20160));
    PFUMX i17831 (.BLUT(n860_adj_2894), .ALUT(n19920), .C0(index_i[5]), 
          .Z(n20161));
    L6MUX21 i18450 (.D0(n20778), .D1(n20779), .SD(index_i[5]), .Z(n20780));
    L6MUX21 i22695 (.D0(n24376), .D1(n24373), .SD(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2126[4]));
    LUT4 n557_bdd_4_lut (.A(n24874), .B(index_i[4]), .C(n23026), .D(index_i[5]), 
         .Z(n24799)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (B (C (D))+!B (C+!(D)))) */ ;
    defparam n557_bdd_4_lut.init = 16'hf099;
    L6MUX21 i18457 (.D0(n20785), .D1(n20786), .SD(index_i[5]), .Z(n20787));
    PFUMX i18460 (.BLUT(n20788), .ALUT(n20789), .C0(index_i[5]), .Z(n20790));
    PFUMX i18463 (.BLUT(n20791), .ALUT(n20792), .C0(index_i[5]), .Z(n20793));
    PFUMX i18466 (.BLUT(n20794), .ALUT(n20795), .C0(index_i[5]), .Z(n20796));
    PFUMX i22690 (.BLUT(n24372), .ALUT(n20175), .C0(index_i[8]), .Z(n24373));
    PFUMX i18469 (.BLUT(n20797), .ALUT(n20798), .C0(index_i[5]), .Z(n20799));
    PFUMX i18472 (.BLUT(n20800), .ALUT(n20801), .C0(index_i[5]), .Z(n20802));
    PFUMX i22693 (.BLUT(n24375), .ALUT(n24374), .C0(index_i[8]), .Z(n24376));
    L6MUX21 i21305 (.D0(n22796), .D1(n24797), .SD(index_i[6]), .Z(n22797));
    PFUMX i18475 (.BLUT(n20803), .ALUT(n20804), .C0(index_i[5]), .Z(n20805));
    L6MUX21 i22670 (.D0(n24350), .D1(n24347), .SD(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2126[9]));
    PFUMX i18478 (.BLUT(n20806), .ALUT(n20807), .C0(index_i[5]), .Z(n20808));
    PFUMX i22668 (.BLUT(n24349), .ALUT(n24348), .C0(index_i[8]), .Z(n24350));
    PFUMX i17850 (.BLUT(n94_adj_2895), .ALUT(n125_adj_2896), .C0(index_i[5]), 
          .Z(n20180));
    PFUMX i17851 (.BLUT(n158_adj_2897), .ALUT(n189_adj_2824), .C0(index_i[5]), 
          .Z(n20181));
    PFUMX i22665 (.BLUT(n24346), .ALUT(n20098), .C0(index_i[8]), .Z(n24347));
    PFUMX i17852 (.BLUT(n221_adj_2898), .ALUT(n252_adj_2821), .C0(index_i[5]), 
          .Z(n20182));
    PFUMX i17853 (.BLUT(n286_adj_2899), .ALUT(n19929), .C0(index_i[5]), 
          .Z(n20183));
    PFUMX i17854 (.BLUT(n349_adj_2900), .ALUT(n19932), .C0(index_i[5]), 
          .Z(n20184));
    PFUMX i17855 (.BLUT(n413_adj_2901), .ALUT(n444_adj_2902), .C0(index_i[5]), 
          .Z(n20185));
    LUT4 n23119_bdd_3_lut (.A(n25274), .B(n444_adj_2903), .C(index_i[5]), 
         .Z(n23120)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n23119_bdd_3_lut.init = 16'hcaca;
    PFUMX i17856 (.BLUT(n476_adj_2904), .ALUT(n507_adj_2905), .C0(index_i[5]), 
          .Z(n20186));
    PFUMX i17857 (.BLUT(n19935), .ALUT(n573_adj_2906), .C0(index_i[5]), 
          .Z(n20187));
    PFUMX i17858 (.BLUT(n11986), .ALUT(n19938), .C0(index_i[5]), .Z(n20188));
    PFUMX i17859 (.BLUT(n669_adj_2907), .ALUT(n700_adj_2908), .C0(index_i[5]), 
          .Z(n20189));
    L6MUX21 i22644 (.D0(n24310), .D1(n24307), .SD(index_i[8]), .Z(n24311));
    LUT4 mux_194_Mux_0_i963_3_lut_3_lut_3_lut_rep_665 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27505)) /* synthesis lut_function=(!(A (B)+!A (B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_0_i963_3_lut_3_lut_3_lut_rep_665.init = 16'h3636;
    L6MUX21 i17860 (.D0(n19941), .D1(n763_adj_2879), .SD(index_i[5]), 
            .Z(n20190));
    PFUMX i17861 (.BLUT(n797_adj_2909), .ALUT(n828), .C0(index_i[5]), 
          .Z(n20191));
    PFUMX i22642 (.BLUT(n24309), .ALUT(n24308), .C0(index_i[7]), .Z(n24310));
    PFUMX i17862 (.BLUT(n860), .ALUT(n891_adj_2910), .C0(index_i[5]), 
          .Z(n20192));
    PFUMX i17863 (.BLUT(n924_adj_2911), .ALUT(n19944), .C0(index_i[5]), 
          .Z(n20193));
    PFUMX i17864 (.BLUT(n19947), .ALUT(n1018), .C0(index_i[5]), .Z(n20194));
    LUT4 mux_194_Mux_6_i844_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n844_adj_2876)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (B (C)+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_6_i844_3_lut_4_lut_4_lut.init = 16'hc1e0;
    PFUMX i22639 (.BLUT(n24306), .ALUT(n21602), .C0(index_i[7]), .Z(n24307));
    PFUMX i17882 (.BLUT(n158_adj_2912), .ALUT(n189_adj_2913), .C0(index_i[5]), 
          .Z(n20212));
    PFUMX i21303 (.BLUT(n24810), .ALUT(n24826), .C0(index_i[7]), .Z(n22796));
    PFUMX i17883 (.BLUT(n221_adj_2914), .ALUT(n19953), .C0(index_i[5]), 
          .Z(n20213));
    PFUMX i17884 (.BLUT(n286_adj_2915), .ALUT(n317_adj_2916), .C0(index_i[5]), 
          .Z(n20214));
    PFUMX i17885 (.BLUT(n349_adj_2917), .ALUT(n19956), .C0(index_i[5]), 
          .Z(n20215));
    PFUMX i17886 (.BLUT(n413_adj_2918), .ALUT(n19959), .C0(index_i[5]), 
          .Z(n20216));
    PFUMX i17887 (.BLUT(n19962), .ALUT(n507_adj_2919), .C0(index_i[5]), 
          .Z(n20217));
    PFUMX i17888 (.BLUT(n19965), .ALUT(n573_adj_2920), .C0(index_i[5]), 
          .Z(n20218));
    PFUMX i17889 (.BLUT(n605_adj_2921), .ALUT(n19968), .C0(index_i[5]), 
          .Z(n20219));
    PFUMX i17890 (.BLUT(n669_adj_2922), .ALUT(n700_adj_2923), .C0(index_i[5]), 
          .Z(n20220));
    PFUMX i17891 (.BLUT(n732_adj_2924), .ALUT(n763_adj_2925), .C0(index_i[5]), 
          .Z(n20221));
    L6MUX21 i17893 (.D0(n860_adj_2869), .D1(n891_adj_2865), .SD(index_i[5]), 
            .Z(n20223));
    L6MUX21 i22619 (.D0(n24283), .D1(n24281), .SD(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2126[7]));
    PFUMX i22617 (.BLUT(n24282), .ALUT(n20111), .C0(index_i[8]), .Z(n24283));
    LUT4 i20310_3_lut_then_4_lut (.A(index_i[0]), .B(index_i[4]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n25261)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)+!C !(D))+!B (C (D)))) */ ;
    defparam i20310_3_lut_then_4_lut.init = 16'hda0e;
    LUT4 i20310_3_lut_else_4_lut (.A(index_i[0]), .B(index_i[4]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n25260)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C))+!A (B (C)+!B (C+(D)))) */ ;
    defparam i20310_3_lut_else_4_lut.init = 16'hf178;
    LUT4 n25101_bdd_4_lut (.A(n141), .B(index_i[5]), .C(index_i[4]), .D(n24996), 
         .Z(n25430)) /* synthesis lut_function=(A (B (D)+!B ((D)+!C))+!A (B (D)+!B (C (D)))) */ ;
    defparam n25101_bdd_4_lut.init = 16'hfe02;
    LUT4 i18700_3_lut (.A(n236), .B(n251), .C(index_i[4]), .Z(n21030)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18700_3_lut.init = 16'hcaca;
    LUT4 i18693_3_lut (.A(n15_adj_2926), .B(n27527), .C(index_i[4]), .Z(n21023)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18693_3_lut.init = 16'hcaca;
    LUT4 n23157_bdd_3_lut (.A(n23157), .B(n476_adj_2882), .C(index_i[5]), 
         .Z(n23158)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n23157_bdd_3_lut.init = 16'hcaca;
    LUT4 i11507_3_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .Z(n11139)) /* synthesis lut_function=(!((B (C))+!A)) */ ;
    defparam i11507_3_lut.init = 16'h2a2a;
    LUT4 i19335_4_lut_4_lut (.A(n24878), .B(n24926), .C(index_i[5]), .D(index_i[4]), 
         .Z(n21665)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C+(D))+!B !(C (D)+!C !(D)))) */ ;
    defparam i19335_4_lut_4_lut.init = 16'hcf50;
    LUT4 n23161_bdd_3_lut (.A(n25265), .B(n23159), .C(index_i[5]), .Z(n23162)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n23161_bdd_3_lut.init = 16'hcaca;
    PFUMX i17578 (.BLUT(n19906), .ALUT(n19907), .C0(index_i[4]), .Z(n476_adj_2882));
    LUT4 i17589_3_lut (.A(n27502), .B(n325), .C(index_i[3]), .Z(n19919)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17589_3_lut.init = 16'hcaca;
    LUT4 i20313_3_lut (.A(n19918), .B(n19919), .C(index_i[4]), .Z(n19920)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20313_3_lut.init = 16'hcaca;
    PFUMX i22615 (.BLUT(n24280), .ALUT(n24279), .C0(index_i[8]), .Z(n24281));
    LUT4 i17576_3_lut (.A(n27508), .B(n25107), .C(index_i[3]), .Z(n19906)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17576_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_6_i653_3_lut (.A(n25141), .B(n85), .C(index_i[3]), 
         .Z(n653_adj_2927)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_6_i653_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_6_i668_3_lut (.A(n108), .B(n27509), .C(index_i[3]), 
         .Z(n668_adj_2928)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_6_i668_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_6_i684_3_lut (.A(n24996), .B(n27508), .C(index_i[3]), 
         .Z(n684_adj_2845)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_6_i684_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_6_i731_3_lut (.A(n25101), .B(n24995), .C(index_i[3]), 
         .Z(n731_adj_2842)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_6_i731_3_lut.init = 16'hcaca;
    PFUMX i21609 (.BLUT(n23162), .ALUT(n23158), .C0(index_i[6]), .Z(n23163));
    LUT4 mux_194_Mux_1_i94_3_lut (.A(index_i[0]), .B(n93_adj_2929), .C(index_i[4]), 
         .Z(n94)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_1_i94_3_lut.init = 16'hcaca;
    PFUMX i23033 (.BLUT(n25260), .ALUT(n25261), .C0(index_i[1]), .Z(n25262));
    LUT4 n20106_bdd_3_lut_23964 (.A(n20106), .B(n20107), .C(index_i[7]), 
         .Z(n24280)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n20106_bdd_3_lut_23964.init = 16'hcaca;
    LUT4 i17585_3_lut (.A(n588), .B(n25121), .C(index_i[3]), .Z(n19915)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17585_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_4_i828_3_lut (.A(n812_adj_2930), .B(n236), .C(index_i[4]), 
         .Z(n828_adj_2893)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_4_i828_3_lut.init = 16'hcaca;
    LUT4 n20106_bdd_3_lut_22614 (.A(n22869), .B(n20109), .C(index_i[7]), 
         .Z(n24279)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n20106_bdd_3_lut_22614.init = 16'hcaca;
    LUT4 n20111_bdd_3_lut (.A(n20102), .B(n25437), .C(index_i[7]), .Z(n24282)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n20111_bdd_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_1_i986_3_lut (.A(n27510), .B(n25143), .C(index_i[3]), 
         .Z(n986_adj_2831)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_1_i986_3_lut.init = 16'hcaca;
    LUT4 i17583_3_lut (.A(n900), .B(n325), .C(index_i[3]), .Z(n19913)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17583_3_lut.init = 16'hcaca;
    LUT4 i20226_3_lut (.A(n716_adj_2931), .B(n731_adj_2932), .C(index_i[4]), 
         .Z(n732_adj_2924)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20226_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_2_i669_3_lut (.A(n653_adj_2933), .B(n475_adj_2934), 
         .C(index_i[4]), .Z(n669_adj_2922)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_2_i669_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_2_i605_3_lut (.A(n142_adj_2935), .B(n604_adj_2936), 
         .C(index_i[4]), .Z(n605_adj_2921)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_2_i605_3_lut.init = 16'hcaca;
    PFUMX i18709 (.BLUT(n21023), .ALUT(n21024), .C0(index_i[5]), .Z(n21039));
    LUT4 mux_194_Mux_8_i892_3_lut_4_lut (.A(n24868), .B(index_i[4]), .C(index_i[5]), 
         .D(n860_adj_2823), .Z(n892_adj_2937)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_8_i892_3_lut_4_lut.init = 16'h4f40;
    LUT4 i20240_3_lut (.A(n25281), .B(n19964), .C(index_i[4]), .Z(n19965)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20240_3_lut.init = 16'hcaca;
    LUT4 i20242_3_lut (.A(n19960), .B(n19961), .C(index_i[4]), .Z(n19962)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20242_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_2_i413_3_lut (.A(n397_adj_2938), .B(n954_adj_2880), 
         .C(index_i[4]), .Z(n413_adj_2918)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_2_i413_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_2_i317_3_lut (.A(n668_adj_2939), .B(n316_adj_2940), 
         .C(index_i[4]), .Z(n317_adj_2916)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_2_i317_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_2_i286_3_lut (.A(n270), .B(n653_adj_2829), .C(index_i[4]), 
         .Z(n286_adj_2915)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_2_i286_3_lut.init = 16'hcaca;
    PFUMX i18710 (.BLUT(n21025), .ALUT(n21026), .C0(index_i[5]), .Z(n21040));
    LUT4 i17571_3_lut (.A(n25144), .B(n25138), .C(index_i[3]), .Z(n19901)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17571_3_lut.init = 16'hcaca;
    LUT4 i17570_3_lut (.A(n25137), .B(n325), .C(index_i[3]), .Z(n19900)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17570_3_lut.init = 16'hcaca;
    LUT4 i20326_3_lut (.A(n19900), .B(n19901), .C(index_i[4]), .Z(n19902)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20326_3_lut.init = 16'hcaca;
    LUT4 i20252_3_lut (.A(n142_adj_2941), .B(n13831), .C(index_i[4]), 
         .Z(n158_adj_2912)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20252_3_lut.init = 16'hcaca;
    L6MUX21 i18711 (.D0(n21027), .D1(n21028), .SD(index_i[5]), .Z(n21041));
    PFUMX i18712 (.BLUT(n21029), .ALUT(n21030), .C0(index_i[5]), .Z(n21042));
    LUT4 i17568_3_lut (.A(n25127), .B(n27515), .C(index_i[3]), .Z(n19898)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17568_3_lut.init = 16'hcaca;
    LUT4 n21602_bdd_3_lut (.A(n21588), .B(n23679), .C(index_i[6]), .Z(n24306)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n21602_bdd_3_lut.init = 16'hacac;
    LUT4 i20329_3_lut (.A(n19897), .B(n19898), .C(index_i[4]), .Z(n19899)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20329_3_lut.init = 16'hcaca;
    LUT4 n22786_bdd_3_lut_22641 (.A(n22786), .B(n21586), .C(index_i[6]), 
         .Z(n24308)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n22786_bdd_3_lut_22641.init = 16'hcaca;
    L6MUX21 i18714 (.D0(n21033), .D1(n21034), .SD(index_i[5]), .Z(n21044));
    LUT4 mux_194_Mux_5_i397_3_lut (.A(n25151), .B(n332), .C(index_i[3]), 
         .Z(n397_adj_2942)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_5_i397_3_lut.init = 16'hcaca;
    L6MUX21 i18715 (.D0(n21035), .D1(n21036), .SD(index_i[5]), .Z(n21045));
    L6MUX21 i18716 (.D0(n21037), .D1(n21038), .SD(index_i[5]), .Z(n21046));
    PFUMX i19396 (.BLUT(n844_adj_2943), .ALUT(n11938), .C0(index_i[4]), 
          .Z(n21726));
    LUT4 mux_194_Mux_5_i506_3_lut (.A(n27515), .B(n25126), .C(index_i[3]), 
         .Z(n506_adj_2944)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_5_i506_3_lut.init = 16'hcaca;
    LUT4 n25430_bdd_3_lut_23847 (.A(n25430), .B(n25429), .C(index_i[6]), 
         .Z(n25431)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n25430_bdd_3_lut_23847.init = 16'hcaca;
    LUT4 mux_194_Mux_11_i638_4_lut_4_lut (.A(n24827), .B(index_i[5]), .C(index_i[6]), 
         .D(n24855), .Z(n638)) /* synthesis lut_function=(A (B (C (D))+!B !(C))+!A (B ((D)+!C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_11_i638_4_lut_4_lut.init = 16'hc707;
    LUT4 mux_194_Mux_5_i15_3_lut (.A(n25146), .B(n25107), .C(index_i[3]), 
         .Z(n15)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_5_i15_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_5_i859_3_lut (.A(n141), .B(n25146), .C(index_i[3]), 
         .Z(n859_adj_2945)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_5_i859_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_5_i875_3_lut (.A(n24996), .B(n27510), .C(index_i[3]), 
         .Z(n875_adj_2946)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_5_i875_3_lut.init = 16'hcaca;
    LUT4 i20266_3_lut (.A(n19945), .B(n25279), .C(index_i[4]), .Z(n19947)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20266_3_lut.init = 16'hcaca;
    LUT4 n22786_bdd_3_lut (.A(n21584), .B(n23740), .C(index_i[6]), .Z(n24309)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n22786_bdd_3_lut.init = 16'hacac;
    LUT4 mux_194_Mux_3_i924_3_lut (.A(n908_adj_2947), .B(index_i[0]), .C(index_i[4]), 
         .Z(n924_adj_2911)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_3_i924_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_3_i891_3_lut (.A(n541_adj_2948), .B(n890_adj_2852), 
         .C(index_i[4]), .Z(n891_adj_2910)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_3_i891_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_3_i797_3_lut (.A(n731_adj_2842), .B(n796_adj_2949), 
         .C(index_i[4]), .Z(n797_adj_2909)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_3_i797_3_lut.init = 16'hcaca;
    LUT4 i12036_3_lut (.A(index_i[3]), .B(index_i[1]), .C(index_i[0]), 
         .Z(n14719)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i12036_3_lut.init = 16'hecec;
    LUT4 mux_194_Mux_3_i669_3_lut (.A(n653_adj_2829), .B(n668_adj_2939), 
         .C(index_i[4]), .Z(n669_adj_2907)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_3_i669_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut_4_lut (.A(n24827), .B(index_i[5]), .C(index_i[8]), .D(n25004), 
         .Z(n19492)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i2_3_lut_4_lut.init = 16'hfff8;
    LUT4 i20281_3_lut (.A(n19933), .B(n19934), .C(index_i[4]), .Z(n19935)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20281_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_3_i476_3_lut (.A(n460_adj_2950), .B(n285), .C(index_i[4]), 
         .Z(n476_adj_2904)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_3_i476_3_lut.init = 16'hcaca;
    LUT4 i11130_3_lut_4_lut (.A(index_i[4]), .B(n25111), .C(index_i[5]), 
         .D(n25098), .Z(n892)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11130_3_lut_4_lut.init = 16'hf8f0;
    LUT4 mux_194_Mux_4_i61_3_lut (.A(n25121), .B(n25154), .C(index_i[3]), 
         .Z(n61)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_4_i61_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_3_i413_3_lut (.A(n397_adj_2951), .B(n25108), .C(index_i[4]), 
         .Z(n413_adj_2901)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_3_i413_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_4_i270_3_lut (.A(n25147), .B(n27515), .C(index_i[3]), 
         .Z(n270_adj_2952)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_4_i270_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_4_i15_3_lut (.A(n25126), .B(n588), .C(index_i[3]), 
         .Z(n15_adj_2854)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_4_i15_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_3_i286_4_lut (.A(n93_adj_2953), .B(index_i[2]), .C(index_i[4]), 
         .D(n14729), .Z(n286_adj_2899)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_3_i286_4_lut.init = 16'h3aca;
    LUT4 mux_194_Mux_4_i348_3_lut (.A(n25125), .B(n25144), .C(index_i[3]), 
         .Z(n348_adj_2954)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_4_i348_3_lut.init = 16'hcaca;
    LUT4 i21607_then_3_lut (.A(index_i[0]), .B(index_i[4]), .C(index_i[3]), 
         .Z(n25264)) /* synthesis lut_function=(A (B)+!A (B (C)+!B !(C))) */ ;
    defparam i21607_then_3_lut.init = 16'hc9c9;
    LUT4 mux_194_Mux_4_i684_3_lut (.A(n85), .B(n108), .C(index_i[3]), 
         .Z(n684_adj_2955)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_4_i684_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_0_i475_3_lut_4_lut (.A(n25030), .B(index_i[1]), .C(index_i[3]), 
         .D(n24952), .Z(n475)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_0_i475_3_lut_4_lut.init = 16'h4f40;
    LUT4 mux_194_Mux_3_i491_3_lut_4_lut (.A(n25030), .B(index_i[1]), .C(index_i[3]), 
         .D(n25143), .Z(n491_adj_2956)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_3_i491_3_lut_4_lut.init = 16'h4f40;
    LUT4 mux_194_Mux_3_i158_3_lut (.A(n142_adj_2935), .B(n157), .C(index_i[4]), 
         .Z(n158_adj_2897)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_3_i158_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_3_i125_3_lut (.A(n46_adj_2867), .B(n526_adj_2957), 
         .C(index_i[4]), .Z(n125_adj_2896)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_3_i125_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_2_i189_3_lut_3_lut_4_lut (.A(index_i[1]), .B(n25111), 
         .C(n173_adj_2958), .D(index_i[4]), .Z(n189_adj_2913)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(C+(D)))) */ ;
    defparam mux_194_Mux_2_i189_3_lut_3_lut_4_lut.init = 16'h77f0;
    LUT4 mux_194_Mux_7_i333_3_lut (.A(n25099), .B(n24996), .C(index_i[3]), 
         .Z(n333_adj_2959)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_7_i333_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_7_i348_3_lut (.A(n27510), .B(n27517), .C(index_i[3]), 
         .Z(n348_adj_2960)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_7_i348_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_7_i397_3_lut (.A(n27510), .B(n25099), .C(index_i[3]), 
         .Z(n397_adj_2961)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_7_i397_3_lut.init = 16'hcaca;
    LUT4 n382_bdd_3_lut (.A(n23004), .B(n26973), .C(index_i[7]), .Z(n24349)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n382_bdd_3_lut.init = 16'hcaca;
    LUT4 n382_bdd_3_lut_22667 (.A(n382_adj_2801), .B(n509_adj_2802), .C(index_i[7]), 
         .Z(n24348)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n382_bdd_3_lut_22667.init = 16'hcaca;
    LUT4 n23032_bdd_3_lut_23915 (.A(n23032), .B(n23037), .C(index_i[7]), 
         .Z(n24346)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n23032_bdd_3_lut_23915.init = 16'hcaca;
    LUT4 i18477_3_lut (.A(n747_adj_2810), .B(n762_adj_2962), .C(index_i[4]), 
         .Z(n20807)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18477_3_lut.init = 16'hcaca;
    LUT4 i18476_3_lut (.A(n716_adj_2963), .B(n14712), .C(index_i[4]), 
         .Z(n20806)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18476_3_lut.init = 16'hcaca;
    LUT4 i18474_3_lut (.A(n93_adj_2964), .B(n699_adj_2816), .C(index_i[4]), 
         .Z(n20804)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18474_3_lut.init = 16'hcaca;
    LUT4 i18473_3_lut (.A(n653), .B(n24844), .C(index_i[4]), .Z(n20803)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18473_3_lut.init = 16'hcaca;
    LUT4 i11061_2_lut_3_lut_4_lut (.A(index_i[1]), .B(n25111), .C(index_i[5]), 
         .D(index_i[4]), .Z(n508)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;
    defparam i11061_2_lut_3_lut_4_lut.init = 16'hf080;
    LUT4 i21607_else_3_lut (.A(index_i[2]), .B(index_i[0]), .C(index_i[4]), 
         .D(index_i[3]), .Z(n25263)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)+!C !(D)))+!A (B (C+!(D))+!B !(C)))) */ ;
    defparam i21607_else_3_lut.init = 16'h1e38;
    LUT4 n20166_bdd_3_lut_23887 (.A(n20165), .B(n20164), .C(index_i[7]), 
         .Z(n24375)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n20166_bdd_3_lut_23887.init = 16'hacac;
    LUT4 i18331_3_lut_4_lut_4_lut (.A(n25093), .B(n24878), .C(index_i[4]), 
         .D(n24994), .Z(n20661)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B (C (D))+!B ((D)+!C)))) */ ;
    defparam i18331_3_lut_4_lut_4_lut.init = 16'h0c5c;
    LUT4 mux_194_Mux_8_i763_3_lut_4_lut_4_lut (.A(n25093), .B(n24960), .C(index_i[4]), 
         .D(n24994), .Z(n14960)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam mux_194_Mux_8_i763_3_lut_4_lut_4_lut.init = 16'hcfca;
    LUT4 n20166_bdd_3_lut_22692 (.A(n20166), .B(n23121), .C(index_i[7]), 
         .Z(n24374)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n20166_bdd_3_lut_22692.init = 16'hcaca;
    LUT4 i9378_3_lut_4_lut_4_lut (.A(n24997), .B(index_i[3]), .C(index_i[5]), 
         .D(n24892), .Z(n11944)) /* synthesis lut_function=(A (B+(C (D)))+!A (B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9378_3_lut_4_lut_4_lut.init = 16'hf8c8;
    LUT4 i18324_3_lut_3_lut_4_lut_4_lut (.A(n24997), .B(index_i[3]), .C(index_i[4]), 
         .D(n24978), .Z(n20654)) /* synthesis lut_function=(!(A (B (C)+!B ((D)+!C))+!A (B+((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18324_3_lut_3_lut_4_lut_4_lut.init = 16'h0838;
    LUT4 n557_bdd_3_lut_22672_4_lut_4_lut (.A(n24997), .B(index_i[3]), .C(index_i[4]), 
         .D(n24952), .Z(n23030)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C))+!A !(B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n557_bdd_3_lut_22672_4_lut_4_lut.init = 16'h838f;
    LUT4 i18467_3_lut (.A(n526_adj_2965), .B(n15_adj_2926), .C(index_i[4]), 
         .Z(n20797)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18467_3_lut.init = 16'hcaca;
    LUT4 i18464_3_lut (.A(n397_adj_2961), .B(n475_adj_2966), .C(index_i[4]), 
         .Z(n20794)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18464_3_lut.init = 16'hcaca;
    LUT4 i18462_3_lut (.A(n348_adj_2960), .B(n443), .C(index_i[4]), .Z(n20792)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18462_3_lut.init = 16'hcaca;
    LUT4 n62_bdd_3_lut_22771_4_lut (.A(n24997), .B(index_i[3]), .C(index_i[4]), 
         .D(n30_adj_2807), .Z(n23002)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n62_bdd_3_lut_22771_4_lut.init = 16'hf808;
    LUT4 i18461_3_lut (.A(n397_adj_2961), .B(n731_adj_2842), .C(index_i[4]), 
         .Z(n20791)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18461_3_lut.init = 16'hcaca;
    LUT4 i18459_3_lut (.A(n364_adj_2967), .B(n379_adj_2968), .C(index_i[4]), 
         .Z(n20789)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18459_3_lut.init = 16'hcaca;
    LUT4 i18458_3_lut (.A(n333_adj_2959), .B(n348_adj_2960), .C(index_i[4]), 
         .Z(n20788)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18458_3_lut.init = 16'hcaca;
    LUT4 i12046_3_lut (.A(index_i[3]), .B(index_i[1]), .C(index_i[0]), 
         .Z(n14729)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i12046_3_lut.init = 16'hc8c8;
    LUT4 mux_194_Mux_3_i348_3_lut (.A(n25143), .B(n25152), .C(index_i[3]), 
         .Z(n348_adj_2969)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_3_i348_3_lut.init = 16'hcaca;
    LUT4 n20168_bdd_3_lut (.A(n20168), .B(n20169), .C(index_i[7]), .Z(n24372)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n20168_bdd_3_lut.init = 16'hcaca;
    LUT4 i17833_4_lut (.A(n25268), .B(n1002_adj_2970), .C(index_i[5]), 
         .D(index_i[4]), .Z(n20163)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;
    defparam i17833_4_lut.init = 16'hfaca;
    LUT4 mux_194_Mux_4_i860_3_lut (.A(n506_adj_2944), .B(n15_adj_2971), 
         .C(index_i[4]), .Z(n860_adj_2894)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_4_i860_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_3_i684_3_lut (.A(n25148), .B(n25136), .C(index_i[3]), 
         .Z(n684_adj_2972)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_3_i684_3_lut.init = 16'hcaca;
    LUT4 i20315_3_lut (.A(n19915), .B(n19916), .C(index_i[4]), .Z(n19917)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20315_3_lut.init = 16'hcaca;
    LUT4 n25101_bdd_3_lut (.A(n25101), .B(n141), .C(index_i[4]), .Z(n25428)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n25101_bdd_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_6_i475_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n475_adj_2934)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A !(B (C+(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_6_i475_3_lut_4_lut_4_lut.init = 16'h9936;
    LUT4 i20317_3_lut (.A(n19912), .B(n19913), .C(index_i[4]), .Z(n19914)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20317_3_lut.init = 16'hcaca;
    LUT4 i9420_3_lut_4_lut (.A(n24952), .B(index_i[4]), .C(index_i[3]), 
         .D(n24998), .Z(n11986)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(C+(D)))) */ ;
    defparam i9420_3_lut_4_lut.init = 16'h7f70;
    CCU2D unary_minus_10_add_3_17 (.A0(\quarter_wave_sample_register_q[15] ), 
          .B0(GND_net), .C0(GND_net), .D0(GND_net), .A1(GND_net), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n17370), .S0(o_val_pipeline_i_0__15__N_2157[15]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam unary_minus_10_add_3_17.INIT0 = 16'hf555;
    defparam unary_minus_10_add_3_17.INIT1 = 16'h0000;
    defparam unary_minus_10_add_3_17.INJECT1_0 = "NO";
    defparam unary_minus_10_add_3_17.INJECT1_1 = "NO";
    LUT4 mux_194_Mux_4_i700_3_lut (.A(n684_adj_2955), .B(index_i[1]), .C(index_i[4]), 
         .Z(n700_adj_2891)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_4_i700_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_4_i669_3_lut (.A(n781_adj_2805), .B(n668_adj_2973), 
         .C(index_i[4]), .Z(n669_adj_2890)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_4_i669_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_4_i542_3_lut (.A(n526_adj_2957), .B(n506), .C(index_i[4]), 
         .Z(n542_adj_2974)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_4_i542_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_3_i908_3_lut (.A(n25131), .B(n25154), .C(index_i[3]), 
         .Z(n908_adj_2947)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_3_i908_3_lut.init = 16'hcaca;
    LUT4 n25100_bdd_4_lut_23850 (.A(n27510), .B(index_i[6]), .C(index_i[4]), 
         .D(n25146), .Z(n25432)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A !(B (C+!(D))+!B !(D))) */ ;
    defparam n25100_bdd_4_lut_23850.init = 16'hbf80;
    LUT4 i17827_4_lut (.A(n24927), .B(n25271), .C(index_i[5]), .D(index_i[4]), 
         .Z(n20157)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam i17827_4_lut.init = 16'hc5ca;
    CCU2D unary_minus_10_add_3_15 (.A0(quarter_wave_sample_register_i[13]), 
          .B0(GND_net), .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[14]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17369), .COUT(n17370), 
          .S0(o_val_pipeline_i_0__15__N_2157[13]), .S1(o_val_pipeline_i_0__15__N_2157[14]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam unary_minus_10_add_3_15.INIT0 = 16'hf555;
    defparam unary_minus_10_add_3_15.INIT1 = 16'hf555;
    defparam unary_minus_10_add_3_15.INJECT1_0 = "NO";
    defparam unary_minus_10_add_3_15.INJECT1_1 = "NO";
    CCU2D unary_minus_10_add_3_13 (.A0(quarter_wave_sample_register_i[11]), 
          .B0(GND_net), .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[12]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17368), .COUT(n17369), 
          .S0(o_val_pipeline_i_0__15__N_2157[11]), .S1(o_val_pipeline_i_0__15__N_2157[12]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam unary_minus_10_add_3_13.INIT0 = 16'hf555;
    defparam unary_minus_10_add_3_13.INIT1 = 16'hf555;
    defparam unary_minus_10_add_3_13.INJECT1_0 = "NO";
    defparam unary_minus_10_add_3_13.INJECT1_1 = "NO";
    LUT4 mux_194_Mux_3_i573_3_lut_3_lut_4_lut (.A(n24998), .B(index_i[3]), 
         .C(n460_adj_2975), .D(index_i[4]), .Z(n573_adj_2906)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_3_i573_3_lut_3_lut_4_lut.init = 16'h11f0;
    LUT4 i18322_3_lut_4_lut (.A(n24998), .B(index_i[3]), .C(index_i[4]), 
         .D(n285_adj_2976), .Z(n20652)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18322_3_lut_4_lut.init = 16'hfe0e;
    LUT4 mux_194_Mux_2_i270_3_lut (.A(n25146), .B(n25142), .C(index_i[3]), 
         .Z(n270)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_2_i270_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_2_i316_3_lut (.A(n25148), .B(n25121), .C(index_i[3]), 
         .Z(n316_adj_2940)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_2_i316_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_4_i286_3_lut (.A(n270_adj_2952), .B(n15_adj_2854), 
         .C(index_i[4]), .Z(n286)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_4_i286_3_lut.init = 16'hcaca;
    CCU2D unary_minus_10_add_3_11 (.A0(quarter_wave_sample_register_i[9]), 
          .B0(GND_net), .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[10]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17367), .COUT(n17368), 
          .S0(o_val_pipeline_i_0__15__N_2157[9]), .S1(o_val_pipeline_i_0__15__N_2157[10]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam unary_minus_10_add_3_11.INIT0 = 16'hf555;
    defparam unary_minus_10_add_3_11.INIT1 = 16'hf555;
    defparam unary_minus_10_add_3_11.INJECT1_0 = "NO";
    defparam unary_minus_10_add_3_11.INJECT1_1 = "NO";
    LUT4 mux_194_Mux_2_i573_3_lut_3_lut_4_lut (.A(n24998), .B(index_i[3]), 
         .C(n557_adj_2977), .D(index_i[4]), .Z(n573_adj_2920)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_2_i573_3_lut_3_lut_4_lut.init = 16'h11f0;
    LUT4 mux_194_Mux_2_i397_3_lut (.A(n27508), .B(n25101), .C(index_i[3]), 
         .Z(n397_adj_2938)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_2_i397_3_lut.init = 16'hcaca;
    LUT4 i18429_3_lut (.A(n491_adj_2978), .B(n506), .C(index_i[4]), .Z(n20759)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18429_3_lut.init = 16'hcaca;
    LUT4 i18428_3_lut (.A(n460_adj_2975), .B(n475_adj_2835), .C(index_i[4]), 
         .Z(n20758)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18428_3_lut.init = 16'hcaca;
    CCU2D unary_minus_10_add_3_9 (.A0(quarter_wave_sample_register_i[7]), 
          .B0(GND_net), .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[8]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17366), .COUT(n17367), 
          .S0(o_val_pipeline_i_0__15__N_2157[7]), .S1(o_val_pipeline_i_0__15__N_2157[8]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam unary_minus_10_add_3_9.INIT0 = 16'hf555;
    defparam unary_minus_10_add_3_9.INIT1 = 16'hf555;
    defparam unary_minus_10_add_3_9.INJECT1_0 = "NO";
    defparam unary_minus_10_add_3_9.INJECT1_1 = "NO";
    LUT4 n124_bdd_3_lut_21457_4_lut (.A(n24998), .B(index_i[3]), .C(index_i[4]), 
         .D(n124), .Z(n22999)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n124_bdd_3_lut_21457_4_lut.init = 16'hf101;
    LUT4 i18426_3_lut (.A(n251_adj_2813), .B(n443_adj_2820), .C(index_i[4]), 
         .Z(n20756)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18426_3_lut.init = 16'hcaca;
    LUT4 i18425_3_lut (.A(n460_adj_2975), .B(n14712), .C(index_i[4]), 
         .Z(n20755)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;
    defparam i18425_3_lut.init = 16'h3a3a;
    LUT4 mux_194_Mux_4_i94_3_lut (.A(n61), .B(n25110), .C(index_i[4]), 
         .Z(n94_adj_2884)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_4_i94_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_4_i573_3_lut_3_lut_4_lut_4_lut (.A(n24998), .B(index_i[3]), 
         .C(index_i[4]), .D(n24978), .Z(n573_adj_2979)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_4_i573_3_lut_3_lut_4_lut_4_lut.init = 16'h1f1c;
    LUT4 mux_194_Mux_5_i731_3_lut (.A(n27501), .B(n27502), .C(index_i[3]), 
         .Z(n731_adj_2883)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_5_i731_3_lut.init = 16'hcaca;
    LUT4 i18413_3_lut (.A(n236_adj_2980), .B(n251_adj_2813), .C(index_i[4]), 
         .Z(n20743)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18413_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_10_i125_3_lut_4_lut_4_lut (.A(n24998), .B(index_i[3]), 
         .C(index_i[4]), .D(n24952), .Z(n125)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B (C (D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_10_i125_3_lut_4_lut_4_lut.init = 16'h3efe;
    LUT4 i18412_3_lut (.A(n205), .B(n15_adj_2887), .C(index_i[4]), .Z(n20742)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18412_3_lut.init = 16'hcaca;
    LUT4 i18409_3_lut (.A(n301_adj_2981), .B(n93_adj_2964), .C(index_i[4]), 
         .Z(n20739)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18409_3_lut.init = 16'hcaca;
    LUT4 i18406_3_lut (.A(n15_adj_2887), .B(n526_adj_2957), .C(index_i[4]), 
         .Z(n20736)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18406_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_10_i574_4_lut_4_lut (.A(n24874), .B(index_i[4]), .C(index_i[5]), 
         .D(n24866), .Z(n574_adj_2826)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_10_i574_4_lut_4_lut.init = 16'h1f1c;
    PFUMX i21576 (.BLUT(n23120), .ALUT(n23117), .C0(index_i[6]), .Z(n23121));
    LUT4 mux_194_Mux_3_i747_3_lut (.A(n25138), .B(n404), .C(index_i[3]), 
         .Z(n747_adj_2878)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_3_i747_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_6_i285_3_lut_4_lut (.A(n25124), .B(index_i[2]), .C(index_i[3]), 
         .D(n25153), .Z(n285)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_6_i285_3_lut_4_lut.init = 16'hf606;
    LUT4 i17643_3_lut_4_lut (.A(n25124), .B(index_i[2]), .C(index_i[3]), 
         .D(n25151), .Z(n19973)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i17643_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_194_Mux_5_i891_3_lut (.A(n875_adj_2946), .B(n379_adj_2968), 
         .C(index_i[4]), .Z(n891_adj_2875)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_5_i891_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_5_i860_3_lut (.A(n15), .B(n859_adj_2945), .C(index_i[4]), 
         .Z(n860_adj_2874)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_5_i860_3_lut.init = 16'hcaca;
    LUT4 i19461_3_lut_4_lut (.A(n25124), .B(index_i[2]), .C(index_i[3]), 
         .D(n27502), .Z(n21791)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19461_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_194_Mux_5_i797_3_lut (.A(n781_adj_2982), .B(n251_adj_2983), 
         .C(index_i[4]), .Z(n797_adj_2872)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_5_i797_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_3_i460_3_lut_4_lut (.A(n25124), .B(index_i[2]), .C(index_i[3]), 
         .D(n25121), .Z(n460_adj_2950)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_3_i460_3_lut_4_lut.init = 16'h6f60;
    LUT4 i20353_3_lut (.A(n21793), .B(n21794), .C(index_i[4]), .Z(n21795)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20353_3_lut.init = 16'hcaca;
    LUT4 i17596_then_4_lut (.A(index_i[0]), .B(index_i[4]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n25267)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C))+!A (B (C)+!B !(C+!(D)))) */ ;
    defparam i17596_then_4_lut.init = 16'hc34a;
    LUT4 n25100_bdd_3_lut_23140 (.A(n12162), .B(n12163), .C(index_i[2]), 
         .Z(n25433)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n25100_bdd_3_lut_23140.init = 16'hacac;
    LUT4 mux_194_Mux_10_i637_3_lut_4_lut_4_lut (.A(n24926), .B(index_i[4]), 
         .C(index_i[5]), .D(n24874), .Z(n637)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_10_i637_3_lut_4_lut_4_lut.init = 16'h1f1c;
    LUT4 mux_194_Mux_5_i636_4_lut (.A(n157_adj_2984), .B(n24928), .C(index_i[4]), 
         .D(index_i[3]), .Z(n636_adj_2863)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_5_i636_4_lut.init = 16'h3aca;
    LUT4 n25100_bdd_3_lut_23372 (.A(n27510), .B(n27509), .C(index_i[4]), 
         .Z(n25434)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n25100_bdd_3_lut_23372.init = 16'hacac;
    LUT4 i20359_3_lut (.A(n17554), .B(n17555), .C(index_i[4]), .Z(n17556)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20359_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_5_i507_3_lut (.A(n491_adj_2985), .B(n506_adj_2944), 
         .C(index_i[4]), .Z(n507)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_5_i507_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_0_i220_3_lut (.A(n24995), .B(n25143), .C(index_i[3]), 
         .Z(n220)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_0_i220_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_5_i476_3_lut (.A(n460_adj_2986), .B(n475_adj_2987), 
         .C(index_i[4]), .Z(n476)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_5_i476_3_lut.init = 16'hcaca;
    LUT4 i11101_2_lut_rep_245_3_lut_4_lut (.A(n24878), .B(index_i[4]), .C(index_i[6]), 
         .D(index_i[5]), .Z(n24805)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11101_2_lut_rep_245_3_lut_4_lut.init = 16'hf080;
    LUT4 i17596_else_4_lut (.A(index_i[0]), .B(index_i[4]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n25266)) /* synthesis lut_function=(A (C)+!A !(B ((D)+!C)+!B !(C))) */ ;
    defparam i17596_else_4_lut.init = 16'hb0f0;
    LUT4 mux_194_Mux_5_i413_3_lut (.A(n397_adj_2942), .B(n251_adj_2847), 
         .C(index_i[4]), .Z(n413_adj_2858)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_5_i413_3_lut.init = 16'hcaca;
    LUT4 i12304_1_lut_2_lut_3_lut_4_lut (.A(n24878), .B(index_i[4]), .C(index_i[6]), 
         .D(index_i[5]), .Z(n382)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i12304_1_lut_2_lut_3_lut_4_lut.init = 16'h0f7f;
    LUT4 i19297_3_lut_4_lut (.A(n24880), .B(n24879), .C(index_i[5]), .D(index_i[6]), 
         .Z(n21627)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (B+((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19297_3_lut_4_lut.init = 16'hffc5;
    LUT4 n25435_bdd_3_lut (.A(n25435), .B(n25432), .C(index_i[5]), .Z(n25436)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n25435_bdd_3_lut.init = 16'hcaca;
    LUT4 i15281_3_lut (.A(n17542), .B(n17543), .C(index_i[4]), .Z(n17544)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15281_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_5_i125_3_lut (.A(n109_adj_2988), .B(n124_adj_2866), 
         .C(index_i[4]), .Z(n125_adj_2851)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_5_i125_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_5_i94_3_lut (.A(n653_adj_2927), .B(n635_adj_2989), 
         .C(index_i[4]), .Z(n94_adj_2850)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_5_i94_3_lut.init = 16'hcaca;
    CCU2D unary_minus_10_add_3_7 (.A0(quarter_wave_sample_register_i[5]), 
          .B0(GND_net), .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[6]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17365), .COUT(n17366), 
          .S0(o_val_pipeline_i_0__15__N_2157[5]), .S1(o_val_pipeline_i_0__15__N_2157[6]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam unary_minus_10_add_3_7.INIT0 = 16'hf555;
    defparam unary_minus_10_add_3_7.INIT1 = 16'hf555;
    defparam unary_minus_10_add_3_7.INJECT1_0 = "NO";
    defparam unary_minus_10_add_3_7.INJECT1_1 = "NO";
    CCU2D unary_minus_10_add_3_5 (.A0(quarter_wave_sample_register_i[3]), 
          .B0(GND_net), .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[4]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17364), .COUT(n17365), 
          .S0(o_val_pipeline_i_0__15__N_2157[3]), .S1(o_val_pipeline_i_0__15__N_2157[4]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam unary_minus_10_add_3_5.INIT0 = 16'hf555;
    defparam unary_minus_10_add_3_5.INIT1 = 16'hf555;
    defparam unary_minus_10_add_3_5.INJECT1_0 = "NO";
    defparam unary_minus_10_add_3_5.INJECT1_1 = "NO";
    LUT4 i17581_then_4_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[4]), 
         .D(index_i[3]), .Z(n25270)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+(D)))+!A !(B (C)+!B !(C+!(D)))) */ ;
    defparam i17581_then_4_lut.init = 16'h9c97;
    LUT4 mux_194_Mux_6_i891_3_lut (.A(n301_adj_2981), .B(n890_adj_2888), 
         .C(index_i[4]), .Z(n891_adj_2839)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_6_i891_3_lut.init = 16'hcaca;
    LUT4 i21155_2_lut (.A(index_i[4]), .B(index_i[3]), .Z(n19821)) /* synthesis lut_function=((B)+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i21155_2_lut.init = 16'hdddd;
    LUT4 mux_194_Mux_6_i828_4_lut (.A(n812_adj_2990), .B(n13817), .C(index_i[4]), 
         .D(index_i[2]), .Z(n828_adj_2837)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_6_i828_4_lut.init = 16'hfaca;
    LUT4 mux_194_Mux_6_i797_3_lut (.A(n781_adj_2805), .B(n24818), .C(index_i[4]), 
         .Z(n797)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_6_i797_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_6_i669_3_lut (.A(n653_adj_2927), .B(n668_adj_2928), 
         .C(index_i[4]), .Z(n669)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_6_i669_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_6_i542_3_lut (.A(n526_adj_2991), .B(n541_adj_2948), 
         .C(index_i[4]), .Z(n542)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_6_i542_3_lut.init = 16'hcaca;
    PFUMX mux_194_Mux_1_i891 (.BLUT(n882), .ALUT(n890_adj_2992), .C0(n19821), 
          .Z(n891)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 mux_194_Mux_6_i252_4_lut (.A(index_i[2]), .B(n251_adj_2847), .C(index_i[4]), 
         .D(n11139), .Z(n252_adj_2993)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_6_i252_4_lut.init = 16'hc5ca;
    LUT4 i20855_3_lut (.A(n23673), .B(n252_adj_2993), .C(index_i[5]), 
         .Z(n21586)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20855_3_lut.init = 16'hcaca;
    PFUMX i23138 (.BLUT(n12163), .ALUT(n25428), .C0(index_i[5]), .Z(n25429));
    LUT4 i10986_2_lut_rep_564 (.A(index_i[0]), .B(index_i[1]), .Z(n25124)) /* synthesis lut_function=((B)+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i10986_2_lut_rep_564.init = 16'hdddd;
    LUT4 i21574_then_4_lut (.A(index_i[0]), .B(index_i[4]), .C(index_i[1]), 
         .D(index_i[3]), .Z(n25273)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam i21574_then_4_lut.init = 16'h3c69;
    PFUMX i23026 (.BLUT(n25248), .ALUT(n25249), .C0(index_i[0]), .Z(n25250));
    L6MUX21 i21563 (.D0(n23107), .D1(n23105), .SD(index_i[6]), .Z(n23108));
    PFUMX i21561 (.BLUT(n924_adj_2994), .ALUT(n23106), .C0(index_i[5]), 
          .Z(n23107));
    LUT4 i21574_else_4_lut (.A(index_i[0]), .B(index_i[4]), .C(index_i[1]), 
         .D(index_i[3]), .Z(n25272)) /* synthesis lut_function=(!(A (B (C)+!B !(C (D)+!C !(D)))+!A (B ((D)+!C)+!B !((D)+!C)))) */ ;
    defparam i21574_else_4_lut.init = 16'h394b;
    PFUMX i21559 (.BLUT(n23104), .ALUT(n24867), .C0(index_i[5]), .Z(n23105));
    LUT4 i21160_2_lut (.A(index_i[5]), .B(index_i[4]), .Z(n19809)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i21160_2_lut.init = 16'heeee;
    LUT4 i18297_3_lut (.A(n20619), .B(n20620), .C(index_i[7]), .Z(n20627)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18297_3_lut.init = 16'hcaca;
    LUT4 i18290_3_lut (.A(n20605), .B(n23710), .C(index_i[6]), .Z(n20620)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18290_3_lut.init = 16'hcaca;
    LUT4 i18299_3_lut (.A(n20623), .B(n20624), .C(index_i[7]), .Z(n20629)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18299_3_lut.init = 16'hcaca;
    PFUMX i18273 (.BLUT(n11999), .ALUT(n62_adj_2995), .C0(index_i[5]), 
          .Z(n20603));
    LUT4 i18293_3_lut (.A(n23716), .B(n20612), .C(index_i[6]), .Z(n20623)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18293_3_lut.init = 16'hcaca;
    LUT4 i17781_3_lut (.A(n20104), .B(n20105), .C(index_i[7]), .Z(n20111)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17781_3_lut.init = 16'hcaca;
    LUT4 i17774_3_lut (.A(n20787), .B(n20790), .C(index_i[6]), .Z(n20104)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17774_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_0_i397_3_lut (.A(n27517), .B(n27502), .C(index_i[3]), 
         .Z(n397)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_0_i397_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_1_i620_3_lut_4_lut (.A(n25061), .B(index_i[1]), .C(index_i[3]), 
         .D(n25147), .Z(n620_adj_2856)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_1_i620_3_lut_4_lut.init = 16'hdfd0;
    LUT4 mux_194_Mux_0_i173_3_lut_4_lut (.A(n25061), .B(index_i[1]), .C(index_i[3]), 
         .D(n25144), .Z(n173)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_0_i173_3_lut_4_lut.init = 16'hdfd0;
    LUT4 i19421_3_lut_4_lut (.A(n25061), .B(index_i[1]), .C(index_i[3]), 
         .D(n404), .Z(n21751)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19421_3_lut_4_lut.init = 16'hdfd0;
    LUT4 mux_194_Mux_0_i581_3_lut_3_lut_rep_677 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27517)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_0_i581_3_lut_3_lut_rep_677.init = 16'hc7c7;
    LUT4 i19299_3_lut (.A(n21622), .B(n21623), .C(index_i[7]), .Z(n21629)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19299_3_lut.init = 16'hcaca;
    LUT4 i19292_3_lut (.A(n23754), .B(n20754), .C(index_i[6]), .Z(n21622)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19292_3_lut.init = 16'hcaca;
    LUT4 i17875_3_lut (.A(n20199), .B(n20200), .C(index_i[7]), .Z(n20205)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17875_3_lut.init = 16'hcaca;
    LUT4 i17870_3_lut (.A(n20189), .B(n20190), .C(index_i[6]), .Z(n20200)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17870_3_lut.init = 16'hcaca;
    LUT4 i17904_3_lut (.A(n23163), .B(n20227), .C(index_i[7]), .Z(n20234)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17904_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_0_i188_3_lut (.A(n27509), .B(n101), .C(index_i[3]), 
         .Z(n188)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_0_i188_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_6_i325_3_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n325)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_6_i325_3_lut_4_lut_3_lut.init = 16'h6d6d;
    LUT4 mux_194_Mux_2_i700_3_lut_4_lut (.A(index_i[1]), .B(n25093), .C(index_i[4]), 
         .D(n684), .Z(n700_adj_2923)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam mux_194_Mux_2_i700_3_lut_4_lut.init = 16'hefe0;
    LUT4 mux_194_Mux_3_i1018_3_lut_4_lut (.A(index_i[1]), .B(n25093), .C(index_i[4]), 
         .D(n19633), .Z(n1018)) /* synthesis lut_function=(A (C+!(D))+!A (B (C+!(D))+!B !(C+(D)))) */ ;
    defparam mux_194_Mux_3_i1018_3_lut_4_lut.init = 16'he0ef;
    L6MUX21 i24333 (.D0(n27043), .D1(n27040), .SD(index_i[4]), .Z(n27044));
    LUT4 i20168_3_lut (.A(n25233), .B(n124_adj_2877), .C(index_i[4]), 
         .Z(n21026)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20168_3_lut.init = 16'hcaca;
    PFUMX i24331 (.BLUT(n27042), .ALUT(n27041), .C0(index_i[5]), .Z(n27043));
    LUT4 mux_194_Mux_1_i747_4_lut_then_4_lut (.A(index_i[0]), .B(index_i[4]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n25276)) /* synthesis lut_function=(A (B ((D)+!C))+!A !(B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_1_i747_4_lut_then_4_lut.init = 16'h9d5d;
    PFUMX i24327 (.BLUT(n27039), .ALUT(n27038), .C0(index_i[3]), .Z(n27040));
    LUT4 mux_194_Mux_0_i635_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n635)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_0_i635_3_lut_4_lut_4_lut.init = 16'hfd0a;
    LUT4 mux_194_Mux_1_i747_4_lut_else_4_lut (.A(index_i[0]), .B(index_i[4]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n25275)) /* synthesis lut_function=(!(A (B (C (D))+!B !(D))+!A ((C (D))+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_1_i747_4_lut_else_4_lut.init = 16'h2ecc;
    LUT4 i19004_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n21334)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (D))+!A !(D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19004_3_lut_4_lut_4_lut_4_lut.init = 16'ha25d;
    LUT4 i17577_3_lut_3_lut (.A(n25099), .B(index_i[3]), .C(n1001), .Z(n19907)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam i17577_3_lut_3_lut.init = 16'h7474;
    LUT4 i9589_3_lut_4_lut (.A(n24994), .B(index_i[2]), .C(index_i[5]), 
         .D(n27516), .Z(n12159)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9589_3_lut_4_lut.init = 16'hfe0e;
    LUT4 i17630_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n19960)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+(D)))+!A !(B (D)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i17630_3_lut_4_lut_4_lut.init = 16'h99c7;
    LUT4 mux_194_Mux_3_i93_3_lut_4_lut (.A(n24994), .B(index_i[2]), .C(index_i[3]), 
         .D(n27516), .Z(n93_adj_2953)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_3_i93_3_lut_4_lut.init = 16'hefe0;
    LUT4 mux_194_Mux_0_i316_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n316_adj_2800)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+(D)))+!A (B (C+(D))+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_0_i316_3_lut_4_lut_4_lut_4_lut.init = 16'h332d;
    LUT4 i11128_2_lut_3_lut_4_lut (.A(n24994), .B(index_i[2]), .C(index_i[5]), 
         .D(n25092), .Z(n764_adj_2799)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11128_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 mux_194_Mux_0_i1002_3_lut_3_lut_4_lut (.A(n24994), .B(index_i[2]), 
         .C(n1001), .D(index_i[3]), .Z(n1002)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_0_i1002_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 i17808_3_lut (.A(n20127), .B(n20128), .C(index_i[6]), .Z(n20138)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17808_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_0_i627_3_lut_rep_565 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n25125)) /* synthesis lut_function=(A (B+!(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_0_i627_3_lut_rep_565.init = 16'hdada;
    LUT4 mux_194_Mux_7_i379_3_lut_3_lut (.A(n25099), .B(index_i[3]), .C(n27517), 
         .Z(n379_adj_2968)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam mux_194_Mux_7_i379_3_lut_3_lut.init = 16'h7474;
    LUT4 mux_194_Mux_4_i668_3_lut_3_lut (.A(n25099), .B(index_i[3]), .C(n27508), 
         .Z(n668_adj_2973)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;
    defparam mux_194_Mux_4_i668_3_lut_3_lut.init = 16'hd1d1;
    PFUMX i21296 (.BLUT(n22785), .ALUT(n25112), .C0(index_i[5]), .Z(n22786));
    LUT4 mux_194_Mux_7_i364_3_lut_3_lut (.A(n25099), .B(index_i[3]), .C(n27510), 
         .Z(n364_adj_2967)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;
    defparam mux_194_Mux_7_i364_3_lut_3_lut.init = 16'hd1d1;
    LUT4 i18438_3_lut_3_lut (.A(n25099), .B(index_i[3]), .C(n27508), .Z(n20768)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam i18438_3_lut_3_lut.init = 16'h7474;
    LUT4 i19285_3_lut_4_lut (.A(n25098), .B(index_i[2]), .C(index_i[3]), 
         .D(n25152), .Z(n21615)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19285_3_lut_4_lut.init = 16'hdfd0;
    PFUMX i24278 (.BLUT(n26971), .ALUT(n26970), .C0(index_i[3]), .Z(n26972));
    PFUMX i24274 (.BLUT(n26967), .ALUT(n26966), .C0(index_i[2]), .Z(n26968));
    LUT4 mux_194_Mux_0_i795_3_lut_3_lut_rep_566 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n25126)) /* synthesis lut_function=(A (B+(C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_0_i795_3_lut_3_lut_rep_566.init = 16'hadad;
    LUT4 mux_194_Mux_12_i254_4_lut (.A(n24826), .B(n24852), .C(index_i[6]), 
         .D(n6), .Z(n254_adj_2827)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_12_i254_4_lut.init = 16'hca0a;
    LUT4 mux_194_Mux_6_i7_3_lut_4_lut_3_lut_rep_567 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n25127)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_6_i7_3_lut_4_lut_3_lut_rep_567.init = 16'hd6d6;
    LUT4 i19464_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21794)) /* synthesis lut_function=(A (B (C)+!B !(C (D)+!C !(D)))+!A (B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19464_3_lut_4_lut_4_lut.init = 16'hd6a5;
    PFUMX i17849 (.BLUT(n31_adj_2860), .ALUT(n62_adj_2996), .C0(index_i[5]), 
          .Z(n20179));
    LUT4 i18694_3_lut_4_lut (.A(n24952), .B(index_i[3]), .C(index_i[4]), 
         .D(n46), .Z(n21024)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18694_3_lut_4_lut.init = 16'h8f80;
    LUT4 index_i_0__bdd_4_lut_23048 (.A(index_i[0]), .B(index_i[3]), .C(index_i[1]), 
         .D(index_i[2]), .Z(n25279)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C))+!A (B (C (D)+!C !(D))+!B !(C+!(D))))) */ ;
    defparam index_i_0__bdd_4_lut_23048.init = 16'h16d3;
    PFUMX i17818 (.BLUT(n31_adj_2855), .ALUT(n62_adj_2853), .C0(index_i[5]), 
          .Z(n20148));
    LUT4 n851_bdd_3_lut_22131_4_lut (.A(n25135), .B(index_i[2]), .C(index_i[3]), 
         .D(n25127), .Z(n23734)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n851_bdd_3_lut_22131_4_lut.init = 16'hf606;
    LUT4 i18718_3_lut (.A(n21041), .B(n21042), .C(index_i[6]), .Z(n21048)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18718_3_lut.init = 16'hcaca;
    LUT4 i18719_3_lut (.A(n27044), .B(n21044), .C(index_i[6]), .Z(n21049)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18719_3_lut.init = 16'hcaca;
    LUT4 index_i_0__bdd_4_lut_23314 (.A(index_i[0]), .B(index_i[3]), .C(index_i[1]), 
         .D(index_i[2]), .Z(n25281)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C (D)))+!A !(B (C+!(D))+!B !(C+(D))))) */ ;
    defparam index_i_0__bdd_4_lut_23314.init = 16'h4ae7;
    PFUMX i17787 (.BLUT(n31), .ALUT(n21749), .C0(index_i[5]), .Z(n20117));
    LUT4 mux_194_Mux_12_i1023_4_lut (.A(n20581), .B(n766_adj_2997), .C(index_i[9]), 
         .D(index_i[8]), .Z(quarter_wave_sample_register_i_15__N_2126[12])) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_12_i1023_4_lut.init = 16'hfaca;
    LUT4 mux_194_Mux_12_i766_4_lut (.A(n24810), .B(n765), .C(index_i[7]), 
         .D(index_i[6]), .Z(n766_adj_2997)) /* synthesis lut_function=(A (B (C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_12_i766_4_lut.init = 16'hc0c5;
    LUT4 i17764_3_lut (.A(n20092), .B(n20093), .C(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2126[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17764_3_lut.init = 16'hcaca;
    LUT4 i17763_4_lut (.A(n20596), .B(n893), .C(index_i[8]), .D(index_i[7]), 
         .Z(n20093)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;
    defparam i17763_4_lut.init = 16'hfaca;
    LUT4 index_i_1__bdd_4_lut_23893 (.A(index_i[1]), .B(index_i[0]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n25283)) /* synthesis lut_function=(!(A (B (D)+!B (C+!(D)))+!A !(B (C (D)+!C !(D))+!B !((D)+!C)))) */ ;
    defparam index_i_1__bdd_4_lut_23893.init = 16'h429c;
    LUT4 i17739_3_lut_4_lut_4_lut (.A(n24997), .B(n25127), .C(index_i[3]), 
         .D(index_i[0]), .Z(n20069)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C))) */ ;
    defparam i17739_3_lut_4_lut_4_lut.init = 16'hcfc5;
    LUT4 i19241_3_lut_3_lut_4_lut (.A(n25098), .B(index_i[2]), .C(n1001), 
         .D(index_i[3]), .Z(n21571)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19241_3_lut_3_lut_4_lut.init = 16'hf077;
    LUT4 mux_194_Mux_3_i668_3_lut_4_lut (.A(n25135), .B(index_i[2]), .C(index_i[3]), 
         .D(n25144), .Z(n668_adj_2939)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_3_i668_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_194_Mux_8_i301_3_lut_4_lut (.A(n25098), .B(index_i[2]), .C(index_i[3]), 
         .D(n27516), .Z(n301_adj_2981)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_8_i301_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_194_Mux_4_i763_3_lut_4_lut (.A(n25135), .B(index_i[2]), .C(index_i[4]), 
         .D(n747_adj_2848), .Z(n763_adj_2892)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_4_i763_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_194_Mux_8_i173_3_lut_3_lut_4_lut (.A(n25098), .B(index_i[2]), 
         .C(n27516), .D(index_i[3]), .Z(n173_adj_2881)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_8_i173_3_lut_3_lut_4_lut.init = 16'hf077;
    LUT4 i9590_3_lut_3_lut_4_lut (.A(n25098), .B(index_i[2]), .C(n15_adj_2887), 
         .D(index_i[4]), .Z(n12160)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9590_3_lut_3_lut_4_lut.init = 16'hf077;
    LUT4 i21125_2_lut_rep_266_3_lut_4_lut (.A(n25098), .B(index_i[2]), .C(index_i[5]), 
         .D(n25092), .Z(n24826)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i21125_2_lut_rep_266_3_lut_4_lut.init = 16'h0f7f;
    LUT4 i11995_3_lut_3_lut_rep_668 (.A(index_i[2]), .B(index_i[0]), .C(index_i[1]), 
         .Z(n27508)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11995_3_lut_3_lut_rep_668.init = 16'hd0d0;
    LUT4 n22_bdd_3_lut_24408_4_lut (.A(index_i[2]), .B(index_i[0]), .C(index_i[1]), 
         .D(index_i[5]), .Z(n27038)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n22_bdd_3_lut_24408_4_lut.init = 16'h0fd0;
    LUT4 mux_194_Mux_6_i15_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n15_adj_2971)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C))+!A !(B (C+!(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_6_i15_3_lut_4_lut_4_lut.init = 16'h5ad6;
    LUT4 n851_bdd_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n23735)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n851_bdd_3_lut_4_lut_4_lut.init = 16'ha5ad;
    PFUMX mux_194_Mux_8_i764 (.BLUT(n716_adj_2808), .ALUT(n732_adj_2849), 
          .C0(n19809), .Z(n764)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    PFUMX mux_194_Mux_8_i574 (.BLUT(n542_adj_2841), .ALUT(n11943), .C0(index_i[5]), 
          .Z(n574)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 i17738_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n20068)) /* synthesis lut_function=(!(A (B (C (D))+!B (C (D)+!C !(D)))+!A !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i17738_3_lut_4_lut_4_lut.init = 16'h5aad;
    LUT4 mux_194_Mux_0_i796_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n796)) /* synthesis lut_function=(A (B (C+(D))+!B (C (D)))+!A !(B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_0_i796_3_lut_4_lut_4_lut.init = 16'hadc0;
    LUT4 i19239_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21569)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C))+!A !(B (C)+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19239_3_lut_4_lut_4_lut.init = 16'h5ad3;
    LUT4 i17607_3_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[0]), .C(index_i[1]), 
         .D(index_i[3]), .Z(n19937)) /* synthesis lut_function=(A (B (C)+!B !(C+!(D)))+!A (B (C)+!B !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i17607_3_lut_4_lut_4_lut.init = 16'hc3d0;
    LUT4 mux_194_Mux_9_i62_3_lut_4_lut_then_4_lut (.A(index_i[4]), .B(index_i[2]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n25300)) /* synthesis lut_function=(!(A (B (C+(D)))+!A (B+(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_9_i62_3_lut_4_lut_then_4_lut.init = 16'h222b;
    LUT4 i1_2_lut_rep_501 (.A(index_i[0]), .B(index_i[2]), .Z(n25061)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i1_2_lut_rep_501.init = 16'heeee;
    LUT4 mux_194_Mux_9_i62_3_lut_4_lut_else_4_lut (.A(index_i[4]), .B(index_i[2]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n25299)) /* synthesis lut_function=((B+(C (D)))+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_9_i62_3_lut_4_lut_else_4_lut.init = 16'hfddd;
    LUT4 i15300_3_lut_4_lut (.A(index_i[0]), .B(index_i[2]), .C(n25062), 
         .D(index_i[4]), .Z(n286_adj_2998)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i15300_3_lut_4_lut.init = 16'hfe00;
    LUT4 i2_2_lut_rep_502 (.A(index_i[1]), .B(index_i[3]), .Z(n25062)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i2_2_lut_rep_502.init = 16'heeee;
    LUT4 i11999_1_lut_2_lut (.A(index_i[1]), .B(index_i[3]), .Z(n541)) /* synthesis lut_function=(!(A+(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11999_1_lut_2_lut.init = 16'h1111;
    LUT4 mux_194_Mux_7_i60_3_lut_4_lut_3_lut_rep_669 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27509)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B+!(C)))) */ ;
    defparam mux_194_Mux_7_i60_3_lut_4_lut_3_lut_rep_669.init = 16'h1818;
    LUT4 mux_194_Mux_2_i557_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n557_adj_2977)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C+!(D))+!B (C (D)+!C !(D))))) */ ;
    defparam mux_194_Mux_2_i557_3_lut_3_lut_4_lut.init = 16'h0f18;
    LUT4 mux_194_Mux_0_i698_3_lut_rep_670 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27510)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B (C)+!B !(C)))) */ ;
    defparam mux_194_Mux_0_i698_3_lut_rep_670.init = 16'h1c1c;
    LUT4 i17588_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n19918)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i17588_3_lut_4_lut_4_lut.init = 16'hda5a;
    LUT4 i11170_2_lut_rep_569 (.A(index_i[0]), .B(index_i[1]), .Z(n25129)) /* synthesis lut_function=(A+!(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11170_2_lut_rep_569.init = 16'hbbbb;
    LUT4 i9429_3_lut_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n875_adj_2864)) /* synthesis lut_function=(A (C (D))+!A !(B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9429_3_lut_3_lut_4_lut_4_lut.init = 16'hb555;
    LUT4 i17604_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n19934)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B (C (D)+!C !(D))))) */ ;
    defparam i17604_3_lut_3_lut_4_lut.init = 16'h0f1c;
    LUT4 i17637_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n19967)) /* synthesis lut_function=(A (C+(D))+!A !(B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i17637_3_lut_4_lut_4_lut.init = 16'haba5;
    LUT4 i1_2_lut_rep_434 (.A(index_i[0]), .B(index_i[1]), .Z(n24994)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i1_2_lut_rep_434.init = 16'h8888;
    LUT4 mux_194_Mux_8_i29_3_lut_rep_671 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27511)) /* synthesis lut_function=(!(A (B (C))+!A !(B+(C)))) */ ;
    defparam mux_194_Mux_8_i29_3_lut_rep_671.init = 16'h7e7e;
    LUT4 mux_194_Mux_7_i526_3_lut_3_lut_4_lut_3_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n526_adj_2965)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(D))+!A !(D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_7_i526_3_lut_3_lut_4_lut_3_lut_4_lut.init = 16'h887f;
    LUT4 mux_194_Mux_3_i1002_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n19633)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (D))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_3_i1002_3_lut_3_lut_4_lut.init = 16'hf708;
    LUT4 mux_194_Mux_6_i332_3_lut_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n332)) /* synthesis lut_function=(!(A (C)+!A !((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_6_i332_3_lut_3_lut_3_lut.init = 16'h5b5b;
    PFUMX i18303 (.BLUT(n20631), .ALUT(n20632), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2126[1]));
    LUT4 mux_194_Mux_6_i812_3_lut_4_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n812_adj_2990)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(D))+!A !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_6_i812_3_lut_4_lut_3_lut_4_lut.init = 16'h7780;
    LUT4 i11057_2_lut_rep_319_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[4]), .D(n25111), .Z(n24879)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11057_2_lut_rep_319_3_lut_4_lut.init = 16'hf8f0;
    LUT4 i10989_2_lut_rep_392_3_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .Z(n24952)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i10989_2_lut_rep_392_3_lut.init = 16'hf8f8;
    LUT4 mux_194_Mux_4_i1002_3_lut_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n1002_adj_2970)) /* synthesis lut_function=(A (B (C (D))+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_4_i1002_3_lut_3_lut_3_lut_4_lut.init = 16'hf007;
    LUT4 mux_194_Mux_4_i900_3_lut_4_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n900)) /* synthesis lut_function=(A ((C)+!B)+!A !(B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_4_i900_3_lut_4_lut_4_lut_3_lut.init = 16'hb2b2;
    LUT4 i12240_2_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(n25094), 
         .D(index_i[2]), .Z(n14932)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i12240_2_lut_3_lut_4_lut.init = 16'hf080;
    LUT4 mux_194_Mux_0_i620_3_lut (.A(n27510), .B(n25147), .C(index_i[3]), 
         .Z(n620)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_0_i620_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_8_i526_3_lut_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n526_adj_2840)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_8_i526_3_lut_3_lut_3_lut_4_lut.init = 16'h0f70;
    LUT4 i20813_3_lut (.A(n20224), .B(n23829), .C(index_i[6]), .Z(n20233)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20813_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_0_i986_3_lut (.A(n27504), .B(n985), .C(index_i[3]), 
         .Z(n986)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_0_i986_3_lut.init = 16'hcaca;
    LUT4 i2_2_lut_rep_307_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(n25092), 
         .D(index_i[2]), .Z(n24867)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i2_2_lut_rep_307_3_lut_4_lut.init = 16'hfff8;
    LUT4 i10990_2_lut_rep_306_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n24866)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i10990_2_lut_rep_306_3_lut_4_lut.init = 16'hf080;
    LUT4 n77_bdd_3_lut_22932_3_lut_4_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n23706)) /* synthesis lut_function=(A (B (C)+!B !(D))+!A !(D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n77_bdd_3_lut_22932_3_lut_4_lut_3_lut_4_lut.init = 16'h80f7;
    LUT4 n72_bdd_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n23672)) /* synthesis lut_function=(!(A (D)+!A !(B (D)+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n72_bdd_4_lut_4_lut_4_lut.init = 16'h54bb;
    LUT4 i12185_2_lut_rep_292_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[4]), .D(index_i[2]), .Z(n24852)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i12185_2_lut_rep_292_3_lut_4_lut.init = 16'hf080;
    LUT4 mux_194_Mux_4_i526_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n526_adj_2957)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A !(B ((D)+!C)+!B (C (D)+!C !(D))))) */ ;
    defparam mux_194_Mux_4_i526_3_lut_3_lut_4_lut.init = 16'h7e0f;
    LUT4 mux_194_Mux_5_i459_3_lut_4_lut_3_lut_rep_571 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n25131)) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_5_i459_3_lut_4_lut_3_lut_rep_571.init = 16'h6b6b;
    LUT4 index_i_6__bdd_3_lut_22005_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(n25111), .D(index_i[6]), .Z(n23035)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam index_i_6__bdd_3_lut_22005_4_lut.init = 16'hf07f;
    LUT4 mux_194_Mux_3_i796_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n796_adj_2949)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C))+!A (B (C+!(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_3_i796_3_lut_4_lut_4_lut_4_lut.init = 16'hf07c;
    LUT4 index_i_6__bdd_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(n25093), 
         .D(index_i[6]), .Z(n23034)) /* synthesis lut_function=(!(A (B (D)+!B (C (D)+!C !(D)))+!A (B (C (D))+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam index_i_6__bdd_4_lut_4_lut.init = 16'h07fc;
    PFUMX i19304 (.BLUT(n21632), .ALUT(n21633), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2126[8]));
    LUT4 mux_194_Mux_0_i364_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n364_adj_2833)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A ((C+!(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_0_i364_3_lut_3_lut_4_lut.init = 16'hdb55;
    LUT4 n699_bdd_4_lut_21492_4_lut (.A(n24978), .B(index_i[3]), .C(n24998), 
         .D(index_i[6]), .Z(n22969)) /* synthesis lut_function=(!(A (B+(C (D)+!C !(D)))+!A (B (D)+!B (C (D)+!C !(D))))) */ ;
    defparam n699_bdd_4_lut_21492_4_lut.init = 16'h0374;
    LUT4 mux_194_Mux_4_i205_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n205_adj_2999)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C (D)+!C !(D))+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_4_i205_3_lut_4_lut_4_lut_4_lut.init = 16'h1fc0;
    LUT4 mux_194_Mux_5_i781_3_lut_4_lut_4_lut (.A(index_i[1]), .B(n25138), 
         .C(index_i[3]), .D(n25030), .Z(n781_adj_2982)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_5_i781_3_lut_4_lut_4_lut.init = 16'hfc5c;
    PFUMX i17761 (.BLUT(n20089), .ALUT(n20090), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2126[11]));
    LUT4 n9595_bdd_3_lut_22148_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n23751)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C (D)+!C !(D))+!B (C)))) */ ;
    defparam n9595_bdd_3_lut_22148_3_lut_4_lut.init = 16'h0fc1;
    LUT4 n19949_bdd_3_lut_3_lut (.A(index_i[1]), .B(n526_adj_2991), .C(index_i[4]), 
         .Z(n23159)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n19949_bdd_3_lut_3_lut.init = 16'h5c5c;
    PFUMX i17611 (.BLUT(n19939), .ALUT(n19940), .C0(index_i[4]), .Z(n19941));
    PFUMX i21494 (.BLUT(n23035), .ALUT(n23034), .C0(index_i[5]), .Z(n23036));
    LUT4 i17634_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n19964)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D))+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i17634_3_lut_4_lut.init = 16'hccdb;
    LUT4 mux_194_Mux_6_i157_3_lut_4_lut_4_lut_4_lut_4_lut (.A(index_i[1]), 
         .B(index_i[2]), .C(index_i[3]), .D(index_i[0]), .Z(n157_adj_2846)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A (B (D)+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_6_i157_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'h19cc;
    LUT4 n476_bdd_3_lut_22270_3_lut (.A(index_i[1]), .B(index_i[4]), .C(n124_adj_2866), 
         .Z(n23157)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n476_bdd_3_lut_22270_3_lut.init = 16'hd1d1;
    LUT4 i11169_2_lut_rep_416_2_lut (.A(index_i[1]), .B(index_i[0]), .Z(n24976)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11169_2_lut_rep_416_2_lut.init = 16'h4444;
    L6MUX21 i21490 (.D0(n23031), .D1(n24799), .SD(index_i[6]), .Z(n23032));
    LUT4 mux_194_Mux_7_i716_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n716_adj_2963)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C+!(D))+!B (C)))) */ ;
    defparam mux_194_Mux_7_i716_3_lut_3_lut_4_lut.init = 16'h0f81;
    PFUMX i21488 (.BLUT(n23030), .ALUT(n23029), .C0(index_i[5]), .Z(n23031));
    LUT4 mux_194_Mux_5_i460_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n460_adj_2986)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A !(B (C)+!B !(C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_5_i460_3_lut_4_lut_4_lut.init = 16'h6b5a;
    LUT4 mux_194_Mux_8_i124_3_lut_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n124_adj_3000)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C+!(D)))+!A (B (C (D)+!C !(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_8_i124_3_lut_3_lut_4_lut_4_lut.init = 16'h07c1;
    PFUMX i17817 (.BLUT(n20145), .ALUT(n20146), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2126[5]));
    LUT4 mux_194_Mux_0_i971_3_lut (.A(n27505), .B(n27511), .C(index_i[3]), 
         .Z(n971)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_0_i971_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_6_i636_4_lut_4_lut (.A(index_i[1]), .B(index_i[4]), 
         .C(n635_adj_2989), .D(n14349), .Z(n636)) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_6_i636_4_lut_4_lut.init = 16'hf3d1;
    LUT4 mux_194_Mux_3_i349_3_lut_3_lut (.A(index_i[1]), .B(index_i[4]), 
         .C(n348_adj_2969), .Z(n349_adj_2900)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_3_i349_3_lut_3_lut.init = 16'hd1d1;
    LUT4 mux_194_Mux_7_i620_3_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .D(index_i[3]), .Z(n620_adj_3001)) /* synthesis lut_function=(A (B (C+!(D)))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_7_i620_3_lut_4_lut_4_lut.init = 16'h9199;
    LUT4 i17567_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n19897)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A !(B (C+!(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i17567_3_lut_4_lut_4_lut.init = 16'ha52b;
    PFUMX i21294 (.BLUT(n25117), .ALUT(n22783), .C0(index_i[2]), .Z(n22784));
    LUT4 mux_194_Mux_7_i262_3_lut_rep_435 (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .Z(n24995)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_7_i262_3_lut_rep_435.init = 16'h6464;
    LUT4 i17753_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[0]), 
         .D(index_i[3]), .Z(n20083)) /* synthesis lut_function=(!(A (B (D)+!B !(C+!(D)))+!A !(B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i17753_3_lut_4_lut.init = 16'h64aa;
    LUT4 i11171_2_lut_rep_437 (.A(index_i[1]), .B(index_i[2]), .Z(n24997)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11171_2_lut_rep_437.init = 16'heeee;
    LUT4 i20664_3_lut (.A(n26429), .B(n25262), .C(index_i[5]), .Z(n20162)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20664_3_lut.init = 16'hcaca;
    LUT4 i10985_2_lut_rep_575 (.A(index_i[0]), .B(index_i[1]), .Z(n25135)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i10985_2_lut_rep_575.init = 16'h4444;
    LUT4 i11112_2_lut_rep_314_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n24874)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11112_2_lut_rep_314_3_lut_4_lut.init = 16'hf0e0;
    LUT4 mux_194_Mux_2_i173_3_lut_3_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n173_adj_2958)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_2_i173_3_lut_3_lut_3_lut_4_lut.init = 16'h0e1e;
    PFUMX i17879 (.BLUT(n20207), .ALUT(n20208), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2126[3]));
    LUT4 mux_194_Mux_5_i954_3_lut_3_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n954_adj_2880)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B (C)+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_5_i954_3_lut_3_lut_4_lut_4_lut.init = 16'h0c1c;
    LUT4 i18699_3_lut_4_lut (.A(n24952), .B(index_i[3]), .C(index_i[4]), 
         .D(n220), .Z(n21029)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18699_3_lut_4_lut.init = 16'hf808;
    LUT4 i20668_3_lut (.A(n542_adj_2974), .B(n573_adj_2979), .C(index_i[5]), 
         .Z(n20156)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20668_3_lut.init = 16'hcaca;
    PFUMX i17910 (.BLUT(n20238), .ALUT(n20239), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2126[2]));
    LUT4 i11153_2_lut_rep_331_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[0]), 
         .Z(n24891)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11153_2_lut_rep_331_3_lut.init = 16'hfefe;
    LUT4 mux_194_Mux_9_i285_3_lut_3_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n285_adj_2976)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_9_i285_3_lut_3_lut_4_lut_4_lut.init = 16'hc0c1;
    LUT4 i11062_2_lut_rep_366_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[3]), 
         .Z(n24926)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11062_2_lut_rep_366_3_lut.init = 16'he0e0;
    LUT4 i11063_2_lut_rep_295_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[4]), .D(index_i[3]), .Z(n24855)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11063_2_lut_rep_295_3_lut_4_lut.init = 16'hfef0;
    LUT4 i7033_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n157_adj_2984)) /* synthesis lut_function=(!(A (C (D))+!A !(B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i7033_3_lut_4_lut_4_lut.init = 16'h4aaa;
    LUT4 mux_194_Mux_0_i954_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n954)) /* synthesis lut_function=(A (D)+!A !(B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_0_i954_3_lut_4_lut_4_lut.init = 16'haf40;
    LUT4 i19469_3_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[3]), 
         .D(index_i[0]), .Z(n21799)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19469_3_lut_3_lut_4_lut.init = 16'h0fe0;
    LUT4 mux_194_Mux_9_i93_3_lut_3_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .Z(n93)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_9_i93_3_lut_3_lut_3_lut.init = 16'hc1c1;
    L6MUX21 i12804359_i1 (.D0(n21053), .D1(n21746), .SD(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2126[0]));
    LUT4 i9407_2_lut_rep_532 (.A(index_i[3]), .B(index_i[4]), .Z(n25092)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9407_2_lut_rep_532.init = 16'heeee;
    LUT4 mux_194_Mux_6_i22_3_lut_3_lut_rep_576 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n25136)) /* synthesis lut_function=(!(A (C)+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_6_i22_3_lut_3_lut_rep_576.init = 16'h4a4a;
    LUT4 i11660_2_lut_rep_281_2_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .Z(n24841)) /* synthesis lut_function=(A (C)+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11660_2_lut_rep_281_2_lut_3_lut.init = 16'hf1f1;
    LUT4 i19306_3_lut_3_lut_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[3]), 
         .Z(n21636)) /* synthesis lut_function=(A (C)+!A (B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19306_3_lut_3_lut_3_lut.init = 16'he5e5;
    LUT4 i9392_3_lut_4_lut (.A(index_i[3]), .B(index_i[4]), .C(n25140), 
         .D(n27508), .Z(n605)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9392_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_194_Mux_7_i506_3_lut_4_lut (.A(n25098), .B(index_i[2]), .C(index_i[3]), 
         .D(n27510), .Z(n506_adj_3002)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_7_i506_3_lut_4_lut.init = 16'h2f20;
    LUT4 mux_194_Mux_0_i953_3_lut_rep_577 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n25137)) /* synthesis lut_function=(A (C)+!A !((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_0_i953_3_lut_rep_577.init = 16'ha4a4;
    LUT4 mux_194_Mux_8_i93_3_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .D(index_i[3]), .Z(n93_adj_2964)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(D))+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_8_i93_3_lut_3_lut_4_lut.init = 16'h3391;
    LUT4 i11113_2_lut_rep_533 (.A(index_i[2]), .B(index_i[3]), .Z(n25093)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11113_2_lut_rep_533.init = 16'heeee;
    LUT4 i11162_2_lut_rep_438 (.A(index_i[1]), .B(index_i[2]), .Z(n24998)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11162_2_lut_rep_438.init = 16'h8888;
    LUT4 i11829_2_lut_rep_391_3_lut (.A(index_i[2]), .B(index_i[3]), .C(index_i[1]), 
         .Z(n24951)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11829_2_lut_rep_391_3_lut.init = 16'hfefe;
    LUT4 i11115_2_lut_rep_367_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[3]), 
         .Z(n24927)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11115_2_lut_rep_367_3_lut.init = 16'hf8f8;
    LUT4 i11049_2_lut_rep_309_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n24869)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11049_2_lut_rep_309_3_lut_4_lut.init = 16'hf8f0;
    LUT4 i12179_2_lut_rep_332_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[0]), 
         .Z(n24892)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i12179_2_lut_rep_332_3_lut.init = 16'h8080;
    LUT4 mux_194_Mux_6_i442_3_lut_4_lut_3_lut_rep_578 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n25138)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_6_i442_3_lut_4_lut_3_lut_rep_578.init = 16'h6464;
    LUT4 i21121_2_lut_rep_308_2_lut_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n24868)) /* synthesis lut_function=(!(A+(B+(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i21121_2_lut_rep_308_2_lut_3_lut_4_lut.init = 16'h0111;
    LUT4 i17622_3_lut_4_lut (.A(n25098), .B(index_i[2]), .C(index_i[3]), 
         .D(n141), .Z(n19952)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i17622_3_lut_4_lut.init = 16'hf202;
    LUT4 mux_194_Mux_8_i491_3_lut_4_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .D(index_i[3]), .Z(n491_adj_2978)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(D))+!A !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_8_i491_3_lut_4_lut_3_lut_4_lut.init = 16'h7780;
    LUT4 mux_194_Mux_3_i221_3_lut_4_lut (.A(n24952), .B(index_i[3]), .C(index_i[4]), 
         .D(n24961), .Z(n221_adj_2898)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_3_i221_3_lut_4_lut.init = 16'h08f8;
    LUT4 i2_3_lut_4_lut_adj_83 (.A(index_i[1]), .B(index_i[2]), .C(index_i[5]), 
         .D(n25092), .Z(n17674)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i2_3_lut_4_lut_adj_83.init = 16'hfff8;
    LUT4 i9417_2_lut_rep_534 (.A(index_i[3]), .B(index_i[4]), .Z(n25094)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9417_2_lut_rep_534.init = 16'h8888;
    LUT4 mux_194_Mux_0_i490_3_lut_4_lut_4_lut_3_lut_rep_579 (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[2]), .Z(n25139)) /* synthesis lut_function=(!(A (B+!(C))+!A ((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_0_i490_3_lut_4_lut_4_lut_3_lut_rep_579.init = 16'h2424;
    LUT4 mux_194_Mux_7_i475_3_lut_3_lut_4_lut (.A(n25098), .B(index_i[2]), 
         .C(n27517), .D(index_i[3]), .Z(n475_adj_2966)) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))+!A !(B ((D)+!C)+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_7_i475_3_lut_3_lut_4_lut.init = 16'h99f0;
    LUT4 i1_2_lut_rep_333_3_lut (.A(index_i[3]), .B(index_i[4]), .C(index_i[5]), 
         .Z(n24893)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i1_2_lut_rep_333_3_lut.init = 16'hf8f8;
    LUT4 i19322_3_lut_3_lut_4_lut (.A(index_i[3]), .B(index_i[4]), .C(n413), 
         .D(index_i[5]), .Z(n21652)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19322_3_lut_3_lut_4_lut.init = 16'h77f0;
    LUT4 mux_194_Mux_0_i557_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n557)) /* synthesis lut_function=(A ((D)+!C)+!A !((D)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_0_i557_3_lut_4_lut.init = 16'haa4e;
    LUT4 mux_194_Mux_0_i939_4_lut (.A(n588), .B(n24976), .C(index_i[3]), 
         .D(index_i[2]), .Z(n939)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_0_i939_4_lut.init = 16'hfaca;
    LUT4 mux_194_Mux_9_i412_3_lut_4_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .Z(n412)) /* synthesis lut_function=(!(A (B (C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_9_i412_3_lut_4_lut_3_lut.init = 16'h7e7e;
    LUT4 mux_194_Mux_0_i491_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n491_adj_2834)) /* synthesis lut_function=(!(A (B (D)+!B !(C+!(D)))+!A ((C+!(D))+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_0_i491_3_lut_4_lut.init = 16'h24aa;
    LUT4 mux_194_Mux_8_i412_3_lut_4_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .Z(n14712)) /* synthesis lut_function=(A (B+!(C))+!A !((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_8_i412_3_lut_4_lut_3_lut.init = 16'h8e8e;
    LUT4 i17582_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n19912)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i17582_3_lut_4_lut.init = 16'h64cc;
    LUT4 i9424_2_lut_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[3]), 
         .Z(n11990)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9424_2_lut_3_lut.init = 16'h8080;
    LUT4 mux_194_Mux_0_i781_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n781)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A (B (C)+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_0_i781_4_lut_4_lut_4_lut.init = 16'h0cb4;
    L6MUX21 i21463 (.D0(n23003), .D1(n23001), .SD(index_i[6]), .Z(n23004));
    LUT4 i18468_3_lut_4_lut_4_lut_4_lut (.A(n25098), .B(index_i[2]), .C(index_i[3]), 
         .D(index_i[4]), .Z(n20798)) /* synthesis lut_function=(A (B)+!A (B (C (D))+!B !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18468_3_lut_4_lut_4_lut_4_lut.init = 16'hc999;
    LUT4 mux_194_Mux_5_i475_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n475_adj_2987)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_5_i475_3_lut_4_lut_4_lut.init = 16'hd4a5;
    LUT4 i20302_3_lut (.A(n620_adj_3001), .B(n13813), .C(index_i[4]), 
         .Z(n20801)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20302_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_0_i157_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n157_adj_2830)) /* synthesis lut_function=(A (B (C+!(D))+!B !(D))+!A (B (D)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_0_i157_3_lut_4_lut.init = 16'hd4aa;
    LUT4 i19242_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21572)) /* synthesis lut_function=(!(A ((D)+!C)+!A !(B ((D)+!C)+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19242_3_lut_3_lut_4_lut.init = 16'h55a4;
    LUT4 i20305_3_lut (.A(n491_adj_2811), .B(n506_adj_3002), .C(index_i[4]), 
         .Z(n20795)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20305_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_4_i812_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n812_adj_2930)) /* synthesis lut_function=(!(A (C+(D))+!A !(B (C+(D))+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_4_i812_3_lut_3_lut_4_lut.init = 16'h554a;
    PFUMX mux_194_Mux_13_i1023 (.BLUT(n511), .ALUT(n19492), .C0(index_i[9]), 
          .Z(quarter_wave_sample_register_i_15__N_2126[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 mux_194_Mux_6_i70_3_lut_rep_675 (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .Z(n27515)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_6_i70_3_lut_rep_675.init = 16'h1c1c;
    LUT4 mux_194_Mux_5_i491_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n491_adj_2985)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A !(B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_5_i491_3_lut_4_lut_4_lut.init = 16'ha54a;
    LUT4 i19001_3_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[0]), 
         .D(index_i[3]), .Z(n21331)) /* synthesis lut_function=(!(A (B (C)+!B !(C (D)))+!A (B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19001_3_lut_4_lut_4_lut.init = 16'h3c1c;
    LUT4 i18454_3_lut (.A(n141), .B(n24995), .C(index_i[3]), .Z(n20784)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18454_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_2_i348_3_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .D(index_i[3]), .Z(n348_adj_3003)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+(D)))+!A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_2_i348_3_lut_4_lut_4_lut.init = 16'h1cc3;
    LUT4 i18453_3_lut (.A(n85), .B(n27510), .C(index_i[3]), .Z(n20783)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18453_3_lut.init = 16'hcaca;
    LUT4 i20990_2_lut_rep_580 (.A(index_i[0]), .B(index_i[1]), .Z(n25140)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20990_2_lut_rep_580.init = 16'h9999;
    LUT4 i18452_3_lut (.A(n25107), .B(n25099), .C(index_i[3]), .Z(n20782)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18452_3_lut.init = 16'hcaca;
    PFUMX i21461 (.BLUT(n23002), .ALUT(n62), .C0(index_i[5]), .Z(n23003));
    LUT4 i11658_2_lut_rep_439 (.A(index_i[1]), .B(index_i[2]), .C(index_i[0]), 
         .Z(n24999)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11658_2_lut_rep_439.init = 16'h7070;
    PFUMX i17647 (.BLUT(n19975), .ALUT(n19976), .C0(index_i[4]), .Z(n19977));
    LUT4 mux_194_Mux_0_i1017_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .D(index_i[3]), .Z(n1017)) /* synthesis lut_function=(A (B (D)+!B !((D)+!C))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_0_i1017_4_lut_4_lut_4_lut.init = 16'hdd70;
    LUT4 i11025_2_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n844_adj_2943)) /* synthesis lut_function=(A (B+!(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11025_2_lut_3_lut_4_lut.init = 16'h9ff9;
    LUT4 i18451_3_lut (.A(n24995), .B(n27517), .C(index_i[3]), .Z(n20781)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18451_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_0_i731_3_lut_4_lut (.A(n24994), .B(index_i[2]), .C(index_i[3]), 
         .D(n27510), .Z(n731)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_0_i731_3_lut_4_lut.init = 16'h4f40;
    LUT4 i18447_3_lut (.A(n25142), .B(n27517), .C(index_i[3]), .Z(n20777)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18447_3_lut.init = 16'hcaca;
    LUT4 i18446_3_lut (.A(n25107), .B(n108), .C(index_i[3]), .Z(n20776)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18446_3_lut.init = 16'hcaca;
    LUT4 i12139_2_lut_rep_538 (.A(index_i[0]), .B(index_i[1]), .Z(n25098)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i12139_2_lut_rep_538.init = 16'heeee;
    LUT4 i19251_3_lut_4_lut (.A(n24994), .B(index_i[2]), .C(index_i[3]), 
         .D(n27504), .Z(n21581)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19251_3_lut_4_lut.init = 16'hf404;
    LUT4 i11163_2_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n635_adj_2857)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A (B (C+!(D))+!B (C+(D)))) */ ;
    defparam i11163_2_lut_4_lut_4_lut.init = 16'hf1fc;
    LUT4 mux_194_Mux_7_i924_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[4]), .D(n25111), .Z(n924_adj_2828)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B ((D)+!C))) */ ;
    defparam mux_194_Mux_7_i924_3_lut_3_lut_4_lut.init = 16'hf10f;
    LUT4 i11117_2_lut_rep_318_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n24878)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i11117_2_lut_rep_318_3_lut_4_lut.init = 16'hfef0;
    LUT4 i17621_3_lut_3_lut_4_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n19951)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B !((D)+!C)))) */ ;
    defparam i17621_3_lut_3_lut_4_lut_3_lut_4_lut.init = 16'h11ef;
    LUT4 mux_194_Mux_0_i923_3_lut (.A(n25101), .B(n27517), .C(index_i[3]), 
         .Z(n923)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_0_i923_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_5_i572_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n572_adj_3004)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A !(B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_5_i572_3_lut_4_lut_4_lut.init = 16'ha9a5;
    LUT4 i18445_3_lut (.A(n85), .B(n25099), .C(index_i[3]), .Z(n20775)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18445_3_lut.init = 16'hcaca;
    LUT4 i18444_3_lut (.A(n24996), .B(n25146), .C(index_i[3]), .Z(n20774)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18444_3_lut.init = 16'hcaca;
    LUT4 i9416_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[4]), .D(n25111), .Z(n189)) /* synthesis lut_function=(A (B (C (D)))+!A !(B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9416_3_lut_4_lut_4_lut_4_lut.init = 16'h9555;
    LUT4 i17663_3_lut_4_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n19993)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))+!A (B (C)+!B ((D)+!C))) */ ;
    defparam i17663_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'hf1e3;
    LUT4 i11098_2_lut_rep_418_3_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .Z(n24978)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i11098_2_lut_rep_418_3_lut.init = 16'he0e0;
    LUT4 i15279_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n17542)) /* synthesis lut_function=(A (B)+!A !(B (C (D))+!B !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i15279_3_lut_4_lut_4_lut.init = 16'h9ccc;
    LUT4 i17664_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n19994)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C+(D)))+!A (B (C (D)+!C !(D))+!B !(C)))) */ ;
    defparam i17664_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h3ef0;
    LUT4 i11006_2_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n668)) /* synthesis lut_function=(!(A ((D)+!B)+!A (B ((D)+!C)+!B (C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11006_2_lut_4_lut_4_lut_4_lut.init = 16'h00c9;
    LUT4 i11120_2_lut_rep_320_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[4]), .D(n25111), .Z(n24880)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i11120_2_lut_rep_320_3_lut_4_lut.init = 16'hfef0;
    LUT4 mux_194_Mux_2_i142_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n142_adj_2941)) /* synthesis lut_function=(!(A (B (D)+!B (C (D)+!C !(D)))+!A (B (D)+!B (C+!(D))))) */ ;
    defparam mux_194_Mux_2_i142_3_lut_4_lut_4_lut_4_lut.init = 16'h03ec;
    LUT4 mux_194_Mux_8_i460_3_lut_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n460_adj_2975)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B ((D)+!C))) */ ;
    defparam mux_194_Mux_8_i460_3_lut_3_lut_3_lut_4_lut.init = 16'hf10f;
    LUT4 mux_194_Mux_8_i236_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n236_adj_2980)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)+!C !(D)))+!A (B (C+!(D))+!B ((D)+!C))) */ ;
    defparam mux_194_Mux_8_i236_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hf1cf;
    LUT4 i19283_3_lut (.A(n24311), .B(n21612), .C(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2126[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19283_3_lut.init = 16'hcaca;
    LUT4 i18440_3_lut (.A(n27517), .B(n27509), .C(index_i[3]), .Z(n20770)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18440_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_2_i716_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n716_adj_2931)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)+!C !(D)))+!A (B (D)+!B !((D)+!C)))) */ ;
    defparam mux_194_Mux_2_i716_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h31cf;
    LUT4 i19282_3_lut (.A(n21609), .B(n21610), .C(index_i[8]), .Z(n21612)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19282_3_lut.init = 16'hcaca;
    LUT4 i18439_3_lut (.A(n1001), .B(n25142), .C(index_i[3]), .Z(n20769)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18439_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_7_i762_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n762_adj_2962)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A (B (C (D)+!C !(D))+!B !(C)))) */ ;
    defparam mux_194_Mux_7_i762_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h1cf0;
    LUT4 n262_bdd_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n27042)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C))+!A (B (C (D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n262_bdd_3_lut_4_lut.init = 16'h0fc7;
    LUT4 mux_194_Mux_3_i157_3_lut_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n157)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B !(C+(D))))) */ ;
    defparam mux_194_Mux_3_i157_3_lut_3_lut_3_lut_4_lut.init = 16'h1ff0;
    LUT4 i9390_3_lut_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n541_adj_2948)) /* synthesis lut_function=(A (B (C (D))+!B !(C (D)))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9390_3_lut_3_lut_4_lut_4_lut.init = 16'h9333;
    LUT4 mux_194_Mux_8_i101_3_lut_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n101)) /* synthesis lut_function=(!(A (B (C))+!A (B (C)+!B !(C)))) */ ;
    defparam mux_194_Mux_8_i101_3_lut_3_lut_3_lut.init = 16'h3e3e;
    LUT4 i17754_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n20084)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)+!C !(D)))+!A (B (C+!(D))+!B ((D)+!C)))) */ ;
    defparam i17754_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h0e30;
    LUT4 i17745_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n20075)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B ((D)+!C)+!B (C))) */ ;
    defparam i17745_3_lut_4_lut_4_lut.init = 16'hfc1c;
    LUT4 i18437_3_lut (.A(n27509), .B(n24996), .C(index_i[3]), .Z(n20767)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18437_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_0_i333_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n333)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B (D))) */ ;
    defparam mux_194_Mux_0_i333_3_lut_3_lut_4_lut.init = 16'hf10e;
    LUT4 mux_194_Mux_7_i572_3_lut_rep_258_3_lut_3_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n24818)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)+!C !(D)))) */ ;
    defparam mux_194_Mux_7_i572_3_lut_rep_258_3_lut_3_lut_4_lut.init = 16'hfe01;
    LUT4 mux_194_Mux_3_i30_3_lut_3_lut_4_lut_3_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n30_adj_2859)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C+!(D)))) */ ;
    defparam mux_194_Mux_3_i30_3_lut_3_lut_4_lut_3_lut_4_lut.init = 16'hfe11;
    LUT4 index_i_0__bdd_4_lut_23046 (.A(index_i[0]), .B(index_i[3]), .C(index_i[1]), 
         .D(index_i[2]), .Z(n25233)) /* synthesis lut_function=(A (B (C)+!B !(C+!(D)))+!A !(B ((D)+!C)+!B !(C (D)+!C !(D)))) */ ;
    defparam index_i_0__bdd_4_lut_23046.init = 16'h92c1;
    LUT4 mux_194_Mux_7_i141_3_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n141)) /* synthesis lut_function=(A ((C)+!B)+!A (B+!(C))) */ ;
    defparam mux_194_Mux_7_i141_3_lut_4_lut_3_lut.init = 16'he7e7;
    LUT4 mux_194_Mux_8_i46_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n46_adj_2867)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (D)+!B !(C (D)+!C !(D)))) */ ;
    defparam mux_194_Mux_8_i46_3_lut_4_lut_4_lut.init = 16'hcf10;
    LUT4 i1_2_lut_rep_444 (.A(index_i[6]), .B(index_i[7]), .Z(n25004)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i1_2_lut_rep_444.init = 16'heeee;
    LUT4 mux_194_Mux_2_i859_3_lut_4_lut (.A(index_i[0]), .B(n24997), .C(index_i[3]), 
         .D(n25137), .Z(n859_adj_2868)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_2_i859_3_lut_4_lut.init = 16'h4f40;
    L6MUX21 i22223 (.D0(n23828), .D1(n23826), .SD(index_i[5]), .Z(n23829));
    LUT4 index_i_5__bdd_3_lut_22292_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n23812)) /* synthesis lut_function=(A (B (C)+!B (C+(D)))+!A (B (C)+!B !(C (D)+!C !(D)))) */ ;
    defparam index_i_5__bdd_3_lut_22292_4_lut_4_lut_4_lut.init = 16'he3f0;
    LUT4 mux_194_Mux_4_i158_3_lut (.A(n142_adj_3005), .B(n157_adj_2984), 
         .C(index_i[4]), .Z(n158)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_4_i158_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_6_i573_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[4]), .D(n572_adj_3006), .Z(n573)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_6_i573_3_lut_4_lut.init = 16'hf909;
    LUT4 mux_194_Mux_7_i92_3_lut_rep_539 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n25099)) /* synthesis lut_function=(A (B+!(C))+!A !((C)+!B)) */ ;
    defparam mux_194_Mux_7_i92_3_lut_rep_539.init = 16'h8e8e;
    LUT4 i19280_3_lut (.A(n21605), .B(n22971), .C(index_i[7]), .Z(n21610)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19280_3_lut.init = 16'hcaca;
    LUT4 i17750_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n20080)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !(B (C+!(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i17750_3_lut_4_lut_4_lut.init = 16'ha5a9;
    LUT4 mux_194_Mux_0_i915_3_lut_rep_541 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n25101)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C)+!B !(C))) */ ;
    defparam mux_194_Mux_0_i915_3_lut_rep_541.init = 16'he3e3;
    PFUMX i22221 (.BLUT(n572_adj_3004), .ALUT(n23827), .C0(index_i[4]), 
          .Z(n23828));
    LUT4 i17646_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n19976)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A (B (D)+!B !(C (D))))) */ ;
    defparam i17646_3_lut_4_lut.init = 16'h18cc;
    LUT4 mux_194_Mux_0_i15_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n15_adj_2926)) /* synthesis lut_function=(A (B (C)+!B ((D)+!C))+!A (B (C)+!B !(C))) */ ;
    defparam mux_194_Mux_0_i15_3_lut_4_lut_4_lut.init = 16'he3c3;
    LUT4 mux_194_Mux_6_i498_3_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n404)) /* synthesis lut_function=(A (B+!(C))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_6_i498_3_lut_4_lut_3_lut.init = 16'h9b9b;
    PFUMX i22219 (.BLUT(n23825), .ALUT(n23824), .C0(index_i[4]), .Z(n23826));
    LUT4 i19250_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21580)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C (D)))+!A (B (C+(D))+!B !(C)))) */ ;
    defparam i19250_4_lut_4_lut_4_lut.init = 16'h301c;
    LUT4 mux_194_Mux_5_i109_3_lut_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .Z(n109_adj_2988)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_5_i109_3_lut_3_lut_3_lut.init = 16'h3939;
    LUT4 mux_194_Mux_0_i699_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n699)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (D))+!A (B (C+!(D))+!B !(C+!(D))))) */ ;
    defparam mux_194_Mux_0_i699_3_lut_3_lut_4_lut.init = 16'h1c33;
    LUT4 i17603_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n19933)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)))+!A !(B (C+!(D))+!B (D)))) */ ;
    defparam i17603_3_lut_3_lut_4_lut.init = 16'h71cc;
    LUT4 i9432_3_lut_4_lut (.A(index_i[0]), .B(n24997), .C(index_i[4]), 
         .D(n588), .Z(n11998)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9432_3_lut_4_lut.init = 16'h4f40;
    PFUMX i21458 (.BLUT(n23000), .ALUT(n22999), .C0(index_i[5]), .Z(n23001));
    LUT4 mux_194_Mux_0_i589_3_lut (.A(n27517), .B(n588), .C(index_i[3]), 
         .Z(n589)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_0_i589_3_lut.init = 16'hcaca;
    PFUMX i21435 (.BLUT(n22969), .ALUT(n22968), .C0(index_i[4]), .Z(n22970));
    LUT4 i11156_3_lut_3_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n13831)) /* synthesis lut_function=(!(A ((C+(D))+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11156_3_lut_3_lut_4_lut_4_lut.init = 16'h555d;
    L6MUX21 i22212 (.D0(n24800), .D1(n23814), .SD(index_i[4]), .Z(n23818));
    LUT4 i11139_3_lut_3_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n13813)) /* synthesis lut_function=(!(A+!(B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11139_3_lut_3_lut_4_lut_4_lut.init = 16'h4555;
    LUT4 mux_194_Mux_3_i142_3_lut_4_lut_3_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[1]), .Z(n142_adj_2935)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_3_i142_3_lut_4_lut_3_lut.init = 16'h6464;
    LUT4 i9592_3_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[4]), 
         .Z(n12162)) /* synthesis lut_function=(A (B)+!A !(B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9592_3_lut_4_lut_3_lut.init = 16'h9898;
    LUT4 i17328_4_lut (.A(n25094), .B(n892), .C(index_i[6]), .D(index_i[5]), 
         .Z(n19630)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D))))) */ ;
    defparam i17328_4_lut.init = 16'h3a35;
    L6MUX21 i18251 (.D0(n20579), .D1(n20580), .SD(index_i[8]), .Z(n20581));
    LUT4 i20901_3_lut (.A(n19630), .B(n17787), .C(index_i[7]), .Z(n20098)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20901_3_lut.init = 16'hcaca;
    LUT4 i17612_3_lut_4_lut (.A(index_i[0]), .B(n24997), .C(index_i[3]), 
         .D(n25131), .Z(n19942)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i17612_3_lut_4_lut.init = 16'hf404;
    LUT4 i12033_3_lut_3_lut (.A(index_i[2]), .B(index_i[0]), .C(index_i[1]), 
         .Z(n1001)) /* synthesis lut_function=(A (C)+!A (B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i12033_3_lut_3_lut.init = 16'hf4f4;
    PFUMX i22208 (.BLUT(n23813), .ALUT(n23812), .C0(index_i[5]), .Z(n23814));
    LUT4 i18695_3_lut_3_lut_4_lut (.A(n24952), .B(index_i[3]), .C(n93_adj_3007), 
         .D(index_i[4]), .Z(n21025)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18695_3_lut_3_lut_4_lut.init = 16'hf077;
    LUT4 mux_194_Mux_5_i924_4_lut_3_lut (.A(index_i[2]), .B(n14719), .C(index_i[4]), 
         .Z(n924_adj_2994)) /* synthesis lut_function=(!(A (B+(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_5_i924_4_lut_3_lut.init = 16'h5656;
    LUT4 mux_194_Mux_5_i251_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .Z(n251_adj_2983)) /* synthesis lut_function=(A (B)+!A (B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_5_i251_3_lut_3_lut.init = 16'hc9c9;
    LUT4 i17485_2_lut_rep_545 (.A(index_i[5]), .B(index_i[4]), .Z(n25105)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i17485_2_lut_rep_545.init = 16'h8888;
    LUT4 i11043_3_lut_4_lut (.A(index_i[5]), .B(index_i[4]), .C(index_i[6]), 
         .D(index_i[3]), .Z(n509)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11043_3_lut_4_lut.init = 16'hf8f0;
    LUT4 i15280_3_lut_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n17543)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i15280_3_lut_3_lut_4_lut_4_lut.init = 16'h3999;
    LUT4 mux_194_Mux_8_i172_3_lut_rep_676 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27516)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_8_i172_3_lut_rep_676.init = 16'h7c7c;
    LUT4 i11673_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[4]), 
         .C(n25111), .D(index_i[1]), .Z(n14348)) /* synthesis lut_function=(!(A (D)+!A !(B (C+!(D))+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11673_3_lut_4_lut_4_lut_4_lut.init = 16'h40ff;
    LUT4 mux_194_Mux_2_i507_3_lut_3_lut (.A(index_i[0]), .B(index_i[4]), 
         .C(n491_adj_3008), .Z(n507_adj_2919)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_2_i507_3_lut_3_lut.init = 16'h7474;
    LUT4 mux_194_Mux_4_i142_3_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[3]), 
         .C(index_i[2]), .Z(n142_adj_3005)) /* synthesis lut_function=(A (B (C))+!A !(B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_4_i142_3_lut_4_lut_3_lut.init = 16'h9595;
    LUT4 n130_bdd_3_lut_22541_4_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .Z(n22783)) /* synthesis lut_function=(A (B)+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n130_bdd_3_lut_22541_4_lut_3_lut.init = 16'hd9d9;
    LUT4 mux_194_Mux_2_i349_3_lut_3_lut (.A(index_i[0]), .B(index_i[4]), 
         .C(n348_adj_3003), .Z(n349_adj_2917)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_2_i349_3_lut_3_lut.init = 16'hd1d1;
    LUT4 mux_194_Mux_6_i645_3_lut_4_lut_3_lut_rep_581 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n25141)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_6_i645_3_lut_4_lut_3_lut_rep_581.init = 16'h1919;
    LUT4 mux_194_Mux_7_i45_3_lut_3_lut_3_lut_rep_582 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n25142)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_7_i45_3_lut_3_lut_3_lut_rep_582.init = 16'h3939;
    LUT4 mux_194_Mux_5_i573_3_lut_3_lut (.A(index_i[0]), .B(index_i[4]), 
         .C(n572_adj_3004), .Z(n573_adj_2861)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_5_i573_3_lut_3_lut.init = 16'hd1d1;
    LUT4 i11670_2_lut_rep_368_3_lut_3_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[1]), .Z(n24928)) /* synthesis lut_function=((B (C))+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11670_2_lut_rep_368_3_lut_3_lut.init = 16'hd5d5;
    LUT4 mux_194_Mux_0_i219_3_lut_3_lut_3_lut_rep_583 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n25143)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_0_i219_3_lut_3_lut_3_lut_rep_583.init = 16'h9393;
    LUT4 mux_194_Mux_0_i165_3_lut_4_lut_4_lut_3_lut_rep_584 (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[2]), .Z(n25144)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_0_i165_3_lut_4_lut_4_lut_3_lut_rep_584.init = 16'h9292;
    LUT4 mux_194_Mux_0_i985_3_lut_4_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[1]), .Z(n985)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_0_i985_3_lut_4_lut_4_lut_3_lut.init = 16'h1919;
    LUT4 mux_194_Mux_7_i77_3_lut_3_lut_rep_586 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n25146)) /* synthesis lut_function=(A (B)+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_7_i77_3_lut_3_lut_rep_586.init = 16'h9c9c;
    LUT4 mux_194_Mux_3_i700_3_lut_3_lut (.A(index_i[0]), .B(index_i[4]), 
         .C(n684_adj_2972), .Z(n700_adj_2908)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_3_i700_3_lut_3_lut.init = 16'h7474;
    LUT4 i9408_3_lut_4_lut_4_lut (.A(index_i[0]), .B(n25121), .C(index_i[4]), 
         .D(index_i[3]), .Z(n605_adj_2862)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A !(B+(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9408_3_lut_4_lut_4_lut.init = 16'h555c;
    LUT4 mux_194_Mux_4_i221_3_lut_3_lut (.A(index_i[0]), .B(index_i[4]), 
         .C(n205_adj_2999), .Z(n221_adj_2885)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_4_i221_3_lut_3_lut.init = 16'h7474;
    LUT4 mux_194_Mux_2_i763_4_lut_4_lut (.A(index_i[0]), .B(n11990), .C(index_i[4]), 
         .D(n157_adj_2846), .Z(n763_adj_2925)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_2_i763_4_lut_4_lut.init = 16'hdfd0;
    LUT4 mux_194_Mux_4_i262_3_lut_3_lut_rep_587 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n25147)) /* synthesis lut_function=(A (B+(C))+!A !(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_4_i262_3_lut_3_lut_rep_587.init = 16'ha9a9;
    L6MUX21 i18300 (.D0(n20625), .D1(n20626), .SD(index_i[7]), .Z(n20630));
    LUT4 i19463_3_lut_4_lut_4_lut (.A(index_i[0]), .B(n25121), .C(index_i[3]), 
         .D(n24998), .Z(n21793)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19463_3_lut_4_lut_4_lut.init = 16'hcfc5;
    LUT4 i11142_3_lut_3_lut_3_lut (.A(index_i[0]), .B(index_i[2]), .C(index_i[1]), 
         .Z(n85)) /* synthesis lut_function=(!(A (C)+!A !(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11142_3_lut_3_lut_3_lut.init = 16'h4f4f;
    LUT4 i11147_3_lut_3_lut_3_lut_rep_547 (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[1]), .Z(n25107)) /* synthesis lut_function=(!(A ((C)+!B)+!A (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11147_3_lut_3_lut_3_lut_rep_547.init = 16'h0d0d;
    LUT4 i17744_3_lut (.A(n25121), .B(n27501), .C(index_i[3]), .Z(n20074)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17744_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_3_i444_3_lut_4_lut (.A(index_i[0]), .B(index_i[3]), 
         .C(n24998), .D(index_i[4]), .Z(n444_adj_2902)) /* synthesis lut_function=(!(A (B (D)+!B (C (D)))+!A !(B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_3_i444_3_lut_4_lut.init = 16'h46aa;
    LUT4 mux_194_Mux_3_i676_3_lut_4_lut_3_lut_rep_588 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n25148)) /* synthesis lut_function=(A (B (C))+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_3_i676_3_lut_4_lut_3_lut_rep_588.init = 16'h9494;
    LUT4 mux_194_Mux_1_i732_3_lut (.A(n716_adj_2819), .B(n491_adj_2985), 
         .C(index_i[4]), .Z(n732)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_1_i732_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_4_i252_4_lut_4_lut (.A(index_i[0]), .B(index_i[3]), 
         .C(n24997), .D(index_i[4]), .Z(n252_adj_2886)) /* synthesis lut_function=(!(A (B (D)+!B !(D))+!A !(B ((D)+!C)+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_4_i252_4_lut_4_lut.init = 16'h669d;
    LUT4 i19238_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[2]), .C(index_i[1]), 
         .D(index_i[3]), .Z(n21568)) /* synthesis lut_function=(!(A ((C (D)+!C !(D))+!B)+!A (B (C (D)+!C !(D))+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19238_3_lut_4_lut_4_lut.init = 16'h0dc0;
    LUT4 i20340_3_lut (.A(n109), .B(n124_adj_3000), .C(index_i[4]), .Z(n20740)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20340_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_6_i134_3_lut_4_lut_3_lut_rep_589 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n25149)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_6_i134_3_lut_4_lut_3_lut_rep_589.init = 16'h9696;
    LUT4 mux_194_Mux_6_i564_3_lut_4_lut_3_lut_rep_590 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n25150)) /* synthesis lut_function=(A (B)+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_6_i564_3_lut_4_lut_3_lut_rep_590.init = 16'hd9d9;
    LUT4 mux_194_Mux_2_i908_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[1]), .D(index_i[3]), .Z(n908_adj_2814)) /* synthesis lut_function=(!(A (B (C)+!B !(C (D)))+!A (B (C)+!B !(C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_2_i908_3_lut_4_lut_4_lut.init = 16'h3c0d;
    LUT4 i1_2_lut_rep_551 (.A(index_i[3]), .B(index_i[2]), .Z(n25111)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i1_2_lut_rep_551.init = 16'h8888;
    L6MUX21 i22151 (.D0(n23753), .D1(n23750), .SD(index_i[5]), .Z(n23754));
    LUT4 mux_194_Mux_6_i356_3_lut_4_lut_3_lut_rep_591 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n25151)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_6_i356_3_lut_4_lut_3_lut_rep_591.init = 16'h4949;
    LUT4 mux_194_Mux_8_i205_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n205)) /* synthesis lut_function=(!(A (B (C)+!B !(C (D)+!C !(D)))+!A !(B ((D)+!C)+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_8_i205_3_lut_3_lut_4_lut.init = 16'h7c0f;
    LUT4 mux_194_Mux_0_i660_3_lut_rep_592 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n25152)) /* synthesis lut_function=(A (B)+!A (B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_0_i660_3_lut_rep_592.init = 16'hc9c9;
    PFUMX i22149 (.BLUT(n23752), .ALUT(n23751), .C0(index_i[4]), .Z(n23753));
    LUT4 i12215_2_lut_rep_400_3_lut_4_lut (.A(index_i[3]), .B(index_i[2]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n24960)) /* synthesis lut_function=(A (B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i12215_2_lut_rep_400_3_lut_4_lut.init = 16'h8880;
    LUT4 i12161_2_lut_rep_365_3_lut (.A(index_i[3]), .B(index_i[2]), .C(index_i[1]), 
         .Z(n24925)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i12161_2_lut_rep_365_3_lut.init = 16'h8080;
    LUT4 mux_194_Mux_0_i134_3_lut_4_lut_3_lut_rep_593 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n25153)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_0_i134_3_lut_4_lut_3_lut_rep_593.init = 16'h6969;
    LUT4 mux_194_Mux_0_i716_3_lut (.A(n25119), .B(n25154), .C(index_i[3]), 
         .Z(n716)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_0_i716_3_lut.init = 16'hcaca;
    LUT4 i18332_3_lut_3_lut_3_lut_4_lut (.A(index_i[3]), .B(index_i[2]), 
         .C(index_i[4]), .D(index_i[1]), .Z(n20662)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18332_3_lut_3_lut_3_lut_4_lut.init = 16'h878f;
    LUT4 mux_194_Mux_0_i715_3_lut_rep_594 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n25154)) /* synthesis lut_function=(A (B (C))+!A !(B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_0_i715_3_lut_rep_594.init = 16'h9595;
    PFUMX i9386 (.BLUT(n12165), .ALUT(n12166), .C0(n19862), .Z(n11952));
    PFUMX i19416 (.BLUT(n21744), .ALUT(n21745), .C0(index_i[8]), .Z(n21746));
    LUT4 i11674_2_lut_2_lut_3_lut (.A(index_i[3]), .B(index_i[2]), .C(index_i[0]), 
         .Z(n14349)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11674_2_lut_2_lut_3_lut.init = 16'h0808;
    LUT4 i17532_1_lut_2_lut (.A(index_i[3]), .B(index_i[2]), .Z(n19862)) /* synthesis lut_function=(!(A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i17532_1_lut_2_lut.init = 16'h7777;
    PFUMX i22146 (.BLUT(n301_adj_2981), .ALUT(n23749), .C0(index_i[4]), 
          .Z(n23750));
    LUT4 mux_194_Mux_1_i93_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n93_adj_2929)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C+(D)))+!A !(B (C (D)+!C !(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_1_i93_3_lut_4_lut_4_lut.init = 16'h955a;
    LUT4 i2_2_lut_rep_401_3_lut_4_lut (.A(index_i[3]), .B(index_i[2]), .C(index_i[1]), 
         .D(index_i[0]), .Z(n24961)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i2_2_lut_rep_401_3_lut_4_lut.init = 16'h8000;
    LUT4 i3044_2_lut_rep_552 (.A(index_i[0]), .B(index_i[2]), .Z(n25112)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i3044_2_lut_rep_552.init = 16'h6666;
    LUT4 mux_194_Mux_1_i62_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[4]), .D(index_i[3]), .Z(n62_adj_2995)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))+!A !(B (C)+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_1_i62_3_lut_4_lut_4_lut.init = 16'ha5a6;
    LUT4 i20736_3_lut (.A(n286_adj_2998), .B(n317), .C(index_i[5]), .Z(n21650)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20736_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_4_i349_3_lut_4_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[4]), .D(n348_adj_2954), .Z(n349_adj_2889)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_4_i349_3_lut_4_lut.init = 16'hf606;
    LUT4 i20848_3_lut (.A(n11945), .B(n892_adj_2937), .C(index_i[6]), 
         .Z(n21626)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20848_3_lut.init = 16'hcaca;
    LUT4 i15292_3_lut_3_lut (.A(index_i[0]), .B(index_i[2]), .C(index_i[3]), 
         .Z(n17555)) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i15292_3_lut_3_lut.init = 16'h6a6a;
    PFUMX i17665 (.BLUT(n19993), .ALUT(n19994), .C0(index_i[4]), .Z(n19995));
    LUT4 mux_194_Mux_0_i142_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n142)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C))+!A !(B (C (D)+!C !(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_0_i142_3_lut_4_lut_4_lut.init = 16'ha569;
    PFUMX i19240 (.BLUT(n21568), .ALUT(n21569), .C0(index_i[4]), .Z(n21570));
    LUT4 i20335_3_lut (.A(n21799), .B(n21800), .C(index_i[4]), .Z(n21801)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20335_3_lut.init = 16'hcaca;
    LUT4 i19288_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21618)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C+(D)))+!A (B (C)+!B !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19288_3_lut_4_lut_4_lut.init = 16'hc95a;
    LUT4 i17741_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n20071)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (D))+!A !(B (C (D))+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i17741_3_lut_3_lut_4_lut.init = 16'h4933;
    LUT4 mux_194_Mux_6_i572_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n572_adj_3006)) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_6_i572_3_lut_4_lut.init = 16'hccd9;
    LUT4 i19466_3_lut (.A(n25138), .B(n27501), .C(index_i[3]), .Z(n21796)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19466_3_lut.init = 16'hcaca;
    PFUMX i19249 (.BLUT(n21577), .ALUT(n21578), .C0(index_i[4]), .Z(n21579));
    L6MUX21 i22137 (.D0(n23739), .D1(n23736), .SD(index_i[5]), .Z(n23740));
    PFUMX i22135 (.BLUT(n15_adj_2971), .ALUT(n23737), .C0(index_i[4]), 
          .Z(n23739));
    PFUMX i19252 (.BLUT(n21580), .ALUT(n21581), .C0(index_i[4]), .Z(n21582));
    LUT4 i17757_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n20087)) /* synthesis lut_function=(A (B (C+(D))+!B ((D)+!C))+!A !(B (C+(D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i17757_3_lut_4_lut.init = 16'haa96;
    LUT4 mux_194_Mux_5_i700_3_lut (.A(n460_adj_2986), .B(n25153), .C(index_i[4]), 
         .Z(n700_adj_2870)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_5_i700_3_lut.init = 16'hcaca;
    LUT4 n676_bdd_3_lut_22927_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n23712)) /* synthesis lut_function=(A (B (C+(D)))+!A (B ((D)+!C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n676_bdd_3_lut_22927_4_lut.init = 16'hcc94;
    LUT4 i19460_3_lut (.A(n325), .B(n27501), .C(index_i[3]), .Z(n21790)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19460_3_lut.init = 16'hcaca;
    PFUMX i22132 (.BLUT(n23735), .ALUT(n23734), .C0(index_i[4]), .Z(n23736));
    LUT4 mux_194_Mux_2_i653_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n653_adj_2933)) /* synthesis lut_function=(A (B (C+!(D))+!B !(D))+!A !(B (C+!(D))+!B !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_2_i653_3_lut_4_lut.init = 16'h94aa;
    LUT4 i19272_3_lut (.A(n21589), .B(n23699), .C(index_i[6]), .Z(n21602)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19272_3_lut.init = 16'hcaca;
    LUT4 i19458_3_lut (.A(n25151), .B(n27502), .C(index_i[3]), .Z(n21788)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19458_3_lut.init = 16'hcaca;
    LUT4 i17609_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n19939)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A !(B (D)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i17609_3_lut_3_lut_4_lut.init = 16'ha955;
    LUT4 i19457_3_lut (.A(n25152), .B(n27505), .C(index_i[3]), .Z(n21787)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19457_3_lut.init = 16'hcaca;
    PFUMX i19286 (.BLUT(n21614), .ALUT(n21615), .C0(index_i[4]), .Z(n21616));
    LUT4 mux_194_Mux_3_i397_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n397_adj_2951)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !(B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_3_i397_3_lut_4_lut_4_lut.init = 16'ha95a;
    LUT4 mux_194_Mux_3_i859_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n859)) /* synthesis lut_function=(!(A (B (D)+!B !(D))+!A (B (C+(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_3_i859_3_lut_3_lut_4_lut.init = 16'h339c;
    LUT4 n781_bdd_3_lut_4_lut_4_lut (.A(index_i[3]), .B(n781_adj_2809), 
         .C(index_i[4]), .D(n24891), .Z(n22867)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B ((D)+!C)+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n781_bdd_3_lut_4_lut_4_lut.init = 16'h5c0c;
    LUT4 i8609_4_lut_4_lut (.A(index_i[3]), .B(index_i[0]), .C(index_i[1]), 
         .D(index_i[2]), .Z(n11113)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (D)+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i8609_4_lut_4_lut.init = 16'h0bf4;
    L6MUX21 i22115 (.D0(n23715), .D1(n23713), .SD(index_i[5]), .Z(n23716));
    LUT4 i11143_2_lut_3_lut_3_lut (.A(index_i[3]), .B(index_i[1]), .C(index_i[0]), 
         .Z(n13817)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11143_2_lut_3_lut_3_lut.init = 16'h4040;
    PFUMX i22113 (.BLUT(n23714), .ALUT(n20087), .C0(index_i[4]), .Z(n23715));
    LUT4 i11026_4_lut_4_lut (.A(index_i[3]), .B(index_i[2]), .C(index_i[0]), 
         .D(index_i[1]), .Z(n875)) /* synthesis lut_function=((B (C)+!B (D))+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11026_4_lut_4_lut.init = 16'hf7d5;
    LUT4 i18330_3_lut_4_lut_3_lut (.A(index_i[3]), .B(index_i[4]), .C(n24952), 
         .Z(n20660)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18330_3_lut_4_lut_3_lut.init = 16'h6464;
    LUT4 mux_194_Mux_1_i890_4_lut_4_lut_4_lut_4_lut (.A(index_i[3]), .B(index_i[4]), 
         .C(n24996), .D(index_i[0]), .Z(n890_adj_2992)) /* synthesis lut_function=(!(A (B (D)+!B !(C))+!A (B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_1_i890_4_lut_4_lut_4_lut_4_lut.init = 16'h31fd;
    PFUMX i22111 (.BLUT(n23712), .ALUT(n23711), .C0(index_i[4]), .Z(n23713));
    LUT4 mux_194_Mux_2_i221_4_lut_4_lut (.A(index_i[3]), .B(index_i[4]), 
         .C(n24892), .D(n24866), .Z(n221_adj_2914)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (B+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_2_i221_4_lut_4_lut.init = 16'hf7c4;
    LUT4 i18483_4_lut_3_lut (.A(index_i[3]), .B(index_i[4]), .C(n24892), 
         .Z(n20813)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18483_4_lut_3_lut.init = 16'h6565;
    LUT4 i9379_3_lut_3_lut (.A(index_i[3]), .B(index_i[4]), .C(n11944), 
         .Z(n11945)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9379_3_lut_3_lut.init = 16'h7474;
    L6MUX21 i22109 (.D0(n23709), .D1(n23707), .SD(index_i[4]), .Z(n23710));
    PFUMX i22107 (.BLUT(n24866), .ALUT(n23708), .C0(index_i[5]), .Z(n23709));
    LUT4 mux_194_Mux_3_i94_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[4]), .D(n93_adj_2953), .Z(n94_adj_2895)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_3_i94_3_lut_4_lut.init = 16'hf606;
    PFUMX i22105 (.BLUT(n23706), .ALUT(n23705), .C0(index_i[5]), .Z(n23707));
    LUT4 mux_194_Mux_3_i62_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[4]), .D(n812_adj_2990), .Z(n62_adj_2996)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_3_i62_3_lut_4_lut.init = 16'h6f60;
    LUT4 i17894_4_lut_4_lut (.A(index_i[4]), .B(index_i[5]), .C(n25250), 
         .D(n908_adj_2814), .Z(n20224)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam i17894_4_lut_4_lut.init = 16'hd1c0;
    PFUMX i19313 (.BLUT(n21641), .ALUT(n21642), .C0(index_i[4]), .Z(n21643));
    L6MUX21 i22097 (.D0(n23698), .D1(n23695), .SD(index_i[5]), .Z(n23699));
    PFUMX i22095 (.BLUT(n23697), .ALUT(n475_adj_2934), .C0(index_i[4]), 
          .Z(n23698));
    PFUMX i22092 (.BLUT(n23694), .ALUT(n23693), .C0(index_i[4]), .Z(n23695));
    LUT4 mux_194_Mux_0_i762_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n762)) /* synthesis lut_function=(A (B+!((D)+!C))+!A !(B (D)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_0_i762_3_lut_4_lut_4_lut.init = 16'h98fc;
    L6MUX21 i22076 (.D0(n23678), .D1(n23676), .SD(index_i[5]), .Z(n23679));
    PFUMX i22074 (.BLUT(n23677), .ALUT(n285), .C0(index_i[4]), .Z(n23678));
    PFUMX i22072 (.BLUT(n23675), .ALUT(n23674), .C0(index_i[4]), .Z(n23676));
    LUT4 i3055_2_lut_rep_557 (.A(index_i[0]), .B(index_i[1]), .Z(n25117)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i3055_2_lut_rep_557.init = 16'h6666;
    PFUMX i22069 (.BLUT(n23672), .ALUT(n25112), .C0(index_i[4]), .Z(n23673));
    LUT4 mux_194_Mux_0_i747_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n747)) /* synthesis lut_function=(!(A (B+!(C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_0_i747_3_lut_4_lut_4_lut_4_lut.init = 16'h6556;
    LUT4 mux_194_Mux_1_i746_3_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n746)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_1_i746_3_lut_4_lut_3_lut.init = 16'h8686;
    LUT4 i20986_2_lut_rep_467 (.A(index_i[1]), .B(index_i[2]), .Z(n25027)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20986_2_lut_rep_467.init = 16'h9999;
    LUT4 i17902_3_lut (.A(n23818), .B(n20223), .C(index_i[6]), .Z(n20232)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17902_3_lut.init = 16'hcaca;
    LUT4 mux_194_Mux_0_i812_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n812)) /* synthesis lut_function=(A (B (C+(D))+!B !(C))+!A (B (D)+!B !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_0_i812_3_lut_4_lut_4_lut_4_lut.init = 16'hcf92;
    LUT4 mux_194_Mux_0_i93_3_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .Z(n93_adj_3007)) /* synthesis lut_function=(A (B)+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_0_i93_3_lut_3_lut.init = 16'h9c9c;
    LUT4 n22_bdd_2_lut_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[3]), 
         .Z(n23824)) /* synthesis lut_function=(A (B+(C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n22_bdd_2_lut_3_lut.init = 16'hf9f9;
    LUT4 mux_194_Mux_5_i828_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[4]), .D(n25093), .Z(n828_adj_2873)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_5_i828_4_lut_4_lut.init = 16'hc66c;
    LUT4 i17624_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n19954)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C))+!A !(B ((D)+!C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i17624_3_lut_4_lut_4_lut.init = 16'h925a;
    LUT4 i21088_2_lut_rep_469 (.A(index_i[4]), .B(index_i[3]), .Z(n25029)) /* synthesis lut_function=(A+!(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i21088_2_lut_rep_469.init = 16'hbbbb;
    LUT4 i9402_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(n25111), .D(index_i[4]), .Z(n221)) /* synthesis lut_function=(!(A (B)+!A (B (C+(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9402_3_lut_4_lut_4_lut_4_lut.init = 16'h3336;
    LUT4 i9418_3_lut_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[4]), .D(index_i[3]), .Z(n444_adj_2903)) /* synthesis lut_function=(!(A (B)+!A !(B (C (D))+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9418_3_lut_3_lut_4_lut_4_lut.init = 16'h6333;
    LUT4 i20729_3_lut_4_lut (.A(index_i[4]), .B(index_i[3]), .C(n25277), 
         .D(n746), .Z(n763)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20729_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_194_Mux_2_i731_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n731_adj_2932)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_2_i731_3_lut_4_lut_4_lut.init = 16'h6cc6;
    LUT4 i19247_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21577)) /* synthesis lut_function=(A (B (C)+!B (C (D)+!C !(D)))+!A !(B (C+!(D))+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19247_3_lut_4_lut_4_lut.init = 16'ha593;
    LUT4 i19423_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21753)) /* synthesis lut_function=(A (B (C (D))+!B !(C (D)))+!A !(B (D)+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19423_3_lut_4_lut_4_lut.init = 16'h9366;
    LUT4 i11996_2_lut_rep_470 (.A(index_i[2]), .B(index_i[0]), .Z(n25030)) /* synthesis lut_function=(A (B)) */ ;
    defparam i11996_2_lut_rep_470.init = 16'h8888;
    LUT4 mux_194_Mux_7_i108_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n108)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_7_i108_3_lut_3_lut.init = 16'hc6c6;
    LUT4 mux_194_Mux_3_i507_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[4]), .D(n491_adj_2956), .Z(n507_adj_2905)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_3_i507_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_194_Mux_2_i604_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n604_adj_2936)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)+!C !(D)))+!A (B (D)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_2_i604_3_lut_4_lut_4_lut_4_lut.init = 16'h39cf;
    LUT4 mux_194_Mux_0_i236_3_lut_3_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[3]), .Z(n236)) /* synthesis lut_function=(A (B+(C))+!A !(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_0_i236_3_lut_3_lut.init = 16'ha9a9;
    LUT4 mux_194_Mux_1_i882_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n882)) /* synthesis lut_function=(A ((C)+!B)+!A !((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_1_i882_3_lut_3_lut.init = 16'ha6a6;
    LUT4 i19417_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21747)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(D))+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19417_3_lut_3_lut_4_lut.init = 16'h3319;
    LUT4 i11050_3_lut_4_lut (.A(n24892), .B(index_i[3]), .C(n25105), .D(index_i[6]), 
         .Z(n765)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11050_3_lut_4_lut.init = 16'hffe0;
    LUT4 i9388_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n526_adj_2991)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+(D)))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9388_3_lut_4_lut_4_lut.init = 16'h666c;
    LUT4 n61_bdd_3_lut_22936_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n23708)) /* synthesis lut_function=(!(A (B)+!A !(B (C+(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n61_bdd_3_lut_22936_3_lut_4_lut_4_lut.init = 16'h6663;
    LUT4 mux_194_Mux_0_i645_3_lut_3_lut_rep_436_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n24996)) /* synthesis lut_function=(!(A (B)+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_0_i645_3_lut_3_lut_rep_436_3_lut.init = 16'h6363;
    LUT4 i9595_3_lut_4_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[4]), .Z(n12165)) /* synthesis lut_function=(!(A (B)+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9595_3_lut_4_lut_4_lut_3_lut.init = 16'h6262;
    PFUMX i18723 (.BLUT(n21051), .ALUT(n21052), .C0(index_i[8]), .Z(n21053));
    LUT4 i9593_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n12163)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B ((D)+!C)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9593_3_lut_4_lut_4_lut.init = 16'h6c3c;
    LUT4 mux_194_Mux_0_i588_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n588)) /* synthesis lut_function=(!(A (B+(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_0_i588_3_lut_3_lut.init = 16'h5656;
    LUT4 mux_194_Mux_5_i754_3_lut_4_lut_4_lut_3_lut_rep_559 (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[2]), .Z(n25119)) /* synthesis lut_function=(!(A (B)+!A ((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_5_i754_3_lut_4_lut_4_lut_3_lut_rep_559.init = 16'h2626;
    LUT4 mux_194_Mux_5_i53_3_lut_4_lut_3_lut_rep_560 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n25120)) /* synthesis lut_function=(A ((C)+!B)+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_5_i53_3_lut_4_lut_3_lut_rep_560.init = 16'he6e6;
    LUT4 mux_194_Mux_0_i525_3_lut_3_lut_rep_561 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n25121)) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_0_i525_3_lut_3_lut_rep_561.init = 16'h6a6a;
    LUT4 mux_194_Mux_2_i491_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n491_adj_3008)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A !(B (C)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_2_i491_3_lut_4_lut_4_lut.init = 16'h6a5a;
    L6MUX21 i21363 (.D0(n22868), .D1(n22866), .SD(index_i[6]), .Z(n22869));
    FD1S3BX quarter_wave_sample_register_i_i14 (.D(quarter_wave_sample_register_i_15__N_2126[14]), 
            .CK(i_ref_clk_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_i[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i14.GSR = "DISABLED";
    PFUMX i17746 (.BLUT(n20074), .ALUT(n20075), .C0(index_i[4]), .Z(n20076));
    LUT4 mux_194_Mux_6_i635_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n635_adj_2989)) /* synthesis lut_function=(A (B (C+(D))+!B !(D))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_194_Mux_6_i635_3_lut_4_lut.init = 16'hcce6;
    LUT4 i17615_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n19945)) /* synthesis lut_function=(!(A (B)+!A (B (C+(D))+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i17615_3_lut_3_lut_4_lut.init = 16'h3326;
    FD1S3BX quarter_wave_sample_register_i_i13 (.D(quarter_wave_sample_register_i_15__N_2126[13]), 
            .CK(i_ref_clk_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_i[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i13.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i12 (.D(quarter_wave_sample_register_i_15__N_2126[12]), 
            .CK(i_ref_clk_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_i[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i12.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i11 (.D(quarter_wave_sample_register_i_15__N_2126[11]), 
            .CK(i_ref_clk_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_i[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i11.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i10 (.D(quarter_wave_sample_register_i_15__N_2126[10]), 
            .CK(i_ref_clk_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_i[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i10.GSR = "DISABLED";
    PFUMX i21359 (.BLUT(n62), .ALUT(n22865), .C0(index_i[5]), .Z(n22866));
    PFUMX i21361 (.BLUT(n22867), .ALUT(n20813), .C0(index_i[5]), .Z(n22868));
    
endmodule
//
// Verilog Description of module \nco(OW=12) 
//

module \nco(OW=12)  (i_ref_clk_c, i_resetb_N_301, increment, o_phase, 
            GND_net) /* synthesis syn_module_defined=1 */ ;
    input i_ref_clk_c;
    input i_resetb_N_301;
    input [30:0]increment;
    output [11:0]o_phase;
    input GND_net;
    
    wire i_ref_clk_c /* synthesis SET_AS_NETWORK=i_ref_clk_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(22[12:21])
    wire [31:0]n233;
    wire [31:0]n133;
    
    wire n17417, n17416, n17415, n17414, n17413, n17412, n17411, 
        n17410, n17409, n17408, n17407, n17406, n17405, n17404, 
        n17403;
    
    FD1S3DX phase_register_507__i0 (.D(n133[0]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(n233[0])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_507__i0.GSR = "DISABLED";
    CCU2D phase_register_507_add_4_32 (.A0(increment[30]), .B0(o_phase[10]), 
          .C0(GND_net), .D0(GND_net), .A1(o_phase[11]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n17417), .S0(n133[30]), .S1(n133[31]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_507_add_4_32.INIT0 = 16'h5666;
    defparam phase_register_507_add_4_32.INIT1 = 16'hfaaa;
    defparam phase_register_507_add_4_32.INJECT1_0 = "NO";
    defparam phase_register_507_add_4_32.INJECT1_1 = "NO";
    CCU2D phase_register_507_add_4_30 (.A0(increment[28]), .B0(o_phase[8]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[29]), .B1(o_phase[9]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17416), .COUT(n17417), .S0(n133[28]), 
          .S1(n133[29]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_507_add_4_30.INIT0 = 16'h5666;
    defparam phase_register_507_add_4_30.INIT1 = 16'h5666;
    defparam phase_register_507_add_4_30.INJECT1_0 = "NO";
    defparam phase_register_507_add_4_30.INJECT1_1 = "NO";
    CCU2D phase_register_507_add_4_28 (.A0(increment[26]), .B0(o_phase[6]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[27]), .B1(o_phase[7]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17415), .COUT(n17416), .S0(n133[26]), 
          .S1(n133[27]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_507_add_4_28.INIT0 = 16'h5666;
    defparam phase_register_507_add_4_28.INIT1 = 16'h5666;
    defparam phase_register_507_add_4_28.INJECT1_0 = "NO";
    defparam phase_register_507_add_4_28.INJECT1_1 = "NO";
    CCU2D phase_register_507_add_4_26 (.A0(increment[24]), .B0(o_phase[4]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[25]), .B1(o_phase[5]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17414), .COUT(n17415), .S0(n133[24]), 
          .S1(n133[25]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_507_add_4_26.INIT0 = 16'h5666;
    defparam phase_register_507_add_4_26.INIT1 = 16'h5666;
    defparam phase_register_507_add_4_26.INJECT1_0 = "NO";
    defparam phase_register_507_add_4_26.INJECT1_1 = "NO";
    CCU2D phase_register_507_add_4_24 (.A0(increment[22]), .B0(o_phase[2]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[23]), .B1(o_phase[3]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17413), .COUT(n17414), .S0(n133[22]), 
          .S1(n133[23]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_507_add_4_24.INIT0 = 16'h5666;
    defparam phase_register_507_add_4_24.INIT1 = 16'h5666;
    defparam phase_register_507_add_4_24.INJECT1_0 = "NO";
    defparam phase_register_507_add_4_24.INJECT1_1 = "NO";
    CCU2D phase_register_507_add_4_22 (.A0(increment[20]), .B0(o_phase[0]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[21]), .B1(o_phase[1]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17412), .COUT(n17413), .S0(n133[20]), 
          .S1(n133[21]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_507_add_4_22.INIT0 = 16'h5666;
    defparam phase_register_507_add_4_22.INIT1 = 16'h5666;
    defparam phase_register_507_add_4_22.INJECT1_0 = "NO";
    defparam phase_register_507_add_4_22.INJECT1_1 = "NO";
    CCU2D phase_register_507_add_4_20 (.A0(increment[18]), .B0(n233[18]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[19]), .B1(n233[19]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17411), .COUT(n17412), .S0(n133[18]), 
          .S1(n133[19]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_507_add_4_20.INIT0 = 16'h5666;
    defparam phase_register_507_add_4_20.INIT1 = 16'h5666;
    defparam phase_register_507_add_4_20.INJECT1_0 = "NO";
    defparam phase_register_507_add_4_20.INJECT1_1 = "NO";
    CCU2D phase_register_507_add_4_18 (.A0(increment[16]), .B0(n233[16]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[17]), .B1(n233[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17410), .COUT(n17411), .S0(n133[16]), 
          .S1(n133[17]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_507_add_4_18.INIT0 = 16'h5666;
    defparam phase_register_507_add_4_18.INIT1 = 16'h5666;
    defparam phase_register_507_add_4_18.INJECT1_0 = "NO";
    defparam phase_register_507_add_4_18.INJECT1_1 = "NO";
    CCU2D phase_register_507_add_4_16 (.A0(increment[14]), .B0(n233[14]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[15]), .B1(n233[15]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17409), .COUT(n17410), .S0(n133[14]), 
          .S1(n133[15]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_507_add_4_16.INIT0 = 16'h5666;
    defparam phase_register_507_add_4_16.INIT1 = 16'h5666;
    defparam phase_register_507_add_4_16.INJECT1_0 = "NO";
    defparam phase_register_507_add_4_16.INJECT1_1 = "NO";
    CCU2D phase_register_507_add_4_14 (.A0(increment[12]), .B0(n233[12]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[13]), .B1(n233[13]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17408), .COUT(n17409), .S0(n133[12]), 
          .S1(n133[13]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_507_add_4_14.INIT0 = 16'h5666;
    defparam phase_register_507_add_4_14.INIT1 = 16'h5666;
    defparam phase_register_507_add_4_14.INJECT1_0 = "NO";
    defparam phase_register_507_add_4_14.INJECT1_1 = "NO";
    CCU2D phase_register_507_add_4_12 (.A0(increment[10]), .B0(n233[10]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[11]), .B1(n233[11]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17407), .COUT(n17408), .S0(n133[10]), 
          .S1(n133[11]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_507_add_4_12.INIT0 = 16'h5666;
    defparam phase_register_507_add_4_12.INIT1 = 16'h5666;
    defparam phase_register_507_add_4_12.INJECT1_0 = "NO";
    defparam phase_register_507_add_4_12.INJECT1_1 = "NO";
    CCU2D phase_register_507_add_4_10 (.A0(increment[8]), .B0(n233[8]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[9]), .B1(n233[9]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17406), .COUT(n17407), .S0(n133[8]), 
          .S1(n133[9]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_507_add_4_10.INIT0 = 16'h5666;
    defparam phase_register_507_add_4_10.INIT1 = 16'h5666;
    defparam phase_register_507_add_4_10.INJECT1_0 = "NO";
    defparam phase_register_507_add_4_10.INJECT1_1 = "NO";
    CCU2D phase_register_507_add_4_8 (.A0(increment[6]), .B0(n233[6]), .C0(GND_net), 
          .D0(GND_net), .A1(increment[7]), .B1(n233[7]), .C1(GND_net), 
          .D1(GND_net), .CIN(n17405), .COUT(n17406), .S0(n133[6]), .S1(n133[7]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_507_add_4_8.INIT0 = 16'h5666;
    defparam phase_register_507_add_4_8.INIT1 = 16'h5666;
    defparam phase_register_507_add_4_8.INJECT1_0 = "NO";
    defparam phase_register_507_add_4_8.INJECT1_1 = "NO";
    CCU2D phase_register_507_add_4_6 (.A0(increment[4]), .B0(n233[4]), .C0(GND_net), 
          .D0(GND_net), .A1(increment[5]), .B1(n233[5]), .C1(GND_net), 
          .D1(GND_net), .CIN(n17404), .COUT(n17405), .S0(n133[4]), .S1(n133[5]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_507_add_4_6.INIT0 = 16'h5666;
    defparam phase_register_507_add_4_6.INIT1 = 16'h5666;
    defparam phase_register_507_add_4_6.INJECT1_0 = "NO";
    defparam phase_register_507_add_4_6.INJECT1_1 = "NO";
    CCU2D phase_register_507_add_4_4 (.A0(increment[2]), .B0(n233[2]), .C0(GND_net), 
          .D0(GND_net), .A1(increment[3]), .B1(n233[3]), .C1(GND_net), 
          .D1(GND_net), .CIN(n17403), .COUT(n17404), .S0(n133[2]), .S1(n133[3]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_507_add_4_4.INIT0 = 16'h5666;
    defparam phase_register_507_add_4_4.INIT1 = 16'h5666;
    defparam phase_register_507_add_4_4.INJECT1_0 = "NO";
    defparam phase_register_507_add_4_4.INJECT1_1 = "NO";
    CCU2D phase_register_507_add_4_2 (.A0(increment[0]), .B0(n233[0]), .C0(GND_net), 
          .D0(GND_net), .A1(increment[1]), .B1(n233[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n17403), .S1(n133[1]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_507_add_4_2.INIT0 = 16'h7000;
    defparam phase_register_507_add_4_2.INIT1 = 16'h5666;
    defparam phase_register_507_add_4_2.INJECT1_0 = "NO";
    defparam phase_register_507_add_4_2.INJECT1_1 = "NO";
    LUT4 i15206_2_lut (.A(increment[0]), .B(n233[0]), .Z(n133[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i15206_2_lut.init = 16'h6666;
    FD1S3DX phase_register_507__i31 (.D(n133[31]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(o_phase[11])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_507__i31.GSR = "DISABLED";
    FD1S3DX phase_register_507__i30 (.D(n133[30]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(o_phase[10])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_507__i30.GSR = "DISABLED";
    FD1S3DX phase_register_507__i29 (.D(n133[29]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(o_phase[9])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_507__i29.GSR = "DISABLED";
    FD1S3DX phase_register_507__i28 (.D(n133[28]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(o_phase[8])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_507__i28.GSR = "DISABLED";
    FD1S3DX phase_register_507__i27 (.D(n133[27]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(o_phase[7])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_507__i27.GSR = "DISABLED";
    FD1S3DX phase_register_507__i26 (.D(n133[26]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(o_phase[6])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_507__i26.GSR = "DISABLED";
    FD1S3DX phase_register_507__i25 (.D(n133[25]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(o_phase[5])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_507__i25.GSR = "DISABLED";
    FD1S3DX phase_register_507__i24 (.D(n133[24]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(o_phase[4])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_507__i24.GSR = "DISABLED";
    FD1S3DX phase_register_507__i23 (.D(n133[23]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(o_phase[3])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_507__i23.GSR = "DISABLED";
    FD1S3DX phase_register_507__i22 (.D(n133[22]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(o_phase[2])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_507__i22.GSR = "DISABLED";
    FD1S3DX phase_register_507__i21 (.D(n133[21]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(o_phase[1])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_507__i21.GSR = "DISABLED";
    FD1S3DX phase_register_507__i20 (.D(n133[20]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(o_phase[0])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_507__i20.GSR = "DISABLED";
    FD1S3DX phase_register_507__i19 (.D(n133[19]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(n233[19])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_507__i19.GSR = "DISABLED";
    FD1S3DX phase_register_507__i18 (.D(n133[18]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(n233[18])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_507__i18.GSR = "DISABLED";
    FD1S3DX phase_register_507__i17 (.D(n133[17]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(n233[17])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_507__i17.GSR = "DISABLED";
    FD1S3DX phase_register_507__i16 (.D(n133[16]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(n233[16])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_507__i16.GSR = "DISABLED";
    FD1S3DX phase_register_507__i15 (.D(n133[15]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(n233[15])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_507__i15.GSR = "DISABLED";
    FD1S3DX phase_register_507__i14 (.D(n133[14]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(n233[14])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_507__i14.GSR = "DISABLED";
    FD1S3DX phase_register_507__i13 (.D(n133[13]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(n233[13])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_507__i13.GSR = "DISABLED";
    FD1S3DX phase_register_507__i12 (.D(n133[12]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(n233[12])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_507__i12.GSR = "DISABLED";
    FD1S3DX phase_register_507__i11 (.D(n133[11]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(n233[11])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_507__i11.GSR = "DISABLED";
    FD1S3DX phase_register_507__i10 (.D(n133[10]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(n233[10])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_507__i10.GSR = "DISABLED";
    FD1S3DX phase_register_507__i9 (.D(n133[9]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(n233[9])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_507__i9.GSR = "DISABLED";
    FD1S3DX phase_register_507__i8 (.D(n133[8]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(n233[8])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_507__i8.GSR = "DISABLED";
    FD1S3DX phase_register_507__i7 (.D(n133[7]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(n233[7])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_507__i7.GSR = "DISABLED";
    FD1S3DX phase_register_507__i6 (.D(n133[6]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(n233[6])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_507__i6.GSR = "DISABLED";
    FD1S3DX phase_register_507__i5 (.D(n133[5]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(n233[5])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_507__i5.GSR = "DISABLED";
    FD1S3DX phase_register_507__i4 (.D(n133[4]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(n233[4])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_507__i4.GSR = "DISABLED";
    FD1S3DX phase_register_507__i3 (.D(n133[3]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(n233[3])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_507__i3.GSR = "DISABLED";
    FD1S3DX phase_register_507__i2 (.D(n133[2]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(n233[2])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_507__i2.GSR = "DISABLED";
    FD1S3DX phase_register_507__i1 (.D(n133[1]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(n233[1])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_507__i1.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module dds_U2
//

module dds_U2 (i_ref_clk_c, i_resetb_N_301, carrier_increment, o_baseband_i_c_15, 
            o_baseband_i_c_14, o_baseband_i_c_13, o_baseband_i_c_12, o_baseband_i_c_11, 
            o_baseband_i_c_10, n3607, i_resetb_c, o_baseband_q_c_7, 
            o_baseband_i_c_7, o_baseband_i_c_8, \quarter_wave_sample_register_q[15] , 
            n27529, o_baseband_q_c_15, o_baseband_q_c_14, o_baseband_q_c_13, 
            o_baseband_q_c_12, o_baseband_q_c_11, o_baseband_q_c_10, n3608, 
            o_baseband_q_c_8, GND_net) /* synthesis syn_module_defined=1 */ ;
    input i_ref_clk_c;
    input i_resetb_N_301;
    input [30:0]carrier_increment;
    output o_baseband_i_c_15;
    output o_baseband_i_c_14;
    output o_baseband_i_c_13;
    output o_baseband_i_c_12;
    output o_baseband_i_c_11;
    output o_baseband_i_c_10;
    output n3607;
    input i_resetb_c;
    output o_baseband_q_c_7;
    output o_baseband_i_c_7;
    output o_baseband_i_c_8;
    output \quarter_wave_sample_register_q[15] ;
    input n27529;
    output o_baseband_q_c_15;
    output o_baseband_q_c_14;
    output o_baseband_q_c_13;
    output o_baseband_q_c_12;
    output o_baseband_q_c_11;
    output o_baseband_q_c_10;
    output n3608;
    output o_baseband_q_c_8;
    input GND_net;
    
    wire i_ref_clk_c /* synthesis SET_AS_NETWORK=i_ref_clk_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(22[12:21])
    wire o_baseband_i_c_15 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[37:47])
    wire o_baseband_i_c_14 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[37:47])
    wire o_baseband_i_c_13 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[37:47])
    wire o_baseband_i_c_12 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[37:47])
    wire o_baseband_i_c_11 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[37:47])
    wire o_baseband_i_c_10 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[37:47])
    wire n3607 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[37:47])
    wire o_baseband_q_c_7 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[49:59])
    wire o_baseband_i_c_7 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[37:47])
    wire o_baseband_i_c_8 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[37:47])
    wire o_baseband_q_c_15 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[49:59])
    wire o_baseband_q_c_14 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[49:59])
    wire o_baseband_q_c_13 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[49:59])
    wire o_baseband_q_c_12 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[49:59])
    wire o_baseband_q_c_11 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[49:59])
    wire o_baseband_q_c_10 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[49:59])
    wire n3608 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[49:59])
    wire o_baseband_q_c_8 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[49:59])
    wire [30:0]increment;   // d:/documents/git_local/fm_modulator/rtl/dds.v(14[31:40])
    wire [11:0]o_phase;   // d:/documents/git_local/fm_modulator/rtl/dds.v(18[26:33])
    
    FD1S3DX increment_i0 (.D(carrier_increment[0]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(increment[0])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=67, LSE_RLINE=67 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i0.GSR = "DISABLED";
    FD1S3DX increment_i30 (.D(carrier_increment[30]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(increment[30])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=67, LSE_RLINE=67 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i30.GSR = "DISABLED";
    FD1S3DX increment_i29 (.D(carrier_increment[29]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(increment[29])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=67, LSE_RLINE=67 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i29.GSR = "DISABLED";
    FD1S3DX increment_i28 (.D(carrier_increment[28]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(increment[28])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=67, LSE_RLINE=67 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i28.GSR = "DISABLED";
    FD1S3DX increment_i27 (.D(carrier_increment[27]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(increment[27])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=67, LSE_RLINE=67 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i27.GSR = "DISABLED";
    FD1S3DX increment_i26 (.D(carrier_increment[26]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(increment[26])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=67, LSE_RLINE=67 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i26.GSR = "DISABLED";
    FD1S3DX increment_i25 (.D(carrier_increment[25]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(increment[25])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=67, LSE_RLINE=67 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i25.GSR = "DISABLED";
    FD1S3DX increment_i24 (.D(carrier_increment[24]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(increment[24])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=67, LSE_RLINE=67 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i24.GSR = "DISABLED";
    FD1S3DX increment_i23 (.D(carrier_increment[23]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(increment[23])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=67, LSE_RLINE=67 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i23.GSR = "DISABLED";
    FD1S3DX increment_i22 (.D(carrier_increment[22]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(increment[22])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=67, LSE_RLINE=67 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i22.GSR = "DISABLED";
    FD1S3DX increment_i21 (.D(carrier_increment[21]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(increment[21])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=67, LSE_RLINE=67 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i21.GSR = "DISABLED";
    FD1S3DX increment_i20 (.D(carrier_increment[20]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(increment[20])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=67, LSE_RLINE=67 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i20.GSR = "DISABLED";
    FD1S3DX increment_i19 (.D(carrier_increment[19]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(increment[19])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=67, LSE_RLINE=67 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i19.GSR = "DISABLED";
    FD1S3DX increment_i18 (.D(carrier_increment[18]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(increment[18])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=67, LSE_RLINE=67 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i18.GSR = "DISABLED";
    FD1S3DX increment_i17 (.D(carrier_increment[17]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(increment[17])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=67, LSE_RLINE=67 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i17.GSR = "DISABLED";
    FD1S3DX increment_i16 (.D(carrier_increment[16]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(increment[16])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=67, LSE_RLINE=67 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i16.GSR = "DISABLED";
    FD1S3DX increment_i15 (.D(carrier_increment[15]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(increment[15])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=67, LSE_RLINE=67 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i15.GSR = "DISABLED";
    FD1S3DX increment_i14 (.D(carrier_increment[14]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(increment[14])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=67, LSE_RLINE=67 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i14.GSR = "DISABLED";
    FD1S3DX increment_i13 (.D(carrier_increment[13]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(increment[13])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=67, LSE_RLINE=67 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i13.GSR = "DISABLED";
    FD1S3DX increment_i12 (.D(carrier_increment[12]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(increment[12])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=67, LSE_RLINE=67 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i12.GSR = "DISABLED";
    FD1S3DX increment_i11 (.D(carrier_increment[11]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(increment[11])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=67, LSE_RLINE=67 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i11.GSR = "DISABLED";
    FD1S3DX increment_i10 (.D(carrier_increment[10]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(increment[10])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=67, LSE_RLINE=67 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i10.GSR = "DISABLED";
    FD1S3DX increment_i9 (.D(carrier_increment[9]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(increment[9])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=67, LSE_RLINE=67 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i9.GSR = "DISABLED";
    FD1S3DX increment_i8 (.D(carrier_increment[8]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(increment[8])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=67, LSE_RLINE=67 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i8.GSR = "DISABLED";
    FD1S3DX increment_i7 (.D(carrier_increment[7]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(increment[7])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=67, LSE_RLINE=67 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i7.GSR = "DISABLED";
    FD1S3DX increment_i6 (.D(carrier_increment[6]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(increment[6])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=67, LSE_RLINE=67 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i6.GSR = "DISABLED";
    FD1S3DX increment_i5 (.D(carrier_increment[5]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(increment[5])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=67, LSE_RLINE=67 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i5.GSR = "DISABLED";
    FD1S3DX increment_i4 (.D(carrier_increment[4]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(increment[4])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=67, LSE_RLINE=67 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i4.GSR = "DISABLED";
    FD1S3DX increment_i3 (.D(carrier_increment[3]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(increment[3])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=67, LSE_RLINE=67 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i3.GSR = "DISABLED";
    FD1S3DX increment_i2 (.D(carrier_increment[2]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(increment[2])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=67, LSE_RLINE=67 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i2.GSR = "DISABLED";
    FD1S3DX increment_i1 (.D(carrier_increment[1]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(increment[1])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=67, LSE_RLINE=67 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i1.GSR = "DISABLED";
    quarter_wave_sine_lookup_U0 qtr_inst (.i_ref_clk_c(i_ref_clk_c), .i_resetb_N_301(i_resetb_N_301), 
            .o_baseband_i_c_15(o_baseband_i_c_15), .o_baseband_i_c_14(o_baseband_i_c_14), 
            .o_baseband_i_c_13(o_baseband_i_c_13), .o_baseband_i_c_12(o_baseband_i_c_12), 
            .o_baseband_i_c_11(o_baseband_i_c_11), .o_baseband_i_c_10(o_baseband_i_c_10), 
            .n3607(n3607), .i_resetb_c(i_resetb_c), .o_phase({o_phase}), 
            .o_baseband_q_c_7(o_baseband_q_c_7), .o_baseband_i_c_7(o_baseband_i_c_7), 
            .o_baseband_i_c_8(o_baseband_i_c_8), .\quarter_wave_sample_register_q[15] (\quarter_wave_sample_register_q[15] ), 
            .n27529(n27529), .o_baseband_q_c_15(o_baseband_q_c_15), .o_baseband_q_c_14(o_baseband_q_c_14), 
            .o_baseband_q_c_13(o_baseband_q_c_13), .o_baseband_q_c_12(o_baseband_q_c_12), 
            .o_baseband_q_c_11(o_baseband_q_c_11), .o_baseband_q_c_10(o_baseband_q_c_10), 
            .n3608(n3608), .o_baseband_q_c_8(o_baseband_q_c_8), .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(21[70:134])
    \nco(OW=12)_U1  nco_inst (.increment({increment}), .o_phase({o_phase}), 
            .GND_net(GND_net), .i_ref_clk_c(i_ref_clk_c), .i_resetb_N_301(i_resetb_N_301)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(20[49:100])
    
endmodule
//
// Verilog Description of module quarter_wave_sine_lookup_U0
//

module quarter_wave_sine_lookup_U0 (i_ref_clk_c, i_resetb_N_301, o_baseband_i_c_15, 
            o_baseband_i_c_14, o_baseband_i_c_13, o_baseband_i_c_12, o_baseband_i_c_11, 
            o_baseband_i_c_10, n3607, i_resetb_c, o_phase, o_baseband_q_c_7, 
            o_baseband_i_c_7, o_baseband_i_c_8, \quarter_wave_sample_register_q[15] , 
            n27529, o_baseband_q_c_15, o_baseband_q_c_14, o_baseband_q_c_13, 
            o_baseband_q_c_12, o_baseband_q_c_11, o_baseband_q_c_10, n3608, 
            o_baseband_q_c_8, GND_net) /* synthesis syn_module_defined=1 */ ;
    input i_ref_clk_c;
    input i_resetb_N_301;
    output o_baseband_i_c_15;
    output o_baseband_i_c_14;
    output o_baseband_i_c_13;
    output o_baseband_i_c_12;
    output o_baseband_i_c_11;
    output o_baseband_i_c_10;
    output n3607;
    input i_resetb_c;
    input [11:0]o_phase;
    output o_baseband_q_c_7;
    output o_baseband_i_c_7;
    output o_baseband_i_c_8;
    output \quarter_wave_sample_register_q[15] ;
    input n27529;
    output o_baseband_q_c_15;
    output o_baseband_q_c_14;
    output o_baseband_q_c_13;
    output o_baseband_q_c_12;
    output o_baseband_q_c_11;
    output o_baseband_q_c_10;
    output n3608;
    output o_baseband_q_c_8;
    input GND_net;
    
    wire i_ref_clk_c /* synthesis SET_AS_NETWORK=i_ref_clk_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(22[12:21])
    wire [15:0]\o_val_pipeline_i[0]  /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(15[24:40])
    wire o_baseband_i_c_15 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[37:47])
    wire o_baseband_i_c_14 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[37:47])
    wire o_baseband_i_c_13 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[37:47])
    wire o_baseband_i_c_12 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[37:47])
    wire o_baseband_i_c_11 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[37:47])
    wire o_baseband_i_c_10 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[37:47])
    wire n3607 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[37:47])
    wire o_baseband_q_c_7 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[49:59])
    wire [15:0]\o_val_pipeline_q[0]  /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(16[24:40])
    wire o_baseband_i_c_7 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[37:47])
    wire o_baseband_i_c_8 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[37:47])
    wire o_baseband_q_c_15 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[49:59])
    wire o_baseband_q_c_14 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[49:59])
    wire o_baseband_q_c_13 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[49:59])
    wire o_baseband_q_c_12 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[49:59])
    wire o_baseband_q_c_11 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[49:59])
    wire o_baseband_q_c_10 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[49:59])
    wire n3608 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[49:59])
    wire o_baseband_q_c_8 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(110[49:59])
    wire [15:0]quarter_wave_sample_register_i;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(22[24:54])
    wire [14:0]quarter_wave_sample_register_i_15__N_2126;
    wire [9:0]index_i;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(31[17:24])
    
    wire n25116, n978, n12126, n25204, n25178;
    wire [9:0]index_q;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(31[26:33])
    
    wire n21201, n24812, n24824, n22855, n875, n890, n21687, o_val_pipeline_i_0__15__N_2156, 
        n25051, n859, o_val_pipeline_i_0__15__N_2158, o_val_pipeline_i_0__15__N_2160, 
        o_val_pipeline_i_0__15__N_2162, n21330, n21323, n20846, o_val_pipeline_i_0__15__N_2164, 
        o_val_pipeline_i_0__15__N_2166, n908, n923, n21688, o_val_pipeline_i_0__15__N_2168, 
        n21267, n21268, n21275, n939, n954, n21689, o_val_pipeline_i_0__15__N_2170, 
        n21298, n21291, n20241, n971, n986, n21690, n1002, n1017, 
        n21691, o_val_pipeline_i_0__15__N_2172, n25050, n21536, n20462, 
        n20463, n20473, n20464, n20465, n20474, n20470, n20471, 
        n20477, n25173, n325, n21200, n21202, n27519, n684, n25085, 
        n21481, n20499, n20500, n20507, n20501, n20502, n20508, 
        n124, n23394, n25176, n25183, n21198, n25122, n20505, 
        n20506, n20510, n348, n349, n20532, n20533, n20539, n20534, 
        n20535, n20540, n21383;
    wire [11:0]phase_q;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(12[17:24])
    
    wire n20536, n20537, n20541;
    wire [1:0]phase_negation_i;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(23[12:28])
    wire [11:0]phase_i;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(11[17:24])
    wire [1:0]phase_negation_q;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(23[30:46])
    wire [9:0]index_i_9__N_2106;
    wire [9:0]index_q_9__N_2116;
    wire [15:0]quarter_wave_sample_register_q;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(22[56:86])
    wire [14:0]quarter_wave_sample_register_q_15__N_2141;
    
    wire n20555, n20556, n20566, n12118, n24909, n20557, n20558, 
        n20567, n20563, n20564, n20570, n21197, n21199, n25096, 
        n24873, n382, n509, n20583, n21343, n382_adj_2251, n509_adj_2252, 
        n20586;
    wire [15:0]o_val_pipeline_i_0__15__N_2157;
    
    wire n21194, n21195, n21196, n25237, n25238, n25239, n21464, 
        n14329, n827, n954_adj_2253;
    wire [14:0]n1807;
    
    wire n21377, n24895, n541, n22817, n24786, n22818, n23437, 
        n23434, n23438, n526, n541_adj_2254, n21756, n20600, n20601, 
        n20602, n25053, n318, n20634, n20635, n20636, n20637, 
        n20638, n20639, n875_adj_2255, n20643, n20644, n20645, n557, 
        n572, n21757, n589, n604, n21758, n17303;
    wire [15:0]o_val_pipeline_q_0__15__N_2189;
    
    wire n17304, n17302, n27520, n25166, n38, n21395;
    wire [11:0]phase_q_11__N_2232;
    
    wire n24945, n24946, n22851, n25052, n17301, n190, n253, n20930, 
        n17300, n20933, n20934, n20939, n25034, n348_adj_2256, n349_adj_2257, 
        n382_adj_2258, n509_adj_2259, n20245, n20267, n20268, n20275, 
        n20269, n20270, n20276, n27503, n668, n17299, n620, n635, 
        n21759, n21145, n21146, n21152, n21191, n21192, n21193, 
        n21147, n21148, n21153, n21167, n21168, n21175, n21171, 
        n21172, n21177, n21173, n21174, n21178, n653, n668_adj_2260, 
        n21760, n20344, n20345, n20352, n20346, n20347, n20353, 
        n526_adj_2261, n541_adj_2262, n21676, n20350, n20351, n20355, 
        n21269, n21270, n21276, n21271, n21272, n21277, n21289, 
        n21290, n21296, n21297, n21299, n21300, n21307, n21303, 
        n21304, n21309, n21305, n21306, n21310, n699, n21761, 
        n20375, n20376, n20383, n20377, n20378, n20384, n716, 
        n731, n21762, n21321, n21322, n21328, n21329, n20408, 
        n20409, n20415, n20410, n20411, n20416, n20412, n20413, 
        n20417, n747, n762, n21763, n20437, n20438, n20445, n781, 
        n796, n21764, n25165, n364, n812, n12132, n21765, n20456, 
        n20457, n30, n875_adj_2263, n890_adj_2264, n21767, n20458, 
        n20459, n24811, n24825, n20466, n20467, n20475, n20483, 
        n20484, n20485, n20486, n20487, n20488, n20489, n20490, 
        n908_adj_2265, n923_adj_2266, n21768, n20491, n20492, n20503, 
        n20495, n20496, n20497, n20498, n939_adj_2267, n21769, n635_adj_2268, 
        n14330, n636, n971_adj_2269, n986_adj_2270, n21770, n20516, 
        n20517, n20531, n20518, n20519, n1002_adj_2271, n1017_adj_2272, 
        n21771, n20520, n20521, n20522, n20523, n20524, n20525, 
        n25159, n732, n763, n25054, n21555, n891, n20545, n20546, 
        n20561, n20549, n20550, n20551, n20552, n20559, n20560, 
        n20568, n620_adj_2273, n25113, n14311, n526_adj_2274, n25160, 
        n620_adj_2275, n635_adj_2276, n636_adj_2277, n25198, n25174, 
        n684_adj_2278, n24887, n24807, n875_adj_2279, n890_adj_2280, 
        n891_adj_2281, n23399, n23395, n23400, n844, n860, n25076, 
        n325_adj_2282, n21185, n379, n21692, n21693, n21700, n21694, 
        n21695, n21701, n21696, n21697, n21702, n27506, n526_adj_2283, 
        n22934, n21698, n21699, n21703, n701, n764, n23388, n23386, 
        n23389, n701_adj_2284, n764_adj_2285, n796_adj_2286, n812_adj_2287, 
        n21446, n924, n23387, n476, n23433, n93, n94, n20948, 
        n812_adj_2288, n62, n21439, n20443, n20444, n20448, n21224, 
        n491, n24044, n475, n25219, n908_adj_2289, n20528, n157, 
        n20441, n20442, n20447, n21545, n21772, n21773, n21780, 
        n21774, n21775, n21781, n21776, n21777, n21782, n21778, 
        n21779, n21783, n25230, n25231, n25232, n20686, n20687, 
        n20688, n20693, n20694, n20695, n204, n747_adj_2290, n762_adj_2291, 
        n763_adj_2292, n20716, n20717, n20723, n20724, n24970, n25040, 
        n20827, n20828, n20831, n20829, n20830, n20832, n620_adj_2293, 
        n635_adj_2294, n636_adj_2295, n20849, n20850, n20853, n20851, 
        n20852, n20854, n412, n23631, n20527, n20856, n20857, 
        n20860, n23385, n24863, n14802, n20858, n20859, n20861, 
        n25163, n506, n20863, n20864, n20867, n21490, n20865, 
        n20866, n20868, n17325, n17324, n20875, n20878, n20932, 
        n20881, n20884, n812_adj_2296, n20450, n20887, n20897, n17323, 
        n20381, n20386, n21434, n251, n12135, n11927, n348_adj_2297, 
        n17322, n251_adj_2298, n21496, n21529, n443, n379_adj_2299, 
        n24938, n24877, n21318, n443_adj_2300, n17788, n24942, n21286, 
        n24985, n20944, n25064, n605, n20913, n20914, n20917, 
        n21524, n27524, n985, n20915, n20916, n20918, n21008, 
        n21009, n21016, n21014, n21015, n21019, n428, n316, n23807, 
        n20251, n20252, n23809, n23919, n23985, n21143, n20253, 
        n20254, n428_adj_2301, n781_adj_2302, n27523, n25189, n747_adj_2303, 
        n20903, n20906, n21428, n20255, n20256, n11930, n20257, 
        n20258, n20259, n20260, n20271, n20263, n20264, n20273, 
        n23225, n20278, n141, n21491, n890_adj_2304, n891_adj_2305, 
        n21070, n21071, n21078, n21076, n21077, n21081, n20439, 
        n20446, n20973, n20976, n20285, n20272, n20277, n747_adj_2306, 
        n20979, n20982, n20286, n781_adj_2307, n762_adj_2308, n844_adj_2309, 
        n859_adj_2310, n860_adj_2311, n23981, n20280, n20985, n20988, 
        n20287, n21374, n21225, n20855, n20862, n20929, n21080, 
        n21083, n21079, n21082, n21135, n21136, n21457, n15, n24838, 
        n251_adj_2312, n157_adj_2313, n21413, n890_adj_2314, n699_adj_2315, 
        n21137, n21138, n24840, n109, n460, n364_adj_2316, n21139, 
        n21140, n21149, n251_adj_2317, n25185, n25201, n716_adj_2318, 
        n254, n25296, n25297, n62_adj_2319, n17321, n20947, n20951, 
        n588, n25181, n25293, n25294, n25295, n25090, n24864, 
        n25156, n653_adj_2320, n924_adj_2321, n956, n85, n23626, 
        n21367, n21433, n25194, n25206, n620_adj_2322, n379_adj_2323, 
        n27521, n589_adj_2324, n21141, n21142, n21150, n252, n21295, 
        n443_adj_2325, n252_adj_2326, n109_adj_2327, n12043, n20909, 
        n20922, n20925, n21170, n574, n20928, n20949, n20950, 
        n20952, n20946, n764_adj_2328, n460_adj_2329, n21553, n699_adj_2330, 
        n21018, n21021, n24884, n252_adj_2331, n716_adj_2332, n21017, 
        n21020, n397, n20297, n20298, n20313, n25184, n21674, 
        n332, n21673, n412_adj_2333, n20954, n20955, n20958, n20299, 
        n20300, n20314, n20301, n20302, n20315, n20305, n20306, 
        n20317, n20307, n20308, n20318, n20309, n20310, n20319, 
        n20311, n20312, n20320, n25047, n25087, n23629, n25290, 
        n25291, n25292, n412_adj_2334, n20956, n20957, n20959, n604_adj_2335, 
        n684_adj_2336, n12168, n12010, n19828, n762_adj_2337, n20328, 
        n20329, n127, n20330, n20331, n20332, n20333, n20334, 
        n20335, n20961, n20962, n20965, n23782, n25459, n25454, 
        n25460, n316_adj_2338, n17320, n20369, n20370, n20380, n20336, 
        n20337, n20348, n23785, n21422, n20340, n20341, n125, 
        n21293, n21259, n21260, n12039, n445, n24959, n445_adj_2339, 
        n684_adj_2340, n716_adj_2341, n21661, n20342, n20343, n21261, 
        n21262, n1001, n21263, n21264, n21273, n254_adj_2342, n21265, 
        n21266, n21274, n25079, n23633, n24948, n924_adj_2343, n956_adj_2344, 
        n23635, n252_adj_2345, n21327, n24876, n24949, n127_adj_2346, 
        n125_adj_2347, n21325, n25082, n23645, n24740, n23186, n20249, 
        n25244, n25284, n25285, n62_adj_2348, n25058, n25068, n23654, 
        n20963, n20964, n20966, n762_adj_2349, n24857, n27494, n12172, 
        n24956, n62_adj_2350, n27496, n860_adj_2351, n14996, n252_adj_2352, 
        n21285, n21287, n21288, n24817, n955, n364_adj_2353, n20685, 
        n21292, n24904, n189, n21294, n24957, n93_adj_2354, n23039, 
        n317, n20817, n20820, n12003, n20823, n20683, n20836, 
        n20839, n21302, n574_adj_2355, n20842, n21639, n20845, n764_adj_2356, 
        n25104, n765, n20844, n25195, n141_adj_2357, n21638, n413, 
        n24832, n24858, n638, n17319, n20359, n20360, n25205, 
        n173, n20361, n20362, n24980, n20363, n20364, n20365, 
        n20366, n20367, n20368, n20379, n20371, n20372, n24738, 
        n24787, n24739, n381, n24737, n24736, n12089, n731_adj_2358, 
        n732_adj_2359, n157_adj_2360, n828, n412_adj_2361, n20689, 
        n574_adj_2362, n637, n574_adj_2363, n637_adj_2364, n381_adj_2365, 
        n653_adj_2366, n21317, n318_adj_2367, n25457, n25456, n25458, 
        n21499, n25208, n17529, n21370, n17528, n21319, n21320, 
        n142, n20996, n638_adj_2368, n766, n173_adj_2369, n188, 
        n20997, n22932, n22933, n254_adj_2370, n20585, n254_adj_2371, 
        n20582, n27495, n21445, n21324, n333, n348_adj_2372, n21002, 
        n21326, n27497, n364_adj_2373, n21003, n27411, n27412, n22937, 
        n24715, n24714, n24716, n21785, n21784, n20385, n397_adj_2374, 
        n21004, n27396, n27397, n23060, n25077, n21559, n21560, 
        n21561, n21005, n20392, n20393, n20407, n21556, n20394, 
        n20395, n21557, n21558, n20396, n20397, n23279, n23276, 
        n23280, n20398, n20399, n20400, n20401, n27522, n21237, 
        n12175, n25451, n25452, n25083, n25065, n21548, n475_adj_2375, 
        n24965, n23184, n20421, n20422, n27498, n124_adj_2376, n20423, 
        n20424, n24969, n24815, n955_adj_2377, n860_adj_2378, n20425, 
        n20426, n27525, n301, n20429, n20430, n475_adj_2379, n21006, 
        n24010, n21705, n21704, n364_adj_2380, n20715, n14998, n252_adj_2381, 
        n27499, n20431, n20432, n20433, n20434, n27526, n20435, 
        n20436, n62_adj_2382, n653_adj_2383, n20587, n766_adj_2384, 
        n14928, n24922, n189_adj_2385, n21541, n491_adj_2386, n11355, 
        n21007, n317_adj_2387, n93_adj_2388, n23064, n890_adj_2389, 
        n22891, n25128, n13921, n20713, n221, n732_adj_2390, n763_adj_2391, 
        n23789, n20945, n21459, n891_adj_2392, n20452, n20453, n20468, 
        n125_adj_2393, n25005, n24955, n20810, n25084, n21533, n23988, 
        n158, n20242, n893, n25114, n24881, n221_adj_2394, n766_adj_2395, 
        n286, n21468, n21155, n21156, n21154, n747_adj_2396, n763_adj_2397, 
        n1002_adj_2398, n22874, n142_adj_2399, n157_adj_2400, n21058, 
        n19504, n20577, n173_adj_2401, n188_adj_2402, n21059, n333_adj_2403, 
        n348_adj_2404, n21064, n21471, n413_adj_2405, n444, n476_adj_2406, 
        n507, n21526, n21474, n573, n413_adj_2407, n157_adj_2408, 
        n828_adj_2409, n21065, n12114, n21477, n24947, n20843, n24802, 
        n25215, n397_adj_2410, n21066, n142_adj_2411, n25214, n669, 
        n700, n20493, n21523, n21525, n20584, n766_adj_2412, n20719, 
        n443_adj_2413, n21067, n21480, n20494, n25202, n23838, n797, 
        n475_adj_2414, n21068, n301_adj_2415, n317_adj_2416, n860_adj_2417, 
        n891_adj_2418, n20847, n924_adj_2419, n21483, n893_adj_2420, 
        n21279, n21280, n21278, n491_adj_2421, n11358, n21069, n21486, 
        n1018, n25164, n23859, n158_adj_2422, n189_adj_2423, n21085, 
        n21086, n21087, n221_adj_2424, n21492, n20449, n286_adj_2425, 
        n317_adj_2426, n349_adj_2427, n21495, n413_adj_2428, n21498, 
        n21501, n507_adj_2429, n21504, n573_adj_2430, n605_adj_2431, 
        n21507, n669_adj_2432, n700_adj_2433, n732_adj_2434, n763_adj_2435, 
        n723, n21514, n21097, n21098, n21099, n20419, n20414, 
        n20418, n21100, n21101, n21102, n12147, n12148, n25010, 
        n21103, n21104, n21105, n12145, n12146, n25032, n21106, 
        n21107, n21108, n94_adj_2436, n21513, n21516, n21519, n20547, 
        n25282, n21512, n20387, n21312, n21308, n21311, n21522, 
        n349_adj_2437, n21528, n21531, n20354, n20357, n21534, n21537, 
        n21112, n21113, n21114, n21543, n20554, n21546, n700_adj_2438, 
        n20356, n236, n21549, n21552, n844_adj_2439, n860_adj_2440, 
        n46, n20902, n21180, n21176, n21179, n498, n21505, n20279, 
        n21506, n25243, n20244, n20248, n23916, n924_adj_2441, n158_adj_2442, 
        n189_adj_2443, n25246, n987, n21500, n21497, n20809, n526_adj_2444, 
        n542, n25171, n21494, n635_adj_2445, n20927, n25025, n700_adj_2446, 
        n25097, n542_adj_2447, n635_adj_2448, n20841, n21164, n21165, 
        n21166, n17535, n17536, n17537, n21493, n508, n21476, 
        n25172, n23835, n17770, n668_adj_2449, n731_adj_2450, n732_adj_2451, 
        n25247, n747_adj_2452, n763_adj_2453, n22856, n20576, n20543, 
        n20538, n20542, n20509, n20512, n20511, n21482, n20940, 
        n20942, n20937, n20938, n20941, n25218, n21677, n844_adj_2454, 
        n860_adj_2455, n46_adj_2456, n20816, n316_adj_2457, n924_adj_2458, 
        n21678, n21679, n21680, n21681, n21682, n21683, n21425, 
        n24941, n124_adj_2459, n21684, n21685, n21686, n21448, n21449, 
        n21450, n508_adj_2460, n20571, n20572, n20574, n27528, n21443, 
        n21444, n20569, n20573, n20478, n20479, n20481, n20476, 
        n20480, n506_adj_2461, n349_adj_2462, n21517, n101, n21424, 
        n21426, n24814, n93_adj_2463, n94_adj_2464, n23625, n142_adj_2465, 
        n23961, n23962, n14105, n25041, n26497, n22895, n20289, 
        n26496, n20284, n26499, n20953, n20960, n26500, n23224, 
        n23222, n26501, n21518, n924_adj_2466, n23223, n24804, n30_adj_2467, 
        n23987, n21414, n1002_adj_2468, n716_adj_2469, n23989, n23986, 
        n23990, n21206, n21207, n476_adj_2470, n506_adj_2471, n23917, 
        n860_adj_2472, n541_adj_2473, n23993, n21403, n21404, n21405, 
        n25088, n23996, n25016, n25074, n24012, n21400, n21401, 
        n21402, n25168, n25169, n25080, n21521, n25217, n684_adj_2474, 
        n700_adj_2475, n635_adj_2476, n781_adj_2477, n669_adj_2478, 
        n716_adj_2479, n24015, n21766, n21248, n25081, n24016, n27518, 
        n24019, n30_adj_2480, n542_adj_2481, n557_adj_2482, n21515, 
        n25255, n285, n21472, n21473, n21550, n23058, n270, n15_adj_2483, 
        n286_adj_2484, n21226, n26637, n23061, n23062, n26638, n882, 
        n890_adj_2485, n19851, n157_adj_2486, n26701, n26700, n26702, 
        n26703, n26704, n26705, n20682, n26706, n26707, n20684, 
        n24043, n61, n94_adj_2487, n684_adj_2488, n812_adj_2489, n491_adj_2490, 
        n26764, n21239, n21240, n21241, n25011, n25199, n491_adj_2491, 
        n26765, n26774, n26775, n24045, n24042, n24046, n781_adj_2492, 
        n26776, n26777, n26778, n25188, n26779, n26780, n26781, 
        n475_adj_2493, n20690, n716_adj_2494, n731_adj_2495, n732_adj_2496, 
        n653_adj_2497, n669_adj_2498, n20880, n20691, n20692, n526_adj_2499, 
        n25207, n24053, n142_adj_2500, n604_adj_2501, n605_adj_2502, 
        n25193, n747_adj_2503, n24452, n24449, n24451, n24450, n882_adj_2504, 
        n475_adj_2505, n25252, n21375, n21371, n21372, n21092, n25091, 
        n828_adj_2506, n397_adj_2507, n954_adj_2508, n413_adj_2509, 
        n444_adj_2510, n12169, n221_adj_2511, n24246, n507_adj_2512, 
        n25221, n108, n25223, n25224, n25225, n25055, n653_adj_2513, 
        n316_adj_2514, n317_adj_2515, n270_adj_2516, n286_adj_2517, 
        n24056, n684_adj_2518, n746, n526_adj_2519, n25177, n142_adj_2520, 
        n14066, n158_adj_2521, n25180, n491_adj_2522, n20882, n25212, 
        n61_adj_2523, n62_adj_2524, n15_adj_2525, n24839, n31, n30_adj_2526, 
        n21212, n460_adj_2527, n24448, n20324, n21110, n781_adj_2528, 
        n30_adj_2529, n31_adj_2530, n15_adj_2531, n15_adj_2532, n30_adj_2533, 
        n31_adj_2534, n205, n157_adj_2535, n124_adj_2536, n900, n25123, 
        n62_adj_2537, n24898, n31_adj_2538, n24073, n348_adj_2539, 
        n12109, n12110, n12171, n23960, n21475, n20712, n31_adj_2540, 
        n404, n25200, n24072, n491_adj_2541, n21245, n25066, n12127, 
        n21657, n859_adj_2542, n24076, n20714, n443_adj_2543, n20720, 
        n20721, n20722, n24875, n23051, n24798, n23092, n875_adj_2544, 
        n891_adj_2545, n859_adj_2546, n860_adj_2547, n24921, n125_adj_2548, 
        n24785, n25045, n285_adj_2549, n25071, n781_adj_2550, n251_adj_2551, 
        n797_adj_2552, n24162, n24816, n21352, n21353, n21354, n21350, 
        n460_adj_2553, n157_adj_2554, n636_adj_2555, n25251, n25057, 
        n21340, n21341, n21342, n21440, n24406, n24403, n511, 
        n21344, n21345, n17538, n17539, n17540, n460_adj_2556, n101_adj_2557, 
        n507_adj_2558, n21346, n21347, n21348, n21458, n460_adj_2559, 
        n476_adj_2560, n24405, n24404, n397_adj_2561, n251_adj_2562, 
        n413_adj_2563, n27395, n21361, n236_adj_2564, n21349, n21351, 
        n24883, n24733, n14882, n22813, n17548, n17549, n17550, 
        n109_adj_2565, n125_adj_2566, n653_adj_2567, n94_adj_2568, n27394, 
        n21355, n21356, n21357, n506_adj_2569, n24402, n20891, n25220, 
        n27409, n27410, n6, n6_adj_2570, n301_adj_2571, n891_adj_2572, 
        n24159, n21247, n13956, n828_adj_2573, n21431, n797_adj_2574, 
        n23610, n908_adj_2575, n924_adj_2576, n173_adj_2577, n189_adj_2578, 
        n653_adj_2579, n668_adj_2580, n669_adj_2581, n541_adj_2582, 
        n890_adj_2583, n891_adj_2584, n25190, n25211, n557_adj_2585, 
        n573_adj_2586, n731_adj_2587, n796_adj_2588, n797_adj_2589, 
        n21421, n542_adj_2590, n285_adj_2591, n573_adj_2592, n669_adj_2593, 
        n25196, n15_adj_2594, n24862, n892, n158_adj_2595, n189_adj_2596, 
        n21419, n27507, n24054, n21454, n124_adj_2597, n23038, n23221, 
        n699_adj_2598, n21234, n573_adj_2599, n21233, n23784, n85_adj_2600, 
        n24160, n716_adj_2601, n20815, n21235, n526_adj_2602, n557_adj_2603, 
        n20818, n20819, n25197, n21394, n572_adj_2604, n573_adj_2605, 
        n511_adj_2606, n20821, n20822, n460_adj_2607, n285_adj_2608, 
        n476_adj_2609, n668_adj_2610, n109_adj_2611, n21436, n124_adj_2612, 
        n844_adj_2613, n397_adj_2614, n25023, n413_adj_2615, n14980, 
        n732_adj_2616, n21091, n25254, n17545, n21236, n491_adj_2617, 
        n23275, n17546, n859_adj_2618, n860_adj_2619, n443_adj_2620, 
        n93_adj_2621, n14811, n286_adj_2622, n25253, n24163, n21640, 
        n25161, n14096, n158_adj_2623, n20833, n572_adj_2624, n125_adj_2625, 
        n20834, n20835, n24170, n24920, n21412, n21658, n20837, 
        n20838, n506_adj_2626, n860_adj_2627, n251_adj_2628, n21215, 
        n21216, n21217, n21213, n21214, n20840, n21418, n21420, 
        n23185, n684_adj_2629, n700_adj_2630, n21423, n25203, n890_adj_2631, 
        n19847, n668_adj_2632, n669_adj_2633, n573_adj_2634, n25070, 
        n684_adj_2635, n25038, n412_adj_2636, n542_adj_2637, n24906, 
        n24172, n25022, n25069, n908_adj_2638, n285_adj_2639, n762_adj_2640, 
        n21427, n20869, n20870, n20871, n20872, n14992, n732_adj_2641, 
        n20873, n20874, n20876, n20877, n124_adj_2642, n23063, n20879, 
        n25072, n25037, n270_adj_2643, n316_adj_2644, n21430, n21432, 
        n21364, n20883, n21435, n812_adj_2645, n20885, n20886, n21094, 
        n21437, n21438, n397_adj_2646, n21441, n21416, n21461, n20895, 
        n20896, n21451, n557_adj_2647, n20901, n270_adj_2648, n286_adj_2649, 
        n20904, n20905, n24897, n20907, n20908, n25256, n491_adj_2650, 
        n25095, n444_adj_2651, n25020, n94_adj_2652, n25258, n21447, 
        n25257, n20919, n251_adj_2653, n78, n890_adj_2654, n891_adj_2655, 
        n14766, n20920, n20921, n14053, n828_adj_2656, n20923, n20924, 
        n21452, n21453, n12093, n797_adj_2657, n21455, n21456, n21368, 
        n668_adj_2658, n669_adj_2659, n20926, n30_adj_2660, n17531, 
        n17673, n20936, n541_adj_2661, n542_adj_2662, n20967, n20968, 
        n20969, n20970, n24861, n892_adj_2663, n20971, n20972, n20974, 
        n20975, n20977, n20978, n270_adj_2664, n285_adj_2665, n21062, 
        n20980, n20981, n236_adj_2666, n21061, n21054, n21362, n20983, 
        n20984, n20986, n20987, n31_adj_2667, n21096, n21479, n94_adj_2668, 
        n125_adj_2669, n20992, n20993, n875_adj_2670, n379_adj_2671, 
        n891_adj_2672, n15_adj_2673, n859_adj_2674, n860_adj_2675, n20994, 
        n20995, n781_adj_2676, n797_adj_2677, n25026, n24243, n21109, 
        n21111, n17547, n636_adj_2678, n17532, n17533, n507_adj_2679, 
        n476_adj_2680, n20999, n413_adj_2681, n397_adj_2682, n24247, 
        n24245, n24248, n986_adj_2683, n21010, n20998, n21011, n21470, 
        n21469, n21467, n21013, n573_adj_2684, n21466, n93_adj_2685, 
        n605_adj_2686, n12047, n24244, n653_adj_2687, n23066, n526_adj_2688, 
        n397_adj_2689, n475_adj_2690, n348_adj_2691, n700_adj_2692, 
        n20261, n21463, n21465, n333_adj_2693, n20262, n21460, n12007, 
        n21462, n23055, n21478, n23041, n491_adj_2694, n475_adj_2695, 
        n205_adj_2696, n93_adj_2697, n397_adj_2698, n348_adj_2699, n364_adj_2700, 
        n333_adj_2701, n24871, n21429, n23788, n908_adj_2702, n317_adj_2703, 
        n21055, n21056, n21057, n21554, n844_adj_2704, n21072, n21060, 
        n21073, n21417, n475_adj_2705, n890_adj_2706, n23994, n173_adj_2707, 
        n21407, n21406, n21408, n21075, n17670, n25073, n747_adj_2708, 
        n444_adj_2709, n828_adj_2710, n205_adj_2711, n21132, n21389, 
        n25259, n573_adj_2712, n21388, n21390, n636_adj_2713, n24870, 
        n700_adj_2714, n732_adj_2715, n21386, n21385, n21387, n142_adj_2716, 
        n221_adj_2717, n252_adj_2718, n21382, n21384, n24872, n21376, 
        n21378, n21369, n21365, n25031, n349_adj_2719, n24173, n24171, 
        n24174, n21366, n716_adj_2720, n19835, n21363, n12046, n24828, 
        n24856, n23057, n700_adj_2721, n23043, n24169, n12071, n828_adj_2722, 
        n21220, n94_adj_2723, n684_adj_2724, n24164, n24161, n24165, 
        n25033, n491_adj_2725, n220, n17305, n221_adj_2726, n14799, 
        n684_adj_2727, n25059, n605_adj_2728, n21229, n220_adj_2729, 
        n25226, n21232, n46_adj_2730, n93_adj_2731, n21249, n21250, 
        n21243, n108_adj_2732, n684_adj_2733, n716_adj_2734, n19824, 
        n21242, n21244, n444_adj_2735, n21238, n12006, n348_adj_2736, 
        n21231, n21230, n21228, n21227, n93_adj_2737, n173_adj_2738, 
        n21659, n21662, n21252, n21219, n25455, n21218, n21675, 
        n17530, n21256, n12015, n21257, n700_adj_2739, n20338, n24859, 
        n668_adj_2740, n46_adj_2741, n23980, n25222, n20339, n23913, 
        n763_adj_2742, n12174, n491_adj_2743, n605_adj_2744, n21551, 
        n19498, n700_adj_2745, n731_adj_2746, n732_adj_2747, n21093, 
        n1018_adj_2748, n14064, n142_adj_2749, n908_adj_2750, n19673, 
        n21527, n21544, n348_adj_2751, n21520, n573_adj_2752, n93_adj_2753, 
        n731_adj_2754, n21095, n653_adj_2755, n475_adj_2756, n604_adj_2757, 
        n25280, n21503, n954_adj_2758, n828_adj_2759, n21484, n25278, 
        n796_adj_2760, n348_adj_2761, n20469, n397_adj_2762, n25035, 
        n20454, n20472, n20460, n20461, n24077, n24074, n24078, 
        n20562, n23650, n23611, n20565, n23656, n23094, n23093, 
        n23095, n986_adj_2763, n20931, n25453, n22878, n62_adj_2764, 
        n20504, n22938, n23068, n21169, n23811, n700_adj_2765, n19655, 
        n20349, n25216, n444_adj_2766, n21301, n23787, n62_adj_2767, 
        n23790, n20404, n62_adj_2768, n24057, n24055, n24058, n20388, 
        n892_adj_2769, n221_adj_2770, n23862, n349_adj_2771, n24853, 
        n24854, n572_adj_2772, n124_adj_2773, n286_adj_2774, n24732, 
        n23054, n23067, n23065, n620_adj_2775, n14014, n507_adj_2776, 
        n23963, n491_adj_2777, n286_adj_2778, n23059, n763_adj_2779, 
        n924_adj_2780, n20403, n25042, n221_adj_2781, n252_adj_2782, 
        n23646, n924_adj_2783, n21530, n173_adj_2784, n21535, n23056, 
        n349_adj_2785, n24847, n23860, n24020, n24017, n24021, n24013, 
        n24011, n24014, n25063, n12177, n23997, n23995, n23998, 
        n572_adj_2786, n21532, n23984, n23982, n23983, n21158, n572_adj_2787, 
        n26502, n26498, n25017, n23651, n23042, n23040, n573_adj_2788, 
        n21547, n987_adj_2789, n985_adj_2790, n205_adj_2791, n157_adj_2792, 
        n23857, n348_adj_2793, n23648, n746_adj_2794, n19638, n25086, 
        n22893, n23918, n23915, n23653, n491_adj_2795, n20990, n25245, 
        n22876, n23914, n20899, n21084, n21706, n12008, n21022, 
        n21786, n21151, n19858, n23396, n23861, n23858, n12048, 
        n23840, n23837, n23841, n23836, n23810, n23808, n21542, 
        n23786, n23783, n23632, n14321, n23637, n635_adj_2796, n21660, 
        n21144, n23655, n23652, n23649, n23647, n23636, n23634, 
        n23627, n22894, n22892, n22877, n22875;
    
    FD1S3BX quarter_wave_sample_register_i_i2 (.D(quarter_wave_sample_register_i_15__N_2126[2]), 
            .CK(i_ref_clk_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_i[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i2.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i1 (.D(quarter_wave_sample_register_i_15__N_2126[1]), 
            .CK(i_ref_clk_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_i[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i1.GSR = "DISABLED";
    LUT4 i9560_3_lut_4_lut (.A(index_i[0]), .B(n25116), .C(index_i[4]), 
         .D(n978), .Z(n12126)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9560_3_lut_4_lut.init = 16'h4f40;
    LUT4 i18871_3_lut (.A(n25204), .B(n25178), .C(index_q[3]), .Z(n21201)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18871_3_lut.init = 16'hcaca;
    PFUMX i21348 (.BLUT(n24812), .ALUT(n24824), .C0(index_i[7]), .Z(n22855));
    PFUMX i19357 (.BLUT(n875), .ALUT(n890), .C0(index_q[4]), .Z(n21687));
    FD1S3DX o_val_pipeline_i_1__i18 (.D(o_val_pipeline_i_0__15__N_2156), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(\o_val_pipeline_i[0] [15])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i18.GSR = "DISABLED";
    LUT4 mux_192_Mux_2_i859_3_lut_4_lut (.A(index_i[0]), .B(n25116), .C(index_i[3]), 
         .D(n25051), .Z(n859)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_2_i859_3_lut_4_lut.init = 16'h4f40;
    FD1S3DX o_val_pipeline_i_1__i17 (.D(o_val_pipeline_i_0__15__N_2158), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(\o_val_pipeline_i[0] [14])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i17.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i16 (.D(o_val_pipeline_i_0__15__N_2160), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(\o_val_pipeline_i[0] [13])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i16.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i15 (.D(o_val_pipeline_i_0__15__N_2162), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(\o_val_pipeline_i[0] [12])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i15.GSR = "DISABLED";
    L6MUX21 i18516 (.D0(n21330), .D1(n21323), .SD(index_q[8]), .Z(n20846));
    FD1S3DX o_val_pipeline_i_1__i14 (.D(o_val_pipeline_i_0__15__N_2164), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(\o_val_pipeline_i[0] [11])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i14.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i13 (.D(o_val_pipeline_i_0__15__N_2166), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(\o_val_pipeline_i[0] [10])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i13.GSR = "DISABLED";
    PFUMX i19358 (.BLUT(n908), .ALUT(n923), .C0(index_q[4]), .Z(n21688));
    FD1S3DX o_val_pipeline_i_1__i12 (.D(o_val_pipeline_i_0__15__N_2168), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(\o_val_pipeline_i[0] [9])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i12.GSR = "DISABLED";
    PFUMX i18945 (.BLUT(n21267), .ALUT(n21268), .C0(index_q[7]), .Z(n21275));
    PFUMX i19359 (.BLUT(n939), .ALUT(n954), .C0(index_q[4]), .Z(n21689));
    FD1S3BX quarter_wave_sample_register_i_i14 (.D(quarter_wave_sample_register_i_15__N_2126[14]), 
            .CK(i_ref_clk_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_i[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i14.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i11 (.D(o_val_pipeline_i_0__15__N_2170), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(\o_val_pipeline_i[0] [8])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i11.GSR = "DISABLED";
    L6MUX21 i17911 (.D0(n21298), .D1(n21291), .SD(index_i[8]), .Z(n20241));
    PFUMX i19360 (.BLUT(n971), .ALUT(n986), .C0(index_q[4]), .Z(n21690));
    PFUMX i19361 (.BLUT(n1002), .ALUT(n1017), .C0(index_q[4]), .Z(n21691));
    FD1S3DX o_val_pipeline_i_1__i10 (.D(o_val_pipeline_i_0__15__N_2172), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(\o_val_pipeline_i[0] [7])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i10.GSR = "DISABLED";
    LUT4 i11346_2_lut_rep_490 (.A(index_i[0]), .B(index_i[1]), .Z(n25050)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11346_2_lut_rep_490.init = 16'h4444;
    LUT4 i19206_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n21536)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)+!C !(D)))+!A (B (C+!(D))+!B ((D)+!C)))) */ ;
    defparam i19206_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h0e30;
    L6MUX21 i18143 (.D0(n20462), .D1(n20463), .SD(index_q[6]), .Z(n20473));
    L6MUX21 i18144 (.D0(n20464), .D1(n20465), .SD(index_q[6]), .Z(n20474));
    L6MUX21 i18147 (.D0(n20470), .D1(n20471), .SD(index_q[7]), .Z(n20477));
    LUT4 i18870_3_lut (.A(n25173), .B(n325), .C(index_q[3]), .Z(n21200)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18870_3_lut.init = 16'hcaca;
    LUT4 i20120_3_lut (.A(n21200), .B(n21201), .C(index_q[4]), .Z(n21202)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20120_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_0_i684_3_lut_4_lut (.A(index_i[0]), .B(n25116), .C(index_i[3]), 
         .D(n27519), .Z(n684)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_0_i684_3_lut_4_lut.init = 16'h4f40;
    FD1S3DX o_val_pipeline_i_1__i9 (.D(\o_val_pipeline_i[0] [15]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(o_baseband_i_c_15)) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i9.GSR = "DISABLED";
    LUT4 i19151_3_lut_4_lut (.A(index_i[0]), .B(n25116), .C(index_i[3]), 
         .D(n25085), .Z(n21481)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19151_3_lut_4_lut.init = 16'hf404;
    FD1S3DX o_val_pipeline_i_1__i8 (.D(\o_val_pipeline_i[0] [14]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(o_baseband_i_c_14)) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i8.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i7 (.D(\o_val_pipeline_i[0] [13]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(o_baseband_i_c_13)) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i7.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i13 (.D(quarter_wave_sample_register_i_15__N_2126[13]), 
            .CK(i_ref_clk_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_i[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i13.GSR = "DISABLED";
    L6MUX21 i18177 (.D0(n20499), .D1(n20500), .SD(index_i[7]), .Z(n20507));
    L6MUX21 i18178 (.D0(n20501), .D1(n20502), .SD(index_i[7]), .Z(n20508));
    FD1S3BX quarter_wave_sample_register_i_i12 (.D(quarter_wave_sample_register_i_15__N_2126[12]), 
            .CK(i_ref_clk_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_i[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i12.GSR = "DISABLED";
    LUT4 n476_bdd_3_lut_21840_3_lut (.A(index_q[1]), .B(index_q[4]), .C(n124), 
         .Z(n23394)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n476_bdd_3_lut_21840_3_lut.init = 16'hd1d1;
    FD1S3DX o_val_pipeline_i_1__i6 (.D(\o_val_pipeline_i[0] [12]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(o_baseband_i_c_12)) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i6.GSR = "DISABLED";
    LUT4 i18868_3_lut (.A(n25176), .B(n25183), .C(index_q[3]), .Z(n21198)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18868_3_lut.init = 16'hcaca;
    LUT4 i8458_2_lut_rep_562 (.A(index_i[1]), .B(index_i[2]), .Z(n25122)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i8458_2_lut_rep_562.init = 16'h8888;
    L6MUX21 i18180 (.D0(n20505), .D1(n20506), .SD(index_i[7]), .Z(n20510));
    FD1S3DX o_val_pipeline_i_1__i5 (.D(\o_val_pipeline_i[0] [11]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(o_baseband_i_c_11)) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i5.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i11 (.D(quarter_wave_sample_register_i_15__N_2126[11]), 
            .CK(i_ref_clk_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_i[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i11.GSR = "DISABLED";
    LUT4 mux_192_Mux_3_i349_3_lut_3_lut (.A(index_i[1]), .B(index_i[4]), 
         .C(n348), .Z(n349)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_3_i349_3_lut_3_lut.init = 16'hd1d1;
    L6MUX21 i18209 (.D0(n20532), .D1(n20533), .SD(index_i[7]), .Z(n20539));
    L6MUX21 i18210 (.D0(n20534), .D1(n20535), .SD(index_i[7]), .Z(n20540));
    FD1S3DX o_val_pipeline_i_1__i4 (.D(\o_val_pipeline_i[0] [10]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(o_baseband_i_c_10)) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i4.GSR = "DISABLED";
    LUT4 i19053_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n21383)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C (D)+!C !(D)))+!A !(B (D)+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19053_3_lut_4_lut_4_lut_4_lut.init = 16'h7c03;
    FD1S3DX o_val_pipeline_i_1__i3 (.D(\o_val_pipeline_i[0] [9]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(n3607)) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i3.GSR = "DISABLED";
    FD1P3AX phase_q__i1 (.D(o_phase[0]), .SP(i_resetb_c), .CK(i_ref_clk_c), 
            .Q(phase_q[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_q__i1.GSR = "DISABLED";
    PFUMX i18211 (.BLUT(n20536), .ALUT(n20537), .C0(index_i[7]), .Z(n20541));
    FD1S3DX o_val_pipeline_q_1__i1 (.D(\o_val_pipeline_q[0] [7]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(o_baseband_q_c_7)) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_q_1__i1.GSR = "DISABLED";
    FD1S3DX phase_negation_i_i0 (.D(phase_i[11]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(phase_negation_i[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_negation_i_i0.GSR = "DISABLED";
    FD1S3DX phase_negation_q_i0 (.D(phase_q[11]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(phase_negation_q[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_negation_q_i0.GSR = "DISABLED";
    FD1S3DX index_i_i0 (.D(index_i_9__N_2106[0]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(index_i[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_i_i0.GSR = "DISABLED";
    FD1S3DX index_q_i0 (.D(index_q_9__N_2116[0]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(index_q[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_q_i0.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i0 (.D(quarter_wave_sample_register_q_15__N_2141[0]), 
            .CK(i_ref_clk_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_q[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_q_i0.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i1 (.D(\o_val_pipeline_i[0] [7]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(o_baseband_i_c_7)) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i1.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i0 (.D(quarter_wave_sample_register_i_15__N_2126[0]), 
            .CK(i_ref_clk_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_i[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i0.GSR = "DISABLED";
    L6MUX21 i18236 (.D0(n20555), .D1(n20556), .SD(index_i[6]), .Z(n20566));
    FD1S3DX o_val_pipeline_i_1__i2 (.D(\o_val_pipeline_i[0] [8]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(o_baseband_i_c_8)) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i2.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i11 (.D(o_phase[11]), .SP(i_resetb_c), .CK(i_ref_clk_c), 
            .Q(phase_i[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i11.GSR = "DISABLED";
    LUT4 i9552_2_lut_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[3]), 
         .Z(n12118)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9552_2_lut_3_lut.init = 16'h8080;
    FD1S3BX quarter_wave_sample_register_i_i10 (.D(quarter_wave_sample_register_i_15__N_2126[10]), 
            .CK(i_ref_clk_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_i[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i10.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i10 (.D(o_phase[10]), .SP(i_resetb_c), .CK(i_ref_clk_c), 
            .Q(phase_i[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i10.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i9 (.D(o_phase[9]), .SP(i_resetb_c), .CK(i_ref_clk_c), 
            .Q(phase_i[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i9.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i8 (.D(o_phase[8]), .SP(i_resetb_c), .CK(i_ref_clk_c), 
            .Q(phase_i[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i8.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i7 (.D(o_phase[7]), .SP(i_resetb_c), .CK(i_ref_clk_c), 
            .Q(phase_i[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i7.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i9 (.D(quarter_wave_sample_register_i_15__N_2126[9]), 
            .CK(i_ref_clk_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_i[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i9.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i6 (.D(o_phase[6]), .SP(i_resetb_c), .CK(i_ref_clk_c), 
            .Q(phase_i[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i6.GSR = "DISABLED";
    LUT4 i11288_2_lut_rep_349_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[3]), 
         .Z(n24909)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11288_2_lut_rep_349_3_lut.init = 16'hf8f8;
    FD1P3AX phase_i_i0_i5 (.D(o_phase[5]), .SP(i_resetb_c), .CK(i_ref_clk_c), 
            .Q(phase_i[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i5.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i8 (.D(quarter_wave_sample_register_i_15__N_2126[8]), 
            .CK(i_ref_clk_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_i[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i8.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i4 (.D(o_phase[4]), .SP(i_resetb_c), .CK(i_ref_clk_c), 
            .Q(phase_i[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i4.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i3 (.D(o_phase[3]), .SP(i_resetb_c), .CK(i_ref_clk_c), 
            .Q(phase_i[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i3.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i2 (.D(o_phase[2]), .SP(i_resetb_c), .CK(i_ref_clk_c), 
            .Q(phase_i[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i2.GSR = "DISABLED";
    L6MUX21 i18237 (.D0(n20557), .D1(n20558), .SD(index_i[6]), .Z(n20567));
    L6MUX21 i18240 (.D0(n20563), .D1(n20564), .SD(index_i[7]), .Z(n20570));
    FD1P3AX phase_i_i0_i1 (.D(o_phase[1]), .SP(i_resetb_c), .CK(i_ref_clk_c), 
            .Q(phase_i[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i1.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i7 (.D(quarter_wave_sample_register_i_15__N_2126[7]), 
            .CK(i_ref_clk_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_i[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i7.GSR = "DISABLED";
    LUT4 i20124_3_lut (.A(n21197), .B(n21198), .C(index_q[4]), .Z(n21199)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20124_3_lut.init = 16'hcaca;
    FD1S3BX quarter_wave_sample_register_i_i6 (.D(quarter_wave_sample_register_i_15__N_2126[6]), 
            .CK(i_ref_clk_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_i[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i6.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i5 (.D(quarter_wave_sample_register_i_15__N_2126[5]), 
            .CK(i_ref_clk_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_i[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i5.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i4 (.D(quarter_wave_sample_register_i_15__N_2126[4]), 
            .CK(i_ref_clk_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_i[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i4.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i3 (.D(quarter_wave_sample_register_i_15__N_2126[3]), 
            .CK(i_ref_clk_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_i[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i3.GSR = "DISABLED";
    LUT4 i11207_2_lut_rep_313_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[4]), .D(n25096), .Z(n24873)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11207_2_lut_rep_313_3_lut_4_lut.init = 16'hf8f0;
    PFUMX i18253 (.BLUT(n382), .ALUT(n509), .C0(index_q[7]), .Z(n20583));
    LUT4 i19013_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21343)) /* synthesis lut_function=(A (B (C (D))+!B !(C (D)))+!A !(B (D)+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19013_3_lut_4_lut_4_lut.init = 16'h9366;
    PFUMX i18256 (.BLUT(n382_adj_2251), .ALUT(n509_adj_2252), .C0(index_i[7]), 
          .Z(n20586));
    LUT4 quarter_wave_sample_register_i_12__I_0_3_lut (.A(quarter_wave_sample_register_i[12]), 
         .B(o_val_pipeline_i_0__15__N_2157[12]), .C(phase_negation_i[1]), 
         .Z(o_val_pipeline_i_0__15__N_2162)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[14] 77[8])
    defparam quarter_wave_sample_register_i_12__I_0_3_lut.init = 16'hcaca;
    LUT4 i20129_3_lut (.A(n21194), .B(n21195), .C(index_q[4]), .Z(n21196)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20129_3_lut.init = 16'hcaca;
    FD1S3BX quarter_wave_sample_register_q_i15 (.D(n27529), .CK(i_ref_clk_c), 
            .PD(i_resetb_N_301), .Q(\quarter_wave_sample_register_q[15] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_q_i15.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i14 (.D(quarter_wave_sample_register_q_15__N_2141[14]), 
            .CK(i_ref_clk_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_q[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_q_i14.GSR = "DISABLED";
    PFUMX i23020 (.BLUT(n25237), .ALUT(n25238), .C0(index_q[0]), .Z(n25239));
    FD1S3BX quarter_wave_sample_register_q_i13 (.D(quarter_wave_sample_register_q_15__N_2141[13]), 
            .CK(i_ref_clk_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_q[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_q_i13.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i12 (.D(quarter_wave_sample_register_q_15__N_2141[12]), 
            .CK(i_ref_clk_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_q[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_q_i12.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i11 (.D(quarter_wave_sample_register_q_15__N_2141[11]), 
            .CK(i_ref_clk_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_q[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_q_i11.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i10 (.D(quarter_wave_sample_register_q_15__N_2141[10]), 
            .CK(i_ref_clk_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_q[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_q_i10.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i9 (.D(quarter_wave_sample_register_q_15__N_2141[9]), 
            .CK(i_ref_clk_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_q[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_q_i9.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i8 (.D(quarter_wave_sample_register_q_15__N_2141[8]), 
            .CK(i_ref_clk_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_q[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_q_i8.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i7 (.D(quarter_wave_sample_register_q_15__N_2141[7]), 
            .CK(i_ref_clk_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_q[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_q_i7.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i6 (.D(quarter_wave_sample_register_q_15__N_2141[6]), 
            .CK(i_ref_clk_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_q[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_q_i6.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i5 (.D(quarter_wave_sample_register_q_15__N_2141[5]), 
            .CK(i_ref_clk_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_q[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_q_i5.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i4 (.D(quarter_wave_sample_register_q_15__N_2141[4]), 
            .CK(i_ref_clk_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_q[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_q_i4.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i3 (.D(quarter_wave_sample_register_q_15__N_2141[3]), 
            .CK(i_ref_clk_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_q[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_q_i3.GSR = "DISABLED";
    LUT4 i19134_3_lut_4_lut_3_lut (.A(index_q[1]), .B(index_q[3]), .C(index_q[2]), 
         .Z(n21464)) /* synthesis lut_function=(A (B)+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19134_3_lut_4_lut_3_lut.init = 16'hd9d9;
    FD1S3BX quarter_wave_sample_register_q_i2 (.D(quarter_wave_sample_register_q_15__N_2141[2]), 
            .CK(i_ref_clk_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_q[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_q_i2.GSR = "DISABLED";
    LUT4 i11654_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[4]), 
         .C(n25096), .D(index_q[0]), .Z(n14329)) /* synthesis lut_function=(!(A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11654_3_lut_4_lut_4_lut_4_lut.init = 16'h55d5;
    FD1S3BX quarter_wave_sample_register_q_i1 (.D(quarter_wave_sample_register_q_15__N_2141[1]), 
            .CK(i_ref_clk_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_q[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_q_i1.GSR = "DISABLED";
    FD1S3DX index_q_i9 (.D(index_q_9__N_2116[9]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(index_q[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_q_i9.GSR = "DISABLED";
    FD1S3DX index_q_i8 (.D(index_q_9__N_2116[8]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(index_q[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_q_i8.GSR = "DISABLED";
    FD1S3DX index_q_i7 (.D(index_q_9__N_2116[7]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(index_q[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_q_i7.GSR = "DISABLED";
    LUT4 mux_192_Mux_4_i827_3_lut_3_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[3]), .Z(n827)) /* synthesis lut_function=(A (B+(C))+!A !(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_4_i827_3_lut_3_lut.init = 16'ha9a9;
    FD1S3DX index_q_i6 (.D(index_q_9__N_2116[6]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(index_q[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_q_i6.GSR = "DISABLED";
    FD1S3DX index_q_i5 (.D(index_q_9__N_2116[5]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(index_q[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_q_i5.GSR = "DISABLED";
    LUT4 mux_192_Mux_0_i954_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n954_adj_2253)) /* synthesis lut_function=(A (D)+!A !(B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_0_i954_3_lut_4_lut_4_lut.init = 16'haf40;
    FD1S3DX index_q_i4 (.D(index_q_9__N_2116[4]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(index_q[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_q_i4.GSR = "DISABLED";
    FD1S3DX index_q_i3 (.D(index_q_9__N_2116[3]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(index_q[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_q_i3.GSR = "DISABLED";
    FD1S3DX index_q_i2 (.D(index_q_9__N_2116[2]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(index_q[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_q_i2.GSR = "DISABLED";
    FD1S3DX index_q_i1 (.D(index_q_9__N_2116[1]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(index_q[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_q_i1.GSR = "DISABLED";
    FD1S3DX index_i_i9 (.D(index_i_9__N_2106[9]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(index_i[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_i_i9.GSR = "DISABLED";
    FD1S3DX index_i_i8 (.D(index_i_9__N_2106[8]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(index_i[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_i_i8.GSR = "DISABLED";
    FD1S3DX index_i_i7 (.D(index_i_9__N_2106[7]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(index_i[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_i_i7.GSR = "DISABLED";
    FD1S3DX index_i_i6 (.D(index_i_9__N_2106[6]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(index_i[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_i_i6.GSR = "DISABLED";
    FD1S3DX index_i_i5 (.D(index_i_9__N_2106[5]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(index_i[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_i_i5.GSR = "DISABLED";
    FD1S3DX index_i_i4 (.D(index_i_9__N_2106[4]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(index_i[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_i_i4.GSR = "DISABLED";
    FD1S3DX index_i_i3 (.D(index_i_9__N_2106[3]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(index_i[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_i_i3.GSR = "DISABLED";
    FD1S3DX index_i_i2 (.D(index_i_9__N_2106[2]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(index_i[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_i_i2.GSR = "DISABLED";
    FD1S3DX index_i_i1 (.D(index_i_9__N_2106[1]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(index_i[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_i_i1.GSR = "DISABLED";
    FD1S3DX phase_negation_q_i1 (.D(phase_negation_q[0]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(phase_negation_q[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_negation_q_i1.GSR = "DISABLED";
    FD1S3DX phase_negation_i_i1 (.D(phase_negation_i[0]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(phase_negation_i[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_negation_i_i1.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i18 (.D(n1807[14]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(\o_val_pipeline_q[0] [15])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_q_1__i18.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i17 (.D(n1807[13]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(\o_val_pipeline_q[0] [14])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_q_1__i17.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i16 (.D(n1807[12]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(\o_val_pipeline_q[0] [13])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_q_1__i16.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i15 (.D(n1807[11]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(\o_val_pipeline_q[0] [12])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_q_1__i15.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i14 (.D(n1807[10]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(\o_val_pipeline_q[0] [11])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_q_1__i14.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i13 (.D(n1807[9]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(\o_val_pipeline_q[0] [10])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_q_1__i13.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i12 (.D(n1807[8]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(\o_val_pipeline_q[0] [9])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_q_1__i12.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i11 (.D(n1807[7]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(\o_val_pipeline_q[0] [8])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_q_1__i11.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i10 (.D(n1807[6]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(\o_val_pipeline_q[0] [7])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_q_1__i10.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i9 (.D(\o_val_pipeline_q[0] [15]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(o_baseband_q_c_15)) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_q_1__i9.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i8 (.D(\o_val_pipeline_q[0] [14]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(o_baseband_q_c_14)) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_q_1__i8.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i7 (.D(\o_val_pipeline_q[0] [13]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(o_baseband_q_c_13)) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_q_1__i7.GSR = "DISABLED";
    LUT4 i19047_3_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[3]), .C(index_q[2]), 
         .D(index_q[0]), .Z(n21377)) /* synthesis lut_function=(A (B (D)+!B (C (D)+!C !(D)))+!A (B (D)+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19047_3_lut_4_lut_4_lut.init = 16'hfc13;
    FD1S3DX o_val_pipeline_q_1__i6 (.D(\o_val_pipeline_q[0] [12]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(o_baseband_q_c_12)) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_q_1__i6.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i5 (.D(\o_val_pipeline_q[0] [11]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(o_baseband_q_c_11)) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_q_1__i5.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i4 (.D(\o_val_pipeline_q[0] [10]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(o_baseband_q_c_10)) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_q_1__i4.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i3 (.D(\o_val_pipeline_q[0] [9]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(n3608)) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_q_1__i3.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i2 (.D(\o_val_pipeline_q[0] [8]), .CK(i_ref_clk_c), 
            .CD(i_resetb_N_301), .Q(o_baseband_q_c_8)) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_q_1__i2.GSR = "DISABLED";
    LUT4 i11631_2_lut_rep_335_2_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .Z(n24895)) /* synthesis lut_function=(A (B+!(C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11631_2_lut_rep_335_2_lut_3_lut.init = 16'h8f8f;
    LUT4 mux_192_Mux_6_i269_3_lut_rep_491 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n25051)) /* synthesis lut_function=(A (C)+!A !((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_6_i269_3_lut_rep_491.init = 16'ha4a4;
    LUT4 mux_192_Mux_4_i541_3_lut_4_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n541)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B ((D)+!C)))) */ ;
    defparam mux_192_Mux_4_i541_3_lut_4_lut_3_lut_4_lut.init = 16'h0ef0;
    L6MUX21 i21322 (.D0(n22817), .D1(n24786), .SD(index_q[6]), .Z(n22818));
    PFUMX i21859 (.BLUT(n23437), .ALUT(n23434), .C0(index_i[6]), .Z(n23438));
    PFUMX i19426 (.BLUT(n526), .ALUT(n541_adj_2254), .C0(index_i[4]), 
          .Z(n21756));
    L6MUX21 i18272 (.D0(n20600), .D1(n20601), .SD(index_q[7]), .Z(n20602));
    LUT4 i11676_3_lut_4_lut (.A(index_i[0]), .B(n25122), .C(n25053), .D(index_i[5]), 
         .Z(n318)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (C (D))) */ ;
    defparam i11676_3_lut_4_lut.init = 16'hf800;
    L6MUX21 i18306 (.D0(n20634), .D1(n20635), .SD(index_q[7]), .Z(n20636));
    L6MUX21 i18309 (.D0(n20637), .D1(n20638), .SD(index_i[7]), .Z(n20639));
    LUT4 i9532_3_lut_4_lut_3_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[0]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n875_adj_2255)) /* synthesis lut_function=(A (B (C (D))+!B !(C (D)))+!A ((C (D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9532_3_lut_4_lut_3_lut_4_lut_4_lut.init = 16'hd333;
    L6MUX21 i18315 (.D0(n20643), .D1(n20644), .SD(index_i[7]), .Z(n20645));
    PFUMX i19427 (.BLUT(n557), .ALUT(n572), .C0(index_i[4]), .Z(n21757));
    PFUMX i19428 (.BLUT(n589), .ALUT(n604), .C0(index_i[4]), .Z(n21758));
    CCU2D add_358_11 (.A0(quarter_wave_sample_register_q[10]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_q[11]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17303), .COUT(n17304), 
          .S0(o_val_pipeline_q_0__15__N_2189[10]), .S1(o_val_pipeline_q_0__15__N_2189[11]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(80[29:60])
    defparam add_358_11.INIT0 = 16'hf555;
    defparam add_358_11.INIT1 = 16'hf555;
    defparam add_358_11.INJECT1_0 = "NO";
    defparam add_358_11.INJECT1_1 = "NO";
    CCU2D add_358_9 (.A0(quarter_wave_sample_register_q[8]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_q[9]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17302), .COUT(n17303), 
          .S0(o_val_pipeline_q_0__15__N_2189[8]), .S1(o_val_pipeline_q_0__15__N_2189[9]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(80[29:60])
    defparam add_358_9.INIT0 = 16'hf555;
    defparam add_358_9.INIT1 = 16'hf555;
    defparam add_358_9.INJECT1_0 = "NO";
    defparam add_358_9.INJECT1_1 = "NO";
    LUT4 mux_192_Mux_0_i589_3_lut (.A(n27520), .B(n978), .C(index_i[3]), 
         .Z(n589)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_0_i589_3_lut.init = 16'hcaca;
    LUT4 i19065_3_lut_3_lut (.A(n25166), .B(index_i[3]), .C(n38), .Z(n21395)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam i19065_3_lut_3_lut.init = 16'h7474;
    FD1P3AX phase_q__i11 (.D(phase_q_11__N_2232[11]), .SP(i_resetb_c), .CK(i_ref_clk_c), 
            .Q(phase_q[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_q__i11.GSR = "DISABLED";
    LUT4 index_i_4__bdd_4_lut_21635 (.A(index_i[4]), .B(n24945), .C(index_i[7]), 
         .D(n24946), .Z(n22851)) /* synthesis lut_function=(A (C+!(D))+!A (B+!(C))) */ ;
    defparam index_i_4__bdd_4_lut_21635.init = 16'he5ef;
    LUT4 mux_192_Mux_6_i22_3_lut_3_lut_rep_492 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n25052)) /* synthesis lut_function=(!(A (C)+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_6_i22_3_lut_3_lut_rep_492.init = 16'h4a4a;
    CCU2D add_358_7 (.A0(quarter_wave_sample_register_q[6]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_q[7]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17301), .COUT(n17302), 
          .S1(o_val_pipeline_q_0__15__N_2189[7]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(80[29:60])
    defparam add_358_7.INIT0 = 16'hf555;
    defparam add_358_7.INIT1 = 16'hf555;
    defparam add_358_7.INJECT1_0 = "NO";
    defparam add_358_7.INJECT1_1 = "NO";
    L6MUX21 i18600 (.D0(n190), .D1(n253), .SD(index_q[6]), .Z(n20930));
    CCU2D add_358_5 (.A0(quarter_wave_sample_register_q[4]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_q[5]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17300), .COUT(n17301));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(80[29:60])
    defparam add_358_5.INIT0 = 16'hf555;
    defparam add_358_5.INIT1 = 16'hf555;
    defparam add_358_5.INJECT1_0 = "NO";
    defparam add_358_5.INJECT1_1 = "NO";
    L6MUX21 i18609 (.D0(n20933), .D1(n20934), .SD(index_q[7]), .Z(n20939));
    LUT4 mux_192_Mux_4_i93_3_lut_4_lut_3_lut_rep_474_4_lut (.A(index_i[1]), 
         .B(index_i[2]), .C(index_i[3]), .D(index_i[0]), .Z(n25034)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_4_i93_3_lut_4_lut_3_lut_rep_474_4_lut.init = 16'h07f0;
    LUT4 mux_193_Mux_3_i349_3_lut_3_lut (.A(index_q[1]), .B(index_q[4]), 
         .C(n348_adj_2256), .Z(n349_adj_2257)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_3_i349_3_lut_3_lut.init = 16'hd1d1;
    L6MUX21 i17915 (.D0(n382_adj_2258), .D1(n509_adj_2259), .SD(index_i[7]), 
            .Z(n20245));
    L6MUX21 i17945 (.D0(n20267), .D1(n20268), .SD(index_q[7]), .Z(n20275));
    L6MUX21 i17946 (.D0(n20269), .D1(n20270), .SD(index_q[7]), .Z(n20276));
    LUT4 mux_192_Mux_4_i668_3_lut_3_lut (.A(n25166), .B(index_i[3]), .C(n27503), 
         .Z(n668)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;
    defparam mux_192_Mux_4_i668_3_lut_3_lut.init = 16'hd1d1;
    CCU2D add_358_3 (.A0(quarter_wave_sample_register_q[2]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_q[3]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17299), .COUT(n17300));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(80[29:60])
    defparam add_358_3.INIT0 = 16'hf555;
    defparam add_358_3.INIT1 = 16'hf555;
    defparam add_358_3.INJECT1_0 = "NO";
    defparam add_358_3.INJECT1_1 = "NO";
    PFUMX i19429 (.BLUT(n620), .ALUT(n635), .C0(index_i[4]), .Z(n21759));
    PFUMX i18822 (.BLUT(n21145), .ALUT(n21146), .C0(index_i[7]), .Z(n21152));
    LUT4 i20135_3_lut (.A(n21191), .B(n21192), .C(index_i[4]), .Z(n21193)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20135_3_lut.init = 16'hcaca;
    L6MUX21 i18823 (.D0(n21147), .D1(n21148), .SD(index_i[7]), .Z(n21153));
    L6MUX21 i18845 (.D0(n21167), .D1(n21168), .SD(index_i[7]), .Z(n21175));
    L6MUX21 i18847 (.D0(n21171), .D1(n21172), .SD(index_i[7]), .Z(n21177));
    PFUMX i18848 (.BLUT(n21173), .ALUT(n21174), .C0(index_i[7]), .Z(n21178));
    PFUMX i19430 (.BLUT(n653), .ALUT(n668_adj_2260), .C0(index_i[4]), 
          .Z(n21760));
    CCU2D add_358_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(quarter_wave_sample_register_q[0]), .B1(quarter_wave_sample_register_q[1]), 
          .C1(GND_net), .D1(GND_net), .COUT(n17299));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(80[29:60])
    defparam add_358_1.INIT0 = 16'hF000;
    defparam add_358_1.INIT1 = 16'ha666;
    defparam add_358_1.INJECT1_0 = "NO";
    defparam add_358_1.INJECT1_1 = "NO";
    L6MUX21 i18022 (.D0(n20344), .D1(n20345), .SD(index_q[7]), .Z(n20352));
    L6MUX21 i18023 (.D0(n20346), .D1(n20347), .SD(index_q[7]), .Z(n20353));
    PFUMX i19346 (.BLUT(n526_adj_2261), .ALUT(n541_adj_2262), .C0(index_q[4]), 
          .Z(n21676));
    L6MUX21 i18025 (.D0(n20350), .D1(n20351), .SD(index_q[7]), .Z(n20355));
    PFUMX i18946 (.BLUT(n21269), .ALUT(n21270), .C0(index_q[7]), .Z(n21276));
    L6MUX21 i18947 (.D0(n21271), .D1(n21272), .SD(index_q[7]), .Z(n21277));
    L6MUX21 i18961 (.D0(n21289), .D1(n21290), .SD(index_i[7]), .Z(n21291));
    L6MUX21 i18968 (.D0(n21296), .D1(n21297), .SD(index_i[7]), .Z(n21298));
    L6MUX21 i18977 (.D0(n21299), .D1(n21300), .SD(index_q[7]), .Z(n21307));
    L6MUX21 i18979 (.D0(n21303), .D1(n21304), .SD(index_q[7]), .Z(n21309));
    PFUMX i18980 (.BLUT(n21305), .ALUT(n21306), .C0(index_q[7]), .Z(n21310));
    PFUMX i19431 (.BLUT(n684), .ALUT(n699), .C0(index_i[4]), .Z(n21761));
    L6MUX21 i18053 (.D0(n20375), .D1(n20376), .SD(index_i[7]), .Z(n20383));
    L6MUX21 i18054 (.D0(n20377), .D1(n20378), .SD(index_i[7]), .Z(n20384));
    PFUMX i19432 (.BLUT(n716), .ALUT(n731), .C0(index_i[4]), .Z(n21762));
    L6MUX21 i18993 (.D0(n21321), .D1(n21322), .SD(index_q[7]), .Z(n21323));
    L6MUX21 i19000 (.D0(n21328), .D1(n21329), .SD(index_q[7]), .Z(n21330));
    L6MUX21 i18085 (.D0(n20408), .D1(n20409), .SD(index_q[7]), .Z(n20415));
    L6MUX21 i18086 (.D0(n20410), .D1(n20411), .SD(index_q[7]), .Z(n20416));
    PFUMX i18087 (.BLUT(n20412), .ALUT(n20413), .C0(index_q[7]), .Z(n20417));
    PFUMX i19433 (.BLUT(n747), .ALUT(n762), .C0(index_i[4]), .Z(n21763));
    L6MUX21 i18115 (.D0(n20437), .D1(n20438), .SD(index_i[7]), .Z(n20445));
    PFUMX i19434 (.BLUT(n781), .ALUT(n796), .C0(index_i[4]), .Z(n21764));
    LUT4 mux_192_Mux_7_i364_3_lut_3_lut (.A(n25166), .B(index_i[3]), .C(n25165), 
         .Z(n364)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;
    defparam mux_192_Mux_7_i364_3_lut_3_lut.init = 16'hd1d1;
    PFUMX i19435 (.BLUT(n812), .ALUT(n12132), .C0(index_i[4]), .Z(n21765));
    L6MUX21 i18140 (.D0(n20456), .D1(n20457), .SD(index_q[6]), .Z(n20470));
    LUT4 mux_192_Mux_9_i30_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .D(index_i[3]), .Z(n30)) /* synthesis lut_function=(A (B (C (D))+!B !(D))+!A !(B+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_9_i30_3_lut_4_lut_4_lut_4_lut.init = 16'h8033;
    PFUMX i19437 (.BLUT(n875_adj_2263), .ALUT(n890_adj_2264), .C0(index_i[4]), 
          .Z(n21767));
    L6MUX21 i18141 (.D0(n20458), .D1(n20459), .SD(index_q[6]), .Z(n20471));
    PFUMX i21320 (.BLUT(n24811), .ALUT(n24825), .C0(index_q[7]), .Z(n22817));
    L6MUX21 i18145 (.D0(n20466), .D1(n20467), .SD(index_q[6]), .Z(n20475));
    L6MUX21 i18169 (.D0(n20483), .D1(n20484), .SD(index_i[6]), .Z(n20499));
    L6MUX21 i18170 (.D0(n20485), .D1(n20486), .SD(index_i[6]), .Z(n20500));
    L6MUX21 i18171 (.D0(n20487), .D1(n20488), .SD(index_i[6]), .Z(n20501));
    L6MUX21 i18172 (.D0(n20489), .D1(n20490), .SD(index_i[6]), .Z(n20502));
    PFUMX i19438 (.BLUT(n908_adj_2265), .ALUT(n923_adj_2266), .C0(index_i[4]), 
          .Z(n21768));
    L6MUX21 i18173 (.D0(n20491), .D1(n20492), .SD(index_i[6]), .Z(n20503));
    L6MUX21 i18175 (.D0(n20495), .D1(n20496), .SD(index_i[6]), .Z(n20505));
    L6MUX21 i18176 (.D0(n20497), .D1(n20498), .SD(index_i[6]), .Z(n20506));
    PFUMX i19439 (.BLUT(n939_adj_2267), .ALUT(n954_adj_2253), .C0(index_i[4]), 
          .Z(n21769));
    LUT4 mux_193_Mux_6_i636_4_lut_4_lut (.A(index_q[1]), .B(index_q[4]), 
         .C(n635_adj_2268), .D(n14330), .Z(n636)) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_6_i636_4_lut_4_lut.init = 16'hf3d1;
    PFUMX i19440 (.BLUT(n971_adj_2269), .ALUT(n986_adj_2270), .C0(index_i[4]), 
          .Z(n21770));
    L6MUX21 i18201 (.D0(n20516), .D1(n20517), .SD(index_i[6]), .Z(n20531));
    L6MUX21 i18202 (.D0(n20518), .D1(n20519), .SD(index_i[6]), .Z(n20532));
    PFUMX i19441 (.BLUT(n1002_adj_2271), .ALUT(n1017_adj_2272), .C0(index_i[4]), 
          .Z(n21771));
    L6MUX21 i18203 (.D0(n20520), .D1(n20521), .SD(index_i[6]), .Z(n20533));
    L6MUX21 i18204 (.D0(n20522), .D1(n20523), .SD(index_i[6]), .Z(n20534));
    L6MUX21 i18205 (.D0(n20524), .D1(n20525), .SD(index_i[6]), .Z(n20535));
    LUT4 i11417_2_lut_rep_599 (.A(index_q[1]), .B(index_q[0]), .Z(n25159)) /* synthesis lut_function=((B)+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11417_2_lut_rep_599.init = 16'hdddd;
    PFUMX i18226 (.BLUT(n732), .ALUT(n763), .C0(index_i[5]), .Z(n20556));
    LUT4 i1_2_lut_rep_494 (.A(index_q[0]), .B(index_q[1]), .Z(n25054)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_2_lut_rep_494.init = 16'h8888;
    L6MUX21 i18228 (.D0(n21555), .D1(n891), .SD(index_i[5]), .Z(n20558));
    L6MUX21 i18231 (.D0(n20545), .D1(n20546), .SD(index_i[6]), .Z(n20561));
    L6MUX21 i18233 (.D0(n20549), .D1(n20550), .SD(index_i[6]), .Z(n20563));
    L6MUX21 i18234 (.D0(n20551), .D1(n20552), .SD(index_i[6]), .Z(n20564));
    L6MUX21 i18238 (.D0(n20559), .D1(n20560), .SD(index_i[6]), .Z(n20568));
    LUT4 mux_193_Mux_7_i620_3_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[0]), .D(index_q[3]), .Z(n620_adj_2273)) /* synthesis lut_function=(A (B (C+!(D)))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_7_i620_3_lut_4_lut_4_lut.init = 16'h9199;
    LUT4 i11636_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(n25113), .C(index_i[4]), 
         .D(index_i[0]), .Z(n14311)) /* synthesis lut_function=(!(A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11636_3_lut_4_lut_4_lut_4_lut.init = 16'h55d5;
    LUT4 mux_193_Mux_8_i526_3_lut_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n526_adj_2274)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_8_i526_3_lut_3_lut_3_lut_4_lut.init = 16'h0f70;
    LUT4 mux_193_Mux_7_i262_3_lut_rep_600 (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[0]), .Z(n25160)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_7_i262_3_lut_rep_600.init = 16'h6464;
    PFUMX mux_192_Mux_1_i636 (.BLUT(n620_adj_2275), .ALUT(n635_adj_2276), 
          .C0(index_i[4]), .Z(n636_adj_2277)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 mux_193_Mux_3_i684_3_lut (.A(n25198), .B(n25174), .C(index_q[3]), 
         .Z(n684_adj_2278)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_3_i684_3_lut.init = 16'hcaca;
    LUT4 i12371_2_lut_rep_247_3_lut_4_lut (.A(n24887), .B(index_i[4]), .C(index_i[6]), 
         .D(index_i[5]), .Z(n24807)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;
    defparam i12371_2_lut_rep_247_3_lut_4_lut.init = 16'hf080;
    PFUMX mux_192_Mux_2_i891 (.BLUT(n875_adj_2279), .ALUT(n890_adj_2280), 
          .C0(index_i[4]), .Z(n891_adj_2281)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    PFUMX i21823 (.BLUT(n23399), .ALUT(n23395), .C0(index_q[6]), .Z(n23400));
    PFUMX mux_192_Mux_2_i860 (.BLUT(n844), .ALUT(n859), .C0(index_i[4]), 
          .Z(n860)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 i18855_3_lut (.A(n25076), .B(n325_adj_2282), .C(index_i[3]), 
         .Z(n21185)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18855_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_7_i379_3_lut_3_lut (.A(n25166), .B(index_i[3]), .C(n27520), 
         .Z(n379)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam mux_192_Mux_7_i379_3_lut_3_lut.init = 16'h7474;
    L6MUX21 i19370 (.D0(n21692), .D1(n21693), .SD(index_q[6]), .Z(n21700));
    L6MUX21 i19371 (.D0(n21694), .D1(n21695), .SD(index_q[6]), .Z(n21701));
    L6MUX21 i19372 (.D0(n21696), .D1(n21697), .SD(index_q[6]), .Z(n21702));
    LUT4 mux_193_Mux_0_i795_3_lut_4_lut_3_lut_rep_666 (.A(index_q[0]), .B(index_q[2]), 
         .C(index_q[1]), .Z(n27506)) /* synthesis lut_function=(A (B+(C))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i795_3_lut_4_lut_3_lut_rep_666.init = 16'hb9b9;
    LUT4 n21488_bdd_3_lut_3_lut (.A(index_i[1]), .B(n526_adj_2283), .C(index_i[4]), 
         .Z(n22934)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n21488_bdd_3_lut_3_lut.init = 16'h5c5c;
    L6MUX21 i19373 (.D0(n21698), .D1(n21699), .SD(index_q[6]), .Z(n21703));
    PFUMX i18305 (.BLUT(n701), .ALUT(n764), .C0(index_q[6]), .Z(n20635));
    L6MUX21 i21815 (.D0(n23388), .D1(n23386), .SD(index_i[6]), .Z(n23389));
    PFUMX i18308 (.BLUT(n701_adj_2284), .ALUT(n764_adj_2285), .C0(index_i[6]), 
          .Z(n20638));
    LUT4 mux_193_Mux_0_i796_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[2]), 
         .C(index_q[1]), .D(index_q[3]), .Z(n796_adj_2286)) /* synthesis lut_function=(A (B (C+(D))+!B (C (D)))+!A !(B ((D)+!C)+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i796_3_lut_4_lut_4_lut.init = 16'hb9c0;
    LUT4 mux_192_Mux_4_i812_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n812_adj_2287)) /* synthesis lut_function=(!(A (C+(D))+!A !(B (C+(D))+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_4_i812_3_lut_3_lut_4_lut.init = 16'h554a;
    LUT4 i19116_3_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[2]), .C(index_q[0]), 
         .D(index_q[3]), .Z(n21446)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A (B (C)+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19116_3_lut_4_lut_4_lut.init = 16'h3c9d;
    PFUMX i21813 (.BLUT(n924), .ALUT(n23387), .C0(index_i[5]), .Z(n23388));
    LUT4 n476_bdd_3_lut_21934 (.A(n476), .B(n23433), .C(index_i[5]), .Z(n23434)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n476_bdd_3_lut_21934.init = 16'hcaca;
    LUT4 mux_192_Mux_3_i94_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[4]), .D(n93), .Z(n94)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_3_i94_3_lut_4_lut.init = 16'hf606;
    LUT4 i18618_3_lut_3_lut (.A(n25166), .B(index_i[3]), .C(n27503), .Z(n20948)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam i18618_3_lut_3_lut.init = 16'h7474;
    LUT4 mux_192_Mux_3_i62_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[4]), .D(n812_adj_2288), .Z(n62)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_3_i62_3_lut_4_lut.init = 16'h6f60;
    LUT4 i19109_3_lut_4_lut (.A(index_q[1]), .B(index_q[2]), .C(index_q[0]), 
         .D(index_q[3]), .Z(n21439)) /* synthesis lut_function=(!(A (B (D)+!B !(C+!(D)))+!A !(B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19109_3_lut_4_lut.init = 16'h64aa;
    LUT4 i18118_3_lut (.A(n20443), .B(n20444), .C(index_i[7]), .Z(n20448)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18118_3_lut.init = 16'hcaca;
    LUT4 i18894_3_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[2]), .C(index_q[0]), 
         .D(index_q[3]), .Z(n21224)) /* synthesis lut_function=(!(A (B+!(C+(D)))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18894_3_lut_4_lut_4_lut.init = 16'h6664;
    LUT4 mux_192_Mux_5_i491_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n491)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A !(B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_5_i491_3_lut_4_lut_4_lut.init = 16'ha54a;
    LUT4 n547_bdd_4_lut_22423_4_lut_4_lut (.A(index_q[1]), .B(index_q[0]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n24044)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B (C)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n547_bdd_4_lut_22423_4_lut_4_lut.init = 16'h3d2d;
    LUT4 mux_192_Mux_5_i475_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n475)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_5_i475_3_lut_4_lut_4_lut.init = 16'hd4a5;
    LUT4 i18198_4_lut_4_lut (.A(index_i[4]), .B(index_i[5]), .C(n25219), 
         .D(n908_adj_2289), .Z(n20528)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam i18198_4_lut_4_lut.init = 16'hd1c0;
    LUT4 mux_192_Mux_0_i157_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n157)) /* synthesis lut_function=(A (B (C+!(D))+!B !(D))+!A (B (D)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_0_i157_3_lut_4_lut.init = 16'hd4aa;
    LUT4 i18117_3_lut (.A(n20441), .B(n20442), .C(index_i[7]), .Z(n20447)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18117_3_lut.init = 16'hcaca;
    LUT4 i19215_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21545)) /* synthesis lut_function=(!(A ((D)+!C)+!A !(B ((D)+!C)+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19215_3_lut_3_lut_4_lut.init = 16'h55a4;
    L6MUX21 i19450 (.D0(n21772), .D1(n21773), .SD(index_i[6]), .Z(n21780));
    L6MUX21 i19451 (.D0(n21774), .D1(n21775), .SD(index_i[6]), .Z(n21781));
    L6MUX21 i19452 (.D0(n21776), .D1(n21777), .SD(index_i[6]), .Z(n21782));
    L6MUX21 i19453 (.D0(n21778), .D1(n21779), .SD(index_i[6]), .Z(n21783));
    PFUMX i23016 (.BLUT(n25230), .ALUT(n25231), .C0(index_q[2]), .Z(n25232));
    L6MUX21 i18358 (.D0(n20686), .D1(n20687), .SD(index_q[6]), .Z(n20688));
    L6MUX21 i18365 (.D0(n20693), .D1(n20694), .SD(index_q[6]), .Z(n20695));
    LUT4 mux_192_Mux_6_i204_3_lut_4_lut_3_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .Z(n204)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_6_i204_3_lut_4_lut_3_lut_3_lut.init = 16'h3d3d;
    PFUMX mux_192_Mux_3_i763 (.BLUT(n747_adj_2290), .ALUT(n762_adj_2291), 
          .C0(index_i[4]), .Z(n763_adj_2292)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    L6MUX21 i18388 (.D0(n20716), .D1(n20717), .SD(index_i[6]), .Z(n382_adj_2258));
    L6MUX21 i18395 (.D0(n20723), .D1(n20724), .SD(index_i[6]), .Z(n509_adj_2259));
    LUT4 i11539_2_lut_rep_410_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[0]), 
         .Z(n24970)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11539_2_lut_rep_410_3_lut.init = 16'h8080;
    LUT4 i11385_2_lut_rep_480 (.A(index_i[1]), .B(index_i[0]), .Z(n25040)) /* synthesis lut_function=((B)+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11385_2_lut_rep_480.init = 16'hdddd;
    PFUMX i18501 (.BLUT(n20827), .ALUT(n20828), .C0(index_q[4]), .Z(n20831));
    PFUMX i18502 (.BLUT(n20829), .ALUT(n20830), .C0(index_q[4]), .Z(n20832));
    PFUMX mux_193_Mux_1_i636 (.BLUT(n620_adj_2293), .ALUT(n635_adj_2294), 
          .C0(index_q[4]), .Z(n636_adj_2295)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    PFUMX i18523 (.BLUT(n20849), .ALUT(n20850), .C0(index_q[4]), .Z(n20853));
    PFUMX i18524 (.BLUT(n20851), .ALUT(n20852), .C0(index_q[4]), .Z(n20854));
    LUT4 mux_192_Mux_9_i412_3_lut_4_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .Z(n412)) /* synthesis lut_function=(!(A (B (C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_9_i412_3_lut_4_lut_3_lut.init = 16'h7e7e;
    LUT4 i18206_3_lut (.A(n23631), .B(n20527), .C(index_i[6]), .Z(n20536)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18206_3_lut.init = 16'hcaca;
    PFUMX i18530 (.BLUT(n20856), .ALUT(n20857), .C0(index_q[4]), .Z(n20860));
    PFUMX i21811 (.BLUT(n23385), .ALUT(n24863), .C0(index_i[5]), .Z(n23386));
    LUT4 mux_192_Mux_0_i781_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n781)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A (B (C)+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_0_i781_4_lut_4_lut_4_lut.init = 16'h0cb4;
    LUT4 mux_192_Mux_8_i412_3_lut_4_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .Z(n14802)) /* synthesis lut_function=(A (B+!(C))+!A !((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_8_i412_3_lut_4_lut_3_lut.init = 16'h8e8e;
    PFUMX i18531 (.BLUT(n20858), .ALUT(n20859), .C0(index_q[4]), .Z(n20861));
    LUT4 mux_192_Mux_7_i506_3_lut_4_lut (.A(n25163), .B(index_i[2]), .C(index_i[3]), 
         .D(n25165), .Z(n506)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_7_i506_3_lut_4_lut.init = 16'h2f20;
    PFUMX i18537 (.BLUT(n20863), .ALUT(n20864), .C0(index_q[4]), .Z(n20867));
    LUT4 i19160_3_lut_3_lut_4_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n21490)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B !((D)+!C)))) */ ;
    defparam i19160_3_lut_3_lut_4_lut_3_lut_4_lut.init = 16'h11ef;
    PFUMX i18538 (.BLUT(n20865), .ALUT(n20866), .C0(index_q[4]), .Z(n20868));
    CCU2D add_357_15 (.A0(quarter_wave_sample_register_i[14]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(\quarter_wave_sample_register_q[15] ), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17325), .S0(o_val_pipeline_i_0__15__N_2157[14]), 
          .S1(o_val_pipeline_i_0__15__N_2157[15]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam add_357_15.INIT0 = 16'hf555;
    defparam add_357_15.INIT1 = 16'hf555;
    defparam add_357_15.INJECT1_0 = "NO";
    defparam add_357_15.INJECT1_1 = "NO";
    CCU2D add_357_13 (.A0(quarter_wave_sample_register_i[12]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[13]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17324), .COUT(n17325), 
          .S0(o_val_pipeline_i_0__15__N_2157[12]), .S1(o_val_pipeline_i_0__15__N_2157[13]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam add_357_13.INIT0 = 16'hf555;
    defparam add_357_13.INIT1 = 16'hf555;
    defparam add_357_13.INJECT1_0 = "NO";
    defparam add_357_13.INJECT1_1 = "NO";
    L6MUX21 i18602 (.D0(n20875), .D1(n20878), .SD(index_q[6]), .Z(n20932));
    L6MUX21 i18603 (.D0(n20881), .D1(n20884), .SD(index_q[6]), .Z(n20933));
    LUT4 i8441_2_lut_rep_493 (.A(index_i[3]), .B(index_i[4]), .Z(n25053)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i8441_2_lut_rep_493.init = 16'heeee;
    LUT4 mux_193_Mux_6_i812_3_lut_4_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n812_adj_2296)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(D))+!A !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_6_i812_3_lut_4_lut_3_lut_4_lut.init = 16'h7780;
    LUT4 i20918_3_lut (.A(n20447), .B(n20448), .C(index_i[8]), .Z(n20450)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20918_3_lut.init = 16'hcaca;
    L6MUX21 i18604 (.D0(n20887), .D1(n20897), .SD(index_q[6]), .Z(n20934));
    CCU2D add_357_11 (.A0(quarter_wave_sample_register_i[10]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[11]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17323), .COUT(n17324), 
          .S0(o_val_pipeline_i_0__15__N_2157[10]), .S1(o_val_pipeline_i_0__15__N_2157[11]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam add_357_11.INIT0 = 16'hf555;
    defparam add_357_11.INIT1 = 16'hf555;
    defparam add_357_11.INJECT1_0 = "NO";
    defparam add_357_11.INJECT1_1 = "NO";
    LUT4 i18056_3_lut (.A(n20381), .B(n23389), .C(index_i[7]), .Z(n20386)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18056_3_lut.init = 16'hcaca;
    LUT4 i18497_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[3]), 
         .C(index_q[2]), .D(index_q[0]), .Z(n20827)) /* synthesis lut_function=(A (B (C (D))+!B (C))+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18497_3_lut_4_lut_4_lut_4_lut.init = 16'hb434;
    LUT4 i19104_3_lut_4_lut_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[0]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n21434)) /* synthesis lut_function=(!(A (B (C)+!B (C+(D)))+!A !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19104_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'h585f;
    LUT4 mux_193_Mux_0_i251_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[0]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n251)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A !(B ((D)+!C)+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i251_3_lut_4_lut_4_lut_4_lut.init = 16'h543c;
    LUT4 i9569_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n12135)) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B ((D)+!C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9569_3_lut_4_lut_4_lut.init = 16'hcdad;
    LUT4 i9361_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[0]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n11927)) /* synthesis lut_function=(A (B (D)+!B !((D)+!C))+!A (((D)+!C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9361_3_lut_4_lut_4_lut_4_lut.init = 16'hdd35;
    LUT4 mux_193_Mux_1_i348_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[3]), 
         .C(index_q[2]), .D(index_q[0]), .Z(n348_adj_2297)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_1_i348_3_lut_4_lut_4_lut_4_lut.init = 16'h7870;
    CCU2D add_357_9 (.A0(quarter_wave_sample_register_i[8]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[9]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17322), .COUT(n17323), 
          .S0(o_val_pipeline_i_0__15__N_2157[8]), .S1(o_val_pipeline_i_0__15__N_2157[9]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam add_357_9.INIT0 = 16'hf555;
    defparam add_357_9.INIT1 = 16'hf555;
    defparam add_357_9.INJECT1_0 = "NO";
    defparam add_357_9.INJECT1_1 = "NO";
    LUT4 mux_192_Mux_0_i251_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n251_adj_2298)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A !(B ((D)+!C)+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_0_i251_3_lut_4_lut_4_lut_4_lut.init = 16'h543c;
    LUT4 i19166_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n21496)) /* synthesis lut_function=(!(A (B (C (D)))+!A !(B+(C+(D))))) */ ;
    defparam i19166_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h7ffe;
    LUT4 i19199_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n21529)) /* synthesis lut_function=(A (B (C (D)))+!A !(B+(C+(D)))) */ ;
    defparam i19199_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h8001;
    LUT4 mux_192_Mux_8_i443_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n443)) /* synthesis lut_function=(A (B (C+!(D))+!B !((D)+!C))+!A !(B (D)+!B ((D)+!C))) */ ;
    defparam mux_192_Mux_8_i443_3_lut_4_lut_4_lut.init = 16'h80fc;
    LUT4 mux_192_Mux_0_i379_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n379_adj_2299)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !((D)+!C))+!A !(B ((D)+!C)+!B (D))) */ ;
    defparam mux_192_Mux_0_i379_3_lut_4_lut_4_lut.init = 16'h8079;
    LUT4 i9566_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n12132)) /* synthesis lut_function=(A (B (D)+!B !((D)+!C))+!A (((D)+!C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9566_3_lut_4_lut_4_lut_4_lut.init = 16'hdd35;
    LUT4 i18988_3_lut_4_lut_4_lut (.A(n24938), .B(index_q[4]), .C(index_q[5]), 
         .D(n24877), .Z(n21318)) /* synthesis lut_function=(A ((C+!(D))+!B)+!A (B (C+!(D))+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18988_3_lut_4_lut_4_lut.init = 16'he3ef;
    LUT4 mux_192_Mux_0_i443_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .D(index_i[3]), .Z(n443_adj_2300)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C (D))+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_0_i443_3_lut_4_lut_4_lut_4_lut.init = 16'h0ed5;
    LUT4 i3_3_lut_4_lut (.A(n24938), .B(index_q[4]), .C(index_q[6]), .D(index_q[5]), 
         .Z(n17788)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i3_3_lut_4_lut.init = 16'hfffe;
    LUT4 i18956_3_lut_4_lut_4_lut (.A(n24942), .B(index_i[4]), .C(index_i[5]), 
         .D(n24887), .Z(n21286)) /* synthesis lut_function=(A ((C+!(D))+!B)+!A (B (C+!(D))+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18956_3_lut_4_lut_4_lut.init = 16'he3ef;
    LUT4 i18614_3_lut_4_lut_4_lut (.A(n24970), .B(index_i[4]), .C(index_i[3]), 
         .D(n24985), .Z(n20944)) /* synthesis lut_function=(A (B (C)+!B !(C+!(D)))+!A (B (C)+!B (C+(D)))) */ ;
    defparam i18614_3_lut_4_lut_4_lut.init = 16'hd3d0;
    LUT4 i9495_3_lut_4_lut (.A(index_i[3]), .B(index_i[4]), .C(n25064), 
         .D(n27503), .Z(n605)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9495_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i18587 (.BLUT(n20913), .ALUT(n20914), .C0(index_i[4]), .Z(n20917));
    LUT4 i19194_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n21524)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(D))+!A (B (D)+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19194_3_lut_4_lut_4_lut_4_lut.init = 16'hd52b;
    LUT4 mux_193_Mux_0_i986_3_lut (.A(n27524), .B(n985), .C(index_q[3]), 
         .Z(n986)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i986_3_lut.init = 16'hcaca;
    PFUMX i18588 (.BLUT(n20915), .ALUT(n20916), .C0(index_i[4]), .Z(n20918));
    L6MUX21 i18686 (.D0(n21008), .D1(n21009), .SD(index_i[6]), .Z(n21016));
    L6MUX21 i18689 (.D0(n21014), .D1(n21015), .SD(index_i[6]), .Z(n21019));
    LUT4 mux_192_Mux_0_i428_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[2]), 
         .B(index_i[0]), .C(index_i[1]), .D(index_i[3]), .Z(n428)) /* synthesis lut_function=(A (B (C+!(D))+!B !((D)+!C))+!A (B (D)+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_0_i428_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hd5a9;
    LUT4 mux_192_Mux_9_i316_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), 
         .B(index_i[2]), .C(index_i[3]), .D(index_i[0]), .Z(n316)) /* synthesis lut_function=(!(A (B (C)+!B !(C+(D)))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_9_i316_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h7e7c;
    LUT4 n78_bdd_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n23807)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A !((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n78_bdd_3_lut_4_lut_4_lut_4_lut.init = 16'h7173;
    L6MUX21 i17937 (.D0(n20251), .D1(n20252), .SD(index_q[6]), .Z(n20267));
    LUT4 n285_bdd_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n23809)) /* synthesis lut_function=(A (B (C)+!B ((D)+!C))+!A (B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n285_bdd_3_lut_4_lut_4_lut_4_lut.init = 16'he7c7;
    LUT4 i18813_3_lut (.A(n23919), .B(n23985), .C(index_i[6]), .Z(n21143)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18813_3_lut.init = 16'hcaca;
    L6MUX21 i17938 (.D0(n20253), .D1(n20254), .SD(index_q[6]), .Z(n20268));
    LUT4 mux_193_Mux_0_i428_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_q[2]), 
         .B(index_q[0]), .C(index_q[1]), .D(index_q[3]), .Z(n428_adj_2301)) /* synthesis lut_function=(A (B (C+!(D))+!B !((D)+!C))+!A (B (D)+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i428_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hd5a9;
    LUT4 mux_192_Mux_7_i781_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), 
         .B(index_i[2]), .C(index_i[3]), .D(index_i[0]), .Z(n781_adj_2302)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_7_i781_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h1e1c;
    LUT4 mux_193_Mux_0_i971_3_lut (.A(n27523), .B(n25189), .C(index_q[3]), 
         .Z(n971)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i971_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_7_i747_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), 
         .B(index_i[2]), .C(index_i[3]), .D(index_i[0]), .Z(n747_adj_2303)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))+!A (B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_7_i747_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'he1e3;
    L6MUX21 i18837 (.D0(n20903), .D1(n20906), .SD(index_i[6]), .Z(n21167));
    LUT4 i19098_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n21428)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(D))+!A (B (D)+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19098_3_lut_4_lut_4_lut_4_lut.init = 16'hd52b;
    L6MUX21 i17939 (.D0(n20255), .D1(n20256), .SD(index_q[6]), .Z(n20269));
    LUT4 i9364_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n11930)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D))+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9364_3_lut_4_lut_4_lut_4_lut.init = 16'hcadd;
    L6MUX21 i17940 (.D0(n20257), .D1(n20258), .SD(index_q[6]), .Z(n20270));
    L6MUX21 i17941 (.D0(n20259), .D1(n20260), .SD(index_q[6]), .Z(n20271));
    L6MUX21 i17943 (.D0(n20263), .D1(n20264), .SD(index_q[6]), .Z(n20273));
    LUT4 i17948_3_lut (.A(n20273), .B(n23225), .C(index_q[7]), .Z(n20278)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17948_3_lut.init = 16'hcaca;
    LUT4 i19161_3_lut_4_lut (.A(n25163), .B(index_i[2]), .C(index_i[3]), 
         .D(n141), .Z(n21491)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19161_3_lut_4_lut.init = 16'hf202;
    PFUMX mux_193_Mux_2_i891 (.BLUT(n875_adj_2255), .ALUT(n890_adj_2304), 
          .C0(index_q[4]), .Z(n891_adj_2305)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    L6MUX21 i18748 (.D0(n21070), .D1(n21071), .SD(index_q[6]), .Z(n21078));
    L6MUX21 i18751 (.D0(n21076), .D1(n21077), .SD(index_q[6]), .Z(n21081));
    LUT4 i18116_3_lut (.A(n20439), .B(n23438), .C(index_i[7]), .Z(n20446)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18116_3_lut.init = 16'hcaca;
    L6MUX21 i17955 (.D0(n20973), .D1(n20976), .SD(index_i[6]), .Z(n20285));
    LUT4 i17947_3_lut (.A(n20271), .B(n20272), .C(index_q[7]), .Z(n20277)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17947_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_7_i747_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), 
         .B(index_q[2]), .C(index_q[3]), .D(index_q[0]), .Z(n747_adj_2306)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))+!A (B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_7_i747_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'he1e3;
    L6MUX21 i17956 (.D0(n20979), .D1(n20982), .SD(index_i[6]), .Z(n20286));
    LUT4 mux_193_Mux_7_i781_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), 
         .B(index_q[2]), .C(index_q[3]), .D(index_q[0]), .Z(n781_adj_2307)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_7_i781_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h1e1c;
    LUT4 quarter_wave_sample_register_i_9__I_0_3_lut (.A(quarter_wave_sample_register_i[9]), 
         .B(o_val_pipeline_i_0__15__N_2157[9]), .C(phase_negation_i[1]), 
         .Z(o_val_pipeline_i_0__15__N_2168)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[14] 77[8])
    defparam quarter_wave_sample_register_i_9__I_0_3_lut.init = 16'hcaca;
    LUT4 i9507_3_lut_3_lut_4_lut_4_lut (.A(index_q[2]), .B(index_q[3]), 
         .C(index_q[0]), .D(index_q[1]), .Z(n762_adj_2308)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C (D)+!C !(D)))+!A !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9507_3_lut_3_lut_4_lut_4_lut.init = 16'h700f;
    PFUMX mux_193_Mux_2_i860 (.BLUT(n844_adj_2309), .ALUT(n859_adj_2310), 
          .C0(index_q[4]), .Z(n860_adj_2311)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 n543_bdd_4_lut_22363_4_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[5]), .D(index_i[2]), .Z(n23981)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n543_bdd_4_lut_22363_4_lut_4_lut.init = 16'hd23d;
    LUT4 i20932_3_lut (.A(n20277), .B(n20278), .C(index_q[8]), .Z(n20280)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20932_3_lut.init = 16'hcaca;
    L6MUX21 i17957 (.D0(n20985), .D1(n20988), .SD(index_i[6]), .Z(n20287));
    LUT4 i19044_3_lut_4_lut (.A(index_q[1]), .B(index_q[0]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21374)) /* synthesis lut_function=(A (B+(C+(D)))+!A !(B (C+(D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19044_3_lut_4_lut.init = 16'haabd;
    LUT4 i12133_2_lut_rep_603 (.A(index_i[0]), .B(index_i[1]), .Z(n25163)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i12133_2_lut_rep_603.init = 16'heeee;
    LUT4 i18895_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n21225)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C))+!A (B (C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18895_3_lut_4_lut_4_lut_4_lut.init = 16'he078;
    L6MUX21 i18599 (.D0(n20855), .D1(n20862), .SD(index_q[6]), .Z(n20929));
    LUT4 i18753_3_lut (.A(n21080), .B(n21081), .C(index_q[7]), .Z(n21083)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18753_3_lut.init = 16'hcaca;
    LUT4 i18499_3_lut_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n20829)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C+!(D))+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18499_3_lut_3_lut_4_lut_4_lut.init = 16'h1f81;
    LUT4 mux_192_Mux_2_i890_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n890_adj_2280)) /* synthesis lut_function=(A (B (C)+!B !(C+!(D)))+!A !(B (C+(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_2_i890_3_lut_4_lut_4_lut.init = 16'h9394;
    LUT4 i18752_3_lut (.A(n21078), .B(n21079), .C(index_q[7]), .Z(n21082)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18752_3_lut.init = 16'hcaca;
    L6MUX21 i18817 (.D0(n21135), .D1(n21136), .SD(index_i[6]), .Z(n21147));
    LUT4 i19127_3_lut_4_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n21457)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B+(C+(D))))) */ ;
    defparam i19127_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'h2aab;
    LUT4 mux_193_Mux_8_i157_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n15)) /* synthesis lut_function=(A (B (C)+!B !(C (D)+!C !(D)))+!A !(B ((D)+!C)+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_8_i157_3_lut_4_lut_4_lut.init = 16'h83e0;
    LUT4 i18585_3_lut_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n20915)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C+!(D))+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18585_3_lut_3_lut_4_lut_4_lut.init = 16'h1f81;
    LUT4 mux_192_Mux_8_i61_3_lut_rep_278_4_lut_4_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[2]), .D(index_i[3]), .Z(n24838)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A (B (C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_8_i61_3_lut_rep_278_4_lut_4_lut_4_lut.init = 16'he0f8;
    LUT4 mux_192_Mux_8_i251_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[2]), .D(index_i[3]), .Z(n251_adj_2312)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_8_i251_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h07e0;
    LUT4 mux_192_Mux_8_i157_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n157_adj_2313)) /* synthesis lut_function=(A (B (C)+!B !(C (D)+!C !(D)))+!A !(B ((D)+!C)+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_8_i157_3_lut_4_lut_4_lut.init = 16'h83e0;
    LUT4 i19083_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n21413)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C))+!A (B (C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19083_3_lut_4_lut_4_lut_4_lut.init = 16'he078;
    LUT4 i18584_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n20914)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18584_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hf81f;
    LUT4 mux_193_Mux_6_i890_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), 
         .B(index_q[1]), .C(index_q[2]), .D(index_q[3]), .Z(n890_adj_2314)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !((D)+!C))+!A !(B ((D)+!C)+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_6_i890_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h7e07;
    LUT4 mux_193_Mux_7_i699_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n699_adj_2315)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C+!(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_7_i699_3_lut_4_lut_4_lut.init = 16'hf07e;
    L6MUX21 i18818 (.D0(n21137), .D1(n21138), .SD(index_i[6]), .Z(n21148));
    LUT4 mux_193_Mux_8_i61_3_lut_rep_280_4_lut_4_lut_4_lut (.A(index_q[0]), 
         .B(index_q[1]), .C(index_q[2]), .D(index_q[3]), .Z(n24840)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A (B (C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_8_i61_3_lut_rep_280_4_lut_4_lut_4_lut.init = 16'he0f8;
    LUT4 i18498_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n20828)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18498_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hf81f;
    LUT4 mux_193_Mux_8_i109_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n109)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C+!(D)))+!A (B (C (D)+!C !(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_8_i109_3_lut_4_lut_4_lut.init = 16'hf83e;
    LUT4 mux_193_Mux_0_i460_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n460)) /* synthesis lut_function=(A (B+(C (D)+!C !(D)))+!A (B (C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i460_3_lut_4_lut_4_lut.init = 16'hf8cb;
    LUT4 mux_193_Mux_0_i364_3_lut_3_lut_4_lut (.A(index_q[1]), .B(index_q[0]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n364_adj_2316)) /* synthesis lut_function=(A (B (D)+!B (C+!(D)))+!A !(B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i364_3_lut_3_lut_4_lut.init = 16'hbd33;
    L6MUX21 i18819 (.D0(n21139), .D1(n21140), .SD(index_i[6]), .Z(n21149));
    LUT4 i18500_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n20830)) /* synthesis lut_function=(A (B (C+!(D))+!B !((D)+!C))+!A !(B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18500_3_lut_4_lut_4_lut.init = 16'h81f8;
    LUT4 mux_193_Mux_8_i251_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), 
         .B(index_q[1]), .C(index_q[2]), .D(index_q[3]), .Z(n251_adj_2317)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_8_i251_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h07e0;
    LUT4 mux_193_Mux_0_i716_3_lut (.A(n25185), .B(n25201), .C(index_q[3]), 
         .Z(n716_adj_2318)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i716_3_lut.init = 16'hcaca;
    LUT4 i11478_2_lut_3_lut_4_lut (.A(n24985), .B(n25053), .C(index_i[6]), 
         .D(index_i[5]), .Z(n254)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11478_2_lut_3_lut_4_lut.init = 16'hfef0;
    LUT4 i9555_3_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[3]), .C(index_i[0]), 
         .D(index_i[1]), .Z(n844)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9555_3_lut_4_lut_4_lut.init = 16'hf00e;
    PFUMX i23058 (.BLUT(n25296), .ALUT(n25297), .C0(index_q[3]), .Z(n62_adj_2319));
    CCU2D add_357_7 (.A0(quarter_wave_sample_register_i[6]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[7]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17321), .COUT(n17322), 
          .S1(o_val_pipeline_i_0__15__N_2157[7]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam add_357_7.INIT0 = 16'hf555;
    defparam add_357_7.INIT1 = 16'hf555;
    defparam add_357_7.INJECT1_0 = "NO";
    defparam add_357_7.INJECT1_1 = "NO";
    PFUMX i18621 (.BLUT(n20947), .ALUT(n20948), .C0(index_i[4]), .Z(n20951));
    LUT4 mux_193_Mux_0_i939_4_lut (.A(n588), .B(n25181), .C(index_q[3]), 
         .D(index_q[2]), .Z(n939)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i939_4_lut.init = 16'hfaca;
    PFUMX i23056 (.BLUT(n25293), .ALUT(n25294), .C0(index_q[1]), .Z(n25295));
    LUT4 i2_2_lut_rep_304_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(n25090), 
         .D(index_q[2]), .Z(n24864)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i2_2_lut_rep_304_3_lut_4_lut.init = 16'hfff8;
    LUT4 mux_193_Mux_0_i653_3_lut (.A(n25156), .B(n25183), .C(index_q[3]), 
         .Z(n653_adj_2320)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i653_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_7_i956_3_lut_3_lut_4_lut (.A(n24945), .B(index_i[4]), 
         .C(n924_adj_2321), .D(index_i[5]), .Z(n956)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_7_i956_3_lut_3_lut_4_lut.init = 16'h11f0;
    LUT4 index_i_5__bdd_4_lut_22661 (.A(n85), .B(index_i[2]), .C(index_i[3]), 
         .D(n25163), .Z(n23626)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (B+!(C (D))))) */ ;
    defparam index_i_5__bdd_4_lut_22661.init = 16'h3a0a;
    LUT4 i19037_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n21367)) /* synthesis lut_function=(!(A (B (C (D)))+!A !(B+(C+(D))))) */ ;
    defparam i19037_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h7ffe;
    LUT4 i19103_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n21433)) /* synthesis lut_function=(A (B (C (D)))+!A !(B+(C+(D)))) */ ;
    defparam i19103_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h8001;
    LUT4 mux_193_Mux_0_i620_3_lut (.A(n25194), .B(n25206), .C(index_q[3]), 
         .Z(n620_adj_2322)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i620_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_0_i379_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n379_adj_2323)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !((D)+!C))+!A !(B ((D)+!C)+!B (D))) */ ;
    defparam mux_193_Mux_0_i379_3_lut_4_lut_4_lut.init = 16'h8079;
    LUT4 mux_193_Mux_0_i589_3_lut (.A(n27521), .B(n588), .C(index_q[3]), 
         .Z(n589_adj_2324)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i589_3_lut.init = 16'hcaca;
    PFUMX i18820 (.BLUT(n21141), .ALUT(n21142), .C0(index_i[6]), .Z(n21150));
    LUT4 i18965_3_lut_3_lut_4_lut (.A(n24945), .B(index_i[4]), .C(n252), 
         .D(index_i[5]), .Z(n21295)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18965_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 mux_193_Mux_8_i443_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n443_adj_2325)) /* synthesis lut_function=(A (B (C+!(D))+!B !((D)+!C))+!A !(B (D)+!B ((D)+!C))) */ ;
    defparam mux_193_Mux_8_i443_3_lut_4_lut_4_lut.init = 16'h80fc;
    LUT4 mux_193_Mux_5_i252_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[4]), .Z(n252_adj_2326)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+(D)))+!A (B (C (D))+!B !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_5_i252_3_lut_4_lut.init = 16'hc993;
    LUT4 mux_192_Mux_8_i109_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n109_adj_2327)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C+!(D)))+!A (B (C (D)+!C !(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_8_i109_3_lut_4_lut_4_lut.init = 16'hf83e;
    L6MUX21 i18838 (.D0(n12043), .D1(n20909), .SD(index_i[6]), .Z(n21168));
    L6MUX21 i18840 (.D0(n20922), .D1(n20925), .SD(index_i[6]), .Z(n21170));
    L6MUX21 i18841 (.D0(n574), .D1(n20928), .SD(index_i[6]), .Z(n21171));
    PFUMX i18622 (.BLUT(n20949), .ALUT(n20950), .C0(index_i[4]), .Z(n20952));
    L6MUX21 i18842 (.D0(n20946), .D1(n764_adj_2328), .SD(index_i[6]), 
            .Z(n21172));
    LUT4 mux_192_Mux_0_i460_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n460_adj_2329)) /* synthesis lut_function=(A (B+(C (D)+!C !(D)))+!A (B (C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_0_i460_3_lut_4_lut_4_lut.init = 16'hf8cb;
    LUT4 i18586_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n20916)) /* synthesis lut_function=(A (B (C+!(D))+!B !((D)+!C))+!A !(B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18586_3_lut_4_lut_4_lut.init = 16'h81f8;
    LUT4 mux_193_Mux_0_i890_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n890)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)+!C !(D)))+!A !(B (C)+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i890_3_lut_4_lut_4_lut.init = 16'h70ca;
    LUT4 mux_192_Mux_0_i604_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n604)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)+!C !(D)))+!A (B (C (D))+!B (C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_0_i604_3_lut_4_lut_4_lut.init = 16'h0e65;
    LUT4 mux_192_Mux_0_i890_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n890_adj_2264)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)+!C !(D)))+!A !(B (C)+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_0_i890_3_lut_4_lut_4_lut.init = 16'h70ca;
    LUT4 i19223_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n21553)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B+(C+(D))))) */ ;
    defparam i19223_3_lut_4_lut_4_lut_4_lut.init = 16'h2aab;
    LUT4 mux_192_Mux_7_i699_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n699_adj_2330)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C+!(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_7_i699_3_lut_4_lut_4_lut.init = 16'hf07e;
    LUT4 i18691_3_lut (.A(n21018), .B(n21019), .C(index_i[7]), .Z(n21021)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18691_3_lut.init = 16'hcaca;
    LUT4 quarter_wave_sample_register_i_8__I_0_3_lut (.A(quarter_wave_sample_register_i[8]), 
         .B(o_val_pipeline_i_0__15__N_2157[8]), .C(phase_negation_i[1]), 
         .Z(o_val_pipeline_i_0__15__N_2170)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[14] 77[8])
    defparam quarter_wave_sample_register_i_8__I_0_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_10_i701_4_lut_4_lut (.A(n24945), .B(index_i[4]), .C(index_i[5]), 
         .D(n24884), .Z(n701_adj_2284)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B (C (D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_10_i701_4_lut_4_lut.init = 16'h3efe;
    LUT4 mux_192_Mux_5_i252_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[4]), .Z(n252_adj_2331)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+(D)))+!A (B (C (D))+!B !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_5_i252_3_lut_4_lut.init = 16'hc993;
    LUT4 mux_192_Mux_1_i716_3_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[1]), .D(index_i[3]), .Z(n716_adj_2332)) /* synthesis lut_function=(!(A (B (D)+!B !(C))+!A !(B (C (D))+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_1_i716_3_lut_4_lut_4_lut.init = 16'h70a9;
    LUT4 i18690_3_lut (.A(n21016), .B(n21017), .C(index_i[7]), .Z(n21020)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18690_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_8_i397_3_lut_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n397)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B ((D)+!C))) */ ;
    defparam mux_192_Mux_8_i397_3_lut_3_lut_3_lut_4_lut.init = 16'hf10f;
    L6MUX21 i17983 (.D0(n20297), .D1(n20298), .SD(index_q[6]), .Z(n20313));
    LUT4 i19344_3_lut (.A(n25204), .B(n25184), .C(index_q[3]), .Z(n21674)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19344_3_lut.init = 16'hcaca;
    LUT4 i19343_3_lut (.A(n325), .B(n332), .C(index_q[3]), .Z(n21673)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19343_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_0_i412_3_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[1]), .D(index_i[3]), .Z(n412_adj_2333)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C (D)))+!A (B (C+!(D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_0_i412_3_lut_4_lut_4_lut.init = 16'hf14c;
    PFUMX i18628 (.BLUT(n20954), .ALUT(n20955), .C0(index_i[4]), .Z(n20958));
    L6MUX21 i17984 (.D0(n20299), .D1(n20300), .SD(index_q[6]), .Z(n20314));
    L6MUX21 i17985 (.D0(n20301), .D1(n20302), .SD(index_q[6]), .Z(n20315));
    PFUMX i17987 (.BLUT(n20305), .ALUT(n20306), .C0(index_q[6]), .Z(n20317));
    L6MUX21 i17988 (.D0(n20307), .D1(n20308), .SD(index_q[6]), .Z(n20318));
    L6MUX21 i17989 (.D0(n20309), .D1(n20310), .SD(index_q[6]), .Z(n20319));
    PFUMX i17990 (.BLUT(n20311), .ALUT(n20312), .C0(index_q[6]), .Z(n20320));
    LUT4 n557_bdd_3_lut_22513 (.A(n25047), .B(n25087), .C(index_i[3]), 
         .Z(n23629)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n557_bdd_3_lut_22513.init = 16'hcaca;
    PFUMX i23054 (.BLUT(n25290), .ALUT(n25291), .C0(index_i[1]), .Z(n25292));
    LUT4 mux_193_Mux_0_i412_3_lut_4_lut_4_lut (.A(index_q[2]), .B(index_q[0]), 
         .C(index_q[1]), .D(index_q[3]), .Z(n412_adj_2334)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C (D)))+!A (B (C+!(D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i412_3_lut_4_lut_4_lut.init = 16'hf14c;
    PFUMX i18629 (.BLUT(n20956), .ALUT(n20957), .C0(index_i[4]), .Z(n20959));
    LUT4 mux_193_Mux_0_i604_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n604_adj_2335)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)+!C !(D)))+!A (B (C (D))+!B (C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i604_3_lut_4_lut_4_lut.init = 16'h0e65;
    LUT4 mux_193_Mux_1_i684_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n684_adj_2336)) /* synthesis lut_function=(A (B ((D)+!C)+!B !((D)+!C))+!A !(B (C+(D))+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_1_i684_3_lut_4_lut_4_lut.init = 16'h992d;
    PFUMX mux_193_Mux_7_i253 (.BLUT(n12168), .ALUT(n12010), .C0(n19828), 
          .Z(n253)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 mux_193_Mux_7_i762_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), 
         .B(index_q[2]), .C(index_q[3]), .D(index_q[0]), .Z(n762_adj_2337)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B ((D)+!C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_7_i762_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h3878;
    L6MUX21 i18014 (.D0(n20328), .D1(n20329), .SD(index_q[6]), .Z(n20344));
    LUT4 i11560_3_lut_4_lut (.A(n24946), .B(index_i[4]), .C(index_i[5]), 
         .D(index_i[6]), .Z(n127)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11560_3_lut_4_lut.init = 16'hf800;
    L6MUX21 i18015 (.D0(n20330), .D1(n20331), .SD(index_q[6]), .Z(n20345));
    L6MUX21 i18016 (.D0(n20332), .D1(n20333), .SD(index_q[6]), .Z(n20346));
    L6MUX21 i18017 (.D0(n20334), .D1(n20335), .SD(index_q[6]), .Z(n20347));
    PFUMX i18635 (.BLUT(n20961), .ALUT(n20962), .C0(index_i[4]), .Z(n20965));
    LUT4 n301_bdd_3_lut_22884_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .D(index_q[0]), .Z(n23782)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A !((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n301_bdd_3_lut_22884_4_lut_4_lut_4_lut.init = 16'h7173;
    PFUMX i23150 (.BLUT(n25459), .ALUT(n25454), .C0(index_i[3]), .Z(n25460));
    LUT4 mux_193_Mux_9_i316_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), 
         .B(index_q[2]), .C(index_q[3]), .D(index_q[0]), .Z(n316_adj_2338)) /* synthesis lut_function=(!(A (B (C)+!B !(C+(D)))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_9_i316_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h7e7c;
    CCU2D add_357_5 (.A0(quarter_wave_sample_register_i[4]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[5]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17320), .COUT(n17321));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam add_357_5.INIT0 = 16'hf555;
    defparam add_357_5.INIT1 = 16'hf555;
    defparam add_357_5.INJECT1_0 = "NO";
    defparam add_357_5.INJECT1_1 = "NO";
    LUT4 i18050_3_lut (.A(n20369), .B(n20370), .C(index_i[6]), .Z(n20380)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18050_3_lut.init = 16'hcaca;
    L6MUX21 i18018 (.D0(n20336), .D1(n20337), .SD(index_q[6]), .Z(n20348));
    LUT4 n10495_bdd_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .D(index_q[0]), .Z(n23785)) /* synthesis lut_function=(A (B (C)+!B ((D)+!C))+!A (B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n10495_bdd_3_lut_4_lut_4_lut_4_lut.init = 16'he7c7;
    LUT4 i19092_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .D(index_q[0]), .Z(n21422)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B (C+(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19092_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h7c78;
    LUT4 i9530_3_lut_4_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n844_adj_2309)) /* synthesis lut_function=(A (B)+!A !(B+!(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9530_3_lut_4_lut_3_lut_4_lut.init = 16'h9998;
    L6MUX21 i18020 (.D0(n20340), .D1(n20341), .SD(index_q[6]), .Z(n20350));
    LUT4 mux_193_Mux_2_i890_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n890_adj_2304)) /* synthesis lut_function=(A (B (C)+!B !(C+!(D)))+!A !(B (C+(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_2_i890_3_lut_4_lut_4_lut.init = 16'h9394;
    LUT4 i18963_3_lut_3_lut_4_lut (.A(n24946), .B(index_i[4]), .C(n125), 
         .D(index_i[5]), .Z(n21293)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18963_3_lut_3_lut_4_lut.init = 16'hf077;
    L6MUX21 i18941 (.D0(n21259), .D1(n21260), .SD(index_q[6]), .Z(n21271));
    LUT4 i9473_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n12039)) /* synthesis lut_function=(!(A (B (C)+!B ((D)+!C))+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9473_3_lut_4_lut_4_lut.init = 16'h4969;
    LUT4 mux_192_Mux_2_i836_3_lut_4_lut_3_lut_rep_679 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27519)) /* synthesis lut_function=(A (B)+!A !(B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_2_i836_3_lut_4_lut_3_lut_rep_679.init = 16'h9898;
    LUT4 mux_192_Mux_11_i445_3_lut_4_lut_4_lut_4_lut (.A(index_i[3]), .B(index_i[4]), 
         .C(index_i[5]), .D(n24985), .Z(n445)) /* synthesis lut_function=(!(A (B (C))+!A !(B+(C+(D))))) */ ;
    defparam mux_192_Mux_11_i445_3_lut_4_lut_4_lut_4_lut.init = 16'h7f7e;
    LUT4 mux_193_Mux_11_i445_3_lut_4_lut_4_lut_4_lut (.A(index_q[3]), .B(index_q[4]), 
         .C(index_q[5]), .D(n24959), .Z(n445_adj_2339)) /* synthesis lut_function=(!(A (B (C))+!A !(B+(C+(D))))) */ ;
    defparam mux_193_Mux_11_i445_3_lut_4_lut_4_lut_4_lut.init = 16'h7f7e;
    LUT4 mux_192_Mux_1_i684_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n684_adj_2340)) /* synthesis lut_function=(A (B ((D)+!C)+!B !((D)+!C))+!A !(B (C+(D))+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_1_i684_3_lut_4_lut_4_lut.init = 16'h992d;
    LUT4 mux_193_Mux_1_i716_3_lut_4_lut_4_lut (.A(index_q[2]), .B(index_q[0]), 
         .C(index_q[1]), .D(index_q[3]), .Z(n716_adj_2341)) /* synthesis lut_function=(!(A (B (D)+!B !(C))+!A !(B (C (D))+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_1_i716_3_lut_4_lut_4_lut.init = 16'h70a9;
    LUT4 i19331_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21661)) /* synthesis lut_function=(A (C)+!A !(B (C)+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19331_3_lut_4_lut_4_lut.init = 16'hb4b5;
    L6MUX21 i18021 (.D0(n20342), .D1(n20343), .SD(index_q[6]), .Z(n20351));
    L6MUX21 i18942 (.D0(n21261), .D1(n21262), .SD(index_q[6]), .Z(n21272));
    LUT4 i12082_3_lut (.A(index_q[2]), .B(index_q[1]), .C(index_q[0]), 
         .Z(n1001)) /* synthesis lut_function=(A (B)+!A (B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12082_3_lut.init = 16'hdcdc;
    L6MUX21 i18943 (.D0(n21263), .D1(n21264), .SD(index_q[6]), .Z(n21273));
    LUT4 i11173_2_lut_3_lut_4_lut (.A(n24959), .B(n25090), .C(index_q[6]), 
         .D(index_q[5]), .Z(n254_adj_2342)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i11173_2_lut_3_lut_4_lut.init = 16'hfef0;
    PFUMX i18944 (.BLUT(n21265), .ALUT(n21266), .C0(index_q[6]), .Z(n21274));
    LUT4 n22_bdd_3_lut_23557 (.A(n27503), .B(n25079), .C(index_i[3]), 
         .Z(n23633)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n22_bdd_3_lut_23557.init = 16'hacac;
    LUT4 mux_193_Mux_7_i956_3_lut_3_lut_4_lut (.A(n24948), .B(index_q[4]), 
         .C(n924_adj_2343), .D(index_q[5]), .Z(n956_adj_2344)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_7_i956_3_lut_3_lut_4_lut.init = 16'h11f0;
    LUT4 n572_bdd_3_lut_22979 (.A(n978), .B(n25047), .C(index_i[3]), .Z(n23635)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n572_bdd_3_lut_22979.init = 16'hcaca;
    LUT4 i18997_3_lut_3_lut_4_lut (.A(n24948), .B(index_q[4]), .C(n252_adj_2345), 
         .D(index_q[5]), .Z(n21327)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18997_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 mux_193_Mux_10_i701_4_lut_4_lut (.A(n24948), .B(index_q[4]), .C(index_q[5]), 
         .D(n24876), .Z(n701)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B (C (D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_10_i701_4_lut_4_lut.init = 16'h3efe;
    LUT4 i11191_3_lut_4_lut (.A(n24949), .B(index_q[4]), .C(index_q[5]), 
         .D(index_q[6]), .Z(n127_adj_2346)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11191_3_lut_4_lut.init = 16'hf800;
    LUT4 i18995_3_lut_3_lut_4_lut (.A(n24949), .B(index_q[4]), .C(n125_adj_2347), 
         .D(index_q[5]), .Z(n21325)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18995_3_lut_3_lut_4_lut.init = 16'hf077;
    LUT4 n123_bdd_3_lut_22042 (.A(n25082), .B(n25087), .C(index_i[3]), 
         .Z(n23645)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n123_bdd_3_lut_22042.init = 16'hacac;
    LUT4 mux_192_Mux_0_i762_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n762)) /* synthesis lut_function=(A (B+!((D)+!C))+!A !(B (D)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_0_i762_3_lut_4_lut_4_lut.init = 16'h98fc;
    LUT4 i20937_3_lut (.A(n24740), .B(n23186), .C(index_i[8]), .Z(n20249)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20937_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_1_i747_4_lut_then_4_lut (.A(index_i[0]), .B(index_i[4]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n25244)) /* synthesis lut_function=(A (B ((D)+!C))+!A !(B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_1_i747_4_lut_then_4_lut.init = 16'h9d5d;
    PFUMX i23050 (.BLUT(n25284), .ALUT(n25285), .C0(index_i[3]), .Z(n62_adj_2348));
    LUT4 i2_2_lut_rep_303_3_lut_4_lut (.A(index_i[3]), .B(index_i[4]), .C(index_i[2]), 
         .D(n25058), .Z(n24863)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i2_2_lut_rep_303_3_lut_4_lut.init = 16'hfffe;
    LUT4 n396_bdd_3_lut_22239 (.A(n25166), .B(n25068), .C(index_i[3]), 
         .Z(n23654)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n396_bdd_3_lut_22239.init = 16'hcaca;
    PFUMX i18636 (.BLUT(n20963), .ALUT(n20964), .C0(index_i[4]), .Z(n20966));
    LUT4 mux_192_Mux_7_i762_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n762_adj_2349)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A (B (C (D)+!C !(D))+!B !(C)))) */ ;
    defparam mux_192_Mux_7_i762_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h1cf0;
    LUT4 i11229_2_lut_rep_297_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n24857)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11229_2_lut_rep_297_3_lut_4_lut.init = 16'hf080;
    LUT4 mux_193_Mux_0_i363_3_lut_4_lut_4_lut_3_lut_rep_654 (.A(index_q[1]), 
         .B(index_q[0]), .C(index_q[2]), .Z(n27494)) /* synthesis lut_function=(A (B+(C))+!A !(B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i363_3_lut_4_lut_4_lut_3_lut_rep_654.init = 16'hbdbd;
    LUT4 i9602_3_lut_3_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[0]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n12172)) /* synthesis lut_function=(!(A (B (D)+!B !(C+(D)))+!A (B (C+(D))+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9602_3_lut_3_lut_4_lut_4_lut.init = 16'h22bd;
    LUT4 mux_193_Mux_10_i62_3_lut_3_lut_4_lut (.A(n24956), .B(index_q[3]), 
         .C(n24938), .D(index_q[4]), .Z(n62_adj_2350)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_10_i62_3_lut_3_lut_4_lut.init = 16'hf077;
    LUT4 mux_192_Mux_6_i459_3_lut_4_lut_3_lut_rep_656 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27496)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_6_i459_3_lut_4_lut_3_lut_rep_656.init = 16'h4d4d;
    LUT4 mux_193_Mux_8_i860_3_lut_4_lut (.A(n24956), .B(index_q[3]), .C(index_q[4]), 
         .D(n24938), .Z(n860_adj_2351)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_8_i860_3_lut_4_lut.init = 16'h08f8;
    LUT4 mux_193_Mux_3_i252_3_lut_4_lut (.A(n24956), .B(index_q[3]), .C(index_q[4]), 
         .D(n14996), .Z(n252_adj_2352)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_3_i252_3_lut_4_lut.init = 16'h08f8;
    PFUMX i18959 (.BLUT(n21285), .ALUT(n21286), .C0(index_i[6]), .Z(n21289));
    PFUMX i18960 (.BLUT(n21287), .ALUT(n21288), .C0(index_i[6]), .Z(n21290));
    LUT4 mux_193_Mux_6_i955_3_lut_4_lut (.A(n24956), .B(index_q[3]), .C(index_q[4]), 
         .D(n24817), .Z(n955)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_6_i955_3_lut_4_lut.init = 16'h8f80;
    LUT4 i18355_3_lut_4_lut (.A(n24956), .B(index_q[3]), .C(index_q[4]), 
         .D(n364_adj_2353), .Z(n20685)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18355_3_lut_4_lut.init = 16'h8f80;
    PFUMX i18966 (.BLUT(n21292), .ALUT(n21293), .C0(index_i[6]), .Z(n21296));
    LUT4 i11181_2_lut_rep_251_3_lut_4_lut (.A(n24956), .B(index_q[3]), .C(index_q[5]), 
         .D(index_q[4]), .Z(n24811)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11181_2_lut_rep_251_3_lut_4_lut.init = 16'hf080;
    LUT4 mux_193_Mux_3_i189_3_lut_3_lut_4_lut (.A(n24956), .B(index_q[3]), 
         .C(index_q[4]), .D(n24904), .Z(n189)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_3_i189_3_lut_3_lut_4_lut.init = 16'h08f8;
    PFUMX i18967 (.BLUT(n21294), .ALUT(n21295), .C0(index_i[6]), .Z(n21297));
    LUT4 n124_bdd_3_lut_22592_4_lut (.A(n24957), .B(index_q[3]), .C(index_q[4]), 
         .D(n93_adj_2354), .Z(n23039)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n124_bdd_3_lut_22592_4_lut.init = 16'hfe0e;
    LUT4 quarter_wave_sample_register_i_7__I_0_3_lut (.A(quarter_wave_sample_register_i[7]), 
         .B(o_val_pipeline_i_0__15__N_2157[7]), .C(phase_negation_i[1]), 
         .Z(o_val_pipeline_i_0__15__N_2172)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[14] 77[8])
    defparam quarter_wave_sample_register_i_7__I_0_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_10_i317_3_lut_3_lut_4_lut (.A(n24957), .B(index_q[3]), 
         .C(n24904), .D(index_q[4]), .Z(n317)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_10_i317_3_lut_3_lut_4_lut.init = 16'hf011;
    L6MUX21 i18969 (.D0(n20817), .D1(n20820), .SD(index_q[6]), .Z(n21299));
    L6MUX21 i18970 (.D0(n12003), .D1(n20823), .SD(index_q[6]), .Z(n21300));
    LUT4 i18353_3_lut_3_lut_4_lut (.A(n24957), .B(index_q[3]), .C(n316_adj_2338), 
         .D(index_q[4]), .Z(n20683)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18353_3_lut_3_lut_4_lut.init = 16'hf011;
    L6MUX21 i18972 (.D0(n20836), .D1(n20839), .SD(index_q[6]), .Z(n21302));
    L6MUX21 i18973 (.D0(n574_adj_2355), .D1(n20842), .SD(index_q[6]), 
            .Z(n21303));
    LUT4 i19309_3_lut (.A(n25194), .B(n25156), .C(index_q[3]), .Z(n21639)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19309_3_lut.init = 16'hcaca;
    L6MUX21 i18974 (.D0(n20845), .D1(n764_adj_2356), .SD(index_q[6]), 
            .Z(n21304));
    LUT4 i11202_3_lut_4_lut (.A(n24957), .B(index_q[3]), .C(n25104), .D(index_q[6]), 
         .Z(n765)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11202_3_lut_4_lut.init = 16'hffe0;
    LUT4 i18514_3_lut_3_lut_4_lut (.A(n24957), .B(index_q[3]), .C(n93_adj_2354), 
         .D(index_q[4]), .Z(n20844)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18514_3_lut_3_lut_4_lut.init = 16'h11f0;
    LUT4 i19308_3_lut (.A(n25195), .B(n141_adj_2357), .C(index_q[3]), 
         .Z(n21638)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19308_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_10_i413_3_lut_4_lut (.A(n24959), .B(index_q[3]), .C(index_q[4]), 
         .D(n24904), .Z(n413)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_10_i413_3_lut_4_lut.init = 16'hf101;
    LUT4 mux_192_Mux_11_i638_4_lut_4_lut (.A(n24832), .B(index_i[5]), .C(index_i[6]), 
         .D(n24858), .Z(n638)) /* synthesis lut_function=(A (B (C (D))+!B !(C))+!A (B ((D)+!C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_11_i638_4_lut_4_lut.init = 16'hc707;
    CCU2D add_357_3 (.A0(quarter_wave_sample_register_i[2]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[3]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17319), .COUT(n17320));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam add_357_3.INIT0 = 16'hf555;
    defparam add_357_3.INIT1 = 16'hf555;
    defparam add_357_3.INJECT1_0 = "NO";
    defparam add_357_3.INJECT1_1 = "NO";
    L6MUX21 i18045 (.D0(n20359), .D1(n20360), .SD(index_i[6]), .Z(n20375));
    LUT4 mux_193_Mux_7_i173_3_lut (.A(n25205), .B(n25156), .C(index_q[3]), 
         .Z(n173)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_7_i173_3_lut.init = 16'hcaca;
    L6MUX21 i18046 (.D0(n20361), .D1(n20362), .SD(index_i[6]), .Z(n20376));
    LUT4 mux_193_Mux_10_i252_3_lut_4_lut_4_lut (.A(n24959), .B(index_q[3]), 
         .C(index_q[4]), .D(n24980), .Z(n252_adj_2345)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B (C (D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_10_i252_3_lut_4_lut_4_lut.init = 16'h3efe;
    L6MUX21 i18047 (.D0(n20363), .D1(n20364), .SD(index_i[6]), .Z(n20377));
    L6MUX21 i18048 (.D0(n20365), .D1(n20366), .SD(index_i[6]), .Z(n20378));
    L6MUX21 i18049 (.D0(n20367), .D1(n20368), .SD(index_i[6]), .Z(n20379));
    L6MUX21 i18051 (.D0(n20371), .D1(n20372), .SD(index_i[6]), .Z(n20381));
    CCU2D add_357_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(quarter_wave_sample_register_i[0]), .B1(quarter_wave_sample_register_i[1]), 
          .C1(GND_net), .D1(GND_net), .COUT(n17319));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam add_357_1.INIT0 = 16'hF000;
    defparam add_357_1.INIT1 = 16'ha666;
    defparam add_357_1.INJECT1_0 = "NO";
    defparam add_357_1.INJECT1_1 = "NO";
    L6MUX21 i22975 (.D0(n24738), .D1(n24787), .SD(index_i[6]), .Z(n24739));
    PFUMX i18313 (.BLUT(n318), .ALUT(n381), .C0(index_i[6]), .Z(n20643));
    PFUMX i22973 (.BLUT(n24737), .ALUT(n24736), .C0(index_i[5]), .Z(n24738));
    PFUMX mux_192_Mux_5_i732 (.BLUT(n12089), .ALUT(n731_adj_2358), .C0(index_i[4]), 
          .Z(n732_adj_2359)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 mux_193_Mux_3_i828_3_lut_3_lut_4_lut (.A(n24959), .B(index_q[3]), 
         .C(n157_adj_2360), .D(index_q[4]), .Z(n828)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_3_i828_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 i18359_3_lut_3_lut_4_lut (.A(n24959), .B(index_q[3]), .C(n412_adj_2361), 
         .D(index_q[4]), .Z(n20689)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18359_3_lut_3_lut_4_lut.init = 16'hf011;
    PFUMX i18307 (.BLUT(n574_adj_2362), .ALUT(n637), .C0(index_i[6]), 
          .Z(n20637));
    PFUMX i18304 (.BLUT(n574_adj_2363), .ALUT(n637_adj_2364), .C0(index_q[6]), 
          .Z(n20634));
    LUT4 i12268_1_lut_2_lut_3_lut_4_lut (.A(n24959), .B(index_q[3]), .C(index_q[5]), 
         .D(index_q[4]), .Z(n381_adj_2365)) /* synthesis lut_function=(!(A (C+(D))+!A (B (C+(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12268_1_lut_2_lut_3_lut_4_lut.init = 16'h010f;
    LUT4 mux_192_Mux_3_i653_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n653_adj_2366)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A !(B (D)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_3_i653_3_lut_4_lut_4_lut.init = 16'h4d99;
    PFUMX i18991 (.BLUT(n21317), .ALUT(n21318), .C0(index_q[6]), .Z(n21321));
    PFUMX i18270 (.BLUT(n318_adj_2367), .ALUT(n381_adj_2365), .C0(index_q[6]), 
          .Z(n20600));
    LUT4 mux_192_Mux_7_i53_3_lut_3_lut_rep_680 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27520)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_7_i53_3_lut_3_lut_rep_680.init = 16'hc7c7;
    PFUMX i23148 (.BLUT(n25457), .ALUT(n25456), .C0(index_i[6]), .Z(n25458));
    LUT4 i19169_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21499)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+(D)))+!A !(B (D)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19169_3_lut_4_lut_4_lut.init = 16'h99c7;
    LUT4 mux_193_Mux_0_i389_3_lut_3_lut_rep_681 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n27521)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i389_3_lut_3_lut_rep_681.init = 16'hc7c7;
    LUT4 i15266_3_lut (.A(n25184), .B(n25208), .C(index_q[3]), .Z(n17529)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15266_3_lut.init = 16'hcaca;
    LUT4 i19040_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21370)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+(D)))+!A !(B (D)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19040_3_lut_4_lut_4_lut.init = 16'h99c7;
    LUT4 i15265_3_lut (.A(n25208), .B(n25204), .C(index_q[3]), .Z(n17528)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15265_3_lut.init = 16'hcaca;
    PFUMX i18992 (.BLUT(n21319), .ALUT(n21320), .C0(index_q[6]), .Z(n21322));
    PFUMX i18666 (.BLUT(n142), .ALUT(n157), .C0(index_i[4]), .Z(n20996));
    LUT4 mux_193_Mux_11_i766_3_lut (.A(n638_adj_2368), .B(n765), .C(index_q[7]), 
         .Z(n766)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_11_i766_3_lut.init = 16'h3a3a;
    PFUMX i18667 (.BLUT(n173_adj_2369), .ALUT(n188), .C0(index_i[4]), 
          .Z(n20997));
    LUT4 n22932_bdd_3_lut (.A(n22932), .B(n476), .C(index_i[5]), .Z(n22933)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n22932_bdd_3_lut.init = 16'hcaca;
    PFUMX i18255 (.BLUT(n127), .ALUT(n254_adj_2370), .C0(index_i[7]), 
          .Z(n20585));
    PFUMX i18252 (.BLUT(n127_adj_2346), .ALUT(n254_adj_2371), .C0(index_q[7]), 
          .Z(n20582));
    LUT4 i11298_3_lut_3_lut_rep_655 (.A(index_q[1]), .B(index_q[0]), .C(index_q[2]), 
         .Z(n27495)) /* synthesis lut_function=(!(A+!((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11298_3_lut_3_lut_rep_655.init = 16'h5151;
    LUT4 i19115_3_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[0]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21445)) /* synthesis lut_function=(!(A ((D)+!C)+!A !(B (C (D))+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19115_3_lut_4_lut_4_lut.init = 16'h51a0;
    PFUMX i18998 (.BLUT(n21324), .ALUT(n21325), .C0(index_q[6]), .Z(n21328));
    PFUMX i18672 (.BLUT(n333), .ALUT(n348_adj_2372), .C0(index_i[4]), 
          .Z(n21002));
    PFUMX i18999 (.BLUT(n21326), .ALUT(n21327), .C0(index_q[6]), .Z(n21329));
    LUT4 mux_192_Mux_6_i38_3_lut_3_lut_rep_657 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27497)) /* synthesis lut_function=(A (B+(C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_6_i38_3_lut_3_lut_rep_657.init = 16'hadad;
    PFUMX i18673 (.BLUT(n364_adj_2373), .ALUT(n379_adj_2299), .C0(index_i[4]), 
          .Z(n21003));
    LUT4 n27411_bdd_3_lut_4_lut (.A(index_i[0]), .B(index_i[2]), .C(index_i[5]), 
         .D(n27411), .Z(n27412)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;
    defparam n27411_bdd_3_lut_4_lut.init = 16'h6f60;
    LUT4 n22936_bdd_3_lut_21935 (.A(n25292), .B(n22934), .C(index_i[5]), 
         .Z(n22937)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n22936_bdd_3_lut_21935.init = 16'hcaca;
    PFUMX i22947 (.BLUT(n24715), .ALUT(n24714), .C0(index_q[4]), .Z(n24716));
    LUT4 i19455_3_lut (.A(n21782), .B(n21783), .C(index_i[7]), .Z(n21785)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19455_3_lut.init = 16'hcaca;
    LUT4 i19454_3_lut (.A(n21780), .B(n21781), .C(index_i[7]), .Z(n21784)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19454_3_lut.init = 16'hcaca;
    LUT4 i18055_3_lut (.A(n20379), .B(n20380), .C(index_i[7]), .Z(n20385)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18055_3_lut.init = 16'hcaca;
    PFUMX i18674 (.BLUT(n397_adj_2374), .ALUT(n412_adj_2333), .C0(index_i[4]), 
          .Z(n21004));
    LUT4 n27396_bdd_3_lut_4_lut (.A(index_q[0]), .B(index_q[2]), .C(index_q[5]), 
         .D(n27396), .Z(n27397)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;
    defparam n27396_bdd_3_lut_4_lut.init = 16'h6f60;
    LUT4 index_q_6__bdd_3_lut_22015_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(n25096), .D(index_q[6]), .Z(n23060)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam index_q_6__bdd_3_lut_22015_4_lut.init = 16'hf07f;
    LUT4 i19229_3_lut (.A(n25077), .B(n25085), .C(index_i[3]), .Z(n21559)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19229_3_lut.init = 16'hcaca;
    LUT4 i20445_3_lut (.A(n21559), .B(n21560), .C(index_i[4]), .Z(n21561)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20445_3_lut.init = 16'hcaca;
    LUT4 i9550_3_lut_3_lut_4_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n762_adj_2291)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A (B))) */ ;
    defparam i9550_3_lut_3_lut_4_lut_3_lut_4_lut.init = 16'h1999;
    PFUMX i18675 (.BLUT(n428), .ALUT(n443_adj_2300), .C0(index_i[4]), 
          .Z(n21005));
    LUT4 i11589_2_lut_rep_382_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n24942)) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;
    defparam i11589_2_lut_rep_382_3_lut_4_lut.init = 16'he000;
    L6MUX21 i18077 (.D0(n20392), .D1(n20393), .SD(index_q[6]), .Z(n20407));
    LUT4 i19226_3_lut (.A(n38), .B(n978), .C(index_i[3]), .Z(n21556)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19226_3_lut.init = 16'hcaca;
    L6MUX21 i18078 (.D0(n20394), .D1(n20395), .SD(index_q[6]), .Z(n20408));
    LUT4 i20447_3_lut (.A(n21556), .B(n21557), .C(index_i[4]), .Z(n21558)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20447_3_lut.init = 16'hcaca;
    L6MUX21 i18079 (.D0(n20396), .D1(n20397), .SD(index_q[6]), .Z(n20409));
    PFUMX i21726 (.BLUT(n23279), .ALUT(n23276), .C0(index_q[6]), .Z(n23280));
    L6MUX21 i18080 (.D0(n20398), .D1(n20399), .SD(index_q[6]), .Z(n20410));
    L6MUX21 i18081 (.D0(n20400), .D1(n20401), .SD(index_q[6]), .Z(n20411));
    LUT4 i11981_3_lut_rep_682 (.A(index_q[2]), .B(index_q[1]), .C(index_q[0]), 
         .Z(n27522)) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11981_3_lut_rep_682.init = 16'hc4c4;
    LUT4 i18907_3_lut_4_lut_4_lut (.A(index_q[2]), .B(index_q[1]), .C(index_q[0]), 
         .D(index_q[3]), .Z(n21237)) /* synthesis lut_function=(A (B (C)+!B !(C+!(D)))+!A (B (C+!(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18907_3_lut_4_lut_4_lut.init = 16'hc3c4;
    PFUMX i23145 (.BLUT(n12175), .ALUT(n25451), .C0(index_i[5]), .Z(n25452));
    LUT4 i19218_3_lut (.A(n25083), .B(n25065), .C(index_i[3]), .Z(n21548)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19218_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_0_i963_3_lut_3_lut_rep_683 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n27523)) /* synthesis lut_function=(!(A (B)+!A (B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i963_3_lut_3_lut_rep_683.init = 16'h3636;
    LUT4 mux_192_Mux_0_i796_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n796)) /* synthesis lut_function=(A (B (C+(D))+!B (C (D)))+!A !(B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_0_i796_3_lut_4_lut_4_lut.init = 16'hadc0;
    LUT4 mux_193_Mux_6_i475_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n475_adj_2375)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A !(B (C+(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_6_i475_3_lut_4_lut_4_lut.init = 16'h9936;
    LUT4 n380_bdd_2_lut_4_lut (.A(n25163), .B(index_i[5]), .C(n24965), 
         .D(index_i[7]), .Z(n23184)) /* synthesis lut_function=(A (B (D)+!B ((D)+!C))+!A ((D)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n380_bdd_2_lut_4_lut.init = 16'hff13;
    L6MUX21 i18107 (.D0(n20421), .D1(n20422), .SD(index_i[6]), .Z(n20437));
    LUT4 mux_193_Mux_0_i123_3_lut_3_lut_rep_684 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n27524)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i123_3_lut_3_lut_rep_684.init = 16'h6c6c;
    LUT4 mux_192_Mux_6_i420_3_lut_4_lut_4_lut_3_lut_rep_658 (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[2]), .Z(n27498)) /* synthesis lut_function=(A (B+!(C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_6_i420_3_lut_4_lut_4_lut_3_lut_rep_658.init = 16'hdbdb;
    LUT4 mux_193_Mux_0_i124_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n124_adj_2376)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A !(B (D)+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i124_3_lut_4_lut_4_lut.init = 16'h6c99;
    L6MUX21 i18108 (.D0(n20423), .D1(n20424), .SD(index_i[6]), .Z(n20438));
    LUT4 mux_192_Mux_6_i955_3_lut_4_lut (.A(n24969), .B(index_i[3]), .C(index_i[4]), 
         .D(n24815), .Z(n955_adj_2377)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_6_i955_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_192_Mux_8_i860_3_lut_4_lut (.A(n24969), .B(index_i[3]), .C(index_i[4]), 
         .D(n24942), .Z(n860_adj_2378)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_8_i860_3_lut_4_lut.init = 16'h08f8;
    L6MUX21 i18109 (.D0(n20425), .D1(n20426), .SD(index_i[6]), .Z(n20439));
    LUT4 mux_193_Mux_0_i396_3_lut_4_lut_4_lut_3_lut_rep_685 (.A(index_q[0]), 
         .B(index_q[1]), .C(index_q[2]), .Z(n27525)) /* synthesis lut_function=(A ((C)+!B)+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i396_3_lut_4_lut_4_lut_3_lut_rep_685.init = 16'hb6b6;
    LUT4 mux_193_Mux_1_i301_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n301)) /* synthesis lut_function=(A (B (C+(D))+!B !(D))+!A !(B (C+(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_1_i301_3_lut_4_lut_4_lut.init = 16'h99b6;
    PFUMX i18111 (.BLUT(n20429), .ALUT(n20430), .C0(index_i[6]), .Z(n20441));
    PFUMX i18676 (.BLUT(n460_adj_2329), .ALUT(n475_adj_2379), .C0(index_i[4]), 
          .Z(n21006));
    LUT4 n420_bdd_3_lut_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n24010)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A !(B (C+(D))+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n420_bdd_3_lut_3_lut_4_lut_4_lut.init = 16'h44db;
    LUT4 i19375_3_lut (.A(n21702), .B(n21703), .C(index_q[7]), .Z(n21705)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19375_3_lut.init = 16'hcaca;
    LUT4 i19374_3_lut (.A(n21700), .B(n21701), .C(index_q[7]), .Z(n21704)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19374_3_lut.init = 16'hcaca;
    LUT4 i18385_3_lut_4_lut (.A(n24969), .B(index_i[3]), .C(index_i[4]), 
         .D(n364_adj_2380), .Z(n20715)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18385_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_192_Mux_3_i252_3_lut_4_lut (.A(n24969), .B(index_i[3]), .C(index_i[4]), 
         .D(n14998), .Z(n252_adj_2381)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_3_i252_3_lut_4_lut.init = 16'h08f8;
    LUT4 i11327_3_lut_3_lut_3_lut_rep_659 (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .Z(n27499)) /* synthesis lut_function=(!(A+!(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11327_3_lut_3_lut_3_lut_rep_659.init = 16'h4545;
    L6MUX21 i18112 (.D0(n20431), .D1(n20432), .SD(index_i[6]), .Z(n20442));
    L6MUX21 i18113 (.D0(n20433), .D1(n20434), .SD(index_i[6]), .Z(n20443));
    LUT4 mux_193_Mux_2_i284_3_lut_4_lut_4_lut_3_lut_rep_686 (.A(index_q[0]), 
         .B(index_q[1]), .C(index_q[2]), .Z(n27526)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_2_i284_3_lut_4_lut_4_lut_3_lut_rep_686.init = 16'h4d4d;
    PFUMX i18114 (.BLUT(n20435), .ALUT(n20436), .C0(index_i[6]), .Z(n20444));
    LUT4 mux_192_Mux_10_i62_3_lut_3_lut_4_lut (.A(n24969), .B(index_i[3]), 
         .C(n24942), .D(index_i[4]), .Z(n62_adj_2382)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_10_i62_3_lut_3_lut_4_lut.init = 16'hf077;
    LUT4 i11485_2_lut_rep_252_3_lut_4_lut (.A(n24969), .B(index_i[3]), .C(index_i[5]), 
         .D(index_i[4]), .Z(n24812)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11485_2_lut_rep_252_3_lut_4_lut.init = 16'hf080;
    LUT4 mux_193_Mux_3_i653_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n653_adj_2383)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A !(B (D)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_3_i653_3_lut_4_lut_4_lut.init = 16'h4d99;
    LUT4 mux_192_Mux_12_i1023_4_lut (.A(n20587), .B(n766_adj_2384), .C(index_i[9]), 
         .D(index_i[8]), .Z(quarter_wave_sample_register_i_15__N_2126[12])) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_12_i1023_4_lut.init = 16'hfaca;
    LUT4 mux_192_Mux_12_i766_4_lut (.A(n24812), .B(n14928), .C(index_i[7]), 
         .D(index_i[6]), .Z(n766_adj_2384)) /* synthesis lut_function=(A (B (C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_12_i766_4_lut.init = 16'hc0c5;
    LUT4 mux_192_Mux_3_i189_3_lut_3_lut_4_lut (.A(n24969), .B(index_i[3]), 
         .C(index_i[4]), .D(n24922), .Z(n189_adj_2385)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_3_i189_3_lut_3_lut_4_lut.init = 16'h08f8;
    LUT4 i19211_3_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[0]), 
         .D(index_i[3]), .Z(n21541)) /* synthesis lut_function=(!(A ((D)+!B)+!A !(B (D)+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19211_3_lut_4_lut_4_lut.init = 16'h4588;
    PFUMX i18677 (.BLUT(n491_adj_2386), .ALUT(n11355), .C0(index_i[4]), 
          .Z(n21007));
    LUT4 mux_192_Mux_10_i317_3_lut_3_lut_4_lut (.A(n24970), .B(index_i[3]), 
         .C(n24922), .D(index_i[4]), .Z(n317_adj_2387)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_10_i317_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 n124_bdd_3_lut_22517_4_lut (.A(n24970), .B(index_i[3]), .C(index_i[4]), 
         .D(n93_adj_2388), .Z(n23064)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n124_bdd_3_lut_22517_4_lut.init = 16'hfe0e;
    LUT4 n62_bdd_3_lut_21524_4_lut (.A(n24970), .B(index_i[3]), .C(index_i[4]), 
         .D(n890_adj_2389), .Z(n22891)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n62_bdd_3_lut_21524_4_lut.init = 16'hfe0e;
    LUT4 i12236_3_lut_4_lut (.A(n24970), .B(index_i[3]), .C(n25128), .D(index_i[6]), 
         .Z(n14928)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i12236_3_lut_4_lut.init = 16'hffe0;
    LUT4 i11246_3_lut_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n13921)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (D))+!A (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11246_3_lut_3_lut_3_lut_4_lut.init = 16'h00f7;
    LUT4 i18383_3_lut_3_lut_4_lut (.A(n24970), .B(index_i[3]), .C(n316), 
         .D(index_i[4]), .Z(n20713)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18383_3_lut_3_lut_4_lut.init = 16'hf011;
    PFUMX i17924 (.BLUT(n221), .ALUT(n252_adj_2326), .C0(index_q[5]), 
          .Z(n20254));
    PFUMX i18133 (.BLUT(n732_adj_2390), .ALUT(n763_adj_2391), .C0(index_q[5]), 
          .Z(n20463));
    LUT4 n953_bdd_3_lut (.A(n27519), .B(n85), .C(index_i[3]), .Z(n23789)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n953_bdd_3_lut.init = 16'hcaca;
    LUT4 i18615_3_lut_3_lut_4_lut (.A(n24970), .B(index_i[3]), .C(n93_adj_2388), 
         .D(index_i[4]), .Z(n20945)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18615_3_lut_3_lut_4_lut.init = 16'h11f0;
    L6MUX21 i18135 (.D0(n21459), .D1(n891_adj_2392), .SD(index_q[5]), 
            .Z(n20465));
    L6MUX21 i18138 (.D0(n20452), .D1(n20453), .SD(index_q[6]), .Z(n20468));
    PFUMX i18154 (.BLUT(n94), .ALUT(n125_adj_2393), .C0(index_i[5]), .Z(n20484));
    LUT4 i20945_3_lut_4_lut (.A(n25005), .B(n24955), .C(index_q[8]), .D(n766), 
         .Z(n20810)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20945_3_lut_4_lut.init = 16'hefe0;
    LUT4 i19203_3_lut (.A(n27497), .B(n25084), .C(index_i[3]), .Z(n21533)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19203_3_lut.init = 16'hcaca;
    LUT4 n543_bdd_4_lut_22367_4_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n23988)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B (C)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n543_bdd_4_lut_22367_4_lut_4_lut.init = 16'h3d2d;
    LUT4 i6359_2_lut (.A(phase_q[0]), .B(phase_i[10]), .Z(index_i_9__N_2106[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i6359_2_lut.init = 16'h6666;
    LUT4 i20966_2_lut (.A(phase_q[0]), .B(phase_i[10]), .Z(index_q_9__N_2116[0])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i20966_2_lut.init = 16'h9999;
    PFUMX i18155 (.BLUT(n158), .ALUT(n189_adj_2385), .C0(index_i[5]), 
          .Z(n20485));
    LUT4 i17913_3_lut (.A(n20241), .B(n20242), .C(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2126[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17913_3_lut.init = 16'hcaca;
    LUT4 i17912_4_lut (.A(n20639), .B(n893), .C(index_i[8]), .D(index_i[7]), 
         .Z(n20242)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;
    defparam i17912_4_lut.init = 16'hfaca;
    LUT4 mux_192_Mux_10_i893_4_lut (.A(n25114), .B(n24881), .C(index_i[6]), 
         .D(index_i[5]), .Z(n893)) /* synthesis lut_function=(A (B (C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_10_i893_4_lut.init = 16'hc0c5;
    LUT4 n1018_bdd_4_lut_4_lut_4_lut (.A(index_i[0]), .B(n25122), .C(index_i[4]), 
         .D(index_i[3]), .Z(n23385)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (D))+!A (B (C (D)+!C !(D))+!B (D)))) */ ;
    defparam n1018_bdd_4_lut_4_lut_4_lut.init = 16'h0c73;
    PFUMX i18156 (.BLUT(n221_adj_2394), .ALUT(n252_adj_2381), .C0(index_i[5]), 
          .Z(n20486));
    LUT4 mux_192_Mux_11_i766_3_lut (.A(n638), .B(n14928), .C(index_i[7]), 
         .Z(n766_adj_2395)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_11_i766_3_lut.init = 16'h3a3a;
    PFUMX i18157 (.BLUT(n286), .ALUT(n21468), .C0(index_i[5]), .Z(n20487));
    LUT4 i18827_3_lut (.A(n21155), .B(n21156), .C(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2126[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18827_3_lut.init = 16'hcaca;
    LUT4 i18826_3_lut (.A(n21153), .B(n21154), .C(index_i[8]), .Z(n21156)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18826_3_lut.init = 16'hcaca;
    LUT4 i18824_3_lut (.A(n21149), .B(n21150), .C(index_i[7]), .Z(n21154)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18824_3_lut.init = 16'hcaca;
    PFUMX mux_193_Mux_3_i763 (.BLUT(n747_adj_2396), .ALUT(n762_adj_2308), 
          .C0(index_q[4]), .Z(n763_adj_2397)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 mux_193_Mux_4_i1002_3_lut_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n1002_adj_2398)) /* synthesis lut_function=(A (B (C (D))+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_4_i1002_3_lut_3_lut_3_lut_4_lut.init = 16'hf007;
    LUT4 n890_bdd_3_lut_4_lut_4_lut (.A(n24980), .B(index_q[3]), .C(n24957), 
         .D(index_q[4]), .Z(n22874)) /* synthesis lut_function=(A (B (C+!(D))+!B !((D)+!C))+!A (B (C+!(D))+!B (C+(D)))) */ ;
    defparam n890_bdd_3_lut_4_lut_4_lut.init = 16'hd1fc;
    PFUMX i18728 (.BLUT(n142_adj_2399), .ALUT(n157_adj_2400), .C0(index_q[4]), 
          .Z(n21058));
    LUT4 i20954_3_lut (.A(n766_adj_2395), .B(n19504), .C(index_i[8]), 
         .Z(n20577)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20954_3_lut.init = 16'hcaca;
    PFUMX i18729 (.BLUT(n173_adj_2401), .ALUT(n188_adj_2402), .C0(index_q[4]), 
          .Z(n21059));
    PFUMX i18734 (.BLUT(n333_adj_2403), .ALUT(n348_adj_2404), .C0(index_q[4]), 
          .Z(n21064));
    PFUMX i18158 (.BLUT(n349), .ALUT(n21471), .C0(index_i[5]), .Z(n20488));
    PFUMX i18159 (.BLUT(n413_adj_2405), .ALUT(n444), .C0(index_i[5]), 
          .Z(n20489));
    PFUMX i18160 (.BLUT(n476_adj_2406), .ALUT(n507), .C0(index_i[5]), 
          .Z(n20490));
    LUT4 i19196_3_lut (.A(n25083), .B(n27498), .C(index_i[3]), .Z(n21526)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19196_3_lut.init = 16'hcaca;
    PFUMX i18161 (.BLUT(n21474), .ALUT(n573), .C0(index_i[5]), .Z(n20491));
    LUT4 mux_192_Mux_10_i413_3_lut_4_lut (.A(n24985), .B(index_i[3]), .C(index_i[4]), 
         .D(n24922), .Z(n413_adj_2407)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_10_i413_3_lut_4_lut.init = 16'hf101;
    LUT4 mux_192_Mux_3_i828_3_lut_3_lut_4_lut (.A(n24985), .B(index_i[3]), 
         .C(n157_adj_2408), .D(index_i[4]), .Z(n828_adj_2409)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_3_i828_3_lut_3_lut_4_lut.init = 16'hf011;
    PFUMX i18735 (.BLUT(n364_adj_2316), .ALUT(n379_adj_2323), .C0(index_q[4]), 
          .Z(n21065));
    PFUMX i18162 (.BLUT(n12114), .ALUT(n21477), .C0(index_i[5]), .Z(n20492));
    LUT4 mux_192_Mux_10_i252_3_lut_4_lut_4_lut (.A(n24985), .B(index_i[3]), 
         .C(index_i[4]), .D(n24947), .Z(n252)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B (C (D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_10_i252_3_lut_4_lut_4_lut.init = 16'h3efe;
    LUT4 i18513_3_lut_4_lut_4_lut (.A(n24957), .B(index_q[4]), .C(index_q[3]), 
         .D(n24959), .Z(n20843)) /* synthesis lut_function=(A (B (C)+!B !(C+!(D)))+!A (B (C)+!B (C+(D)))) */ ;
    defparam i18513_3_lut_4_lut_4_lut.init = 16'hd3d0;
    LUT4 n557_bdd_3_lut_4_lut (.A(n24985), .B(index_i[3]), .C(index_i[5]), 
         .D(n23629), .Z(n24802)) /* synthesis lut_function=(!(A (C+!(D))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n557_bdd_3_lut_4_lut.init = 16'h1f10;
    LUT4 i21857_then_4_lut (.A(index_i[0]), .B(index_i[4]), .C(index_i[1]), 
         .D(index_i[3]), .Z(n25215)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam i21857_then_4_lut.init = 16'h3c69;
    PFUMX i18736 (.BLUT(n397_adj_2410), .ALUT(n412_adj_2334), .C0(index_q[4]), 
          .Z(n21066));
    LUT4 mux_192_Mux_3_i142_3_lut_3_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .Z(n142_adj_2411)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_3_i142_3_lut_3_lut_3_lut.init = 16'h3838;
    LUT4 i21857_else_4_lut (.A(index_i[0]), .B(index_i[4]), .C(index_i[1]), 
         .D(index_i[3]), .Z(n25214)) /* synthesis lut_function=(!(A (B (C)+!B !(C (D)+!C !(D)))+!A (B ((D)+!C)+!B !((D)+!C)))) */ ;
    defparam i21857_else_4_lut.init = 16'h394b;
    PFUMX i18163 (.BLUT(n669), .ALUT(n700), .C0(index_i[5]), .Z(n20493));
    LUT4 i20465_3_lut (.A(n21523), .B(n21524), .C(index_i[4]), .Z(n21525)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20465_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_12_i1023_4_lut (.A(n20584), .B(n766_adj_2412), .C(index_q[9]), 
         .D(index_q[8]), .Z(quarter_wave_sample_register_q_15__N_2141[12])) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_12_i1023_4_lut.init = 16'hfaca;
    LUT4 i18389_3_lut_3_lut_4_lut (.A(n24985), .B(index_i[3]), .C(n412), 
         .D(index_i[4]), .Z(n20719)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18389_3_lut_3_lut_4_lut.init = 16'hf011;
    PFUMX i18737 (.BLUT(n428_adj_2301), .ALUT(n443_adj_2413), .C0(index_q[4]), 
          .Z(n21067));
    L6MUX21 i18164 (.D0(n21480), .D1(n763_adj_2292), .SD(index_i[5]), 
            .Z(n20494));
    LUT4 mux_193_Mux_12_i766_4_lut (.A(n24811), .B(n765), .C(index_q[7]), 
         .D(index_q[6]), .Z(n766_adj_2412)) /* synthesis lut_function=(A (B (C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_12_i766_4_lut.init = 16'hc0c5;
    LUT4 n7_bdd_3_lut_22231 (.A(n25202), .B(n25174), .C(index_q[3]), .Z(n23838)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n7_bdd_3_lut_22231.init = 16'hacac;
    PFUMX i18165 (.BLUT(n797), .ALUT(n828_adj_2409), .C0(index_i[5]), 
          .Z(n20495));
    PFUMX i18738 (.BLUT(n460), .ALUT(n475_adj_2414), .C0(index_q[4]), 
          .Z(n21068));
    LUT4 i12367_1_lut_2_lut_3_lut_4_lut (.A(n24985), .B(index_i[3]), .C(index_i[5]), 
         .D(index_i[4]), .Z(n381)) /* synthesis lut_function=(!(A (C+(D))+!A (B (C+(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i12367_1_lut_2_lut_3_lut_4_lut.init = 16'h010f;
    LUT4 mux_192_Mux_1_i317_3_lut (.A(n301_adj_2415), .B(n908_adj_2289), 
         .C(index_i[4]), .Z(n317_adj_2416)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_1_i317_3_lut.init = 16'hcaca;
    PFUMX i18166 (.BLUT(n860_adj_2417), .ALUT(n891_adj_2418), .C0(index_i[5]), 
          .Z(n20496));
    LUT4 i18518_3_lut (.A(n20846), .B(n20847), .C(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_2141[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18518_3_lut.init = 16'hcaca;
    PFUMX i18167 (.BLUT(n924_adj_2419), .ALUT(n21483), .C0(index_i[5]), 
          .Z(n20497));
    LUT4 i18517_4_lut (.A(n20636), .B(n893_adj_2420), .C(index_q[8]), 
         .D(index_q[7]), .Z(n20847)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;
    defparam i18517_4_lut.init = 16'hfaca;
    LUT4 i18951_3_lut (.A(n21279), .B(n21280), .C(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_2141[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18951_3_lut.init = 16'hcaca;
    LUT4 i18950_3_lut (.A(n21277), .B(n21278), .C(index_q[8]), .Z(n21280)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18950_3_lut.init = 16'hcaca;
    LUT4 i18948_3_lut (.A(n21273), .B(n21274), .C(index_q[7]), .Z(n21278)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18948_3_lut.init = 16'hcaca;
    PFUMX i18739 (.BLUT(n491_adj_2421), .ALUT(n11358), .C0(index_q[4]), 
          .Z(n21069));
    LUT4 i20968_2_lut (.A(phase_i[9]), .B(phase_i[10]), .Z(index_q_9__N_2116[9])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i20968_2_lut.init = 16'h9999;
    LUT4 i20970_2_lut (.A(phase_i[8]), .B(phase_i[10]), .Z(index_q_9__N_2116[8])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i20970_2_lut.init = 16'h9999;
    PFUMX i18168 (.BLUT(n21486), .ALUT(n1018), .C0(index_i[5]), .Z(n20498));
    LUT4 n269_bdd_3_lut_22254 (.A(n25164), .B(n27503), .C(index_i[3]), 
         .Z(n23859)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n269_bdd_3_lut_22254.init = 16'hcaca;
    PFUMX i18186 (.BLUT(n158_adj_2422), .ALUT(n189_adj_2423), .C0(index_i[5]), 
          .Z(n20516));
    LUT4 i20972_2_lut (.A(phase_i[7]), .B(phase_i[10]), .Z(index_q_9__N_2116[7])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i20972_2_lut.init = 16'h9999;
    PFUMX i18757 (.BLUT(n21085), .ALUT(n21086), .C0(index_q[4]), .Z(n21087));
    LUT4 i20974_2_lut (.A(phase_i[6]), .B(phase_i[10]), .Z(index_q_9__N_2116[6])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i20974_2_lut.init = 16'h9999;
    LUT4 i20976_2_lut (.A(phase_i[5]), .B(phase_i[10]), .Z(index_q_9__N_2116[5])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i20976_2_lut.init = 16'h9999;
    LUT4 i20978_2_lut (.A(phase_i[4]), .B(phase_i[10]), .Z(index_q_9__N_2116[4])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i20978_2_lut.init = 16'h9999;
    PFUMX i18187 (.BLUT(n221_adj_2424), .ALUT(n21492), .C0(index_i[5]), 
          .Z(n20517));
    LUT4 i20980_2_lut (.A(phase_i[3]), .B(phase_i[10]), .Z(index_q_9__N_2116[3])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i20980_2_lut.init = 16'h9999;
    LUT4 i20982_2_lut (.A(phase_i[2]), .B(phase_i[10]), .Z(index_q_9__N_2116[2])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i20982_2_lut.init = 16'h9999;
    LUT4 i18119_3_lut (.A(n20445), .B(n20446), .C(index_i[8]), .Z(n20449)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18119_3_lut.init = 16'hcaca;
    PFUMX i18188 (.BLUT(n286_adj_2425), .ALUT(n317_adj_2426), .C0(index_i[5]), 
          .Z(n20518));
    PFUMX i18189 (.BLUT(n349_adj_2427), .ALUT(n21495), .C0(index_i[5]), 
          .Z(n20519));
    LUT4 i20984_2_lut (.A(phase_i[1]), .B(phase_i[10]), .Z(index_q_9__N_2116[1])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i20984_2_lut.init = 16'h9999;
    PFUMX i18190 (.BLUT(n413_adj_2428), .ALUT(n21498), .C0(index_i[5]), 
          .Z(n20520));
    PFUMX i18191 (.BLUT(n21501), .ALUT(n507_adj_2429), .C0(index_i[5]), 
          .Z(n20521));
    LUT4 i6380_2_lut (.A(phase_i[9]), .B(phase_i[10]), .Z(index_i_9__N_2106[9])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i6380_2_lut.init = 16'h6666;
    LUT4 i6381_2_lut (.A(phase_i[8]), .B(phase_i[10]), .Z(index_i_9__N_2106[8])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i6381_2_lut.init = 16'h6666;
    PFUMX i18192 (.BLUT(n21504), .ALUT(n573_adj_2430), .C0(index_i[5]), 
          .Z(n20522));
    PFUMX i18193 (.BLUT(n605_adj_2431), .ALUT(n21507), .C0(index_i[5]), 
          .Z(n20523));
    PFUMX i18194 (.BLUT(n669_adj_2432), .ALUT(n700_adj_2433), .C0(index_i[5]), 
          .Z(n20524));
    LUT4 i6382_2_lut (.A(phase_i[7]), .B(phase_i[10]), .Z(index_i_9__N_2106[7])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i6382_2_lut.init = 16'h6666;
    LUT4 i6383_2_lut (.A(phase_i[6]), .B(phase_i[10]), .Z(index_i_9__N_2106[6])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i6383_2_lut.init = 16'h6666;
    LUT4 i6384_2_lut (.A(phase_i[5]), .B(phase_i[10]), .Z(index_i_9__N_2106[5])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i6384_2_lut.init = 16'h6666;
    PFUMX i18195 (.BLUT(n732_adj_2434), .ALUT(n763_adj_2435), .C0(index_i[5]), 
          .Z(n20525));
    LUT4 i6385_2_lut (.A(phase_i[4]), .B(phase_i[10]), .Z(index_i_9__N_2106[4])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i6385_2_lut.init = 16'h6666;
    LUT4 i6386_2_lut (.A(phase_i[3]), .B(phase_i[10]), .Z(index_i_9__N_2106[3])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i6386_2_lut.init = 16'h6666;
    LUT4 i19184_3_lut (.A(n723), .B(n25065), .C(index_i[3]), .Z(n21514)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19184_3_lut.init = 16'hcaca;
    PFUMX i18769 (.BLUT(n21097), .ALUT(n21098), .C0(index_q[4]), .Z(n21099));
    L6MUX21 i18197 (.D0(n860), .D1(n891_adj_2281), .SD(index_i[5]), .Z(n20527));
    LUT4 i18089_3_lut (.A(n20416), .B(n20417), .C(index_q[8]), .Z(n20419)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18089_3_lut.init = 16'hcaca;
    LUT4 i18088_3_lut (.A(n20414), .B(n20415), .C(index_q[8]), .Z(n20418)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18088_3_lut.init = 16'hcaca;
    LUT4 i6387_2_lut (.A(phase_i[2]), .B(phase_i[10]), .Z(index_i_9__N_2106[2])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i6387_2_lut.init = 16'h6666;
    LUT4 i6388_2_lut (.A(phase_i[1]), .B(phase_i[10]), .Z(index_i_9__N_2106[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i6388_2_lut.init = 16'h6666;
    LUT4 mux_398_i9_3_lut (.A(\quarter_wave_sample_register_q[15] ), .B(o_val_pipeline_q_0__15__N_2189[15]), 
         .C(phase_negation_q[1]), .Z(n1807[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(80[29:60])
    defparam mux_398_i9_3_lut.init = 16'hcaca;
    PFUMX i18772 (.BLUT(n21100), .ALUT(n21101), .C0(index_q[4]), .Z(n21102));
    LUT4 mux_398_i8_3_lut (.A(quarter_wave_sample_register_q[14]), .B(o_val_pipeline_q_0__15__N_2189[14]), 
         .C(phase_negation_q[1]), .Z(n1807[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(80[29:60])
    defparam mux_398_i8_3_lut.init = 16'hcaca;
    PFUMX i9437 (.BLUT(n12147), .ALUT(n12148), .C0(n25010), .Z(n12003));
    LUT4 mux_398_i7_3_lut (.A(quarter_wave_sample_register_q[13]), .B(o_val_pipeline_q_0__15__N_2189[13]), 
         .C(phase_negation_q[1]), .Z(n1807[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(80[29:60])
    defparam mux_398_i7_3_lut.init = 16'hcaca;
    LUT4 mux_398_i6_3_lut (.A(quarter_wave_sample_register_q[12]), .B(o_val_pipeline_q_0__15__N_2189[12]), 
         .C(phase_negation_q[1]), .Z(n1807[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(80[29:60])
    defparam mux_398_i6_3_lut.init = 16'hcaca;
    LUT4 mux_398_i5_3_lut (.A(quarter_wave_sample_register_q[11]), .B(o_val_pipeline_q_0__15__N_2189[11]), 
         .C(phase_negation_q[1]), .Z(n1807[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(80[29:60])
    defparam mux_398_i5_3_lut.init = 16'hcaca;
    PFUMX i18775 (.BLUT(n21103), .ALUT(n21104), .C0(index_q[4]), .Z(n21105));
    LUT4 mux_398_i4_3_lut (.A(quarter_wave_sample_register_q[10]), .B(o_val_pipeline_q_0__15__N_2189[10]), 
         .C(phase_negation_q[1]), .Z(n1807[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(80[29:60])
    defparam mux_398_i4_3_lut.init = 16'hcaca;
    PFUMX i9477 (.BLUT(n12145), .ALUT(n12146), .C0(n25032), .Z(n12043));
    PFUMX i18778 (.BLUT(n21106), .ALUT(n21107), .C0(index_q[4]), .Z(n21108));
    LUT4 mux_398_i3_3_lut (.A(quarter_wave_sample_register_q[9]), .B(o_val_pipeline_q_0__15__N_2189[9]), 
         .C(phase_negation_q[1]), .Z(n1807[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(80[29:60])
    defparam mux_398_i3_3_lut.init = 16'hcaca;
    LUT4 mux_398_i2_3_lut (.A(quarter_wave_sample_register_q[8]), .B(o_val_pipeline_q_0__15__N_2189[8]), 
         .C(phase_negation_q[1]), .Z(n1807[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(80[29:60])
    defparam mux_398_i2_3_lut.init = 16'hcaca;
    LUT4 mux_398_i1_3_lut (.A(quarter_wave_sample_register_q[7]), .B(o_val_pipeline_q_0__15__N_2189[7]), 
         .C(phase_negation_q[1]), .Z(n1807[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(80[29:60])
    defparam mux_398_i1_3_lut.init = 16'hcaca;
    PFUMX i18216 (.BLUT(n94_adj_2436), .ALUT(n21513), .C0(index_i[5]), 
          .Z(n20546));
    L6MUX21 i18217 (.D0(n21516), .D1(n21519), .SD(index_i[5]), .Z(n20547));
    LUT4 i20472_3_lut (.A(n25282), .B(n21512), .C(index_i[4]), .Z(n21513)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20472_3_lut.init = 16'hcaca;
    LUT4 i18057_3_lut (.A(n20383), .B(n20384), .C(index_i[8]), .Z(n20387)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18057_3_lut.init = 16'hcaca;
    LUT4 i18982_3_lut (.A(n21309), .B(n21310), .C(index_q[8]), .Z(n21312)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18982_3_lut.init = 16'hcaca;
    LUT4 i18981_3_lut (.A(n21307), .B(n21308), .C(index_q[8]), .Z(n21311)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18981_3_lut.init = 16'hcaca;
    PFUMX i18219 (.BLUT(n21522), .ALUT(n317_adj_2416), .C0(index_i[5]), 
          .Z(n20549));
    PFUMX i18220 (.BLUT(n349_adj_2437), .ALUT(n21525), .C0(index_i[5]), 
          .Z(n20550));
    L6MUX21 i18221 (.D0(n21528), .D1(n21531), .SD(index_i[5]), .Z(n20551));
    LUT4 i18027_3_lut (.A(n20354), .B(n20355), .C(index_q[8]), .Z(n20357)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18027_3_lut.init = 16'hcaca;
    L6MUX21 i18222 (.D0(n21534), .D1(n21537), .SD(index_i[5]), .Z(n20552));
    PFUMX i18784 (.BLUT(n21112), .ALUT(n21113), .C0(index_q[4]), .Z(n21114));
    L6MUX21 i18224 (.D0(n21543), .D1(n636_adj_2277), .SD(index_i[5]), 
            .Z(n20554));
    PFUMX i18225 (.BLUT(n21546), .ALUT(n700_adj_2438), .C0(index_i[5]), 
          .Z(n20555));
    LUT4 i18026_3_lut (.A(n20352), .B(n20353), .C(index_q[8]), .Z(n20356)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18026_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_8_i236_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n236)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)+!C !(D)))+!A (B (C+!(D))+!B ((D)+!C))) */ ;
    defparam mux_192_Mux_8_i236_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hf1cf;
    L6MUX21 i18227 (.D0(n21549), .D1(n21552), .SD(index_i[5]), .Z(n20557));
    LUT4 mux_192_Mux_6_i860_3_lut_3_lut (.A(n24838), .B(index_i[4]), .C(n844_adj_2439), 
         .Z(n860_adj_2440)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam mux_192_Mux_6_i860_3_lut_3_lut.init = 16'h7474;
    LUT4 i18572_3_lut_3_lut (.A(n24838), .B(index_i[4]), .C(n46), .Z(n20902)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam i18572_3_lut_3_lut.init = 16'h7474;
    LUT4 i18850_3_lut (.A(n21177), .B(n21178), .C(index_i[8]), .Z(n21180)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18850_3_lut.init = 16'hcaca;
    LUT4 i18849_3_lut (.A(n21175), .B(n21176), .C(index_i[8]), .Z(n21179)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18849_3_lut.init = 16'hcaca;
    LUT4 i19175_3_lut (.A(n498), .B(n25051), .C(index_i[3]), .Z(n21505)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19175_3_lut.init = 16'hcaca;
    LUT4 i17949_3_lut (.A(n20275), .B(n20276), .C(index_q[8]), .Z(n20279)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17949_3_lut.init = 16'hcaca;
    LUT4 i20484_3_lut (.A(n21505), .B(n21506), .C(index_i[4]), .Z(n21507)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20484_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_1_i747_4_lut_else_4_lut (.A(index_i[0]), .B(index_i[4]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n25243)) /* synthesis lut_function=(!(A (B (C (D))+!B !(D))+!A ((C (D))+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_1_i747_4_lut_else_4_lut.init = 16'h2ecc;
    LUT4 i17918_3_lut (.A(n20244), .B(n20245), .C(index_i[8]), .Z(n20248)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17918_3_lut.init = 16'hcaca;
    LUT4 n483_bdd_3_lut_22309 (.A(n25052), .B(n25082), .C(index_i[3]), 
         .Z(n23916)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n483_bdd_3_lut_22309.init = 16'hcaca;
    LUT4 quarter_wave_sample_register_i_15__I_0_3_lut (.A(\quarter_wave_sample_register_q[15] ), 
         .B(o_val_pipeline_i_0__15__N_2157[15]), .C(phase_negation_i[1]), 
         .Z(o_val_pipeline_i_0__15__N_2156)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[14] 77[8])
    defparam quarter_wave_sample_register_i_15__I_0_3_lut.init = 16'hcaca;
    PFUMX i18229 (.BLUT(n924_adj_2441), .ALUT(n21558), .C0(index_i[5]), 
          .Z(n20559));
    PFUMX i17969 (.BLUT(n158_adj_2442), .ALUT(n189_adj_2443), .C0(index_q[5]), 
          .Z(n20299));
    LUT4 index_q_0__bdd_4_lut_23028 (.A(index_q[0]), .B(index_q[3]), .C(index_q[1]), 
         .D(index_q[2]), .Z(n25246)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C))+!A (B (C (D)+!C !(D))+!B !(C+!(D))))) */ ;
    defparam index_q_0__bdd_4_lut_23028.init = 16'h16d3;
    PFUMX i18230 (.BLUT(n987), .ALUT(n21561), .C0(index_i[5]), .Z(n20560));
    LUT4 i19170_3_lut (.A(n498), .B(n27496), .C(index_i[3]), .Z(n21500)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19170_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut (.A(o_phase[11]), .B(o_phase[10]), .Z(phase_q_11__N_2232[11])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i1_2_lut.init = 16'h9999;
    LUT4 i20490_3_lut (.A(n21496), .B(n21497), .C(index_i[4]), .Z(n21498)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20490_3_lut.init = 16'hcaca;
    LUT4 i18479_3_lut (.A(n22818), .B(n20602), .C(index_q[8]), .Z(n20809)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18479_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_8_i542_3_lut_4_lut (.A(n25116), .B(index_i[3]), .C(index_i[4]), 
         .D(n526_adj_2444), .Z(n542)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_8_i542_3_lut_4_lut.init = 16'h6f60;
    LUT4 i19164_3_lut (.A(n27496), .B(n25171), .C(index_i[3]), .Z(n21494)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19164_3_lut.init = 16'hcaca;
    LUT4 i18597_3_lut_4_lut (.A(n25116), .B(index_i[3]), .C(index_i[4]), 
         .D(n635_adj_2445), .Z(n20927)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18597_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_193_Mux_1_i700_3_lut_4_lut (.A(n25025), .B(index_q[3]), .C(index_q[4]), 
         .D(n684_adj_2336), .Z(n700_adj_2446)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_1_i700_3_lut_4_lut.init = 16'hefe0;
    LUT4 mux_193_Mux_8_i542_3_lut_4_lut (.A(n25097), .B(index_q[3]), .C(index_q[4]), 
         .D(n526_adj_2274), .Z(n542_adj_2447)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_8_i542_3_lut_4_lut.init = 16'h6f60;
    LUT4 i18511_3_lut_4_lut (.A(n25097), .B(index_q[3]), .C(index_q[4]), 
         .D(n635_adj_2448), .Z(n20841)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18511_3_lut_4_lut.init = 16'hf606;
    PFUMX i18836 (.BLUT(n21164), .ALUT(n21165), .C0(index_i[4]), .Z(n21166));
    PFUMX i15274 (.BLUT(n17535), .ALUT(n17536), .C0(index_i[4]), .Z(n17537));
    LUT4 i20492_3_lut (.A(n21493), .B(n21494), .C(index_i[4]), .Z(n21495)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20492_3_lut.init = 16'hcaca;
    PFUMX i18271 (.BLUT(n445_adj_2339), .ALUT(n508), .C0(index_q[6]), 
          .Z(n20601));
    LUT4 i11376_3_lut_3_lut_rep_663 (.A(index_i[2]), .B(index_i[0]), .C(index_i[1]), 
         .Z(n27503)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11376_3_lut_3_lut_rep_663.init = 16'hd0d0;
    LUT4 i19146_3_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[0]), .C(index_i[1]), 
         .D(index_i[3]), .Z(n21476)) /* synthesis lut_function=(A (B (C)+!B !(C+!(D)))+!A (B (C)+!B !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19146_3_lut_4_lut_4_lut.init = 16'hc3d0;
    LUT4 n851_bdd_3_lut_22228_4_lut (.A(n25172), .B(index_q[2]), .C(index_q[3]), 
         .D(n25176), .Z(n23835)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n851_bdd_3_lut_22228_4_lut.init = 16'hf606;
    LUT4 i3_4_lut (.A(n24812), .B(index_i[6]), .C(index_i[8]), .D(index_i[7]), 
         .Z(n17770)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i3_4_lut.init = 16'hfffe;
    LUT4 mux_193_Mux_3_i668_3_lut_4_lut (.A(n25172), .B(index_q[2]), .C(index_q[3]), 
         .D(n25204), .Z(n668_adj_2449)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_3_i668_3_lut_4_lut.init = 16'h6f60;
    PFUMX mux_193_Mux_5_i732 (.BLUT(n12039), .ALUT(n731_adj_2450), .C0(index_q[4]), 
          .Z(n732_adj_2451)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 index_q_2__bdd_4_lut_23165 (.A(index_q[2]), .B(index_q[1]), .C(index_q[3]), 
         .D(index_q[0]), .Z(n25247)) /* synthesis lut_function=(A (B ((D)+!C))+!A !(B+!(C+!(D)))) */ ;
    defparam index_q_2__bdd_4_lut_23165.init = 16'h9819;
    LUT4 mux_193_Mux_4_i763_3_lut_4_lut (.A(n25172), .B(index_q[2]), .C(index_q[4]), 
         .D(n747_adj_2452), .Z(n763_adj_2453)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_4_i763_3_lut_4_lut.init = 16'h6f60;
    LUT4 i18246_3_lut (.A(n22856), .B(n20645), .C(index_i[8]), .Z(n20576)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18246_3_lut.init = 16'hcaca;
    LUT4 i20495_3_lut (.A(n21490), .B(n21491), .C(index_i[4]), .Z(n21492)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20495_3_lut.init = 16'hcaca;
    LUT4 i18213_3_lut (.A(n20540), .B(n20541), .C(index_i[8]), .Z(n20543)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18213_3_lut.init = 16'hcaca;
    LUT4 i18212_3_lut (.A(n20538), .B(n20539), .C(index_i[8]), .Z(n20542)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18212_3_lut.init = 16'hcaca;
    LUT4 i18182_3_lut (.A(n20509), .B(n20510), .C(index_i[8]), .Z(n20512)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18182_3_lut.init = 16'hcaca;
    LUT4 i18181_3_lut (.A(n20507), .B(n20508), .C(index_i[8]), .Z(n20511)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18181_3_lut.init = 16'hcaca;
    LUT4 i19152_3_lut (.A(n325_adj_2282), .B(n25065), .C(index_i[3]), 
         .Z(n21482)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19152_3_lut.init = 16'hcaca;
    LUT4 i18612_3_lut (.A(n20939), .B(n20940), .C(index_q[8]), .Z(n20942)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18612_3_lut.init = 16'hcaca;
    LUT4 i20501_3_lut (.A(n21481), .B(n21482), .C(index_i[4]), .Z(n21483)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20501_3_lut.init = 16'hcaca;
    LUT4 i18611_3_lut (.A(n20937), .B(n20938), .C(index_q[8]), .Z(n20941)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18611_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_2_i955_then_4_lut (.A(index_i[4]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n25218)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B (C+!(D))+!B !(C (D)))) */ ;
    defparam mux_192_Mux_2_i955_then_4_lut.init = 16'he95d;
    L6MUX21 i19362 (.D0(n21676), .D1(n21677), .SD(index_q[5]), .Z(n21692));
    LUT4 mux_193_Mux_6_i860_3_lut_3_lut (.A(n24840), .B(index_q[4]), .C(n844_adj_2454), 
         .Z(n860_adj_2455)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam mux_193_Mux_6_i860_3_lut_3_lut.init = 16'h7474;
    LUT4 i18486_3_lut_3_lut (.A(n24840), .B(index_q[4]), .C(n46_adj_2456), 
         .Z(n20816)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam i18486_3_lut_3_lut.init = 16'h7474;
    LUT4 mux_193_Mux_1_i924_3_lut (.A(n316_adj_2457), .B(n412_adj_2361), 
         .C(index_q[4]), .Z(n924_adj_2458)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_1_i924_3_lut.init = 16'hcaca;
    L6MUX21 i19363 (.D0(n21678), .D1(n21679), .SD(index_q[5]), .Z(n21693));
    L6MUX21 i19364 (.D0(n21680), .D1(n21681), .SD(index_q[5]), .Z(n21694));
    L6MUX21 i19365 (.D0(n21682), .D1(n21683), .SD(index_q[5]), .Z(n21695));
    LUT4 i19095_3_lut_4_lut_4_lut (.A(n25097), .B(n25176), .C(index_q[3]), 
         .D(index_q[0]), .Z(n21425)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C))) */ ;
    defparam i19095_3_lut_4_lut_4_lut.init = 16'hcfc5;
    LUT4 mux_192_Mux_5_i124_3_lut (.A(n24941), .B(n25171), .C(index_i[3]), 
         .Z(n124_adj_2459)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_5_i124_3_lut.init = 16'hcaca;
    L6MUX21 i19366 (.D0(n21684), .D1(n21685), .SD(index_q[5]), .Z(n21696));
    L6MUX21 i19367 (.D0(n21686), .D1(n21687), .SD(index_q[5]), .Z(n21697));
    LUT4 i19953_3_lut (.A(n21448), .B(n21449), .C(index_q[4]), .Z(n21450)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19953_3_lut.init = 16'hcaca;
    L6MUX21 i19368 (.D0(n21688), .D1(n21689), .SD(index_q[5]), .Z(n21698));
    L6MUX21 i19369 (.D0(n21690), .D1(n21691), .SD(index_q[5]), .Z(n21699));
    PFUMX i18314 (.BLUT(n445), .ALUT(n508_adj_2460), .C0(index_i[6]), 
          .Z(n20644));
    LUT4 i18244_3_lut (.A(n20571), .B(n20572), .C(index_i[8]), .Z(n20574)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18244_3_lut.init = 16'hcaca;
    LUT4 i19956_3_lut (.A(n27528), .B(n21443), .C(index_q[4]), .Z(n21444)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19956_3_lut.init = 16'hcaca;
    LUT4 i18243_3_lut (.A(n20569), .B(n20570), .C(index_i[8]), .Z(n20573)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18243_3_lut.init = 16'hcaca;
    LUT4 i18151_3_lut (.A(n20478), .B(n20479), .C(index_q[8]), .Z(n20481)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18151_3_lut.init = 16'hcaca;
    LUT4 i18150_3_lut (.A(n20476), .B(n20477), .C(index_q[8]), .Z(n20480)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18150_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_1_i349_3_lut (.A(n506_adj_2461), .B(n348_adj_2297), 
         .C(index_q[4]), .Z(n349_adj_2462)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_1_i349_3_lut.init = 16'hcaca;
    LUT4 i19187_3_lut_4_lut_4_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n21517)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))+!A (B (C)+!B ((D)+!C))) */ ;
    defparam i19187_3_lut_4_lut_4_lut_4_lut_4_lut_4_lut.init = 16'hf1e3;
    LUT4 mux_192_Mux_8_i101_3_lut_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n101)) /* synthesis lut_function=(!(A (B (C))+!A (B (C)+!B !(C)))) */ ;
    defparam mux_192_Mux_8_i101_3_lut_3_lut_3_lut.init = 16'h3e3e;
    LUT4 i19962_3_lut (.A(n21424), .B(n21425), .C(index_q[4]), .Z(n21426)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19962_3_lut.init = 16'hcaca;
    LUT4 i11440_2_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n635_adj_2276)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A (B (C+!(D))+!B (C+(D)))) */ ;
    defparam i11440_2_lut_4_lut_4_lut.init = 16'hf1fc;
    LUT4 mux_192_Mux_3_i157_3_lut_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n157_adj_2408)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B !(C+(D))))) */ ;
    defparam mux_192_Mux_3_i157_3_lut_3_lut_3_lut_4_lut.init = 16'h1ff0;
    LUT4 mux_192_Mux_7_i572_3_lut_rep_254_3_lut_3_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n24814)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)+!C !(D)))) */ ;
    defparam mux_192_Mux_7_i572_3_lut_rep_254_3_lut_3_lut_4_lut.init = 16'hfe01;
    LUT4 mux_193_Mux_1_i94_3_lut (.A(index_q[0]), .B(n93_adj_2463), .C(index_q[4]), 
         .Z(n94_adj_2464)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_1_i94_3_lut.init = 16'hcaca;
    LUT4 index_i_5__bdd_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n23625)) /* synthesis lut_function=(A (B (C)+!B (C+(D)))+!A (B (C)+!B !(C (D)+!C !(D)))) */ ;
    defparam index_i_5__bdd_3_lut_4_lut_4_lut_4_lut.init = 16'he3f0;
    LUT4 mux_192_Mux_2_i142_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n142_adj_2465)) /* synthesis lut_function=(!(A (B (D)+!B (C (D)+!C !(D)))+!A (B (D)+!B (C+!(D))))) */ ;
    defparam mux_192_Mux_2_i142_3_lut_4_lut_4_lut_4_lut.init = 16'h03ec;
    LUT4 n23961_bdd_3_lut (.A(n23961), .B(n316_adj_2457), .C(index_q[4]), 
         .Z(n23962)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n23961_bdd_3_lut.init = 16'hcaca;
    LUT4 i11430_3_lut_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n14105)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B !(C+!(D))))) */ ;
    defparam i11430_3_lut_3_lut_3_lut_4_lut.init = 16'h10ff;
    LUT4 i11293_2_lut_rep_327_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n24887)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i11293_2_lut_rep_327_3_lut_4_lut.init = 16'hfef0;
    LUT4 mux_192_Mux_7_i540_3_lut_rep_481_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n25041)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C)+!B !(C))) */ ;
    defparam mux_192_Mux_7_i540_3_lut_rep_481_3_lut.init = 16'he3e3;
    LUT4 n22895_bdd_3_lut (.A(n20287), .B(n20286), .C(index_i[7]), .Z(n26497)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n22895_bdd_3_lut.init = 16'hacac;
    LUT4 n22895_bdd_3_lut_23952 (.A(n22895), .B(n20289), .C(index_i[7]), 
         .Z(n26496)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n22895_bdd_3_lut_23952.init = 16'hcaca;
    LUT4 n25460_bdd_3_lut_23955 (.A(n20284), .B(n20285), .C(index_i[7]), 
         .Z(n26499)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n25460_bdd_3_lut_23955.init = 16'hcaca;
    LUT4 n25460_bdd_3_lut_24162 (.A(n20953), .B(n20960), .C(index_i[6]), 
         .Z(n26500)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n25460_bdd_3_lut_24162.init = 16'hcaca;
    L6MUX21 i21669 (.D0(n23224), .D1(n23222), .SD(index_q[6]), .Z(n23225));
    LUT4 n26500_bdd_3_lut (.A(n26500), .B(n25460), .C(index_i[7]), .Z(n26501)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n26500_bdd_3_lut.init = 16'hcaca;
    LUT4 i19188_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n21518)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C+(D)))+!A (B (C (D)+!C !(D))+!B !(C)))) */ ;
    defparam i19188_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h3ef0;
    PFUMX i21667 (.BLUT(n924_adj_2466), .ALUT(n23223), .C0(index_q[5]), 
          .Z(n23224));
    L6MUX21 i19442 (.D0(n21756), .D1(n21757), .SD(index_i[5]), .Z(n21772));
    L6MUX21 i19443 (.D0(n21758), .D1(n21759), .SD(index_i[5]), .Z(n21773));
    LUT4 i11188_3_lut_4_lut (.A(n24804), .B(index_q[7]), .C(index_q[8]), 
         .D(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_2141[14])) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (D))) */ ;
    defparam i11188_3_lut_4_lut.init = 16'hffe0;
    LUT4 mux_192_Mux_8_i46_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n46)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (B (C)+!B !(C (D)+!C !(D)))) */ ;
    defparam mux_192_Mux_8_i46_3_lut_4_lut_4_lut_4_lut.init = 16'hc1f0;
    LUT4 mux_192_Mux_3_i30_3_lut_4_lut_4_lut_4_lut_3_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n30_adj_2467)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C+!(D)))) */ ;
    defparam mux_192_Mux_3_i30_3_lut_4_lut_4_lut_4_lut_3_lut_4_lut.init = 16'hfe11;
    L6MUX21 i19444 (.D0(n21760), .D1(n21761), .SD(index_i[5]), .Z(n21774));
    LUT4 n543_bdd_4_lut_22364 (.A(index_i[2]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[0]), .Z(n23987)) /* synthesis lut_function=(A (B (C+!(D))+!B !(D))+!A !(B (C+!(D))+!B !(D))) */ ;
    defparam n543_bdd_4_lut_22364.init = 16'h95aa;
    LUT4 i18106_4_lut (.A(n21414), .B(n1002_adj_2468), .C(index_i[5]), 
         .D(index_i[4]), .Z(n20436)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;
    defparam i18106_4_lut.init = 16'hfaca;
    LUT4 mux_192_Mux_2_i716_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n716_adj_2469)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)+!C !(D)))+!A (B (D)+!B !((D)+!C)))) */ ;
    defparam mux_192_Mux_2_i716_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h31cf;
    LUT4 n23989_bdd_3_lut (.A(n23989), .B(n23986), .C(index_i[4]), .Z(n23990)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n23989_bdd_3_lut.init = 16'hcaca;
    PFUMX i18878 (.BLUT(n21206), .ALUT(n21207), .C0(index_q[4]), .Z(n476_adj_2470));
    LUT4 mux_192_Mux_4_i860_3_lut (.A(n506_adj_2471), .B(n23917), .C(index_i[4]), 
         .Z(n860_adj_2472)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_4_i860_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_7_i541_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n541_adj_2473)) /* synthesis lut_function=(A (B (D)+!B (C+!(D)))+!A (B (D)+!B !(D))) */ ;
    defparam mux_192_Mux_7_i541_3_lut_4_lut_4_lut_4_lut.init = 16'hec33;
    LUT4 n85_bdd_3_lut_22370 (.A(n25084), .B(n25051), .C(index_i[3]), 
         .Z(n23993)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n85_bdd_3_lut_22370.init = 16'hcaca;
    LUT4 i19977_3_lut (.A(n21403), .B(n21404), .C(index_i[4]), .Z(n21405)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19977_3_lut.init = 16'hcaca;
    LUT4 n262_bdd_3_lut_22475 (.A(n25088), .B(n25051), .C(index_i[3]), 
         .Z(n23996)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n262_bdd_3_lut_22475.init = 16'hcaca;
    LUT4 mux_192_Mux_8_i29_3_lut_rep_604 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n25164)) /* synthesis lut_function=(!(A (B (C))+!A !(B+(C)))) */ ;
    defparam mux_192_Mux_8_i29_3_lut_rep_604.init = 16'h7e7e;
    LUT4 mux_192_Mux_1_i700_3_lut_4_lut (.A(n25016), .B(index_i[3]), .C(index_i[4]), 
         .D(n684_adj_2340), .Z(n700_adj_2438)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_1_i700_3_lut_4_lut.init = 16'hefe0;
    LUT4 mux_192_Mux_7_i243_3_lut_rep_605 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n25165)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B (C)+!B !(C)))) */ ;
    defparam mux_192_Mux_7_i243_3_lut_rep_605.init = 16'h1c1c;
    LUT4 n498_bdd_3_lut_22392 (.A(n498), .B(n25074), .C(index_i[3]), .Z(n24012)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n498_bdd_3_lut_22392.init = 16'hcaca;
    LUT4 mux_192_Mux_7_i29_3_lut_rep_606 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n25166)) /* synthesis lut_function=(A (B+!(C))+!A !((C)+!B)) */ ;
    defparam mux_192_Mux_7_i29_3_lut_rep_606.init = 16'h8e8e;
    L6MUX21 i19445 (.D0(n21762), .D1(n21763), .SD(index_i[5]), .Z(n21775));
    LUT4 i19979_3_lut (.A(n21400), .B(n21401), .C(index_i[4]), .Z(n21402)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19979_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_7_i7_3_lut_3_lut_4_lut_3_lut_rep_608 (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[2]), .Z(n25168)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B+!(C)))) */ ;
    defparam mux_192_Mux_7_i7_3_lut_3_lut_4_lut_3_lut_rep_608.init = 16'h1818;
    LUT4 mux_192_Mux_6_i645_3_lut_3_lut_4_lut_3_lut_rep_609 (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[2]), .Z(n25169)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B))) */ ;
    defparam mux_192_Mux_6_i645_3_lut_3_lut_4_lut_3_lut_rep_609.init = 16'h1919;
    LUT4 i19191_3_lut_4_lut (.A(index_i[0]), .B(n25116), .C(index_i[3]), 
         .D(n25080), .Z(n21521)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19191_3_lut_4_lut.init = 16'hfb0b;
    LUT4 mux_192_Mux_2_i955_else_4_lut (.A(index_i[4]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n25217)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+(D)))+!A !(B (C+!(D))+!B !(C+!(D))))) */ ;
    defparam mux_192_Mux_2_i955_else_4_lut.init = 16'h49c6;
    LUT4 mux_192_Mux_5_i53_3_lut_4_lut_3_lut_rep_611 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n25171)) /* synthesis lut_function=(A ((C)+!B)+!A (B)) */ ;
    defparam mux_192_Mux_5_i53_3_lut_4_lut_3_lut_rep_611.init = 16'he6e6;
    LUT4 mux_192_Mux_4_i700_3_lut (.A(n684_adj_2474), .B(index_i[1]), .C(index_i[4]), 
         .Z(n700_adj_2475)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_4_i700_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_0_i557_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n557)) /* synthesis lut_function=(A ((D)+!C)+!A !((D)+!B)) */ ;
    defparam mux_192_Mux_0_i557_3_lut_4_lut.init = 16'haa4e;
    LUT4 mux_192_Mux_6_i635_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n635_adj_2476)) /* synthesis lut_function=(A (B (C+(D))+!B !(D))+!A (B)) */ ;
    defparam mux_192_Mux_6_i635_3_lut_4_lut.init = 16'hcce6;
    L6MUX21 i19446 (.D0(n21764), .D1(n21765), .SD(index_i[5]), .Z(n21776));
    LUT4 mux_192_Mux_4_i669_3_lut (.A(n781_adj_2477), .B(n668), .C(index_i[4]), 
         .Z(n669_adj_2478)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_4_i669_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_7_i716_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n716_adj_2479)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C+!(D))+!B (C)))) */ ;
    defparam mux_192_Mux_7_i716_3_lut_3_lut_4_lut.init = 16'h0f81;
    LUT4 n498_bdd_3_lut_22393 (.A(n498), .B(n25065), .C(index_i[3]), .Z(n24015)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n498_bdd_3_lut_22393.init = 16'hcaca;
    L6MUX21 i19447 (.D0(n21766), .D1(n21767), .SD(index_i[5]), .Z(n21777));
    L6MUX21 i19448 (.D0(n21768), .D1(n21769), .SD(index_i[5]), .Z(n21778));
    LUT4 i18918_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21248)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(D))+!A (B))) */ ;
    defparam i18918_3_lut_3_lut_4_lut.init = 16'h3319;
    LUT4 n498_bdd_3_lut_22554 (.A(n25081), .B(n25087), .C(index_i[3]), 
         .Z(n24016)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n498_bdd_3_lut_22554.init = 16'hcaca;
    LUT4 n452_bdd_3_lut_22558 (.A(n27518), .B(n27496), .C(index_i[3]), 
         .Z(n24019)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n452_bdd_3_lut_22558.init = 16'hcaca;
    LUT4 mux_192_Mux_4_i542_3_lut (.A(n30_adj_2480), .B(n541), .C(index_i[4]), 
         .Z(n542_adj_2481)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_4_i542_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_2_i557_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n557_adj_2482)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C+!(D))+!B (C (D)+!C !(D))))) */ ;
    defparam mux_192_Mux_2_i557_3_lut_3_lut_4_lut.init = 16'h0f18;
    LUT4 i19185_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21515)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A (B (D)+!B !(C (D))))) */ ;
    defparam i19185_3_lut_4_lut.init = 16'h18cc;
    L6MUX21 i19449 (.D0(n21770), .D1(n21771), .SD(index_i[5]), .Z(n21779));
    LUT4 i18100_4_lut (.A(n24909), .B(n25255), .C(index_i[5]), .D(index_i[4]), 
         .Z(n20430)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam i18100_4_lut.init = 16'hc5ca;
    LUT4 mux_192_Mux_8_i285_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n285)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C (D)+!C !(D))+!B (C)))) */ ;
    defparam mux_192_Mux_8_i285_3_lut_3_lut_4_lut.init = 16'h0fc1;
    LUT4 i19142_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21472)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)))+!A !(B (C+!(D))+!B (D)))) */ ;
    defparam i19142_3_lut_3_lut_4_lut.init = 16'h71cc;
    LUT4 i19143_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21473)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B (C (D)+!C !(D))))) */ ;
    defparam i19143_3_lut_3_lut_4_lut.init = 16'h0f1c;
    LUT4 i19220_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21550)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C (D)))+!A (B (C+(D))+!B !(C)))) */ ;
    defparam i19220_4_lut_4_lut_4_lut.init = 16'h301c;
    LUT4 mux_192_Mux_0_i699_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n699)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (D))+!A (B (C+!(D))+!B !(C+!(D))))) */ ;
    defparam mux_192_Mux_0_i699_3_lut_3_lut_4_lut.init = 16'h1c33;
    LUT4 mux_192_Mux_8_i30_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n30_adj_2480)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A !(B ((D)+!C)+!B (C (D)+!C !(D))))) */ ;
    defparam mux_192_Mux_8_i30_3_lut_3_lut_4_lut.init = 16'h7e0f;
    LUT4 n699_bdd_4_lut_22545 (.A(n24876), .B(index_q[6]), .C(n24938), 
         .D(index_q[5]), .Z(n23058)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C+!(D))+!B (D))) */ ;
    defparam n699_bdd_4_lut_22545.init = 16'hd1cc;
    LUT4 mux_192_Mux_4_i286_3_lut (.A(n270), .B(n15_adj_2483), .C(index_i[4]), 
         .Z(n286_adj_2484)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_4_i286_3_lut.init = 16'hcaca;
    PFUMX i18896 (.BLUT(n21224), .ALUT(n21225), .C0(index_q[4]), .Z(n21226));
    LUT4 index_q_1__bdd_4_lut_24616 (.A(index_q[1]), .B(index_q[3]), .C(index_q[0]), 
         .D(index_q[2]), .Z(n26637)) /* synthesis lut_function=(A (B (C+(D))+!B (C (D)))+!A !(B (C)+!B !(C+(D)))) */ ;
    defparam index_q_1__bdd_4_lut_24616.init = 16'hbd94;
    LUT4 i10928_2_lut_rep_612 (.A(index_q[0]), .B(index_q[1]), .Z(n25172)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i10928_2_lut_rep_612.init = 16'h4444;
    LUT4 n23061_bdd_3_lut (.A(n23061), .B(n23058), .C(index_q[4]), .Z(n23062)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n23061_bdd_3_lut.init = 16'hcaca;
    LUT4 n26637_bdd_3_lut (.A(n26637), .B(index_q[1]), .C(index_q[4]), 
         .Z(n26638)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n26637_bdd_3_lut.init = 16'hcaca;
    PFUMX mux_192_Mux_1_i891 (.BLUT(n882), .ALUT(n890_adj_2485), .C0(n19851), 
          .Z(n891)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 i7660_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n157_adj_2486)) /* synthesis lut_function=(!(A (C (D))+!A !(B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i7660_3_lut_4_lut_4_lut.init = 16'h4aaa;
    LUT4 index_i_6__bdd_4_lut_24114 (.A(index_i[6]), .B(index_i[5]), .C(index_i[1]), 
         .D(index_i[0]), .Z(n26701)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C))+!A (B (C)+!B !(C)))) */ ;
    defparam index_i_6__bdd_4_lut_24114.init = 16'h3cbc;
    LUT4 index_i_6__bdd_1_lut (.A(index_i[5]), .Z(n26700)) /* synthesis lut_function=(!(A)) */ ;
    defparam index_i_6__bdd_1_lut.init = 16'h5555;
    LUT4 index_i_5__bdd_3_lut_24120 (.A(index_i[5]), .B(n26702), .C(index_i[3]), 
         .Z(n26703)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam index_i_5__bdd_3_lut_24120.init = 16'hcaca;
    LUT4 n25163_bdd_4_lut_24111 (.A(n24887), .B(n24970), .C(index_i[6]), 
         .D(index_i[5]), .Z(n26704)) /* synthesis lut_function=(!(A (B (C)+!B (D))+!A !(B (D)+!B (C)))) */ ;
    defparam n25163_bdd_4_lut_24111.init = 16'h5c3a;
    LUT4 n25163_bdd_4_lut_24490 (.A(n25163), .B(index_i[6]), .C(index_i[2]), 
         .D(index_i[5]), .Z(n26705)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A !(B (C+(D))+!B (D)))) */ ;
    defparam n25163_bdd_4_lut_24490.init = 16'h5fe0;
    PFUMX i18356 (.BLUT(n20682), .ALUT(n20683), .C0(index_q[5]), .Z(n20686));
    LUT4 n26706_bdd_3_lut (.A(n26706), .B(n26703), .C(index_i[4]), .Z(n26707)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n26706_bdd_3_lut.init = 16'hcaca;
    PFUMX i18357 (.BLUT(n20684), .ALUT(n20685), .C0(index_q[5]), .Z(n20687));
    LUT4 n547_bdd_4_lut_22420 (.A(index_q[2]), .B(index_q[1]), .C(index_q[3]), 
         .D(index_q[0]), .Z(n24043)) /* synthesis lut_function=(A (B (C+!(D))+!B !(D))+!A !(B (C+!(D))+!B !(D))) */ ;
    defparam n547_bdd_4_lut_22420.init = 16'h95aa;
    LUT4 mux_193_Mux_0_i954_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n954)) /* synthesis lut_function=(A (D)+!A !(B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i954_3_lut_4_lut_4_lut.init = 16'haf40;
    LUT4 mux_192_Mux_4_i94_3_lut (.A(n61), .B(n25034), .C(index_i[4]), 
         .Z(n94_adj_2487)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_4_i94_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_0_i684_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n684_adj_2488)) /* synthesis lut_function=(!(A ((D)+!B)+!A !(B (D)+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i684_3_lut_4_lut_4_lut_4_lut.init = 16'h5498;
    LUT4 mux_193_Mux_0_i953_3_lut_rep_613 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n25173)) /* synthesis lut_function=(A (C)+!A !((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i953_3_lut_rep_613.init = 16'ha4a4;
    LUT4 mux_193_Mux_6_i22_3_lut_3_lut_rep_614 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n25174)) /* synthesis lut_function=(!(A (C)+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_6_i22_3_lut_3_lut_rep_614.init = 16'h4a4a;
    LUT4 mux_193_Mux_4_i812_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n812_adj_2489)) /* synthesis lut_function=(!(A (C+(D))+!A !(B (C+(D))+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_4_i812_3_lut_3_lut_4_lut.init = 16'h554a;
    LUT4 mux_193_Mux_5_i491_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n491_adj_2490)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A !(B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_5_i491_3_lut_4_lut_4_lut.init = 16'ha54a;
    LUT4 index_i_1__bdd_4_lut (.A(index_i[1]), .B(index_i[3]), .C(index_i[0]), 
         .D(index_i[2]), .Z(n26764)) /* synthesis lut_function=(A (B (C+(D))+!B (C (D)))+!A !(B (C)+!B !(C+(D)))) */ ;
    defparam index_i_1__bdd_4_lut.init = 16'hbd94;
    PFUMX i18911 (.BLUT(n21239), .ALUT(n21240), .C0(index_q[4]), .Z(n21241));
    LUT4 mux_193_Mux_0_i475_3_lut_4_lut (.A(n25011), .B(index_q[1]), .C(index_q[3]), 
         .D(n24980), .Z(n475_adj_2414)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i475_3_lut_4_lut.init = 16'h4f40;
    LUT4 mux_193_Mux_3_i491_3_lut_4_lut (.A(n25011), .B(index_q[1]), .C(index_q[3]), 
         .D(n25199), .Z(n491_adj_2491)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_3_i491_3_lut_4_lut.init = 16'h4f40;
    LUT4 n26764_bdd_3_lut (.A(n26764), .B(index_i[1]), .C(index_i[4]), 
         .Z(n26765)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n26764_bdd_3_lut.init = 16'hcaca;
    LUT4 index_q_6__bdd_1_lut (.A(index_q[5]), .Z(n26774)) /* synthesis lut_function=(!(A)) */ ;
    defparam index_q_6__bdd_1_lut.init = 16'h5555;
    LUT4 index_q_6__bdd_4_lut_24177 (.A(index_q[6]), .B(index_q[5]), .C(index_q[1]), 
         .D(index_q[0]), .Z(n26775)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C))+!A (B (C)+!B !(C)))) */ ;
    defparam index_q_6__bdd_4_lut_24177.init = 16'h3cbc;
    LUT4 i19119_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21449)) /* synthesis lut_function=(!(A ((D)+!C)+!A !(B ((D)+!C)+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19119_3_lut_3_lut_4_lut.init = 16'h55a4;
    LUT4 n24045_bdd_3_lut (.A(n24045), .B(n24042), .C(index_q[4]), .Z(n24046)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n24045_bdd_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_0_i781_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n781_adj_2492)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A (B (C)+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i781_4_lut_4_lut_4_lut.init = 16'h0cb4;
    LUT4 index_q_5__bdd_3_lut (.A(index_q[5]), .B(n26776), .C(index_q[3]), 
         .Z(n26777)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam index_q_5__bdd_3_lut.init = 16'hcaca;
    LUT4 n25188_bdd_4_lut_24156 (.A(n24877), .B(n24957), .C(index_q[6]), 
         .D(index_q[5]), .Z(n26778)) /* synthesis lut_function=(!(A (B (C)+!B (D))+!A !(B (D)+!B (C)))) */ ;
    defparam n25188_bdd_4_lut_24156.init = 16'h5c3a;
    LUT4 n25188_bdd_4_lut (.A(n25188), .B(index_q[6]), .C(index_q[2]), 
         .D(index_q[5]), .Z(n26779)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A !(B (C+(D))+!B (D)))) */ ;
    defparam n25188_bdd_4_lut.init = 16'h5fe0;
    LUT4 n26780_bdd_3_lut (.A(n26780), .B(n26777), .C(index_q[4]), .Z(n26781)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n26780_bdd_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_5_i475_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n475_adj_2493)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_5_i475_3_lut_4_lut_4_lut.init = 16'hd4a5;
    LUT4 mux_193_Mux_0_i157_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n157_adj_2400)) /* synthesis lut_function=(A (B (C+!(D))+!B !(D))+!A (B (D)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i157_3_lut_4_lut.init = 16'hd4aa;
    PFUMX i18363 (.BLUT(n20689), .ALUT(n20690), .C0(index_q[5]), .Z(n20693));
    LUT4 i20003_3_lut (.A(n716_adj_2494), .B(n731_adj_2495), .C(index_q[4]), 
         .Z(n732_adj_2496)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20003_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_2_i669_3_lut (.A(n653_adj_2497), .B(n475_adj_2375), 
         .C(index_q[4]), .Z(n669_adj_2498)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_2_i669_3_lut.init = 16'hcaca;
    LUT4 i18550_3_lut_4_lut_4_lut_4_lut (.A(n25188), .B(index_q[2]), .C(index_q[3]), 
         .D(index_q[4]), .Z(n20880)) /* synthesis lut_function=(A (B)+!A (B (C (D))+!B !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18550_3_lut_4_lut_4_lut_4_lut.init = 16'hc999;
    PFUMX i18364 (.BLUT(n20691), .ALUT(n20692), .C0(index_q[5]), .Z(n20694));
    LUT4 mux_193_Mux_6_i325_3_lut_4_lut_4_lut_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n325)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_6_i325_3_lut_4_lut_4_lut_3_lut.init = 16'h6d6d;
    LUT4 i9451_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n526_adj_2499)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+(D)))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9451_3_lut_4_lut_4_lut.init = 16'h666c;
    LUT4 n347_bdd_3_lut_22429 (.A(n25207), .B(n25173), .C(index_q[3]), 
         .Z(n24053)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n347_bdd_3_lut_22429.init = 16'hcaca;
    LUT4 mux_193_Mux_2_i605_3_lut (.A(n142_adj_2500), .B(n604_adj_2501), 
         .C(index_q[4]), .Z(n605_adj_2502)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_2_i605_3_lut.init = 16'hcaca;
    LUT4 i18520_3_lut_3_lut (.A(n25193), .B(index_q[3]), .C(n27522), .Z(n20850)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam i18520_3_lut_3_lut.init = 16'h7474;
    LUT4 mux_193_Mux_0_i747_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n747_adj_2503)) /* synthesis lut_function=(!(A (B+!(C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i747_3_lut_4_lut_4_lut_4_lut.init = 16'h6556;
    L6MUX21 i22754 (.D0(n24452), .D1(n24449), .SD(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_2141[4]));
    LUT4 i9465_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(n25096), .D(index_q[4]), .Z(n221)) /* synthesis lut_function=(!(A (B)+!A (B (C+(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9465_3_lut_4_lut_4_lut_4_lut.init = 16'h3336;
    PFUMX i22752 (.BLUT(n24451), .ALUT(n24450), .C0(index_q[8]), .Z(n24452));
    LUT4 mux_193_Mux_1_i882_3_lut_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n882_adj_2504)) /* synthesis lut_function=(A ((C)+!B)+!A !((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_1_i882_3_lut_3_lut.init = 16'ha6a6;
    LUT4 mux_193_Mux_7_i475_3_lut_3_lut_4_lut (.A(n25188), .B(index_q[2]), 
         .C(n27521), .D(index_q[3]), .Z(n475_adj_2505)) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))+!A !(B ((D)+!C)+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_7_i475_3_lut_3_lut_4_lut.init = 16'h99f0;
    LUT4 i20011_3_lut (.A(n25252), .B(n21374), .C(index_q[4]), .Z(n21375)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20011_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_0_i645_3_lut_3_lut_rep_596_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n25156)) /* synthesis lut_function=(!(A (B)+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i645_3_lut_3_lut_rep_596_3_lut.init = 16'h6363;
    LUT4 i20013_3_lut (.A(n21370), .B(n21371), .C(index_q[4]), .Z(n21372)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20013_3_lut.init = 16'hcaca;
    LUT4 i18762_3_lut_4_lut (.A(n25188), .B(index_q[2]), .C(index_q[3]), 
         .D(n25160), .Z(n21092)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18762_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_193_Mux_5_i828_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[4]), .D(n25091), .Z(n828_adj_2506)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_5_i828_4_lut_4_lut.init = 16'hc66c;
    LUT4 mux_193_Mux_2_i413_3_lut (.A(n397_adj_2507), .B(n954_adj_2508), 
         .C(index_q[4]), .Z(n413_adj_2509)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_2_i413_3_lut.init = 16'hcaca;
    LUT4 i9503_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[4]), .Z(n444_adj_2510)) /* synthesis lut_function=(!(A (B)+!A !(B (C (D))+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9503_3_lut_4_lut_4_lut_4_lut.init = 16'h6333;
    LUT4 i9599_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n12169)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B ((D)+!C)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9599_3_lut_4_lut_4_lut.init = 16'h6c3c;
    PFUMX i18032 (.BLUT(n221_adj_2511), .ALUT(n252_adj_2331), .C0(index_i[5]), 
          .Z(n20362));
    LUT4 n61_bdd_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n24246)) /* synthesis lut_function=(!(A (B)+!A !(B (C+(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n61_bdd_3_lut_4_lut_4_lut_4_lut.init = 16'h6663;
    LUT4 mux_193_Mux_3_i507_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[4]), .D(n491_adj_2491), .Z(n507_adj_2512)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_3_i507_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_193_Mux_6_i844_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n844_adj_2454)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (B (C)+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_6_i844_3_lut_4_lut_4_lut.init = 16'hc1e0;
    LUT4 i21821_then_3_lut (.A(index_q[0]), .B(index_q[4]), .C(index_q[3]), 
         .Z(n25221)) /* synthesis lut_function=(A (B)+!A (B (C)+!B !(C))) */ ;
    defparam i21821_then_3_lut.init = 16'hc9c9;
    LUT4 mux_193_Mux_7_i108_3_lut_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n108)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_7_i108_3_lut_3_lut.init = 16'hc6c6;
    PFUMX i23012 (.BLUT(n25223), .ALUT(n25224), .C0(index_q[0]), .Z(n25225));
    LUT4 mux_193_Mux_7_i653_3_lut_4_lut (.A(n25188), .B(index_q[2]), .C(index_q[3]), 
         .D(n25055), .Z(n653_adj_2513)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_7_i653_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_193_Mux_0_i908_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n908)) /* synthesis lut_function=(!(A (B (C (D))+!B !(D))+!A (B+((D)+!C)))) */ ;
    defparam mux_193_Mux_0_i908_3_lut_4_lut_4_lut.init = 16'h2a98;
    LUT4 mux_193_Mux_5_i731_3_lut (.A(n27494), .B(n27525), .C(index_q[3]), 
         .Z(n731_adj_2450)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_5_i731_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_2_i731_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n731_adj_2495)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_2_i731_3_lut_4_lut_4_lut.init = 16'h6cc6;
    LUT4 mux_193_Mux_2_i317_3_lut (.A(n668_adj_2449), .B(n316_adj_2514), 
         .C(index_q[4]), .Z(n317_adj_2515)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_2_i317_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_2_i286_3_lut (.A(n270_adj_2516), .B(n653_adj_2383), 
         .C(index_q[4]), .Z(n286_adj_2517)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_2_i286_3_lut.init = 16'hcaca;
    LUT4 n396_bdd_3_lut_22459 (.A(n27525), .B(n25173), .C(index_q[3]), 
         .Z(n24056)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n396_bdd_3_lut_22459.init = 16'hcaca;
    LUT4 mux_193_Mux_0_i588_3_lut_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n588)) /* synthesis lut_function=(!(A (B+(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i588_3_lut_3_lut.init = 16'h5656;
    LUT4 mux_193_Mux_2_i684_3_lut_4_lut (.A(n25188), .B(index_q[2]), .C(index_q[3]), 
         .D(n27495), .Z(n684_adj_2518)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_2_i684_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_193_Mux_1_i746_3_lut_4_lut_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n746)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_1_i746_3_lut_4_lut_3_lut.init = 16'h8686;
    LUT4 mux_193_Mux_7_i526_3_lut_3_lut_4_lut_4_lut_3_lut_4_lut (.A(index_q[0]), 
         .B(index_q[1]), .C(index_q[3]), .D(index_q[2]), .Z(n526_adj_2519)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(D))+!A !(D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_7_i526_3_lut_3_lut_4_lut_4_lut_3_lut_4_lut.init = 16'h887f;
    LUT4 mux_193_Mux_6_i7_3_lut_4_lut_4_lut_3_lut_rep_616 (.A(index_q[0]), 
         .B(index_q[1]), .C(index_q[2]), .Z(n25176)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_6_i7_3_lut_4_lut_4_lut_3_lut_rep_616.init = 16'hd6d6;
    LUT4 mux_193_Mux_5_i459_3_lut_4_lut_4_lut_3_lut_rep_617 (.A(index_q[0]), 
         .B(index_q[1]), .C(index_q[2]), .Z(n25177)) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_5_i459_3_lut_4_lut_4_lut_3_lut_rep_617.init = 16'h6b6b;
    LUT4 mux_193_Mux_6_i442_3_lut_4_lut_3_lut_rep_618 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n25178)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_6_i442_3_lut_4_lut_3_lut_rep_618.init = 16'h6464;
    LUT4 i20025_3_lut (.A(n142_adj_2520), .B(n14066), .C(index_q[4]), 
         .Z(n158_adj_2521)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20025_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_0_i525_3_lut_3_lut_rep_620 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n25180)) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i525_3_lut_3_lut_rep_620.init = 16'h6a6a;
    LUT4 mux_193_Mux_2_i491_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n491_adj_2522)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A !(B (C)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_2_i491_3_lut_4_lut_4_lut.init = 16'h6a5a;
    LUT4 i18552_4_lut_4_lut_4_lut (.A(n25188), .B(index_q[2]), .C(index_q[4]), 
         .D(index_q[3]), .Z(n20882)) /* synthesis lut_function=(A (B)+!A !(B (C+(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18552_4_lut_4_lut_4_lut.init = 16'h999c;
    LUT4 mux_192_Mux_6_i844_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n844_adj_2439)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (B (C)+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_6_i844_3_lut_4_lut_4_lut.init = 16'hc1e0;
    LUT4 mux_193_Mux_4_i62_4_lut (.A(n25212), .B(n61_adj_2523), .C(index_q[4]), 
         .D(index_q[3]), .Z(n62_adj_2524)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_4_i62_4_lut.init = 16'hc5ca;
    LUT4 mux_193_Mux_4_i31_4_lut (.A(n15_adj_2525), .B(n24839), .C(index_q[4]), 
         .D(index_q[3]), .Z(n31)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_4_i31_4_lut.init = 16'h3aca;
    LUT4 mux_193_Mux_5_i30_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n30_adj_2526)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A (B+!(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_5_i30_3_lut_4_lut.init = 16'hcc67;
    LUT4 i18882_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21212)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18882_3_lut_4_lut.init = 16'h64cc;
    LUT4 mux_193_Mux_5_i460_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n460_adj_2527)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A !(B (C)+!B !(C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_5_i460_3_lut_4_lut_4_lut.init = 16'h6b5a;
    PFUMX i22749 (.BLUT(n24448), .ALUT(n20324), .C0(index_q[8]), .Z(n24449));
    LUT4 i18780_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21110)) /* synthesis lut_function=(A (B (C)+!B !(C (D)+!C !(D)))+!A (B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18780_3_lut_4_lut_4_lut.init = 16'hd6a5;
    LUT4 mux_193_Mux_3_i31_3_lut (.A(n781_adj_2528), .B(n30_adj_2529), .C(index_q[4]), 
         .Z(n31_adj_2530)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_3_i31_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_6_i15_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n15_adj_2531)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C))+!A !(B (C+!(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_6_i15_3_lut_4_lut_4_lut.init = 16'h5ad6;
    LUT4 i11416_2_lut_rep_621 (.A(index_q[0]), .B(index_q[1]), .Z(n25181)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11416_2_lut_rep_621.init = 16'h2222;
    LUT4 mux_192_Mux_5_i31_3_lut (.A(n15_adj_2532), .B(n30_adj_2533), .C(index_i[4]), 
         .Z(n31_adj_2534)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_5_i31_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_4_i205_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n205)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_4_i205_3_lut_4_lut_4_lut.init = 16'h5a2a;
    LUT4 mux_193_Mux_6_i157_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n157_adj_2535)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (D))+!A !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_6_i157_3_lut_4_lut_4_lut_4_lut.init = 16'h5d22;
    LUT4 mux_193_Mux_8_i124_3_lut_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n124_adj_2536)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C+!(D)))+!A (B (C (D)+!C !(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_8_i124_3_lut_3_lut_4_lut_4_lut.init = 16'h07c1;
    LUT4 mux_193_Mux_4_i900_3_lut_4_lut_4_lut_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n900)) /* synthesis lut_function=(A ((C)+!B)+!A !(B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_4_i900_3_lut_4_lut_4_lut_3_lut.init = 16'hb2b2;
    LUT4 mux_192_Mux_4_i62_4_lut (.A(n25123), .B(n61), .C(index_i[4]), 
         .D(index_i[3]), .Z(n62_adj_2537)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_4_i62_4_lut.init = 16'hc5ca;
    LUT4 mux_192_Mux_4_i31_4_lut (.A(n15_adj_2483), .B(n24898), .C(index_i[4]), 
         .D(index_i[3]), .Z(n31_adj_2538)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_4_i31_4_lut.init = 16'h3aca;
    LUT4 n404_bdd_3_lut_22456 (.A(n27524), .B(n27523), .C(index_q[3]), 
         .Z(n24073)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n404_bdd_3_lut_22456.init = 16'hcaca;
    LUT4 mux_193_Mux_2_i348_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n348_adj_2539)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)+!C !(D)))+!A !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_2_i348_3_lut_4_lut_4_lut_4_lut.init = 16'h5a25;
    LUT4 i18861_3_lut_3_lut_4_lut (.A(n25058), .B(index_i[2]), .C(n25041), 
         .D(index_i[3]), .Z(n21191)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18861_3_lut_3_lut_4_lut.init = 16'hf099;
    LUT4 i9544_3_lut (.A(n12109), .B(n25206), .C(index_q[3]), .Z(n12110)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9544_3_lut.init = 16'hcaca;
    LUT4 i9601_3_lut_4_lut_3_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[4]), 
         .Z(n12171)) /* synthesis lut_function=(!(A (B)+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9601_3_lut_4_lut_3_lut.init = 16'h6262;
    LUT4 n547_bdd_3_lut_22419_3_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .Z(n23960)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A ((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n547_bdd_3_lut_22419_3_lut.init = 16'h2c2c;
    LUT4 i19145_3_lut_3_lut_4_lut (.A(n25058), .B(index_i[2]), .C(n24941), 
         .D(index_i[3]), .Z(n21475)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19145_3_lut_3_lut_4_lut.init = 16'hf099;
    PFUMX i18386 (.BLUT(n20712), .ALUT(n20713), .C0(index_i[5]), .Z(n20716));
    LUT4 mux_192_Mux_3_i31_3_lut (.A(n781_adj_2477), .B(n30_adj_2467), .C(index_i[4]), 
         .Z(n31_adj_2540)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_3_i31_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_0_i985_3_lut_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n985)) /* synthesis lut_function=(!(A (B+!(C))+!A (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i985_3_lut_3_lut.init = 16'h2525;
    LUT4 mux_193_Mux_6_i70_3_lut_3_lut_rep_623 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n25183)) /* synthesis lut_function=(!(A (B+(C))+!A !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_6_i70_3_lut_3_lut_rep_623.init = 16'h5252;
    LUT4 mux_193_Mux_0_i490_3_lut_4_lut_3_lut_rep_624 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n25184)) /* synthesis lut_function=(!(A (B+!(C))+!A ((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i490_3_lut_4_lut_3_lut_rep_624.init = 16'h2424;
    LUT4 mux_193_Mux_5_i754_3_lut_4_lut_3_lut_rep_625 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n25185)) /* synthesis lut_function=(!(A (B)+!A ((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_5_i754_3_lut_4_lut_3_lut_rep_625.init = 16'h2626;
    LUT4 n404_bdd_3_lut_22448 (.A(n404), .B(n25200), .C(index_q[3]), .Z(n24072)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n404_bdd_3_lut_22448.init = 16'hcaca;
    LUT4 n476_bdd_3_lut_21856_4_lut (.A(n25058), .B(index_i[2]), .C(index_i[4]), 
         .D(n491_adj_2541), .Z(n23433)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n476_bdd_3_lut_21856_4_lut.init = 16'h9f90;
    LUT4 i18915_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21245)) /* synthesis lut_function=(!(A (B)+!A (B (C+(D))+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18915_3_lut_3_lut_4_lut.init = 16'h3326;
    LUT4 mux_193_Mux_0_i491_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n491_adj_2421)) /* synthesis lut_function=(!(A (B (D)+!B !(C+!(D)))+!A ((C+!(D))+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i491_3_lut_4_lut.init = 16'h24aa;
    LUT4 i9561_3_lut (.A(n12126), .B(n25066), .C(index_i[3]), .Z(n12127)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9561_3_lut.init = 16'hcaca;
    LUT4 i19327_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21657)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C))+!A !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19327_3_lut_4_lut_4_lut.init = 16'h5a52;
    LUT4 i18867_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21197)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A !(B (C+!(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18867_3_lut_4_lut_4_lut.init = 16'ha52b;
    LUT4 mux_192_Mux_3_i860_3_lut_4_lut (.A(n25058), .B(index_i[2]), .C(index_i[4]), 
         .D(n859_adj_2542), .Z(n860_adj_2417)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_3_i860_3_lut_4_lut.init = 16'hf606;
    LUT4 n308_bdd_3_lut_22496 (.A(n27526), .B(n25199), .C(index_q[3]), 
         .Z(n24076)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n308_bdd_3_lut_22496.init = 16'hacac;
    PFUMX i18387 (.BLUT(n20714), .ALUT(n20715), .C0(index_i[5]), .Z(n20717));
    LUT4 mux_192_Mux_7_i443_3_lut_4_lut (.A(n25058), .B(index_i[2]), .C(index_i[3]), 
         .D(n25041), .Z(n443_adj_2543)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_7_i443_3_lut_4_lut.init = 16'h6f60;
    PFUMX i18393 (.BLUT(n20719), .ALUT(n20720), .C0(index_i[5]), .Z(n20723));
    PFUMX i18394 (.BLUT(n20721), .ALUT(n20722), .C0(index_i[5]), .Z(n20724));
    LUT4 n46_bdd_4_lut (.A(n24875), .B(index_q[4]), .C(n23051), .D(index_q[5]), 
         .Z(n24798)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (B (C (D))+!B (C+!(D)))) */ ;
    defparam n46_bdd_4_lut.init = 16'hf099;
    LUT4 n78_bdd_4_lut_22479 (.A(n24884), .B(index_i[6]), .C(n24942), 
         .D(index_i[5]), .Z(n23092)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C+!(D))+!B (D))) */ ;
    defparam n78_bdd_4_lut_22479.init = 16'hd1cc;
    LUT4 mux_192_Mux_5_i891_3_lut (.A(n875_adj_2544), .B(n379), .C(index_i[4]), 
         .Z(n891_adj_2545)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_5_i891_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_5_i860_3_lut (.A(n15_adj_2532), .B(n859_adj_2546), 
         .C(index_i[4]), .Z(n860_adj_2547)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_5_i860_3_lut.init = 16'hcaca;
    LUT4 i18996_4_lut_4_lut (.A(n24877), .B(n24921), .C(index_q[5]), .D(index_q[4]), 
         .Z(n21326)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C+(D))+!B !(C (D)+!C !(D)))) */ ;
    defparam i18996_4_lut_4_lut.init = 16'hcf50;
    LUT4 i12135_2_lut_rep_628 (.A(index_q[0]), .B(index_q[1]), .Z(n25188)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i12135_2_lut_rep_628.init = 16'heeee;
    LUT4 index_i_7__bdd_4_lut (.A(index_i[7]), .B(n125_adj_2548), .C(n22851), 
         .D(index_i[5]), .Z(n24785)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(B (C+(D))+!B !((D)+!C)))) */ ;
    defparam index_i_7__bdd_4_lut.init = 16'h66f0;
    LUT4 mux_192_Mux_6_i285_3_lut_4_lut (.A(n25045), .B(index_i[2]), .C(index_i[3]), 
         .D(n25082), .Z(n285_adj_2549)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_6_i285_3_lut_4_lut.init = 16'hf606;
    LUT4 i19182_3_lut_4_lut (.A(n25045), .B(index_i[2]), .C(index_i[3]), 
         .D(n25071), .Z(n21512)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19182_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_192_Mux_5_i797_3_lut (.A(n781_adj_2550), .B(n251_adj_2551), 
         .C(index_i[4]), .Z(n797_adj_2552)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_5_i797_3_lut.init = 16'hcaca;
    LUT4 n627_bdd_1_lut_2_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n24162)) /* synthesis lut_function=(!(A (C+(D))+!A (B (C+(D))+!B (C)))) */ ;
    defparam n627_bdd_1_lut_2_lut_3_lut_4_lut.init = 16'h010f;
    LUT4 mux_193_Mux_7_i572_3_lut_rep_256_3_lut_3_lut_4_lut (.A(index_q[0]), 
         .B(index_q[1]), .C(index_q[3]), .D(index_q[2]), .Z(n24816)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)+!C !(D)))) */ ;
    defparam mux_193_Mux_7_i572_3_lut_rep_256_3_lut_3_lut_4_lut.init = 16'hfe01;
    LUT4 i20048_3_lut (.A(n21352), .B(n21353), .C(index_i[4]), .Z(n21354)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20048_3_lut.init = 16'hcaca;
    LUT4 i11223_2_lut_rep_317_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n24877)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i11223_2_lut_rep_317_3_lut_4_lut.init = 16'hfef0;
    LUT4 i19020_3_lut_4_lut (.A(n25045), .B(index_i[2]), .C(index_i[3]), 
         .D(n25088), .Z(n21350)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19020_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_192_Mux_3_i460_3_lut_4_lut (.A(n25045), .B(index_i[2]), .C(index_i[3]), 
         .D(n25083), .Z(n460_adj_2553)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_3_i460_3_lut_4_lut.init = 16'h6f60;
    LUT4 i11182_2_lut_rep_399_3_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .Z(n24959)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i11182_2_lut_rep_399_3_lut.init = 16'he0e0;
    LUT4 mux_192_Mux_5_i636_4_lut (.A(n157_adj_2554), .B(n24895), .C(index_i[4]), 
         .D(index_i[3]), .Z(n636_adj_2555)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_5_i636_4_lut.init = 16'h3aca;
    LUT4 index_i_1__bdd_4_lut_23049 (.A(index_i[1]), .B(index_i[0]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n25251)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A !(B ((D)+!C)+!B (D))) */ ;
    defparam index_i_1__bdd_4_lut_23049.init = 16'h8a51;
    LUT4 i20580_3_lut_4_lut (.A(n25057), .B(index_i[4]), .C(index_i[5]), 
         .D(n62_adj_2382), .Z(n21292)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20580_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_193_Mux_0_i333_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n333_adj_2403)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B (D))) */ ;
    defparam mux_193_Mux_0_i333_3_lut_3_lut_4_lut.init = 16'hf10e;
    LUT4 mux_193_Mux_2_i142_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n142_adj_2520)) /* synthesis lut_function=(!(A (B (D)+!B (C (D)+!C !(D)))+!A (B (D)+!B (C+!(D))))) */ ;
    defparam mux_193_Mux_2_i142_3_lut_4_lut_4_lut_4_lut.init = 16'h03ec;
    PFUMX i19012 (.BLUT(n21340), .ALUT(n21341), .C0(index_i[4]), .Z(n21342));
    LUT4 i19110_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n21440)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)+!C !(D)))+!A (B (C+!(D))+!B ((D)+!C)))) */ ;
    defparam i19110_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h0e30;
    LUT4 mux_193_Mux_3_i157_3_lut_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n157_adj_2360)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B !(C+(D))))) */ ;
    defparam mux_193_Mux_3_i157_3_lut_3_lut_3_lut_4_lut.init = 16'h1ff0;
    L6MUX21 i22715 (.D0(n24406), .D1(n24403), .SD(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_2141[9]));
    LUT4 mux_193_Mux_14_i511_4_lut_4_lut (.A(n24804), .B(index_q[7]), .C(index_q[8]), 
         .D(n254_adj_2342), .Z(n511)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (B (C+!(D))+!B !(C)))) */ ;
    defparam mux_193_Mux_14_i511_4_lut_4_lut.init = 16'h1c10;
    PFUMX i19015 (.BLUT(n21343), .ALUT(n21344), .C0(index_i[4]), .Z(n21345));
    LUT4 i20052_3_lut (.A(n17538), .B(n17539), .C(index_i[4]), .Z(n17540)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20052_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_8_i460_3_lut_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n460_adj_2556)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B ((D)+!C))) */ ;
    defparam mux_193_Mux_8_i460_3_lut_3_lut_3_lut_4_lut.init = 16'hf10f;
    LUT4 mux_193_Mux_8_i101_3_lut_3_lut_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n101_adj_2557)) /* synthesis lut_function=(!(A (B (C))+!A (B (C)+!B !(C)))) */ ;
    defparam mux_193_Mux_8_i101_3_lut_3_lut_3_lut.init = 16'h3e3e;
    LUT4 mux_192_Mux_5_i507_3_lut (.A(n491), .B(n506_adj_2471), .C(index_i[4]), 
         .Z(n507_adj_2558)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_5_i507_3_lut.init = 16'hcaca;
    PFUMX i19018 (.BLUT(n21346), .ALUT(n21347), .C0(index_i[4]), .Z(n21348));
    LUT4 i19128_3_lut_4_lut_4_lut (.A(n25188), .B(n25200), .C(index_q[3]), 
         .D(index_q[2]), .Z(n21458)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B+(C))) */ ;
    defparam i19128_3_lut_4_lut_4_lut.init = 16'hfc5c;
    LUT4 mux_192_Mux_5_i476_3_lut (.A(n460_adj_2559), .B(n475), .C(index_i[4]), 
         .Z(n476_adj_2560)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_5_i476_3_lut.init = 16'hcaca;
    PFUMX i22713 (.BLUT(n24405), .ALUT(n24404), .C0(index_q[8]), .Z(n24406));
    LUT4 mux_192_Mux_5_i413_3_lut (.A(n397_adj_2561), .B(n251_adj_2562), 
         .C(index_i[4]), .Z(n413_adj_2563)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_5_i413_3_lut.init = 16'hcaca;
    LUT4 index_q_0__bdd_2_lut (.A(index_q[0]), .B(index_q[2]), .Z(n27395)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam index_q_0__bdd_2_lut.init = 16'h6666;
    LUT4 i19031_3_lut_3_lut_4_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n21361)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B !((D)+!C)))) */ ;
    defparam i19031_3_lut_3_lut_4_lut_3_lut_4_lut.init = 16'h11ef;
    LUT4 mux_193_Mux_8_i236_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), 
         .B(index_q[1]), .C(index_q[3]), .D(index_q[2]), .Z(n236_adj_2564)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)+!C !(D)))+!A (B (C+!(D))+!B ((D)+!C))) */ ;
    defparam mux_193_Mux_8_i236_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hf1cf;
    PFUMX i19021 (.BLUT(n21349), .ALUT(n21350), .C0(index_i[4]), .Z(n21351));
    LUT4 n604_bdd_4_lut (.A(n24883), .B(index_i[4]), .C(n24733), .D(index_i[5]), 
         .Z(n24787)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (B (C (D))+!B (C+!(D)))) */ ;
    defparam n604_bdd_4_lut.init = 16'hf099;
    LUT4 index_q_0__bdd_4_lut_23112 (.A(index_q[0]), .B(index_q[3]), .C(index_q[1]), 
         .D(index_q[2]), .Z(n25252)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C (D)))+!A !(B (C+!(D))+!B !(C+(D))))) */ ;
    defparam index_q_0__bdd_4_lut_23112.init = 16'h4ae7;
    LUT4 index_q_7__bdd_4_lut_23170 (.A(index_q[7]), .B(n14882), .C(n22813), 
         .D(index_q[5]), .Z(n24786)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(B (C+(D))+!B !((D)+!C)))) */ ;
    defparam index_q_7__bdd_4_lut_23170.init = 16'h66f0;
    LUT4 i15287_3_lut (.A(n17548), .B(n17549), .C(index_i[4]), .Z(n17550)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15287_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_5_i125_3_lut (.A(n109_adj_2565), .B(n124_adj_2459), 
         .C(index_i[4]), .Z(n125_adj_2566)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_5_i125_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_8_i46_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n46_adj_2456)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (D)+!B !(C (D)+!C !(D)))) */ ;
    defparam mux_193_Mux_8_i46_3_lut_4_lut_4_lut.init = 16'hcf10;
    LUT4 mux_192_Mux_5_i94_3_lut (.A(n653_adj_2567), .B(n635_adj_2476), 
         .C(index_i[4]), .Z(n94_adj_2568)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_5_i94_3_lut.init = 16'hcaca;
    LUT4 index_q_0__bdd_4_lut (.A(index_q[0]), .B(index_q[4]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n27394)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(D))+!A !(B (D)+!B (C+!(D))))) */ ;
    defparam index_q_0__bdd_4_lut.init = 16'h7e11;
    PFUMX i19027 (.BLUT(n21355), .ALUT(n21356), .C0(index_i[4]), .Z(n21357));
    LUT4 mux_193_Mux_7_i506_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n506_adj_2569)) /* synthesis lut_function=(!(A (B (D)+!B ((D)+!C))+!A (B (D)+!B (C+!(D))))) */ ;
    defparam mux_193_Mux_7_i506_3_lut_4_lut_4_lut_4_lut.init = 16'h01ec;
    LUT4 i11211_2_lut_3_lut_4_lut (.A(index_q[1]), .B(n25096), .C(index_q[5]), 
         .D(index_q[4]), .Z(n508)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;
    defparam i11211_2_lut_3_lut_4_lut.init = 16'hf080;
    PFUMX i22710 (.BLUT(n24402), .ALUT(n20891), .C0(index_q[8]), .Z(n24403));
    LUT4 i21821_else_3_lut (.A(index_q[2]), .B(index_q[0]), .C(index_q[4]), 
         .D(index_q[3]), .Z(n25220)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)+!C !(D)))+!A (B (C+!(D))+!B !(C)))) */ ;
    defparam i21821_else_3_lut.init = 16'h1e38;
    LUT4 i11551_3_lut_4_lut (.A(n24807), .B(index_i[7]), .C(index_i[8]), 
         .D(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2126[14])) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (D))) */ ;
    defparam i11551_3_lut_4_lut.init = 16'hffe0;
    LUT4 index_i_0__bdd_4_lut (.A(index_i[0]), .B(index_i[4]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n27409)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(D))+!A !(B (D)+!B (C+!(D))))) */ ;
    defparam index_i_0__bdd_4_lut.init = 16'h7e11;
    LUT4 index_i_0__bdd_2_lut (.A(index_i[0]), .B(index_i[2]), .Z(n27410)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam index_i_0__bdd_2_lut.init = 16'h6666;
    LUT4 i2_2_lut (.A(index_i[3]), .B(index_i[5]), .Z(n6)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2_2_lut.init = 16'h8888;
    LUT4 i2_2_lut_adj_77 (.A(index_q[3]), .B(index_q[5]), .Z(n6_adj_2570)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2_2_lut_adj_77.init = 16'h8888;
    LUT4 i11410_2_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n635_adj_2294)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A (B (C+!(D))+!B (C+(D)))) */ ;
    defparam i11410_2_lut_4_lut_4_lut.init = 16'hf1fc;
    LUT4 i11391_3_lut_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n14066)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B !(C+!(D))))) */ ;
    defparam i11391_3_lut_3_lut_3_lut_4_lut.init = 16'h10ff;
    LUT4 mux_193_Mux_6_i891_3_lut (.A(n301_adj_2571), .B(n890_adj_2314), 
         .C(index_q[4]), .Z(n891_adj_2572)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_6_i891_3_lut.init = 16'hcaca;
    LUT4 i12165_2_lut_rep_378_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n24938)) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;
    defparam i12165_2_lut_rep_378_3_lut_4_lut.init = 16'he000;
    LUT4 index_q_5__bdd_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n24159)) /* synthesis lut_function=(A (B (D)+!B (C+(D)))+!A (B (D)+!B !(C (D)+!C !(D)))) */ ;
    defparam index_q_5__bdd_3_lut_4_lut_4_lut.init = 16'hef30;
    LUT4 i20064_3_lut (.A(n21245), .B(n25246), .C(index_q[4]), .Z(n21247)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20064_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_6_i828_4_lut (.A(n812_adj_2296), .B(n13956), .C(index_q[4]), 
         .D(index_q[2]), .Z(n828_adj_2573)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_6_i828_4_lut.init = 16'hfaca;
    LUT4 i19101_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n21431)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (B (C+!(D))+!B (D))) */ ;
    defparam i19101_3_lut_4_lut_4_lut_4_lut.init = 16'hf1cc;
    LUT4 mux_193_Mux_6_i797_3_lut (.A(n781_adj_2528), .B(n24816), .C(index_q[4]), 
         .Z(n797_adj_2574)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_6_i797_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_8_i506_3_lut_4_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n506_adj_2461)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B ((D)+!C)))) */ ;
    defparam mux_193_Mux_8_i506_3_lut_4_lut_3_lut_4_lut.init = 16'h0ef0;
    LUT4 mux_193_Mux_3_i30_3_lut_4_lut_4_lut_4_lut_3_lut_4_lut (.A(index_q[0]), 
         .B(index_q[1]), .C(index_q[2]), .D(index_q[3]), .Z(n30_adj_2529)) /* synthesis lut_function=(A (C)+!A (B (C)+!B ((D)+!C))) */ ;
    defparam mux_193_Mux_3_i30_3_lut_4_lut_4_lut_4_lut_3_lut_4_lut.init = 16'hf1e1;
    LUT4 n183_bdd_3_lut_22823_4_lut_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n23610)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)+!B !(C)))) */ ;
    defparam n183_bdd_3_lut_22823_4_lut_3_lut.init = 16'h6161;
    LUT4 mux_193_Mux_3_i924_3_lut (.A(n908_adj_2575), .B(index_q[0]), .C(index_q[4]), 
         .Z(n924_adj_2576)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_3_i924_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_2_i189_3_lut_3_lut_4_lut (.A(index_q[1]), .B(n25096), 
         .C(n173_adj_2577), .D(index_q[4]), .Z(n189_adj_2578)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(C+(D)))) */ ;
    defparam mux_193_Mux_2_i189_3_lut_3_lut_4_lut.init = 16'h77f0;
    LUT4 mux_193_Mux_6_i669_3_lut (.A(n653_adj_2579), .B(n668_adj_2580), 
         .C(index_q[4]), .Z(n669_adj_2581)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_6_i669_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_7_i141_3_lut_4_lut_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n141_adj_2357)) /* synthesis lut_function=(A ((C)+!B)+!A (B+!(C))) */ ;
    defparam mux_193_Mux_7_i141_3_lut_4_lut_3_lut.init = 16'he7e7;
    LUT4 mux_193_Mux_3_i891_3_lut (.A(n541_adj_2582), .B(n890_adj_2583), 
         .C(index_q[4]), .Z(n891_adj_2584)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_3_i891_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_5_i124_3_lut (.A(n25156), .B(n25190), .C(index_q[3]), 
         .Z(n124)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_5_i124_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_2_i573_3_lut_3_lut_4_lut (.A(n25211), .B(index_q[3]), 
         .C(n557_adj_2585), .D(index_q[4]), .Z(n573_adj_2586)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_2_i573_3_lut_3_lut_4_lut.init = 16'h11f0;
    LUT4 mux_193_Mux_3_i797_3_lut (.A(n731_adj_2587), .B(n796_adj_2588), 
         .C(index_q[4]), .Z(n797_adj_2589)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_3_i797_3_lut.init = 16'hcaca;
    LUT4 i19091_3_lut_4_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n21421)) /* synthesis lut_function=(A (B (D)+!B ((D)+!C))+!A (B (D)+!B (C+!(D)))) */ ;
    defparam i19091_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'hfe13;
    LUT4 mux_193_Mux_2_i716_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), 
         .B(index_q[1]), .C(index_q[3]), .D(index_q[2]), .Z(n716_adj_2494)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)+!C !(D)))+!A (B (D)+!B !((D)+!C)))) */ ;
    defparam mux_193_Mux_2_i716_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h31cf;
    LUT4 mux_193_Mux_8_i29_3_lut_rep_629 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n25189)) /* synthesis lut_function=(!(A (B (C))+!A !(B+(C)))) */ ;
    defparam mux_193_Mux_8_i29_3_lut_rep_629.init = 16'h7e7e;
    LUT4 mux_193_Mux_6_i542_3_lut (.A(n526_adj_2499), .B(n541_adj_2582), 
         .C(index_q[4]), .Z(n542_adj_2590)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_6_i542_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_5_i53_3_lut_4_lut_3_lut_rep_630 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n25190)) /* synthesis lut_function=(A ((C)+!B)+!A (B)) */ ;
    defparam mux_193_Mux_5_i53_3_lut_4_lut_3_lut_rep_630.init = 16'he6e6;
    LUT4 index_q_1__bdd_4_lut (.A(index_q[1]), .B(index_q[0]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n27528)) /* synthesis lut_function=(A (B+(C (D)+!C !(D)))+!A !(B (C+(D))+!B !(C))) */ ;
    defparam index_q_1__bdd_4_lut.init = 16'hb89e;
    LUT4 mux_193_Mux_7_i92_3_lut_rep_633 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n25193)) /* synthesis lut_function=(A (B+!(C))+!A !((C)+!B)) */ ;
    defparam mux_193_Mux_7_i92_3_lut_rep_633.init = 16'h8e8e;
    LUT4 i18352_3_lut_4_lut (.A(n25211), .B(index_q[3]), .C(index_q[4]), 
         .D(n285_adj_2591), .Z(n20682)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18352_3_lut_4_lut.init = 16'hfe0e;
    LUT4 mux_193_Mux_4_i573_3_lut_3_lut_4_lut_4_lut (.A(n25211), .B(index_q[3]), 
         .C(index_q[4]), .D(n24959), .Z(n573_adj_2592)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_4_i573_3_lut_3_lut_4_lut_4_lut.init = 16'h1f1c;
    LUT4 mux_193_Mux_0_i698_3_lut_rep_634 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n25194)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B (C)+!B !(C)))) */ ;
    defparam mux_193_Mux_0_i698_3_lut_rep_634.init = 16'h1c1c;
    LUT4 mux_193_Mux_7_i7_3_lut_4_lut_3_lut_rep_635 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n25195)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B+!(C)))) */ ;
    defparam mux_193_Mux_7_i7_3_lut_4_lut_3_lut_rep_635.init = 16'h1818;
    LUT4 mux_193_Mux_3_i669_3_lut (.A(n653_adj_2383), .B(n668_adj_2449), 
         .C(index_q[4]), .Z(n669_adj_2593)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_3_i669_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_0_i915_3_lut_rep_636 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n25196)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C)+!B !(C))) */ ;
    defparam mux_193_Mux_0_i915_3_lut_rep_636.init = 16'he3e3;
    LUT4 mux_193_Mux_0_i15_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n15_adj_2594)) /* synthesis lut_function=(A (B (C)+!B ((D)+!C))+!A (B (C)+!B !(C))) */ ;
    defparam mux_193_Mux_0_i15_3_lut_4_lut_4_lut.init = 16'he3c3;
    LUT4 mux_193_Mux_8_i892_3_lut_4_lut (.A(n24862), .B(index_q[4]), .C(index_q[5]), 
         .D(n860_adj_2351), .Z(n892)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_8_i892_3_lut_4_lut.init = 16'h4f40;
    PFUMX i18093 (.BLUT(n158_adj_2595), .ALUT(n189_adj_2596), .C0(index_i[5]), 
          .Z(n20423));
    LUT4 i19089_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21419)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A (B (D)+!B !(C (D))))) */ ;
    defparam i19089_3_lut_4_lut.init = 16'h18cc;
    LUT4 mux_193_Mux_2_i557_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n557_adj_2585)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C+!(D))+!B (C (D)+!C !(D))))) */ ;
    defparam mux_193_Mux_2_i557_3_lut_3_lut_4_lut.init = 16'h0f18;
    LUT4 n347_bdd_3_lut_22506_4_lut (.A(n25159), .B(index_q[2]), .C(index_q[3]), 
         .D(n27507), .Z(n24054)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n347_bdd_3_lut_22506_4_lut.init = 16'hf606;
    LUT4 i19124_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21454)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C (D)))+!A (B (C+(D))+!B !(C)))) */ ;
    defparam i19124_4_lut_4_lut_4_lut.init = 16'h301c;
    LUT4 n124_bdd_3_lut_21496_4_lut (.A(n25211), .B(index_q[3]), .C(index_q[4]), 
         .D(n124_adj_2597), .Z(n23038)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n124_bdd_3_lut_21496_4_lut.init = 16'hf101;
    PFUMX i21665 (.BLUT(n23221), .ALUT(n24864), .C0(index_q[5]), .Z(n23222));
    LUT4 mux_193_Mux_3_i890_3_lut_4_lut (.A(n25159), .B(index_q[2]), .C(index_q[3]), 
         .D(n325), .Z(n890_adj_2583)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_3_i890_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_193_Mux_0_i699_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n699_adj_2598)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (D))+!A (B (C+!(D))+!B !(C+!(D))))) */ ;
    defparam mux_193_Mux_0_i699_3_lut_3_lut_4_lut.init = 16'h1c33;
    LUT4 i18904_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21234)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B (C (D)+!C !(D))))) */ ;
    defparam i18904_3_lut_3_lut_4_lut.init = 16'h0f1c;
    LUT4 mux_193_Mux_3_i573_3_lut_3_lut_4_lut (.A(n25211), .B(index_q[3]), 
         .C(n460_adj_2556), .D(index_q[4]), .Z(n573_adj_2599)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_3_i573_3_lut_3_lut_4_lut.init = 16'h11f0;
    LUT4 i18903_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21233)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)))+!A !(B (C+!(D))+!B (D)))) */ ;
    defparam i18903_3_lut_3_lut_4_lut.init = 16'h71cc;
    LUT4 n10495_bdd_3_lut_22178_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n23784)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C (D)+!C !(D))+!B (C)))) */ ;
    defparam n10495_bdd_3_lut_22178_3_lut_4_lut.init = 16'h0fc1;
    LUT4 index_q_5__bdd_4_lut_24074 (.A(n85_adj_2600), .B(index_q[2]), .C(index_q[3]), 
         .D(n25188), .Z(n24160)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (B+!(C (D))))) */ ;
    defparam index_q_5__bdd_4_lut_24074.init = 16'h3a0a;
    LUT4 mux_193_Mux_7_i716_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n716_adj_2601)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C+!(D))+!B (C)))) */ ;
    defparam mux_193_Mux_7_i716_3_lut_3_lut_4_lut.init = 16'h0f81;
    LUT4 mux_193_Mux_6_i635_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n635_adj_2268)) /* synthesis lut_function=(A (B (C+(D))+!B !(D))+!A (B)) */ ;
    defparam mux_193_Mux_6_i635_3_lut_4_lut.init = 16'hcce6;
    PFUMX i18487 (.BLUT(n20815), .ALUT(n20816), .C0(index_q[5]), .Z(n20817));
    LUT4 mux_193_Mux_10_i125_3_lut_4_lut_4_lut (.A(n25211), .B(index_q[3]), 
         .C(index_q[4]), .D(n24980), .Z(n125_adj_2347)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B (C (D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_10_i125_3_lut_4_lut_4_lut.init = 16'h3efe;
    LUT4 i20088_3_lut (.A(n21233), .B(n21234), .C(index_q[4]), .Z(n21235)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20088_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_4_i526_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n526_adj_2602)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A !(B ((D)+!C)+!B (C (D)+!C !(D))))) */ ;
    defparam mux_193_Mux_4_i526_3_lut_3_lut_4_lut.init = 16'h7e0f;
    LUT4 mux_193_Mux_0_i557_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n557_adj_2603)) /* synthesis lut_function=(A ((D)+!C)+!A !((D)+!B)) */ ;
    defparam mux_193_Mux_0_i557_3_lut_4_lut.init = 16'haa4e;
    PFUMX i18490 (.BLUT(n20818), .ALUT(n20819), .C0(index_q[5]), .Z(n20820));
    LUT4 i21008_2_lut_rep_637 (.A(index_q[0]), .B(index_q[1]), .Z(n25197)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21008_2_lut_rep_637.init = 16'h9999;
    PFUMX i19066 (.BLUT(n21394), .ALUT(n21395), .C0(index_i[4]), .Z(n476));
    LUT4 i19074_3_lut_4_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n21404)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19074_3_lut_4_lut_3_lut_4_lut.init = 16'hf80f;
    LUT4 mux_193_Mux_6_i573_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[4]), .D(n572_adj_2604), .Z(n573_adj_2605)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_6_i573_3_lut_4_lut.init = 16'hf909;
    LUT4 mux_192_Mux_14_i511_4_lut_4_lut (.A(n24807), .B(index_i[7]), .C(index_i[8]), 
         .D(n254), .Z(n511_adj_2606)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (B (C+!(D))+!B !(C)))) */ ;
    defparam mux_192_Mux_14_i511_4_lut_4_lut.init = 16'h1c10;
    PFUMX i18493 (.BLUT(n20821), .ALUT(n20822), .C0(index_q[5]), .Z(n20823));
    LUT4 mux_193_Mux_3_i476_3_lut (.A(n460_adj_2607), .B(n285_adj_2608), 
         .C(index_q[4]), .Z(n476_adj_2609)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_3_i476_3_lut.init = 16'hcaca;
    LUT4 i10974_2_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n668_adj_2610)) /* synthesis lut_function=(!(A ((D)+!B)+!A (B ((D)+!C)+!B (C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i10974_2_lut_4_lut_4_lut_4_lut.init = 16'h00c9;
    LUT4 mux_193_Mux_5_i109_3_lut_3_lut_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .Z(n109_adj_2611)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_5_i109_3_lut_3_lut_3_lut.init = 16'h3939;
    LUT4 mux_193_Mux_2_i604_3_lut_4_lut_4_lut_4_lut_4_lut (.A(index_q[0]), 
         .B(index_q[1]), .C(index_q[3]), .D(index_q[2]), .Z(n604_adj_2501)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)+!C !(D)))+!A (B (C)+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_2_i604_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'h3c9f;
    LUT4 i19106_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n21436)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !(B (C+!(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19106_3_lut_4_lut_4_lut.init = 16'ha5a9;
    LUT4 mux_192_Mux_8_i124_3_lut_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n124_adj_2612)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C+!(D)))+!A (B (C (D)+!C !(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_8_i124_3_lut_3_lut_4_lut_4_lut.init = 16'h07c1;
    LUT4 i10978_2_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n844_adj_2613)) /* synthesis lut_function=(A (B+!(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i10978_2_lut_3_lut_4_lut.init = 16'h9ff9;
    LUT4 mux_193_Mux_3_i413_3_lut (.A(n397_adj_2614), .B(n25023), .C(index_q[4]), 
         .Z(n413_adj_2615)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_3_i413_3_lut.init = 16'hcaca;
    LUT4 i18783_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21113)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A (B (C (D)+!C !(D))+!B (D))) */ ;
    defparam i18783_3_lut_4_lut.init = 16'hd926;
    LUT4 mux_193_Mux_8_i732_3_lut (.A(index_q[3]), .B(n14980), .C(index_q[5]), 
         .Z(n732_adj_2616)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_8_i732_3_lut.init = 16'h3a3a;
    LUT4 i18761_3_lut_3_lut_4_lut (.A(n25054), .B(index_q[2]), .C(n25196), 
         .D(index_q[3]), .Z(n21091)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18761_3_lut_3_lut_4_lut.init = 16'hf099;
    LUT4 i19069_then_4_lut (.A(index_i[2]), .B(index_i[1]), .C(index_i[4]), 
         .D(index_i[3]), .Z(n25254)) /* synthesis lut_function=(A (B (C+(D))+!B !(C))+!A !(B (C+(D))+!B !(C+!(D)))) */ ;
    defparam i19069_then_4_lut.init = 16'h9a97;
    LUT4 i19026_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21356)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A (B (C (D)+!C !(D))+!B (D))) */ ;
    defparam i19026_3_lut_4_lut.init = 16'hd926;
    LUT4 i15282_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n17545)) /* synthesis lut_function=(A (B)+!A !(B (C (D))+!B !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i15282_3_lut_4_lut_4_lut.init = 16'h9ccc;
    LUT4 i18906_3_lut_3_lut_4_lut (.A(n25054), .B(index_q[2]), .C(n25156), 
         .D(index_q[3]), .Z(n21236)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18906_3_lut_3_lut_4_lut.init = 16'hf099;
    LUT4 n476_bdd_3_lut_21723_4_lut (.A(n25054), .B(index_q[2]), .C(index_q[4]), 
         .D(n491_adj_2617), .Z(n23275)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n476_bdd_3_lut_21723_4_lut.init = 16'h9f90;
    LUT4 i15283_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n17546)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i15283_3_lut_4_lut_4_lut_4_lut.init = 16'h3999;
    LUT4 i20597_3_lut (.A(n12169), .B(n24716), .C(index_q[5]), .Z(n12010)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20597_3_lut.init = 16'hcaca;
    LUT4 i9453_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n541_adj_2582)) /* synthesis lut_function=(A (B (C (D))+!B !(C (D)))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9453_3_lut_4_lut_4_lut_4_lut.init = 16'h9333;
    LUT4 mux_193_Mux_3_i860_3_lut_4_lut (.A(n25054), .B(index_q[2]), .C(index_q[4]), 
         .D(n859_adj_2618), .Z(n860_adj_2619)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_3_i860_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_193_Mux_7_i443_3_lut_4_lut (.A(n25054), .B(index_q[2]), .C(index_q[3]), 
         .D(n25196), .Z(n443_adj_2620)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_7_i443_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_193_Mux_3_i286_4_lut (.A(n93_adj_2621), .B(index_q[2]), .C(index_q[4]), 
         .D(n14811), .Z(n286_adj_2622)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_3_i286_4_lut.init = 16'h3aca;
    LUT4 i19069_else_4_lut (.A(index_i[2]), .B(index_i[1]), .C(index_i[4]), 
         .D(index_i[3]), .Z(n25253)) /* synthesis lut_function=(!(A (B (C)+!B (C+(D)))+!A !(B (C (D)+!C !(D))+!B (C+!(D))))) */ ;
    defparam i19069_else_4_lut.init = 16'h581f;
    LUT4 n627_bdd_3_lut_22534 (.A(n27507), .B(n27523), .C(index_q[3]), 
         .Z(n24163)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n627_bdd_3_lut_22534.init = 16'hcaca;
    LUT4 i20101_3_lut (.A(n21638), .B(n21639), .C(index_q[4]), .Z(n21640)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20101_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_7_i45_3_lut_3_lut_rep_601_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n25161)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_7_i45_3_lut_3_lut_rep_601_3_lut.init = 16'h3939;
    LUT4 mux_193_Mux_2_i955_then_4_lut (.A(index_q[4]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n25224)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B (C+!(D))+!B !(C (D)))) */ ;
    defparam mux_193_Mux_2_i955_then_4_lut.init = 16'he95d;
    LUT4 i11421_3_lut (.A(index_i[3]), .B(index_i[1]), .C(index_i[0]), 
         .Z(n14096)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11421_3_lut.init = 16'hc8c8;
    LUT4 mux_193_Mux_0_i348_3_lut_4_lut (.A(n25159), .B(index_q[2]), .C(index_q[3]), 
         .D(n27495), .Z(n348_adj_2404)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i348_3_lut_4_lut.init = 16'h6f60;
    LUT4 i9598_3_lut_4_lut_3_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[4]), 
         .Z(n12168)) /* synthesis lut_function=(A (B)+!A !(B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9598_3_lut_4_lut_3_lut.init = 16'h9898;
    LUT4 mux_193_Mux_3_i158_3_lut (.A(n142_adj_2500), .B(n157_adj_2360), 
         .C(index_q[4]), .Z(n158_adj_2623)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_3_i158_3_lut.init = 16'hcaca;
    L6MUX21 i18503 (.D0(n20831), .D1(n20832), .SD(index_q[5]), .Z(n20833));
    LUT4 mux_193_Mux_5_i572_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n572_adj_2624)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A !(B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_5_i572_3_lut_4_lut_4_lut.init = 16'ha9a5;
    LUT4 i9501_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[4]), .D(n25096), .Z(n189_adj_2443)) /* synthesis lut_function=(A (B (C (D)))+!A !(B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9501_3_lut_4_lut_4_lut_4_lut.init = 16'h9555;
    LUT4 mux_193_Mux_3_i125_3_lut (.A(n46_adj_2456), .B(n526_adj_2602), 
         .C(index_q[4]), .Z(n125_adj_2625)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_3_i125_3_lut.init = 16'hcaca;
    PFUMX i18506 (.BLUT(n20834), .ALUT(n20835), .C0(index_q[5]), .Z(n20836));
    LUT4 mux_193_Mux_2_i955_else_4_lut (.A(index_q[4]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n25223)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+(D)))+!A !(B (C+!(D))+!B !(C+!(D))))) */ ;
    defparam mux_193_Mux_2_i955_else_4_lut.init = 16'h49c6;
    LUT4 n262_bdd_3_lut_22540 (.A(n25178), .B(n27522), .C(index_q[3]), 
         .Z(n24170)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n262_bdd_3_lut_22540.init = 16'hcaca;
    LUT4 i18964_4_lut_4_lut (.A(n24887), .B(n24920), .C(index_i[5]), .D(index_i[4]), 
         .Z(n21294)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C+(D))+!B !(C (D)+!C !(D)))) */ ;
    defparam i18964_4_lut_4_lut.init = 16'hcf50;
    PFUMX i19084 (.BLUT(n21412), .ALUT(n21413), .C0(index_i[4]), .Z(n21414));
    LUT4 mux_193_Mux_6_i498_3_lut_4_lut_4_lut_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n404)) /* synthesis lut_function=(A (B+!(C))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_6_i498_3_lut_4_lut_4_lut_3_lut.init = 16'h9b9b;
    LUT4 i19328_3_lut_4_lut (.A(n25159), .B(index_q[2]), .C(index_q[3]), 
         .D(n25202), .Z(n21658)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19328_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_192_Mux_3_i348_3_lut (.A(n27518), .B(n25065), .C(index_i[3]), 
         .Z(n348)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_3_i348_3_lut.init = 16'hcaca;
    PFUMX i18509 (.BLUT(n20837), .ALUT(n20838), .C0(index_q[5]), .Z(n20839));
    LUT4 i17982_4_lut (.A(n21226), .B(n1002_adj_2398), .C(index_q[5]), 
         .D(index_q[4]), .Z(n20312)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;
    defparam i17982_4_lut.init = 16'hfaca;
    LUT4 mux_193_Mux_4_i860_3_lut (.A(n506_adj_2626), .B(n15_adj_2531), 
         .C(index_q[4]), .Z(n860_adj_2627)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_4_i860_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_5_i251_3_lut_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .Z(n251_adj_2628)) /* synthesis lut_function=(A (B)+!A (B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_5_i251_3_lut_3_lut.init = 16'hc9c9;
    LUT4 i20110_3_lut (.A(n21215), .B(n21216), .C(index_q[4]), .Z(n21217)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20110_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_3_i676_3_lut_4_lut_3_lut_rep_638 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n25198)) /* synthesis lut_function=(A (B (C))+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_3_i676_3_lut_4_lut_3_lut_rep_638.init = 16'h9494;
    LUT4 i20112_3_lut (.A(n21212), .B(n21213), .C(index_q[4]), .Z(n21214)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20112_3_lut.init = 16'hcaca;
    LUT4 i12372_1_lut_2_lut_3_lut_4_lut (.A(n24887), .B(index_i[4]), .C(index_i[6]), 
         .D(index_i[5]), .Z(n382_adj_2251)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A (C (D)))) */ ;
    defparam i12372_1_lut_2_lut_3_lut_4_lut.init = 16'h0f7f;
    PFUMX i18512 (.BLUT(n20840), .ALUT(n20841), .C0(index_q[5]), .Z(n20842));
    LUT4 mux_193_Mux_0_i219_3_lut_3_lut_3_lut_rep_639 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n25199)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i219_3_lut_3_lut_3_lut_rep_639.init = 16'h9393;
    LUT4 mux_193_Mux_0_i660_3_lut_rep_640 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n25200)) /* synthesis lut_function=(A (B)+!A (B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i660_3_lut_rep_640.init = 16'hc9c9;
    PFUMX i19090 (.BLUT(n21418), .ALUT(n21419), .C0(index_q[4]), .Z(n21420));
    PFUMX i21628 (.BLUT(n23185), .ALUT(n23184), .C0(index_i[6]), .Z(n23186));
    LUT4 mux_193_Mux_0_i715_3_lut_3_lut_rep_641 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n25201)) /* synthesis lut_function=(A (B (C))+!A !(B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i715_3_lut_3_lut_rep_641.init = 16'h9595;
    LUT4 mux_193_Mux_4_i700_3_lut (.A(n684_adj_2629), .B(index_q[1]), .C(index_q[4]), 
         .Z(n700_adj_2630)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_4_i700_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_0_i134_3_lut_4_lut_3_lut_rep_642 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n25202)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i134_3_lut_4_lut_3_lut_rep_642.init = 16'h6969;
    PFUMX i19093 (.BLUT(n21421), .ALUT(n21422), .C0(index_q[4]), .Z(n21423));
    LUT4 mux_193_Mux_6_i645_3_lut_3_lut_4_lut_3_lut_rep_643 (.A(index_q[0]), 
         .B(index_q[1]), .C(index_q[2]), .Z(n25203)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_6_i645_3_lut_3_lut_4_lut_3_lut_rep_643.init = 16'h1919;
    PFUMX mux_193_Mux_1_i891 (.BLUT(n882_adj_2504), .ALUT(n890_adj_2631), 
          .C0(n19847), .Z(n891_adj_2392)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 mux_193_Mux_4_i669_3_lut (.A(n781_adj_2528), .B(n668_adj_2632), 
         .C(index_q[4]), .Z(n669_adj_2633)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_4_i669_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_4_i573_3_lut_3_lut_4_lut_4_lut (.A(n25122), .B(index_i[3]), 
         .C(index_i[4]), .D(n24985), .Z(n573_adj_2634)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_4_i573_3_lut_3_lut_4_lut_4_lut.init = 16'h1f1c;
    LUT4 mux_193_Mux_0_i518_3_lut_4_lut_3_lut_rep_644 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n25204)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i518_3_lut_4_lut_3_lut_rep_644.init = 16'h9292;
    LUT4 mux_193_Mux_7_i77_3_lut_3_lut_rep_645 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n25205)) /* synthesis lut_function=(A (B)+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_7_i77_3_lut_3_lut_rep_645.init = 16'h9c9c;
    PFUMX i18515 (.BLUT(n20843), .ALUT(n20844), .C0(index_q[5]), .Z(n20845));
    LUT4 mux_192_Mux_3_i684_3_lut (.A(n25070), .B(n25052), .C(index_i[3]), 
         .Z(n684_adj_2635)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_3_i684_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_4_i262_3_lut_3_lut_rep_646 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n25206)) /* synthesis lut_function=(A (B+(C))+!A !(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_4_i262_3_lut_3_lut_rep_646.init = 16'ha9a9;
    LUT4 mux_193_Mux_6_i134_3_lut_4_lut_3_lut_rep_647 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n25207)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_6_i134_3_lut_4_lut_3_lut_rep_647.init = 16'h9696;
    LUT4 mux_192_Mux_7_i412_3_lut (.A(n25041), .B(n25038), .C(index_i[3]), 
         .Z(n412_adj_2636)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_7_i412_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_6_i356_3_lut_4_lut_3_lut_rep_648 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n25208)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_6_i356_3_lut_4_lut_3_lut_rep_648.init = 16'h4949;
    LUT4 mux_193_Mux_4_i542_3_lut (.A(n526_adj_2602), .B(n506_adj_2461), 
         .C(index_q[4]), .Z(n542_adj_2637)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_4_i542_3_lut.init = 16'hcaca;
    LUT4 i17976_4_lut (.A(n24906), .B(n25239), .C(index_q[5]), .D(index_q[4]), 
         .Z(n20306)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam i17976_4_lut.init = 16'hc5ca;
    LUT4 n627_bdd_3_lut (.A(n27507), .B(n588), .C(index_q[3]), .Z(n24172)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n627_bdd_3_lut.init = 16'hacac;
    LUT4 i18777_3_lut_4_lut (.A(n25022), .B(index_q[2]), .C(index_q[3]), 
         .D(n27525), .Z(n21107)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18777_3_lut_4_lut.init = 16'h6f60;
    L6MUX21 i18525 (.D0(n20853), .D1(n20854), .SD(index_q[5]), .Z(n20855));
    LUT4 mux_192_Mux_3_i908_3_lut (.A(n25085), .B(n25069), .C(index_i[3]), 
         .Z(n908_adj_2638)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_3_i908_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_6_i572_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n572_adj_2604)) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_6_i572_3_lut_4_lut.init = 16'hccd9;
    LUT4 i18382_3_lut_4_lut (.A(n25122), .B(index_i[3]), .C(index_i[4]), 
         .D(n285_adj_2639), .Z(n20712)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18382_3_lut_4_lut.init = 16'hfe0e;
    L6MUX21 i18532 (.D0(n20860), .D1(n20861), .SD(index_q[5]), .Z(n20862));
    LUT4 mux_193_Mux_0_i762_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n762_adj_2640)) /* synthesis lut_function=(A (B+!((D)+!C))+!A !(B (D)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i762_3_lut_4_lut_4_lut.init = 16'h98fc;
    LUT4 i19097_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21427)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (D))+!A !(B (C (D))+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19097_3_lut_3_lut_4_lut.init = 16'h4933;
    L6MUX21 i18539 (.D0(n20867), .D1(n20868), .SD(index_q[5]), .Z(n20869));
    PFUMX i18542 (.BLUT(n20870), .ALUT(n20871), .C0(index_q[5]), .Z(n20872));
    LUT4 mux_192_Mux_8_i732_3_lut (.A(index_i[3]), .B(n14992), .C(index_i[5]), 
         .Z(n732_adj_2641)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_8_i732_3_lut.init = 16'h3a3a;
    PFUMX i18545 (.BLUT(n20873), .ALUT(n20874), .C0(index_q[5]), .Z(n20875));
    LUT4 i19113_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21443)) /* synthesis lut_function=(A (B (C+(D))+!B ((D)+!C))+!A !(B (C+(D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19113_3_lut_4_lut.init = 16'haa96;
    PFUMX i18548 (.BLUT(n20876), .ALUT(n20877), .C0(index_q[5]), .Z(n20878));
    LUT4 n124_bdd_3_lut_21521_4_lut (.A(n25122), .B(index_i[3]), .C(index_i[4]), 
         .D(n124_adj_2642), .Z(n23063)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n124_bdd_3_lut_21521_4_lut.init = 16'hf101;
    LUT4 mux_193_Mux_3_i397_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n397_adj_2614)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !(B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_3_i397_3_lut_4_lut_4_lut.init = 16'ha95a;
    PFUMX i18551 (.BLUT(n20879), .ALUT(n20880), .C0(index_q[5]), .Z(n20881));
    LUT4 i18909_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21239)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A !(B (D)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18909_3_lut_3_lut_4_lut.init = 16'ha955;
    LUT4 mux_192_Mux_2_i270_3_lut (.A(n25072), .B(n25037), .C(index_i[3]), 
         .Z(n270_adj_2643)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_2_i270_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_2_i316_3_lut (.A(n25070), .B(n25083), .C(index_i[3]), 
         .Z(n316_adj_2644)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_2_i316_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_2_i573_3_lut_3_lut_4_lut (.A(n25122), .B(index_i[3]), 
         .C(n557_adj_2482), .D(index_i[4]), .Z(n573_adj_2430)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_2_i573_3_lut_3_lut_4_lut.init = 16'h11f0;
    PFUMX i19102 (.BLUT(n21430), .ALUT(n21431), .C0(index_q[4]), .Z(n21432));
    LUT4 mux_193_Mux_3_i859_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n859_adj_2618)) /* synthesis lut_function=(!(A (B (D)+!B !(D))+!A (B (C+(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_3_i859_3_lut_3_lut_4_lut.init = 16'h339c;
    LUT4 i19034_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21364)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C))+!A !(B ((D)+!C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19034_3_lut_4_lut_4_lut.init = 16'h925a;
    PFUMX i18554 (.BLUT(n20882), .ALUT(n20883), .C0(index_q[5]), .Z(n20884));
    LUT4 i19167_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .D(index_i[3]), .Z(n21497)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(D))+!A (B+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19167_3_lut_4_lut_4_lut_4_lut.init = 16'h3380;
    PFUMX i19105 (.BLUT(n21433), .ALUT(n21434), .C0(index_q[4]), .Z(n21435));
    LUT4 mux_192_Mux_3_i573_3_lut_3_lut_4_lut (.A(n25122), .B(index_i[3]), 
         .C(n397), .D(index_i[4]), .Z(n573)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_3_i573_3_lut_3_lut_4_lut.init = 16'h11f0;
    LUT4 mux_193_Mux_0_i812_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n812_adj_2645)) /* synthesis lut_function=(A (B (C+(D))+!B !(C))+!A (B (D)+!B !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i812_3_lut_4_lut_4_lut_4_lut.init = 16'hcf92;
    PFUMX i18557 (.BLUT(n20885), .ALUT(n20886), .C0(index_q[5]), .Z(n20887));
    LUT4 i18764_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21094)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(D))+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18764_3_lut_3_lut_4_lut.init = 16'h3319;
    LUT4 mux_193_Mux_0_i142_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n142_adj_2399)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C))+!A !(B (C (D)+!C !(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i142_3_lut_4_lut_4_lut.init = 16'ha569;
    PFUMX i19108 (.BLUT(n21436), .ALUT(n21437), .C0(index_q[4]), .Z(n21438));
    LUT4 mux_193_Mux_1_i93_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n93_adj_2463)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C+(D)))+!A !(B (C (D)+!C !(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_1_i93_3_lut_4_lut_4_lut.init = 16'h955a;
    LUT4 mux_192_Mux_4_i491_3_lut_4_lut_4_lut (.A(index_i[2]), .B(n25165), 
         .C(index_i[3]), .D(n25058), .Z(n491_adj_2541)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_4_i491_3_lut_4_lut_4_lut.init = 16'hfc5c;
    LUT4 i18936_3_lut_4_lut (.A(n24906), .B(n24876), .C(index_q[4]), .D(index_q[5]), 
         .Z(n21266)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (B+((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18936_3_lut_4_lut.init = 16'hffc5;
    LUT4 mux_192_Mux_2_i397_3_lut (.A(n27503), .B(n25041), .C(index_i[3]), 
         .Z(n397_adj_2646)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_2_i397_3_lut.init = 16'hcaca;
    PFUMX i19111 (.BLUT(n21439), .ALUT(n21440), .C0(index_q[4]), .Z(n21441));
    LUT4 mux_192_Mux_10_i125_3_lut_4_lut_4_lut (.A(n25122), .B(index_i[3]), 
         .C(index_i[4]), .D(n24947), .Z(n125)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B (C (D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_10_i125_3_lut_4_lut_4_lut.init = 16'h3efe;
    LUT4 i19086_3_lut_4_lut (.A(n25022), .B(index_q[2]), .C(index_q[3]), 
         .D(n25208), .Z(n21416)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19086_3_lut_4_lut.init = 16'hf606;
    LUT4 i19131_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21461)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C+(D)))+!A (B (C)+!B !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19131_3_lut_4_lut_4_lut.init = 16'hc95a;
    PFUMX i18567 (.BLUT(n20895), .ALUT(n20896), .C0(index_q[5]), .Z(n20897));
    LUT4 i18770_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21100)) /* synthesis lut_function=(A (B (C (D))+!B !(C (D)))+!A !(B (D)+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18770_3_lut_4_lut_4_lut.init = 16'h9366;
    LUT4 i19121_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21451)) /* synthesis lut_function=(A (B (C)+!B (C (D)+!C !(D)))+!A !(B (C+!(D))+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19121_3_lut_4_lut_4_lut.init = 16'ha593;
    LUT4 mux_193_Mux_1_i557_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n557_adj_2647)) /* synthesis lut_function=(A (B (C+(D)))+!A (B ((D)+!C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_1_i557_3_lut_4_lut.init = 16'hcc94;
    PFUMX i18573 (.BLUT(n20901), .ALUT(n20902), .C0(index_i[5]), .Z(n20903));
    LUT4 mux_193_Mux_4_i286_3_lut (.A(n270_adj_2648), .B(n15_adj_2525), 
         .C(index_q[4]), .Z(n286_adj_2649)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_4_i286_3_lut.init = 16'hcaca;
    PFUMX i18576 (.BLUT(n20904), .ALUT(n20905), .C0(index_i[5]), .Z(n20906));
    LUT4 mux_193_Mux_2_i653_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n653_adj_2497)) /* synthesis lut_function=(A (B (C+!(D))+!B !(D))+!A !(B (C+!(D))+!B !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_2_i653_3_lut_4_lut.init = 16'h94aa;
    LUT4 i11409_2_lut_rep_651 (.A(index_q[1]), .B(index_q[2]), .Z(n25211)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11409_2_lut_rep_651.init = 16'h8888;
    LUT4 i11652_2_lut_rep_337_2_lut_3_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[0]), .Z(n24897)) /* synthesis lut_function=(A (B+!(C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11652_2_lut_rep_337_2_lut_3_lut.init = 16'h8f8f;
    PFUMX i18579 (.BLUT(n20907), .ALUT(n20908), .C0(index_i[5]), .Z(n20909));
    LUT4 index_q_1__bdd_4_lut_23356 (.A(index_q[1]), .B(index_q[0]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n25256)) /* synthesis lut_function=(!(A (B (D)+!B (C+!(D)))+!A !(B (C (D)+!C !(D))+!B !((D)+!C)))) */ ;
    defparam index_q_1__bdd_4_lut_23356.init = 16'h429c;
    LUT4 i20551_3_lut_4_lut (.A(n25091), .B(index_q[4]), .C(index_q[5]), 
         .D(n62_adj_2350), .Z(n21324)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20551_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_193_Mux_8_i491_3_lut_3_lut_3_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .D(index_q[0]), .Z(n491_adj_2650)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_8_i491_3_lut_3_lut_3_lut_4_lut.init = 16'h7870;
    LUT4 i9467_3_lut_4_lut (.A(n25181), .B(index_q[2]), .C(n25095), .D(n25207), 
         .Z(n444_adj_2651)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9467_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_193_Mux_4_i94_3_lut (.A(n61_adj_2523), .B(n25020), .C(index_q[4]), 
         .Z(n94_adj_2652)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_4_i94_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_8_i635_3_lut_4_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n635_adj_2448)) /* synthesis lut_function=(!(A (B (C (D))+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_8_i635_3_lut_4_lut_3_lut_4_lut.init = 16'h0ff8;
    LUT4 mux_193_Mux_1_i747_4_lut_then_4_lut (.A(index_q[0]), .B(index_q[4]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n25258)) /* synthesis lut_function=(A (B ((D)+!C))+!A !(B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_1_i747_4_lut_then_4_lut.init = 16'h9d5d;
    PFUMX i19117 (.BLUT(n21445), .ALUT(n21446), .C0(index_q[4]), .Z(n21447));
    LUT4 mux_193_Mux_4_i747_3_lut_4_lut (.A(n25181), .B(index_q[2]), .C(index_q[3]), 
         .D(n27525), .Z(n747_adj_2452)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_4_i747_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_193_Mux_1_i747_4_lut_else_4_lut (.A(index_q[0]), .B(index_q[4]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n25257)) /* synthesis lut_function=(!(A (B (C (D))+!B !(D))+!A ((C (D))+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_1_i747_4_lut_else_4_lut.init = 16'h2ecc;
    LUT4 mux_193_Mux_6_i285_3_lut_4_lut (.A(n25022), .B(index_q[2]), .C(index_q[3]), 
         .D(n25202), .Z(n285_adj_2608)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_6_i285_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_193_Mux_3_i460_3_lut_4_lut (.A(n25022), .B(index_q[2]), .C(index_q[3]), 
         .D(n25180), .Z(n460_adj_2607)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_3_i460_3_lut_4_lut.init = 16'h6f60;
    LUT4 i11568_2_lut_rep_397_3_lut (.A(index_q[1]), .B(index_q[2]), .C(index_q[0]), 
         .Z(n24957)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11568_2_lut_rep_397_3_lut.init = 16'h8080;
    L6MUX21 i18589 (.D0(n20917), .D1(n20918), .SD(index_i[5]), .Z(n20919));
    LUT4 mux_193_Mux_6_i251_3_lut_4_lut (.A(n25181), .B(index_q[2]), .C(index_q[3]), 
         .D(n25207), .Z(n251_adj_2653)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_6_i251_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_192_Mux_6_i891_3_lut (.A(n78), .B(n890_adj_2654), .C(index_i[4]), 
         .Z(n891_adj_2655)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_6_i891_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_8_i412_3_lut_4_lut_3_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .Z(n14766)) /* synthesis lut_function=(A (B+!(C))+!A !((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_8_i412_3_lut_4_lut_3_lut.init = 16'h8e8e;
    PFUMX i18592 (.BLUT(n20920), .ALUT(n20921), .C0(index_i[5]), .Z(n20922));
    LUT4 mux_192_Mux_6_i828_4_lut (.A(n812_adj_2288), .B(n14053), .C(index_i[4]), 
         .D(index_i[2]), .Z(n828_adj_2656)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_6_i828_4_lut.init = 16'hfaca;
    PFUMX i18595 (.BLUT(n20923), .ALUT(n20924), .C0(index_i[5]), .Z(n20925));
    PFUMX i19123 (.BLUT(n21451), .ALUT(n21452), .C0(index_q[4]), .Z(n21453));
    LUT4 i9527_2_lut_3_lut (.A(index_q[1]), .B(index_q[2]), .C(index_q[3]), 
         .Z(n12093)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9527_2_lut_3_lut.init = 16'h8080;
    LUT4 mux_192_Mux_6_i797_3_lut (.A(n781_adj_2477), .B(n24814), .C(index_i[4]), 
         .Z(n797_adj_2657)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_6_i797_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_4_i93_3_lut_4_lut_3_lut_rep_460_4_lut (.A(index_q[1]), 
         .B(index_q[2]), .C(index_q[3]), .D(index_q[0]), .Z(n25020)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_4_i93_3_lut_4_lut_3_lut_rep_460_4_lut.init = 16'h07f0;
    LUT4 mux_193_Mux_9_i412_3_lut_3_lut_4_lut_3_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .Z(n412_adj_2361)) /* synthesis lut_function=(!(A (B (C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_9_i412_3_lut_3_lut_4_lut_3_lut.init = 16'h7e7e;
    PFUMX i19126 (.BLUT(n21454), .ALUT(n21455), .C0(index_q[4]), .Z(n21456));
    LUT4 i19038_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[0]), .D(index_q[3]), .Z(n21368)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(D))+!A (B+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19038_3_lut_4_lut_4_lut_4_lut.init = 16'h3380;
    LUT4 i11221_2_lut_rep_346_3_lut (.A(index_q[1]), .B(index_q[2]), .C(index_q[3]), 
         .Z(n24906)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11221_2_lut_rep_346_3_lut.init = 16'hf8f8;
    LUT4 mux_192_Mux_6_i669_3_lut (.A(n653_adj_2567), .B(n668_adj_2658), 
         .C(index_i[4]), .Z(n669_adj_2659)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_6_i669_3_lut.init = 16'hcaca;
    PFUMX i18598 (.BLUT(n20926), .ALUT(n20927), .C0(index_i[5]), .Z(n20928));
    LUT4 mux_193_Mux_9_i30_3_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .D(index_q[0]), .Z(n30_adj_2660)) /* synthesis lut_function=(A (B (C (D))+!B !(C))+!A !(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_9_i30_3_lut_4_lut_4_lut.init = 16'h8303;
    LUT4 i15268_3_lut_4_lut_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .D(index_q[0]), .Z(n17531)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C (D)+!C !(D)))+!A !(B (D)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i15268_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'h83fc;
    PFUMX i18606 (.BLUT(n956_adj_2344), .ALUT(n17673), .C0(index_q[6]), 
          .Z(n20936));
    LUT4 i11201_2_lut_rep_316_3_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .D(index_q[0]), .Z(n24876)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11201_2_lut_rep_316_3_lut_4_lut.init = 16'hf8f0;
    PFUMX i19129 (.BLUT(n21457), .ALUT(n21458), .C0(index_q[4]), .Z(n21459));
    LUT4 mux_192_Mux_6_i542_3_lut (.A(n526_adj_2283), .B(n541_adj_2661), 
         .C(index_i[4]), .Z(n542_adj_2662)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_6_i542_3_lut.init = 16'hcaca;
    LUT4 i18886_3_lut_4_lut_3_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .D(index_q[0]), .Z(n21216)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18886_3_lut_4_lut_3_lut_4_lut.init = 16'hf80f;
    LUT4 i18865_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .D(index_q[0]), .Z(n21195)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C (D)+!C !(D)))+!A !(B (D)+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18865_3_lut_4_lut_4_lut_4_lut.init = 16'h7c03;
    PFUMX i18616 (.BLUT(n20944), .ALUT(n20945), .C0(index_i[5]), .Z(n20946));
    LUT4 mux_193_Mux_3_i142_3_lut_3_lut_3_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .Z(n142_adj_2500)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_3_i142_3_lut_3_lut_3_lut.init = 16'h3838;
    LUT4 i11565_2_lut_rep_652 (.A(index_q[1]), .B(index_q[2]), .C(index_q[0]), 
         .Z(n25212)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11565_2_lut_rep_652.init = 16'h7070;
    LUT4 mux_193_Mux_0_i1017_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[0]), .D(index_q[3]), .Z(n1017)) /* synthesis lut_function=(A (B (D)+!B !((D)+!C))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i1017_4_lut_4_lut_4_lut.init = 16'hdd70;
    L6MUX21 i18623 (.D0(n20951), .D1(n20952), .SD(index_i[5]), .Z(n20953));
    L6MUX21 i18630 (.D0(n20958), .D1(n20959), .SD(index_i[5]), .Z(n20960));
    L6MUX21 i18637 (.D0(n20965), .D1(n20966), .SD(index_i[5]), .Z(n20967));
    PFUMX i18640 (.BLUT(n20968), .ALUT(n20969), .C0(index_i[5]), .Z(n20970));
    LUT4 mux_192_Mux_8_i892_3_lut_4_lut (.A(n24861), .B(index_i[4]), .C(index_i[5]), 
         .D(n860_adj_2378), .Z(n892_adj_2663)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_8_i892_3_lut_4_lut.init = 16'h4f40;
    PFUMX i18643 (.BLUT(n20971), .ALUT(n20972), .C0(index_i[5]), .Z(n20973));
    PFUMX i18646 (.BLUT(n20974), .ALUT(n20975), .C0(index_i[5]), .Z(n20976));
    PFUMX i18649 (.BLUT(n20977), .ALUT(n20978), .C0(index_i[5]), .Z(n20979));
    LUT4 i18812_3_lut_4_lut (.A(n24909), .B(n24884), .C(index_i[4]), .D(index_i[5]), 
         .Z(n21142)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (B+((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18812_3_lut_4_lut.init = 16'hffc5;
    LUT4 i20152_3_lut (.A(n270_adj_2664), .B(n285_adj_2665), .C(index_q[4]), 
         .Z(n21062)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20152_3_lut.init = 16'hcaca;
    PFUMX i18652 (.BLUT(n20980), .ALUT(n20981), .C0(index_i[5]), .Z(n20982));
    LUT4 i18731_3_lut (.A(n236_adj_2666), .B(n251), .C(index_q[4]), .Z(n21061)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18731_3_lut.init = 16'hcaca;
    LUT4 i18724_3_lut (.A(n15_adj_2594), .B(n25247), .C(index_q[4]), .Z(n21054)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18724_3_lut.init = 16'hcaca;
    LUT4 i19032_3_lut_4_lut (.A(n25188), .B(index_q[2]), .C(index_q[3]), 
         .D(n141_adj_2357), .Z(n21362)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19032_3_lut_4_lut.init = 16'hf202;
    PFUMX i18655 (.BLUT(n20983), .ALUT(n20984), .C0(index_i[5]), .Z(n20985));
    PFUMX i18658 (.BLUT(n20986), .ALUT(n20987), .C0(index_i[5]), .Z(n20988));
    PFUMX i17921 (.BLUT(n31_adj_2667), .ALUT(n21096), .C0(index_q[5]), 
          .Z(n20251));
    LUT4 i19149_3_lut (.A(n25070), .B(n25088), .C(index_i[3]), .Z(n21479)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19149_3_lut.init = 16'hcaca;
    PFUMX i17922 (.BLUT(n94_adj_2668), .ALUT(n125_adj_2669), .C0(index_q[5]), 
          .Z(n20252));
    PFUMX i18678 (.BLUT(n20992), .ALUT(n20993), .C0(index_i[5]), .Z(n21008));
    LUT4 mux_193_Mux_5_i891_3_lut (.A(n875_adj_2670), .B(n379_adj_2671), 
         .C(index_q[4]), .Z(n891_adj_2672)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_5_i891_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_5_i860_3_lut (.A(n15_adj_2673), .B(n859_adj_2674), 
         .C(index_q[4]), .Z(n860_adj_2675)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_5_i860_3_lut.init = 16'hcaca;
    PFUMX i18679 (.BLUT(n20994), .ALUT(n20995), .C0(index_i[5]), .Z(n21009));
    LUT4 mux_193_Mux_5_i797_3_lut (.A(n781_adj_2676), .B(n251_adj_2628), 
         .C(index_q[4]), .Z(n797_adj_2677)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_5_i797_3_lut.init = 16'hcaca;
    LUT4 i18768_3_lut_4_lut (.A(n25026), .B(index_q[1]), .C(index_q[3]), 
         .D(n404), .Z(n21098)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18768_3_lut_4_lut.init = 16'hdfd0;
    LUT4 i20507_3_lut (.A(n21475), .B(n21476), .C(index_i[4]), .Z(n21477)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20507_3_lut.init = 16'hcaca;
    LUT4 n250_bdd_3_lut_22582 (.A(n25202), .B(n27523), .C(index_q[3]), 
         .Z(n24243)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n250_bdd_3_lut_22582.init = 16'hacac;
    LUT4 i20175_3_lut (.A(n21109), .B(n21110), .C(index_q[4]), .Z(n21111)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20175_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_0_i173_3_lut_4_lut (.A(n25026), .B(index_q[1]), .C(index_q[3]), 
         .D(n25204), .Z(n173_adj_2401)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i173_3_lut_4_lut.init = 16'hdfd0;
    PFUMX i17923 (.BLUT(n17547), .ALUT(n14329), .C0(index_q[5]), .Z(n20253));
    LUT4 mux_193_Mux_1_i620_3_lut_4_lut (.A(n25026), .B(index_q[1]), .C(index_q[3]), 
         .D(n25206), .Z(n620_adj_2293)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_1_i620_3_lut_4_lut.init = 16'hdfd0;
    LUT4 mux_193_Mux_5_i636_4_lut (.A(n157_adj_2486), .B(n24897), .C(index_q[4]), 
         .D(index_q[3]), .Z(n636_adj_2678)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_5_i636_4_lut.init = 16'h3aca;
    L6MUX21 i17925 (.D0(n21099), .D1(n21102), .SD(index_q[5]), .Z(n20255));
    L6MUX21 i17926 (.D0(n21105), .D1(n21108), .SD(index_q[5]), .Z(n20256));
    LUT4 i20178_3_lut (.A(n17531), .B(n17532), .C(index_q[4]), .Z(n17533)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20178_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_5_i507_3_lut (.A(n491_adj_2490), .B(n506_adj_2626), 
         .C(index_q[4]), .Z(n507_adj_2679)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_5_i507_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_5_i476_3_lut (.A(n460_adj_2527), .B(n475_adj_2493), 
         .C(index_q[4]), .Z(n476_adj_2680)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_5_i476_3_lut.init = 16'hcaca;
    LUT4 i18669_3_lut (.A(n827), .B(n251_adj_2298), .C(index_i[4]), .Z(n20999)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18669_3_lut.init = 16'hcaca;
    LUT4 i18391_3_lut_4_lut_4_lut (.A(n25057), .B(n24887), .C(index_i[4]), 
         .D(n25058), .Z(n20721)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B (C (D))+!B ((D)+!C)))) */ ;
    defparam i18391_3_lut_4_lut_4_lut.init = 16'h0c5c;
    PFUMX i17927 (.BLUT(n413_adj_2681), .ALUT(n444_adj_2651), .C0(index_q[5]), 
          .Z(n20257));
    LUT4 mux_193_Mux_5_i413_3_lut (.A(n397_adj_2682), .B(n251_adj_2653), 
         .C(index_q[4]), .Z(n413_adj_2681)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_5_i413_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_8_i763_3_lut_4_lut_4_lut (.A(n25057), .B(n24942), .C(index_i[4]), 
         .D(n25058), .Z(n14992)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam mux_192_Mux_8_i763_3_lut_4_lut_4_lut.init = 16'hcfca;
    L6MUX21 i22587 (.D0(n24247), .D1(n24245), .SD(index_q[4]), .Z(n24248));
    LUT4 mux_192_Mux_1_i986_3_lut (.A(n25165), .B(n27518), .C(index_i[3]), 
         .Z(n986_adj_2683)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_1_i986_3_lut.init = 16'hcaca;
    LUT4 i15284_3_lut (.A(n17545), .B(n17546), .C(index_q[4]), .Z(n17547)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15284_3_lut.init = 16'hcaca;
    L6MUX21 i18680 (.D0(n20996), .D1(n20997), .SD(index_i[5]), .Z(n21010));
    PFUMX i18681 (.BLUT(n20998), .ALUT(n20999), .C0(index_i[5]), .Z(n21011));
    LUT4 i19140_3_lut (.A(n27498), .B(n25077), .C(index_i[3]), .Z(n21470)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19140_3_lut.init = 16'hcaca;
    LUT4 i19139_3_lut (.A(n25087), .B(n25071), .C(index_i[3]), .Z(n21469)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19139_3_lut.init = 16'hcaca;
    LUT4 i20513_3_lut (.A(n21469), .B(n21470), .C(index_i[4]), .Z(n21471)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20513_3_lut.init = 16'hcaca;
    LUT4 i19137_3_lut (.A(n27503), .B(n25169), .C(index_i[3]), .Z(n21467)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19137_3_lut.init = 16'hcaca;
    LUT4 i18662_3_lut (.A(n541_adj_2473), .B(n25251), .C(index_i[4]), 
         .Z(n20992)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18662_3_lut.init = 16'hcaca;
    PFUMX i22585 (.BLUT(n24857), .ALUT(n24246), .C0(index_q[5]), .Z(n24247));
    PFUMX i17928 (.BLUT(n476_adj_2680), .ALUT(n507_adj_2679), .C0(index_q[5]), 
          .Z(n20258));
    L6MUX21 i18683 (.D0(n21002), .D1(n21003), .SD(index_i[5]), .Z(n21013));
    LUT4 mux_193_Mux_5_i125_3_lut (.A(n109_adj_2611), .B(n124), .C(index_q[4]), 
         .Z(n125_adj_2669)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_5_i125_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_5_i94_3_lut (.A(n653_adj_2579), .B(n635_adj_2268), 
         .C(index_q[4]), .Z(n94_adj_2668)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_5_i94_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_5_i31_3_lut (.A(n15_adj_2673), .B(n30_adj_2526), .C(index_q[4]), 
         .Z(n31_adj_2667)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_5_i31_3_lut.init = 16'hcaca;
    L6MUX21 i18684 (.D0(n21004), .D1(n21005), .SD(index_i[5]), .Z(n21014));
    LUT4 i18657_3_lut (.A(n747_adj_2303), .B(n762_adj_2349), .C(index_i[4]), 
         .Z(n20987)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18657_3_lut.init = 16'hcaca;
    L6MUX21 i18685 (.D0(n21006), .D1(n21007), .SD(index_i[5]), .Z(n21015));
    PFUMX i17929 (.BLUT(n17533), .ALUT(n573_adj_2684), .C0(index_q[5]), 
          .Z(n20259));
    LUT4 i18656_3_lut (.A(n716_adj_2479), .B(n14802), .C(index_i[4]), 
         .Z(n20986)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18656_3_lut.init = 16'hcaca;
    LUT4 i19136_3_lut (.A(n25166), .B(n85), .C(index_i[3]), .Z(n21466)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19136_3_lut.init = 16'hcaca;
    LUT4 i20515_3_lut (.A(n21466), .B(n21467), .C(index_i[4]), .Z(n21468)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20515_3_lut.init = 16'hcaca;
    LUT4 i18654_3_lut (.A(n93_adj_2685), .B(n699_adj_2330), .C(index_i[4]), 
         .Z(n20984)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18654_3_lut.init = 16'hcaca;
    PFUMX i17930 (.BLUT(n605_adj_2686), .ALUT(n636_adj_2678), .C0(index_q[5]), 
          .Z(n20260));
    LUT4 i9481_3_lut_4_lut_4_lut (.A(n25116), .B(index_i[3]), .C(index_i[5]), 
         .D(n24970), .Z(n12047)) /* synthesis lut_function=(A (B+(C (D)))+!A (B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9481_3_lut_4_lut_4_lut.init = 16'hf8c8;
    PFUMX i22583 (.BLUT(n24244), .ALUT(n24243), .C0(index_q[5]), .Z(n24245));
    LUT4 n604_bdd_3_lut_4_lut_4_lut (.A(n25116), .B(index_i[3]), .C(index_i[4]), 
         .D(n24947), .Z(n24737)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C))+!A !(B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n604_bdd_3_lut_4_lut_4_lut.init = 16'h838f;
    LUT4 i18653_3_lut (.A(n653_adj_2687), .B(n24838), .C(index_i[4]), 
         .Z(n20983)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18653_3_lut.init = 16'hcaca;
    LUT4 i18384_3_lut_3_lut_4_lut_4_lut (.A(n25116), .B(index_i[3]), .C(index_i[4]), 
         .D(n24985), .Z(n20714)) /* synthesis lut_function=(!(A (B (C)+!B ((D)+!C))+!A (B+((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18384_3_lut_3_lut_4_lut_4_lut.init = 16'h0838;
    LUT4 n62_bdd_3_lut_22521_4_lut (.A(n25116), .B(index_i[3]), .C(index_i[4]), 
         .D(n30), .Z(n23066)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n62_bdd_3_lut_22521_4_lut.init = 16'hf808;
    LUT4 i18647_3_lut (.A(n526_adj_2688), .B(n541_adj_2473), .C(index_i[4]), 
         .Z(n20977)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18647_3_lut.init = 16'hcaca;
    LUT4 i18644_3_lut (.A(n397_adj_2689), .B(n475_adj_2690), .C(index_i[4]), 
         .Z(n20974)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18644_3_lut.init = 16'hcaca;
    LUT4 i18642_3_lut (.A(n348_adj_2691), .B(n443_adj_2543), .C(index_i[4]), 
         .Z(n20972)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18642_3_lut.init = 16'hcaca;
    LUT4 i18641_3_lut (.A(n397_adj_2689), .B(n412_adj_2636), .C(index_i[4]), 
         .Z(n20971)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18641_3_lut.init = 16'hcaca;
    LUT4 i19125_3_lut_4_lut (.A(n25054), .B(index_q[2]), .C(index_q[3]), 
         .D(n27524), .Z(n21455)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19125_3_lut_4_lut.init = 16'hf404;
    PFUMX i17931 (.BLUT(n21111), .ALUT(n700_adj_2692), .C0(index_q[5]), 
          .Z(n20261));
    LUT4 i19133_3_lut (.A(n25183), .B(n25177), .C(index_q[3]), .Z(n21463)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19133_3_lut.init = 16'hcaca;
    LUT4 i19948_3_lut (.A(n21463), .B(n21464), .C(index_q[4]), .Z(n21465)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19948_3_lut.init = 16'hcaca;
    LUT4 i18639_3_lut (.A(n364), .B(n379), .C(index_i[4]), .Z(n20969)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18639_3_lut.init = 16'hcaca;
    LUT4 i18638_3_lut (.A(n333_adj_2693), .B(n348_adj_2691), .C(index_i[4]), 
         .Z(n20968)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18638_3_lut.init = 16'hcaca;
    LUT4 i12191_2_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(n25095), 
         .D(index_q[2]), .Z(n14882)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12191_2_lut_3_lut_4_lut.init = 16'hf080;
    LUT4 i18361_3_lut_4_lut_4_lut (.A(n25091), .B(n24877), .C(index_q[4]), 
         .D(n25054), .Z(n20691)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B (C (D))+!B ((D)+!C)))) */ ;
    defparam i18361_3_lut_4_lut_4_lut.init = 16'h0c5c;
    L6MUX21 i17932 (.D0(n732_adj_2451), .D1(n21114), .SD(index_q[5]), 
            .Z(n20262));
    LUT4 mux_193_Mux_8_i763_3_lut_4_lut_4_lut (.A(n25091), .B(n24938), .C(index_q[4]), 
         .D(n25054), .Z(n14980)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam mux_193_Mux_8_i763_3_lut_4_lut_4_lut.init = 16'hcfca;
    PFUMX i17933 (.BLUT(n797_adj_2677), .ALUT(n828_adj_2506), .C0(index_q[5]), 
          .Z(n20263));
    LUT4 i11285_2_lut_rep_324_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n24884)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11285_2_lut_rep_324_3_lut_4_lut.init = 16'hf8f0;
    LUT4 i19130_3_lut (.A(n1001), .B(n588), .C(index_q[3]), .Z(n21460)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19130_3_lut.init = 16'hcaca;
    LUT4 i18354_3_lut_3_lut_4_lut_4_lut (.A(n25097), .B(index_q[3]), .C(index_q[4]), 
         .D(n24959), .Z(n20684)) /* synthesis lut_function=(!(A (B (C)+!B ((D)+!C))+!A (B+((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18354_3_lut_3_lut_4_lut_4_lut.init = 16'h0838;
    LUT4 i9441_3_lut_4_lut_4_lut (.A(n25097), .B(index_q[3]), .C(index_q[5]), 
         .D(n24957), .Z(n12007)) /* synthesis lut_function=(A (B+(C (D)))+!A (B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9441_3_lut_4_lut_4_lut.init = 16'hf8c8;
    LUT4 i19950_3_lut (.A(n21460), .B(n21461), .C(index_q[4]), .Z(n21462)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19950_3_lut.init = 16'hcaca;
    LUT4 n46_bdd_3_lut_21796_4_lut_4_lut (.A(n25097), .B(index_q[3]), .C(index_q[4]), 
         .D(n24980), .Z(n23055)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C))+!A !(B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n46_bdd_3_lut_21796_4_lut_4_lut.init = 16'h838f;
    PFUMX i17934 (.BLUT(n860_adj_2675), .ALUT(n891_adj_2672), .C0(index_q[5]), 
          .Z(n20264));
    LUT4 i19122_3_lut (.A(n25180), .B(n25200), .C(index_q[3]), .Z(n21452)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19122_3_lut.init = 16'hcaca;
    PFUMX i19150 (.BLUT(n21478), .ALUT(n21479), .C0(index_i[4]), .Z(n21480));
    LUT4 n62_bdd_3_lut_22596_4_lut (.A(n25097), .B(index_q[3]), .C(index_q[4]), 
         .D(n30_adj_2660), .Z(n23041)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n62_bdd_3_lut_22596_4_lut.init = 16'hf808;
    LUT4 i18594_3_lut (.A(n491_adj_2694), .B(n541), .C(index_i[4]), .Z(n20924)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18594_3_lut.init = 16'hcaca;
    LUT4 i18593_3_lut (.A(n397), .B(n475_adj_2695), .C(index_i[4]), .Z(n20923)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18593_3_lut.init = 16'hcaca;
    LUT4 i18591_3_lut (.A(n251_adj_2312), .B(n443), .C(index_i[4]), .Z(n20921)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18591_3_lut.init = 16'hcaca;
    LUT4 i18590_3_lut (.A(n397), .B(n14802), .C(index_i[4]), .Z(n20920)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;
    defparam i18590_3_lut.init = 16'h3a3a;
    LUT4 i18578_3_lut (.A(n236), .B(n251_adj_2312), .C(index_i[4]), .Z(n20908)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18578_3_lut.init = 16'hcaca;
    LUT4 i18577_3_lut (.A(n205_adj_2696), .B(n157_adj_2313), .C(index_i[4]), 
         .Z(n20907)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18577_3_lut.init = 16'hcaca;
    LUT4 i18877_3_lut_3_lut (.A(n25193), .B(index_q[3]), .C(n1001), .Z(n21207)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam i18877_3_lut_3_lut.init = 16'h7474;
    LUT4 i18574_3_lut (.A(n78), .B(n93_adj_2685), .C(index_i[4]), .Z(n20904)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18574_3_lut.init = 16'hcaca;
    LUT4 i18571_3_lut (.A(n157_adj_2313), .B(n30_adj_2480), .C(index_i[4]), 
         .Z(n20901)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18571_3_lut.init = 16'hcaca;
    LUT4 i18566_3_lut (.A(n747_adj_2306), .B(n762_adj_2337), .C(index_q[4]), 
         .Z(n20896)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18566_3_lut.init = 16'hcaca;
    LUT4 i18565_3_lut (.A(n716_adj_2601), .B(n14766), .C(index_q[4]), 
         .Z(n20895)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18565_3_lut.init = 16'hcaca;
    LUT4 i15273_3_lut (.A(n25074), .B(n25071), .C(index_i[3]), .Z(n17536)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15273_3_lut.init = 16'hcaca;
    LUT4 i19107_3_lut (.A(n27506), .B(n25207), .C(index_q[3]), .Z(n21437)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19107_3_lut.init = 16'hcaca;
    LUT4 i21102_2_lut (.A(index_i[4]), .B(index_i[3]), .Z(n19851)) /* synthesis lut_function=((B)+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i21102_2_lut.init = 16'hdddd;
    LUT4 i18556_3_lut (.A(n93_adj_2697), .B(n699_adj_2315), .C(index_q[4]), 
         .Z(n20886)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18556_3_lut.init = 16'hcaca;
    LUT4 i18555_3_lut (.A(n653_adj_2513), .B(n24840), .C(index_q[4]), 
         .Z(n20885)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18555_3_lut.init = 16'hcaca;
    LUT4 i19100_3_lut (.A(n25180), .B(n27494), .C(index_q[3]), .Z(n21430)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19100_3_lut.init = 16'hcaca;
    LUT4 i18549_3_lut (.A(n526_adj_2519), .B(n15_adj_2594), .C(index_q[4]), 
         .Z(n20879)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18549_3_lut.init = 16'hcaca;
    LUT4 i18546_3_lut (.A(n397_adj_2698), .B(n475_adj_2505), .C(index_q[4]), 
         .Z(n20876)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18546_3_lut.init = 16'hcaca;
    LUT4 i18544_3_lut (.A(n348_adj_2699), .B(n443_adj_2620), .C(index_q[4]), 
         .Z(n20874)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18544_3_lut.init = 16'hcaca;
    LUT4 i18543_3_lut (.A(n397_adj_2698), .B(n731_adj_2587), .C(index_q[4]), 
         .Z(n20873)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18543_3_lut.init = 16'hcaca;
    LUT4 i18541_3_lut (.A(n364_adj_2700), .B(n379_adj_2671), .C(index_q[4]), 
         .Z(n20871)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18541_3_lut.init = 16'hcaca;
    LUT4 i18540_3_lut (.A(n333_adj_2701), .B(n348_adj_2699), .C(index_q[4]), 
         .Z(n20870)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18540_3_lut.init = 16'hcaca;
    PFUMX i19356 (.BLUT(n844_adj_2613), .ALUT(n11930), .C0(index_q[4]), 
          .Z(n21686));
    LUT4 n380_bdd_4_lut (.A(n24871), .B(index_i[7]), .C(n25114), .D(index_i[5]), 
         .Z(n23185)) /* synthesis lut_function=(A (B+(C (D)+!C !(D)))+!A (B (D)+!B (C (D)+!C !(D)))) */ ;
    defparam n380_bdd_4_lut.init = 16'hfc8b;
    LUT4 i19960_3_lut (.A(n21427), .B(n21428), .C(index_q[4]), .Z(n21429)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19960_3_lut.init = 16'hcaca;
    LUT4 n953_bdd_3_lut_22183_4_lut_4_lut (.A(n25163), .B(n25166), .C(index_i[3]), 
         .D(index_i[2]), .Z(n23788)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B+(C))) */ ;
    defparam n953_bdd_3_lut_22183_4_lut_4_lut.init = 16'hfc5c;
    LUT4 mux_193_Mux_1_i317_3_lut (.A(n301), .B(n908_adj_2702), .C(index_q[4]), 
         .Z(n317_adj_2703)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_1_i317_3_lut.init = 16'hcaca;
    PFUMX i18740 (.BLUT(n21054), .ALUT(n21055), .C0(index_q[5]), .Z(n21070));
    LUT4 quarter_wave_sample_register_i_14__I_0_3_lut (.A(quarter_wave_sample_register_i[14]), 
         .B(o_val_pipeline_i_0__15__N_2157[14]), .C(phase_negation_i[1]), 
         .Z(o_val_pipeline_i_0__15__N_2158)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[14] 77[8])
    defparam quarter_wave_sample_register_i_14__I_0_3_lut.init = 16'hcaca;
    PFUMX i18741 (.BLUT(n21056), .ALUT(n21057), .C0(index_q[5]), .Z(n21071));
    LUT4 i19224_3_lut_4_lut_4_lut (.A(n25163), .B(n25065), .C(index_i[3]), 
         .D(index_i[2]), .Z(n21554)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B+(C))) */ ;
    defparam i19224_3_lut_4_lut_4_lut.init = 16'hfc5c;
    PFUMX i19436 (.BLUT(n844_adj_2704), .ALUT(n12135), .C0(index_i[4]), 
          .Z(n21766));
    L6MUX21 i18742 (.D0(n21058), .D1(n21059), .SD(index_q[5]), .Z(n21072));
    LUT4 i19088_3_lut (.A(n900), .B(n25200), .C(index_q[3]), .Z(n21418)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19088_3_lut.init = 16'hcaca;
    PFUMX i18743 (.BLUT(n21060), .ALUT(n21061), .C0(index_q[5]), .Z(n21073));
    LUT4 i11722_2_lut_3_lut_4_lut (.A(index_i[1]), .B(n25113), .C(index_i[5]), 
         .D(index_i[4]), .Z(n508_adj_2460)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;
    defparam i11722_2_lut_3_lut_4_lut.init = 16'hf080;
    LUT4 i19967_3_lut (.A(n25256), .B(n21416), .C(index_q[4]), .Z(n21417)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19967_3_lut.init = 16'hcaca;
    LUT4 i18508_3_lut (.A(n491_adj_2650), .B(n506_adj_2461), .C(index_q[4]), 
         .Z(n20838)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18508_3_lut.init = 16'hcaca;
    LUT4 i18507_3_lut (.A(n460_adj_2556), .B(n475_adj_2705), .C(index_q[4]), 
         .Z(n20837)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18507_3_lut.init = 16'hcaca;
    LUT4 i18505_3_lut (.A(n251_adj_2317), .B(n443_adj_2325), .C(index_q[4]), 
         .Z(n20835)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18505_3_lut.init = 16'hcaca;
    LUT4 i18504_3_lut (.A(n460_adj_2556), .B(n14766), .C(index_q[4]), 
         .Z(n20834)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;
    defparam i18504_3_lut.init = 16'h3a3a;
    LUT4 mux_192_Mux_3_i890_3_lut_4_lut (.A(n25040), .B(index_i[2]), .C(index_i[3]), 
         .D(n325_adj_2282), .Z(n890_adj_2706)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_3_i890_3_lut_4_lut.init = 16'h6f60;
    LUT4 n85_bdd_3_lut_22562_4_lut (.A(n25040), .B(index_i[2]), .C(index_i[3]), 
         .D(n25047), .Z(n23994)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n85_bdd_3_lut_22562_4_lut.init = 16'hf606;
    LUT4 mux_192_Mux_2_i189_3_lut_3_lut_4_lut (.A(index_i[1]), .B(n25113), 
         .C(n173_adj_2707), .D(index_i[4]), .Z(n189_adj_2423)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(C+(D)))) */ ;
    defparam mux_192_Mux_2_i189_3_lut_3_lut_4_lut.init = 16'h77f0;
    LUT4 i19077_3_lut (.A(n25088), .B(n325_adj_2282), .C(index_i[3]), 
         .Z(n21407)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19077_3_lut.init = 16'hcaca;
    LUT4 i19975_3_lut (.A(n21406), .B(n21407), .C(index_i[4]), .Z(n21408)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19975_3_lut.init = 16'hcaca;
    L6MUX21 i18745 (.D0(n21064), .D1(n21065), .SD(index_q[5]), .Z(n21075));
    L6MUX21 i18746 (.D0(n21066), .D1(n21067), .SD(index_q[5]), .Z(n21076));
    L6MUX21 i18747 (.D0(n21068), .D1(n21069), .SD(index_q[5]), .Z(n21077));
    PFUMX i17959 (.BLUT(n956), .ALUT(n17670), .C0(index_i[6]), .Z(n20289));
    LUT4 mux_192_Mux_4_i747_3_lut_4_lut (.A(n25073), .B(index_i[2]), .C(index_i[3]), 
         .D(n25088), .Z(n747_adj_2708)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_4_i747_3_lut_4_lut.init = 16'hf606;
    LUT4 i9517_3_lut_4_lut (.A(n25073), .B(index_i[2]), .C(n25114), .D(n25084), 
         .Z(n444_adj_2709)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9517_3_lut_4_lut.init = 16'h6f60;
    LUT4 i19073_3_lut (.A(n978), .B(n25083), .C(index_i[3]), .Z(n21403)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19073_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_4_i828_3_lut (.A(n812_adj_2287), .B(n827), .C(index_i[4]), 
         .Z(n828_adj_2710)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_4_i828_3_lut.init = 16'hcaca;
    LUT4 i19071_3_lut (.A(n723), .B(n325_adj_2282), .C(index_i[3]), .Z(n21401)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19071_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_6_i251_3_lut_4_lut (.A(n25073), .B(index_i[2]), .C(index_i[3]), 
         .D(n25084), .Z(n251_adj_2562)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_6_i251_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_192_Mux_0_i348_3_lut_4_lut (.A(n25040), .B(index_i[2]), .C(index_i[3]), 
         .D(n27499), .Z(n348_adj_2372)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_0_i348_3_lut_4_lut.init = 16'h6f60;
    LUT4 i18492_3_lut (.A(n236_adj_2564), .B(n251_adj_2317), .C(index_q[4]), 
         .Z(n20822)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18492_3_lut.init = 16'hcaca;
    LUT4 i18491_3_lut (.A(n205_adj_2711), .B(n15), .C(index_q[4]), .Z(n20821)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18491_3_lut.init = 16'hcaca;
    L6MUX21 i18802 (.D0(n21166), .D1(n17537), .SD(index_i[5]), .Z(n21132));
    LUT4 i19064_3_lut (.A(n27503), .B(n27499), .C(index_i[3]), .Z(n21394)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19064_3_lut.init = 16'hcaca;
    LUT4 i18488_3_lut (.A(n301_adj_2571), .B(n93_adj_2697), .C(index_q[4]), 
         .Z(n20818)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18488_3_lut.init = 16'hcaca;
    LUT4 i18485_3_lut (.A(n15), .B(n526_adj_2602), .C(index_q[4]), .Z(n20815)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18485_3_lut.init = 16'hcaca;
    LUT4 i19059_3_lut (.A(n25076), .B(n25079), .C(index_i[3]), .Z(n21389)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19059_3_lut.init = 16'hcaca;
    PFUMX i23031 (.BLUT(n25257), .ALUT(n25258), .C0(index_q[1]), .Z(n25259));
    PFUMX i18805 (.BLUT(n542_adj_2662), .ALUT(n573_adj_2712), .C0(index_i[5]), 
          .Z(n21135));
    LUT4 i19058_3_lut (.A(n25051), .B(n325_adj_2282), .C(index_i[3]), 
         .Z(n21388)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19058_3_lut.init = 16'hcaca;
    LUT4 i19985_3_lut (.A(n21388), .B(n21389), .C(index_i[4]), .Z(n21390)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19985_3_lut.init = 16'hcaca;
    PFUMX i18806 (.BLUT(n605), .ALUT(n636_adj_2713), .C0(index_i[5]), 
          .Z(n21136));
    LUT4 i18976_3_lut_4_lut (.A(n24870), .B(n24873), .C(index_q[5]), .D(index_q[6]), 
         .Z(n21306)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (B+((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18976_3_lut_4_lut.init = 16'hffc5;
    PFUMX i18807 (.BLUT(n669_adj_2659), .ALUT(n700_adj_2714), .C0(index_i[5]), 
          .Z(n21137));
    LUT4 i2_3_lut_4_lut (.A(index_i[3]), .B(index_i[4]), .C(index_i[5]), 
         .D(n25122), .Z(n17670)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i2_3_lut_4_lut.init = 16'hfffe;
    PFUMX i18808 (.BLUT(n732_adj_2715), .ALUT(n21193), .C0(index_i[5]), 
          .Z(n21138));
    LUT4 i19056_3_lut (.A(n25080), .B(n25077), .C(index_i[3]), .Z(n21386)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19056_3_lut.init = 16'hcaca;
    PFUMX i18809 (.BLUT(n797_adj_2657), .ALUT(n828_adj_2656), .C0(index_i[5]), 
          .Z(n21139));
    LUT4 i15272_3_lut (.A(n25071), .B(n25076), .C(index_i[3]), .Z(n17535)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15272_3_lut.init = 16'hcaca;
    PFUMX i18810 (.BLUT(n860_adj_2440), .ALUT(n891_adj_2655), .C0(index_i[5]), 
          .Z(n21140));
    LUT4 i19987_3_lut (.A(n21385), .B(n21386), .C(index_i[4]), .Z(n21387)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19987_3_lut.init = 16'hcaca;
    PFUMX i17968 (.BLUT(n94_adj_2652), .ALUT(n21196), .C0(index_q[5]), 
          .Z(n20298));
    LUT4 mux_192_Mux_4_i158_3_lut (.A(n142_adj_2716), .B(n157_adj_2554), 
         .C(index_i[4]), .Z(n158_adj_2595)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_4_i158_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_8_i491_3_lut_3_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n491_adj_2694)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_8_i491_3_lut_3_lut_3_lut_4_lut.init = 16'h7870;
    PFUMX i17970 (.BLUT(n221_adj_2717), .ALUT(n252_adj_2718), .C0(index_q[5]), 
          .Z(n20300));
    LUT4 i19996_3_lut (.A(n21382), .B(n21383), .C(index_i[4]), .Z(n21384)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19996_3_lut.init = 16'hcaca;
    LUT4 i18844_3_lut_4_lut (.A(n24871), .B(n24872), .C(index_i[5]), .D(index_i[6]), 
         .Z(n21174)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (B+((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18844_3_lut_4_lut.init = 16'hffc5;
    LUT4 i19046_3_lut (.A(n404), .B(n25173), .C(index_q[3]), .Z(n21376)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19046_3_lut.init = 16'hcaca;
    LUT4 i20006_3_lut (.A(n21376), .B(n21377), .C(index_q[4]), .Z(n21378)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20006_3_lut.init = 16'hcaca;
    PFUMX i17971 (.BLUT(n286_adj_2649), .ALUT(n21199), .C0(index_q[5]), 
          .Z(n20301));
    LUT4 i19041_3_lut (.A(n404), .B(n27526), .C(index_q[3]), .Z(n21371)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19041_3_lut.init = 16'hcaca;
    LUT4 i20015_3_lut (.A(n21367), .B(n21368), .C(index_q[4]), .Z(n21369)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20015_3_lut.init = 16'hcaca;
    LUT4 i19035_3_lut (.A(n27526), .B(n25190), .C(index_q[3]), .Z(n21365)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19035_3_lut.init = 16'hcaca;
    LUT4 i19011_3_lut_4_lut (.A(n25031), .B(index_i[1]), .C(index_i[3]), 
         .D(n498), .Z(n21341)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19011_3_lut_4_lut.init = 16'hdfd0;
    PFUMX i17972 (.BLUT(n349_adj_2719), .ALUT(n21202), .C0(index_q[5]), 
          .Z(n20302));
    L6MUX21 i22537 (.D0(n24173), .D1(n24171), .SD(index_q[5]), .Z(n24174));
    LUT4 i20020_3_lut (.A(n21364), .B(n21365), .C(index_q[4]), .Z(n21366)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20020_3_lut.init = 16'hcaca;
    LUT4 i21104_2_lut (.A(index_q[4]), .B(index_q[3]), .Z(n19847)) /* synthesis lut_function=((B)+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21104_2_lut.init = 16'hdddd;
    LUT4 mux_192_Mux_0_i173_3_lut_4_lut (.A(n25031), .B(index_i[1]), .C(index_i[3]), 
         .D(n25076), .Z(n173_adj_2369)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_0_i173_3_lut_4_lut.init = 16'hdfd0;
    LUT4 mux_193_Mux_7_i333_3_lut (.A(n25193), .B(n25156), .C(index_q[3]), 
         .Z(n333_adj_2701)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_7_i333_3_lut.init = 16'hcaca;
    PFUMX mux_192_Mux_8_i764 (.BLUT(n716_adj_2720), .ALUT(n732_adj_2641), 
          .C0(n19835), .Z(n764_adj_2328)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 mux_192_Mux_1_i620_3_lut_4_lut (.A(n25031), .B(index_i[1]), .C(index_i[3]), 
         .D(n25066), .Z(n620_adj_2275)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_1_i620_3_lut_4_lut.init = 16'hdfd0;
    PFUMX i22535 (.BLUT(n572_adj_2624), .ALUT(n24172), .C0(index_q[4]), 
          .Z(n24173));
    LUT4 i20023_3_lut (.A(n21361), .B(n21362), .C(index_q[4]), .Z(n21363)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20023_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_7_i348_3_lut (.A(n25194), .B(n27521), .C(index_q[3]), 
         .Z(n348_adj_2699)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_7_i348_3_lut.init = 16'hcaca;
    PFUMX mux_192_Mux_8_i574 (.BLUT(n542), .ALUT(n12046), .C0(index_i[5]), 
          .Z(n574)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 mux_193_Mux_11_i638_4_lut_4_lut (.A(n24828), .B(index_q[5]), .C(index_q[6]), 
         .D(n24856), .Z(n638_adj_2368)) /* synthesis lut_function=(A (B (C (D))+!B !(C))+!A (B ((D)+!C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_11_i638_4_lut_4_lut.init = 16'hc707;
    LUT4 n23057_bdd_3_lut_23867 (.A(n23057), .B(n23062), .C(index_q[7]), 
         .Z(n24402)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n23057_bdd_3_lut_23867.init = 16'hcaca;
    LUT4 mux_193_Mux_7_i397_3_lut (.A(n25194), .B(n25193), .C(index_q[3]), 
         .Z(n397_adj_2698)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_7_i397_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_6_i731_3_lut (.A(n25196), .B(n25160), .C(index_q[3]), 
         .Z(n731_adj_2587)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_6_i731_3_lut.init = 16'hcaca;
    LUT4 i19025_3_lut (.A(n25079), .B(n27498), .C(index_i[3]), .Z(n21355)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19025_3_lut.init = 16'hcaca;
    LUT4 n20688_bdd_3_lut_22712 (.A(n20688), .B(n20695), .C(index_q[7]), 
         .Z(n24404)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n20688_bdd_3_lut_22712.init = 16'hcaca;
    LUT4 mux_192_Mux_5_i700_3_lut (.A(n460_adj_2559), .B(n25082), .C(index_i[4]), 
         .Z(n700_adj_2721)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_5_i700_3_lut.init = 16'hcaca;
    LUT4 n20688_bdd_3_lut (.A(n23043), .B(n26781), .C(index_q[7]), .Z(n24405)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n20688_bdd_3_lut.init = 16'hcaca;
    PFUMX i22532 (.BLUT(n24170), .ALUT(n24169), .C0(index_q[4]), .Z(n24171));
    LUT4 i19019_3_lut (.A(n325_adj_2282), .B(n27498), .C(index_i[3]), 
         .Z(n21349)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19019_3_lut.init = 16'hcaca;
    LUT4 i19017_3_lut (.A(n25071), .B(n25088), .C(index_i[3]), .Z(n21347)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19017_3_lut.init = 16'hcaca;
    LUT4 i19016_3_lut (.A(n25065), .B(n25087), .C(index_i[3]), .Z(n21346)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19016_3_lut.init = 16'hcaca;
    LUT4 i19014_3_lut (.A(n27496), .B(n25087), .C(index_i[3]), .Z(n21344)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19014_3_lut.init = 16'hcaca;
    LUT4 i19010_3_lut (.A(n25079), .B(n25087), .C(index_i[3]), .Z(n21340)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19010_3_lut.init = 16'hcaca;
    PFUMX i17977 (.BLUT(n669_adj_2633), .ALUT(n700_adj_2630), .C0(index_q[5]), 
          .Z(n20307));
    PFUMX i17978 (.BLUT(n21214), .ALUT(n763_adj_2453), .C0(index_q[5]), 
          .Z(n20308));
    LUT4 i9505_3_lut_4_lut (.A(n24980), .B(index_q[4]), .C(index_q[3]), 
         .D(n25211), .Z(n12071)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(C+(D)))) */ ;
    defparam i9505_3_lut_4_lut.init = 16'h7f70;
    PFUMX i17979 (.BLUT(n21217), .ALUT(n828_adj_2722), .C0(index_q[5]), 
          .Z(n20309));
    PFUMX i23029 (.BLUT(n25253), .ALUT(n25254), .C0(index_i[0]), .Z(n25255));
    LUT4 mux_192_Mux_7_i333_3_lut (.A(n25166), .B(n24941), .C(index_i[3]), 
         .Z(n333_adj_2693)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_7_i333_3_lut.init = 16'hcaca;
    PFUMX i17980 (.BLUT(n860_adj_2627), .ALUT(n21220), .C0(index_q[5]), 
          .Z(n20310));
    LUT4 mux_192_Mux_7_i348_3_lut (.A(n25165), .B(n27520), .C(index_i[3]), 
         .Z(n348_adj_2691)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_7_i348_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_7_i397_3_lut (.A(n25165), .B(n25166), .C(index_i[3]), 
         .Z(n397_adj_2689)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_7_i397_3_lut.init = 16'hcaca;
    LUT4 i9548_3_lut_4_lut (.A(n24947), .B(index_i[4]), .C(index_i[3]), 
         .D(n25122), .Z(n12114)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(C+(D)))) */ ;
    defparam i9548_3_lut_4_lut.init = 16'h7f70;
    LUT4 i18990_3_lut_4_lut_4_lut (.A(n24904), .B(index_q[4]), .C(index_q[5]), 
         .D(n24862), .Z(n21320)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A (B (C+(D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18990_3_lut_4_lut_4_lut.init = 16'h101c;
    LUT4 mux_193_Mux_10_i574_4_lut_4_lut (.A(n24875), .B(index_q[4]), .C(index_q[5]), 
         .D(n24857), .Z(n574_adj_2363)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_10_i574_4_lut_4_lut.init = 16'h1f1c;
    LUT4 mux_193_Mux_2_i908_3_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[0]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n908_adj_2702)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C)+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_2_i908_3_lut_4_lut_4_lut.init = 16'h5a51;
    PFUMX i17999 (.BLUT(n94_adj_2723), .ALUT(n125_adj_2625), .C0(index_q[5]), 
          .Z(n20329));
    LUT4 mux_193_Mux_6_i668_3_lut (.A(n108), .B(n25195), .C(index_q[3]), 
         .Z(n668_adj_2580)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_6_i668_3_lut.init = 16'hcaca;
    PFUMX i18000 (.BLUT(n158_adj_2623), .ALUT(n189), .C0(index_q[5]), 
          .Z(n20330));
    LUT4 mux_193_Mux_6_i684_3_lut (.A(n25156), .B(n27522), .C(index_q[3]), 
         .Z(n684_adj_2724)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_6_i684_3_lut.init = 16'hcaca;
    L6MUX21 i22528 (.D0(n24164), .D1(n24161), .SD(index_q[4]), .Z(n24165));
    LUT4 mux_193_Mux_5_i15_3_lut (.A(n25205), .B(n27495), .C(index_q[3]), 
         .Z(n15_adj_2673)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_5_i15_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_0_i475_3_lut_4_lut (.A(n25033), .B(index_i[1]), .C(index_i[3]), 
         .D(n24947), .Z(n475_adj_2379)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_0_i475_3_lut_4_lut.init = 16'h4f40;
    LUT4 mux_192_Mux_3_i491_3_lut_4_lut (.A(n25033), .B(index_i[1]), .C(index_i[3]), 
         .D(n27518), .Z(n491_adj_2725)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_3_i491_3_lut_4_lut.init = 16'h4f40;
    LUT4 mux_193_Mux_6_i653_3_lut (.A(n25203), .B(n85_adj_2600), .C(index_q[3]), 
         .Z(n653_adj_2579)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_6_i653_3_lut.init = 16'hcaca;
    PFUMX mux_193_Mux_7_i190 (.BLUT(n21640), .ALUT(n173), .C0(index_q[5]), 
          .Z(n190)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 mux_193_Mux_5_i397_3_lut (.A(n25208), .B(n332), .C(index_q[3]), 
         .Z(n397_adj_2682)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_5_i397_3_lut.init = 16'hcaca;
    LUT4 i18862_3_lut_4_lut (.A(n25163), .B(index_i[2]), .C(index_i[3]), 
         .D(n25038), .Z(n21192)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;
    defparam i18862_3_lut_4_lut.init = 16'h6f60;
    LUT4 i18648_3_lut_4_lut_4_lut_4_lut (.A(n25163), .B(index_i[2]), .C(index_i[3]), 
         .D(index_i[4]), .Z(n20978)) /* synthesis lut_function=(A (B)+!A (B (C (D))+!B !(C (D)))) */ ;
    defparam i18648_3_lut_4_lut_4_lut_4_lut.init = 16'hc999;
    LUT4 mux_192_Mux_7_i475_3_lut_3_lut_4_lut (.A(n25163), .B(index_i[2]), 
         .C(n27520), .D(index_i[3]), .Z(n475_adj_2690)) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))+!A !(B ((D)+!C)+!B !(C+(D)))) */ ;
    defparam mux_192_Mux_7_i475_3_lut_3_lut_4_lut.init = 16'h99f0;
    LUT4 mux_192_Mux_0_i220_3_lut (.A(n25038), .B(n27518), .C(index_i[3]), 
         .Z(n220)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_0_i220_3_lut.init = 16'hcaca;
    PFUMX i22526 (.BLUT(n24163), .ALUT(n24162), .C0(index_q[5]), .Z(n24164));
    LUT4 mux_193_Mux_10_i637_3_lut_4_lut_4_lut (.A(n24921), .B(index_q[4]), 
         .C(index_q[5]), .D(n24875), .Z(n637_adj_2364)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_10_i637_3_lut_4_lut_4_lut.init = 16'h1f1c;
    LUT4 i11185_2_lut_rep_244_3_lut_4_lut (.A(n24877), .B(index_q[4]), .C(index_q[6]), 
         .D(index_q[5]), .Z(n24804)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11185_2_lut_rep_244_3_lut_4_lut.init = 16'hf080;
    LUT4 mux_193_Mux_5_i506_3_lut (.A(n25183), .B(n27506), .C(index_q[3]), 
         .Z(n506_adj_2626)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_5_i506_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_5_i859_3_lut (.A(n141_adj_2357), .B(n25205), .C(index_q[3]), 
         .Z(n859_adj_2674)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_5_i859_3_lut.init = 16'hcaca;
    CCU2D add_358_15 (.A0(quarter_wave_sample_register_q[14]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(\quarter_wave_sample_register_q[15] ), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17305), .S0(o_val_pipeline_q_0__15__N_2189[14]), 
          .S1(o_val_pipeline_q_0__15__N_2189[15]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(80[29:60])
    defparam add_358_15.INIT0 = 16'hf555;
    defparam add_358_15.INIT1 = 16'hf555;
    defparam add_358_15.INJECT1_0 = "NO";
    defparam add_358_15.INJECT1_1 = "NO";
    LUT4 mux_193_Mux_3_i221_3_lut_4_lut (.A(n24980), .B(index_q[3]), .C(index_q[4]), 
         .D(n24948), .Z(n221_adj_2726)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_3_i221_3_lut_4_lut.init = 16'h08f8;
    LUT4 mux_193_Mux_5_i875_3_lut (.A(n25156), .B(n25194), .C(index_q[3]), 
         .Z(n875_adj_2670)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_5_i875_3_lut.init = 16'hcaca;
    LUT4 i12111_3_lut (.A(index_q[3]), .B(index_q[1]), .C(index_q[0]), 
         .Z(n14799)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12111_3_lut.init = 16'hecec;
    PFUMX i18001 (.BLUT(n221_adj_2726), .ALUT(n252_adj_2352), .C0(index_q[5]), 
          .Z(n20331));
    LUT4 mux_192_Mux_2_i684_3_lut_4_lut (.A(n25163), .B(index_i[2]), .C(index_i[3]), 
         .D(n27499), .Z(n684_adj_2727)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;
    defparam mux_192_Mux_2_i684_3_lut_4_lut.init = 16'h6f60;
    LUT4 i12352_1_lut_2_lut_3_lut_4_lut (.A(n24877), .B(index_q[4]), .C(index_q[6]), 
         .D(index_q[5]), .Z(n382)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12352_1_lut_2_lut_3_lut_4_lut.init = 16'h0f7f;
    LUT4 mux_192_Mux_7_i653_3_lut_4_lut (.A(n25163), .B(index_i[2]), .C(index_i[3]), 
         .D(n25059), .Z(n653_adj_2687)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam mux_192_Mux_7_i653_3_lut_4_lut.init = 16'hf606;
    LUT4 n20313_bdd_3_lut_22751 (.A(n20315), .B(n23280), .C(index_q[7]), 
         .Z(n24450)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n20313_bdd_3_lut_22751.init = 16'hcaca;
    LUT4 i9519_3_lut_3_lut_4_lut (.A(index_i[3]), .B(index_i[4]), .C(n25083), 
         .D(index_i[0]), .Z(n605_adj_2728)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9519_3_lut_3_lut_4_lut.init = 16'h10fe;
    PFUMX i18002 (.BLUT(n286_adj_2622), .ALUT(n21229), .C0(index_q[5]), 
          .Z(n20332));
    LUT4 i18730_3_lut_4_lut (.A(n24980), .B(index_q[3]), .C(index_q[4]), 
         .D(n220_adj_2729), .Z(n21060)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18730_3_lut_4_lut.init = 16'hf808;
    PFUMX i22524 (.BLUT(n24160), .ALUT(n24159), .C0(index_q[5]), .Z(n24161));
    LUT4 i18650_4_lut_4_lut_4_lut (.A(n25163), .B(index_i[2]), .C(index_i[4]), 
         .D(index_i[3]), .Z(n20980)) /* synthesis lut_function=(A (B)+!A !(B (C+(D))+!B !(C+(D)))) */ ;
    defparam i18650_4_lut_4_lut_4_lut.init = 16'h999c;
    LUT4 index_i_0__bdd_4_lut_23045 (.A(index_i[0]), .B(index_i[3]), .C(index_i[1]), 
         .D(index_i[2]), .Z(n25226)) /* synthesis lut_function=(A (B (C)+!B !(C+!(D)))+!A !(B ((D)+!C)+!B !(C (D)+!C !(D)))) */ ;
    defparam index_i_0__bdd_4_lut_23045.init = 16'h92c1;
    PFUMX i18003 (.BLUT(n349_adj_2257), .ALUT(n21232), .C0(index_q[5]), 
          .Z(n20333));
    LUT4 mux_193_Mux_0_i220_3_lut (.A(n25160), .B(n25199), .C(index_q[3]), 
         .Z(n220_adj_2729)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i220_3_lut.init = 16'hcaca;
    LUT4 i18725_3_lut_4_lut (.A(n24980), .B(index_q[3]), .C(index_q[4]), 
         .D(n46_adj_2730), .Z(n21055)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18725_3_lut_4_lut.init = 16'h8f80;
    LUT4 i18726_3_lut_3_lut_4_lut (.A(n24980), .B(index_q[3]), .C(n93_adj_2731), 
         .D(index_q[4]), .Z(n21056)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18726_3_lut_3_lut_4_lut.init = 16'hf077;
    LUT4 i18919_3_lut (.A(n25171), .B(n27503), .C(index_i[3]), .Z(n21249)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18919_3_lut.init = 16'hcaca;
    LUT4 n20324_bdd_3_lut (.A(n20317), .B(n20318), .C(index_q[7]), .Z(n24448)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n20324_bdd_3_lut.init = 16'hcaca;
    LUT4 n20313_bdd_3_lut (.A(n20313), .B(n20314), .C(index_q[7]), .Z(n24451)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n20313_bdd_3_lut.init = 16'hcaca;
    LUT4 i20029_3_lut (.A(n21248), .B(n21249), .C(index_i[4]), .Z(n21250)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20029_3_lut.init = 16'hcaca;
    LUT4 i18913_3_lut (.A(n325), .B(n25200), .C(index_q[3]), .Z(n21243)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18913_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_6_i653_3_lut (.A(n25169), .B(n85), .C(index_i[3]), 
         .Z(n653_adj_2567)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_6_i653_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_6_i668_3_lut (.A(n108_adj_2732), .B(n25168), .C(index_i[3]), 
         .Z(n668_adj_2658)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_6_i668_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_6_i684_3_lut (.A(n24941), .B(n27503), .C(index_i[3]), 
         .Z(n684_adj_2733)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_6_i684_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_8_i93_3_lut_3_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[0]), .D(index_q[3]), .Z(n93_adj_2697)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(D))+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_8_i93_3_lut_3_lut_4_lut.init = 16'h3391;
    PFUMX mux_193_Mux_8_i764 (.BLUT(n716_adj_2734), .ALUT(n732_adj_2616), 
          .C0(n19824), .Z(n764_adj_2356)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 i20067_3_lut (.A(n21242), .B(n21243), .C(index_q[4]), .Z(n21244)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20067_3_lut.init = 16'hcaca;
    LUT4 i18910_3_lut (.A(n25198), .B(n27525), .C(index_q[3]), .Z(n21240)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18910_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_4_i61_3_lut (.A(n25180), .B(n25201), .C(index_q[3]), 
         .Z(n61_adj_2523)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_4_i61_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_10_i637_3_lut_4_lut_4_lut (.A(n24920), .B(index_i[4]), 
         .C(index_i[5]), .D(n24883), .Z(n637)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B !(C+(D))))) */ ;
    defparam mux_192_Mux_10_i637_3_lut_4_lut_4_lut.init = 16'h1f1c;
    PFUMX i18004 (.BLUT(n413_adj_2615), .ALUT(n444_adj_2735), .C0(index_q[5]), 
          .Z(n20334));
    LUT4 mux_193_Mux_4_i270_3_lut (.A(n25206), .B(n25183), .C(index_q[3]), 
         .Z(n270_adj_2648)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_4_i270_3_lut.init = 16'hcaca;
    LUT4 i20086_3_lut (.A(n21236), .B(n21237), .C(index_q[4]), .Z(n21238)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20086_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_4_i15_3_lut (.A(n27506), .B(n588), .C(index_q[3]), 
         .Z(n15_adj_2525)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_4_i15_3_lut.init = 16'hcaca;
    PFUMX mux_193_Mux_8_i574 (.BLUT(n542_adj_2447), .ALUT(n12006), .C0(index_q[5]), 
          .Z(n574_adj_2355)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 mux_193_Mux_4_i348_3_lut (.A(n27507), .B(n25204), .C(index_q[3]), 
         .Z(n348_adj_2736)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_4_i348_3_lut.init = 16'hcaca;
    PFUMX i18005 (.BLUT(n476_adj_2609), .ALUT(n507_adj_2512), .C0(index_q[5]), 
          .Z(n20335));
    LUT4 i21116_2_lut (.A(index_i[5]), .B(index_i[4]), .Z(n19835)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i21116_2_lut.init = 16'heeee;
    LUT4 i18901_3_lut (.A(n27494), .B(n25183), .C(index_q[3]), .Z(n21231)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18901_3_lut.init = 16'hcaca;
    LUT4 i18900_3_lut (.A(n27523), .B(n25208), .C(index_q[3]), .Z(n21230)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18900_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_0_i908_3_lut_4_lut (.A(index_i[0]), .B(n25122), .C(index_i[3]), 
         .D(n27519), .Z(n908_adj_2265)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (C+!(D)))) */ ;
    defparam mux_192_Mux_0_i908_3_lut_4_lut.init = 16'h2f20;
    PFUMX i18006 (.BLUT(n21235), .ALUT(n573_adj_2599), .C0(index_q[5]), 
          .Z(n20336));
    LUT4 i20096_3_lut (.A(n21230), .B(n21231), .C(index_q[4]), .Z(n21232)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20096_3_lut.init = 16'hcaca;
    LUT4 i18898_3_lut (.A(n27522), .B(n25203), .C(index_q[3]), .Z(n21228)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18898_3_lut.init = 16'hcaca;
    LUT4 i18897_3_lut (.A(n25193), .B(n85_adj_2600), .C(index_q[3]), .Z(n21227)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18897_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_4_i684_3_lut (.A(n85_adj_2600), .B(n108), .C(index_q[3]), 
         .Z(n684_adj_2629)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_4_i684_3_lut.init = 16'hcaca;
    LUT4 i20098_3_lut (.A(n21227), .B(n21228), .C(index_q[4]), .Z(n21229)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20098_3_lut.init = 16'hcaca;
    LUT4 i18664_3_lut_3_lut_4_lut (.A(n24947), .B(index_i[3]), .C(n93_adj_2737), 
         .D(index_i[4]), .Z(n20994)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18664_3_lut_3_lut_4_lut.init = 16'hf077;
    PFUMX i18007 (.BLUT(n12071), .ALUT(n21238), .C0(index_q[5]), .Z(n20337));
    LUT4 n954_bdd_3_lut (.A(n954_adj_2508), .B(n173_adj_2738), .C(index_q[4]), 
         .Z(n23223)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n954_bdd_3_lut.init = 16'hacac;
    L6MUX21 i18922 (.D0(n21659), .D1(n21662), .SD(index_q[5]), .Z(n21252));
    LUT4 i18889_3_lut (.A(n27525), .B(n325), .C(index_q[3]), .Z(n21219)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18889_3_lut.init = 16'hcaca;
    LUT4 n25165_bdd_4_lut_23485 (.A(n25165), .B(index_i[6]), .C(index_i[4]), 
         .D(n25072), .Z(n25455)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A !(B (C+!(D))+!B !(D))) */ ;
    defparam n25165_bdd_4_lut_23485.init = 16'hbf80;
    LUT4 i20108_3_lut (.A(n21218), .B(n21219), .C(index_q[4]), .Z(n21220)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20108_3_lut.init = 16'hcaca;
    LUT4 i12120_3_lut (.A(index_q[3]), .B(index_q[1]), .C(index_q[0]), 
         .Z(n14811)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12120_3_lut.init = 16'hc8c8;
    LUT4 mux_193_Mux_3_i348_3_lut (.A(n25199), .B(n25200), .C(index_q[3]), 
         .Z(n348_adj_2256)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_3_i348_3_lut.init = 16'hcaca;
    LUT4 i18885_3_lut (.A(n588), .B(n25180), .C(index_q[3]), .Z(n21215)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18885_3_lut.init = 16'hcaca;
    L6MUX21 i18926 (.D0(n21675), .D1(n17530), .SD(index_q[5]), .Z(n21256));
    L6MUX21 i18927 (.D0(n21087), .D1(n12015), .SD(index_q[5]), .Z(n21257));
    LUT4 mux_193_Mux_4_i828_3_lut (.A(n812_adj_2489), .B(n236_adj_2666), 
         .C(index_q[4]), .Z(n828_adj_2722)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_4_i828_3_lut.init = 16'hcaca;
    LUT4 i18883_3_lut (.A(n900), .B(n325), .C(index_q[3]), .Z(n21213)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18883_3_lut.init = 16'hcaca;
    PFUMX i18008 (.BLUT(n669_adj_2593), .ALUT(n700_adj_2739), .C0(index_q[5]), 
          .Z(n20338));
    LUT4 mux_192_Mux_10_i574_4_lut_4_lut (.A(n24883), .B(index_i[4]), .C(index_i[5]), 
         .D(n24859), .Z(n574_adj_2362)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_10_i574_4_lut_4_lut.init = 16'h1f1c;
    LUT4 mux_192_Mux_3_i668_3_lut_4_lut (.A(n25050), .B(index_i[2]), .C(index_i[3]), 
         .D(n25076), .Z(n668_adj_2740)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_3_i668_3_lut_4_lut.init = 16'h6f60;
    LUT4 i18663_3_lut_4_lut (.A(n24947), .B(index_i[3]), .C(index_i[4]), 
         .D(n46_adj_2741), .Z(n20993)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18663_3_lut_4_lut.init = 16'h8f80;
    LUT4 n543_bdd_3_lut_22362_4_lut (.A(n25050), .B(index_i[2]), .C(n25082), 
         .D(index_i[5]), .Z(n23980)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(B (C+(D))+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n543_bdd_3_lut_22362_4_lut.init = 16'h66f0;
    LUT4 i21149_2_lut (.A(index_q[5]), .B(index_q[4]), .Z(n19824)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21149_2_lut.init = 16'heeee;
    PFUMX i23010 (.BLUT(n25220), .ALUT(n25221), .C0(index_q[1]), .Z(n25222));
    L6MUX21 i18009 (.D0(n21241), .D1(n763_adj_2397), .SD(index_q[5]), 
            .Z(n20339));
    PFUMX i18929 (.BLUT(n542_adj_2590), .ALUT(n573_adj_2605), .C0(index_q[5]), 
          .Z(n21259));
    LUT4 i18668_3_lut_4_lut (.A(n24947), .B(index_i[3]), .C(index_i[4]), 
         .D(n220), .Z(n20998)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18668_3_lut_4_lut.init = 16'hf808;
    LUT4 n277_bdd_3_lut_22306_4_lut (.A(n25050), .B(index_i[2]), .C(index_i[3]), 
         .D(n25080), .Z(n23913)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n277_bdd_3_lut_22306_4_lut.init = 16'hf606;
    LUT4 mux_192_Mux_4_i763_3_lut_4_lut (.A(n25050), .B(index_i[2]), .C(index_i[4]), 
         .D(n747_adj_2708), .Z(n763_adj_2742)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_4_i763_3_lut_4_lut.init = 16'h6f60;
    PFUMX i18010 (.BLUT(n797_adj_2589), .ALUT(n828), .C0(index_q[5]), 
          .Z(n20340));
    LUT4 n25165_bdd_3_lut_23147 (.A(n12174), .B(n12175), .C(index_i[2]), 
         .Z(n25456)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n25165_bdd_3_lut_23147.init = 16'hacac;
    LUT4 mux_192_Mux_3_i221_3_lut_4_lut (.A(n24947), .B(index_i[3]), .C(index_i[4]), 
         .D(n24945), .Z(n221_adj_2394)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_3_i221_3_lut_4_lut.init = 16'h08f8;
    LUT4 i18876_3_lut (.A(n27522), .B(n27495), .C(index_q[3]), .Z(n21206)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18876_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_7_i491_3_lut_4_lut (.A(n25054), .B(index_q[2]), .C(index_q[3]), 
         .D(n25160), .Z(n491_adj_2743)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_7_i491_3_lut_4_lut.init = 16'hf404;
    PFUMX i18930 (.BLUT(n605_adj_2744), .ALUT(n636), .C0(index_q[5]), 
          .Z(n21260));
    LUT4 i18958_3_lut_4_lut_4_lut (.A(n24922), .B(index_i[4]), .C(index_i[5]), 
         .D(n24861), .Z(n21288)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A (B (C+(D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18958_3_lut_4_lut_4_lut.init = 16'h101c;
    LUT4 mux_192_Mux_0_i731_3_lut_4_lut (.A(n25058), .B(index_i[2]), .C(index_i[3]), 
         .D(n25165), .Z(n731)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_0_i731_3_lut_4_lut.init = 16'h4f40;
    LUT4 i19221_3_lut_4_lut (.A(n25058), .B(index_i[2]), .C(index_i[3]), 
         .D(n25081), .Z(n21551)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19221_3_lut_4_lut.init = 16'hf404;
    PFUMX i18011 (.BLUT(n860_adj_2619), .ALUT(n891_adj_2584), .C0(index_q[5]), 
          .Z(n20341));
    LUT4 i2_3_lut_4_lut_adj_78 (.A(n24828), .B(index_q[5]), .C(index_q[8]), 
         .D(n25005), .Z(n19498)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i2_3_lut_4_lut_adj_78.init = 16'hfff8;
    LUT4 n25165_bdd_3_lut_23486 (.A(n25165), .B(n25168), .C(index_i[4]), 
         .Z(n25457)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n25165_bdd_3_lut_23486.init = 16'hacac;
    LUT4 i18835_3_lut (.A(n25076), .B(n25074), .C(index_i[3]), .Z(n21165)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18835_3_lut.init = 16'hcaca;
    LUT4 i18834_3_lut (.A(n325_adj_2282), .B(n204), .C(index_i[3]), .Z(n21164)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18834_3_lut.init = 16'hcaca;
    PFUMX i18931 (.BLUT(n669_adj_2581), .ALUT(n700_adj_2745), .C0(index_q[5]), 
          .Z(n21261));
    LUT4 mux_193_Mux_3_i908_3_lut (.A(n25177), .B(n25201), .C(index_q[3]), 
         .Z(n908_adj_2575)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_3_i908_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_7_i379_3_lut_3_lut (.A(n25193), .B(index_q[3]), .C(n27521), 
         .Z(n379_adj_2671)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam mux_193_Mux_7_i379_3_lut_3_lut.init = 16'h7474;
    LUT4 mux_193_Mux_0_i731_3_lut_4_lut (.A(n25054), .B(index_q[2]), .C(index_q[3]), 
         .D(n25194), .Z(n731_adj_2746)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i731_3_lut_4_lut.init = 16'h4f40;
    PFUMX i18932 (.BLUT(n732_adj_2747), .ALUT(n21093), .C0(index_q[5]), 
          .Z(n21262));
    PFUMX i18012 (.BLUT(n924_adj_2576), .ALUT(n21244), .C0(index_q[5]), 
          .Z(n20342));
    LUT4 mux_192_Mux_5_i397_3_lut (.A(n25071), .B(n204), .C(index_i[3]), 
         .Z(n397_adj_2561)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_5_i397_3_lut.init = 16'hcaca;
    PFUMX i18933 (.BLUT(n797_adj_2574), .ALUT(n828_adj_2573), .C0(index_q[5]), 
          .Z(n21263));
    LUT4 mux_193_Mux_7_i364_3_lut_3_lut (.A(n25193), .B(index_q[3]), .C(n25194), 
         .Z(n364_adj_2700)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;
    defparam mux_193_Mux_7_i364_3_lut_3_lut.init = 16'hd1d1;
    LUT4 mux_192_Mux_5_i506_3_lut (.A(n25077), .B(n27497), .C(index_i[3]), 
         .Z(n506_adj_2471)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_5_i506_3_lut.init = 16'hcaca;
    PFUMX i18013 (.BLUT(n21247), .ALUT(n1018_adj_2748), .C0(index_q[5]), 
          .Z(n20343));
    LUT4 mux_192_Mux_5_i15_3_lut (.A(n25072), .B(n27499), .C(index_i[3]), 
         .Z(n15_adj_2532)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_5_i15_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_4_i668_3_lut_3_lut (.A(n25193), .B(index_q[3]), .C(n27522), 
         .Z(n668_adj_2632)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;
    defparam mux_193_Mux_4_i668_3_lut_3_lut.init = 16'hd1d1;
    LUT4 mux_192_Mux_5_i859_3_lut (.A(n141), .B(n25072), .C(index_i[3]), 
         .Z(n859_adj_2546)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_5_i859_3_lut.init = 16'hcaca;
    LUT4 i15275_3_lut_4_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n17538)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C (D)+!C !(D)))+!A !(B (D)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i15275_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'h83fc;
    LUT4 mux_192_Mux_5_i875_3_lut (.A(n24941), .B(n25165), .C(index_i[3]), 
         .Z(n875_adj_2544)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_5_i875_3_lut.init = 16'hcaca;
    PFUMX i18934 (.BLUT(n860_adj_2455), .ALUT(n891_adj_2572), .C0(index_q[5]), 
          .Z(n21264));
    LUT4 i11389_3_lut (.A(index_i[3]), .B(index_i[1]), .C(index_i[0]), 
         .Z(n14064)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11389_3_lut.init = 16'hecec;
    LUT4 i11554_2_lut_rep_563 (.A(index_i[1]), .B(index_i[2]), .C(index_i[0]), 
         .Z(n25123)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11554_2_lut_rep_563.init = 16'h7070;
    LUT4 mux_193_Mux_4_i158_3_lut (.A(n142_adj_2749), .B(n157_adj_2486), 
         .C(index_q[4]), .Z(n158_adj_2442)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_4_i158_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_1_i924_3_lut (.A(n908_adj_2750), .B(n412), .C(index_i[4]), 
         .Z(n924_adj_2441)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_1_i924_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_2_i700_3_lut_4_lut (.A(index_i[1]), .B(n25057), .C(index_i[4]), 
         .D(n684_adj_2727), .Z(n700_adj_2433)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_2_i700_3_lut_4_lut.init = 16'hefe0;
    LUT4 mux_192_Mux_4_i15_3_lut (.A(n27497), .B(n978), .C(index_i[3]), 
         .Z(n15_adj_2483)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_4_i15_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_3_i1018_3_lut_4_lut (.A(index_i[1]), .B(n25057), .C(index_i[4]), 
         .D(n19673), .Z(n1018)) /* synthesis lut_function=(A (C+!(D))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_3_i1018_3_lut_4_lut.init = 16'he0ef;
    PFUMX i24574 (.BLUT(n27410), .ALUT(n27409), .C0(index_i[1]), .Z(n27411));
    LUT4 i19094_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[2]), .C(index_q[1]), 
         .D(index_q[3]), .Z(n21424)) /* synthesis lut_function=(!(A (B (D)+!B !(C+(D)))+!A !(B (D)+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19094_3_lut_4_lut_4_lut.init = 16'h66b9;
    LUT4 mux_192_Mux_4_i61_3_lut (.A(n25083), .B(n25069), .C(index_i[3]), 
         .Z(n61)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_4_i61_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_0_i1017_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .D(index_i[3]), .Z(n1017_adj_2272)) /* synthesis lut_function=(A (B (D)+!B !((D)+!C))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_0_i1017_4_lut_4_lut_4_lut.init = 16'hdd70;
    LUT4 i19197_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n21527)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (B (C+!(D))+!B (D))) */ ;
    defparam i19197_3_lut_4_lut_4_lut_4_lut.init = 16'hf1cc;
    LUT4 mux_193_Mux_0_i627_3_lut_rep_667 (.A(index_q[0]), .B(index_q[2]), 
         .C(index_q[1]), .Z(n27507)) /* synthesis lut_function=(A ((C)+!B)+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i627_3_lut_rep_667.init = 16'he6e6;
    PFUMX i24563 (.BLUT(n27395), .ALUT(n27394), .C0(index_q[1]), .Z(n27396));
    LUT4 i20458_3_lut (.A(n21544), .B(n21545), .C(index_i[4]), .Z(n21546)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20458_3_lut.init = 16'hcaca;
    PFUMX i18030 (.BLUT(n94_adj_2568), .ALUT(n125_adj_2566), .C0(index_i[5]), 
          .Z(n20360));
    LUT4 i18782_3_lut (.A(n25178), .B(n27494), .C(index_q[3]), .Z(n21112)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18782_3_lut.init = 16'hcaca;
    PFUMX i18031 (.BLUT(n17550), .ALUT(n14311), .C0(index_i[5]), .Z(n20361));
    L6MUX21 i18033 (.D0(n21342), .D1(n21345), .SD(index_i[5]), .Z(n20363));
    L6MUX21 i18034 (.D0(n21348), .D1(n21351), .SD(index_i[5]), .Z(n20364));
    PFUMX i18035 (.BLUT(n413_adj_2563), .ALUT(n444_adj_2709), .C0(index_i[5]), 
          .Z(n20365));
    LUT4 mux_192_Mux_6_i890_3_lut_3_lut_4_lut (.A(n25058), .B(index_i[2]), 
         .C(n25164), .D(index_i[3]), .Z(n890_adj_2654)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_6_i890_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 n476_bdd_3_lut_21820 (.A(n476_adj_2470), .B(n23275), .C(index_q[5]), 
         .Z(n23276)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n476_bdd_3_lut_21820.init = 16'hcaca;
    LUT4 mux_192_Mux_1_i349_3_lut (.A(n541), .B(n348_adj_2751), .C(index_i[4]), 
         .Z(n349_adj_2437)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_1_i349_3_lut.init = 16'hcaca;
    PFUMX i18036 (.BLUT(n476_adj_2560), .ALUT(n507_adj_2558), .C0(index_i[5]), 
          .Z(n20366));
    LUT4 i20467_3_lut (.A(n21520), .B(n21521), .C(index_i[4]), .Z(n21522)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20467_3_lut.init = 16'hcaca;
    PFUMX i18037 (.BLUT(n17540), .ALUT(n573_adj_2752), .C0(index_i[5]), 
          .Z(n20367));
    LUT4 mux_193_Mux_5_i700_3_lut (.A(n460_adj_2527), .B(n25202), .C(index_q[4]), 
         .Z(n700_adj_2692)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_5_i700_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_2_i270_3_lut (.A(n25205), .B(n25161), .C(index_q[3]), 
         .Z(n270_adj_2516)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_2_i270_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_1_i94_3_lut (.A(index_i[0]), .B(n93_adj_2753), .C(index_i[4]), 
         .Z(n94_adj_2436)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_1_i94_3_lut.init = 16'hcaca;
    LUT4 i18776_3_lut (.A(n325), .B(n27494), .C(index_q[3]), .Z(n21106)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18776_3_lut.init = 16'hcaca;
    LUT4 i18774_3_lut (.A(n25208), .B(n27525), .C(index_q[3]), .Z(n21104)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18774_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_2_i316_3_lut (.A(n25198), .B(n25180), .C(index_q[3]), 
         .Z(n316_adj_2514)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_2_i316_3_lut.init = 16'hcaca;
    LUT4 i18773_3_lut (.A(n25200), .B(n27523), .C(index_q[3]), .Z(n21103)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18773_3_lut.init = 16'hcaca;
    LUT4 i18771_3_lut (.A(n27526), .B(n27523), .C(index_q[3]), .Z(n21101)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18771_3_lut.init = 16'hcaca;
    LUT4 i18767_3_lut (.A(n25178), .B(n27523), .C(index_q[3]), .Z(n21097)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18767_3_lut.init = 16'hcaca;
    LUT4 i20481_3_lut (.A(n716_adj_2469), .B(n731_adj_2754), .C(index_i[4]), 
         .Z(n732_adj_2434)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20481_3_lut.init = 16'hcaca;
    LUT4 i18765_3_lut (.A(n25190), .B(n27522), .C(index_q[3]), .Z(n21095)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18765_3_lut.init = 16'hcaca;
    PFUMX i18038 (.BLUT(n605_adj_2728), .ALUT(n636_adj_2555), .C0(index_i[5]), 
          .Z(n20368));
    LUT4 i20196_3_lut (.A(n21094), .B(n21095), .C(index_q[4]), .Z(n21096)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20196_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_2_i669_3_lut (.A(n653_adj_2755), .B(n475_adj_2756), 
         .C(index_i[4]), .Z(n669_adj_2432)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_2_i669_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_3_i93_3_lut_4_lut (.A(n25058), .B(index_i[2]), .C(index_i[3]), 
         .D(n25059), .Z(n93)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_3_i93_3_lut_4_lut.init = 16'hefe0;
    LUT4 mux_192_Mux_2_i605_3_lut (.A(n142_adj_2411), .B(n604_adj_2757), 
         .C(index_i[4]), .Z(n605_adj_2431)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_2_i605_3_lut.init = 16'hcaca;
    LUT4 i20069_3_lut (.A(n21091), .B(n21092), .C(index_q[4]), .Z(n21093)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20069_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_2_i397_3_lut (.A(n27522), .B(n25196), .C(index_q[3]), 
         .Z(n397_adj_2507)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_2_i397_3_lut.init = 16'hcaca;
    LUT4 i20486_3_lut (.A(n25280), .B(n21503), .C(index_i[4]), .Z(n21504)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20486_3_lut.init = 16'hcaca;
    PFUMX i18039 (.BLUT(n21354), .ALUT(n700_adj_2721), .C0(index_i[5]), 
          .Z(n20369));
    LUT4 i20488_3_lut (.A(n21499), .B(n21500), .C(index_i[4]), .Z(n21501)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20488_3_lut.init = 16'hcaca;
    L6MUX21 i18040 (.D0(n732_adj_2359), .D1(n21357), .SD(index_i[5]), 
            .Z(n20370));
    LUT4 mux_192_Mux_2_i413_3_lut (.A(n397_adj_2646), .B(n954_adj_2758), 
         .C(index_i[4]), .Z(n413_adj_2428)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_2_i413_3_lut.init = 16'hcaca;
    PFUMX i18041 (.BLUT(n797_adj_2552), .ALUT(n828_adj_2759), .C0(index_i[5]), 
          .Z(n20371));
    LUT4 mux_192_Mux_2_i317_3_lut (.A(n668_adj_2740), .B(n316_adj_2644), 
         .C(index_i[4]), .Z(n317_adj_2426)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_2_i317_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_2_i286_3_lut (.A(n270_adj_2643), .B(n653_adj_2366), 
         .C(index_i[4]), .Z(n286_adj_2425)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_2_i286_3_lut.init = 16'hcaca;
    LUT4 i9577_3_lut_4_lut (.A(n25058), .B(index_i[2]), .C(index_i[5]), 
         .D(n25059), .Z(n12145)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9577_3_lut_4_lut.init = 16'hfe0e;
    LUT4 i18756_3_lut (.A(n404), .B(n25184), .C(index_q[3]), .Z(n21086)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18756_3_lut.init = 16'hcaca;
    LUT4 i18755_3_lut (.A(n25204), .B(n325), .C(index_q[3]), .Z(n21085)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18755_3_lut.init = 16'hcaca;
    LUT4 i20497_3_lut (.A(n142_adj_2465), .B(n14105), .C(index_i[4]), 
         .Z(n158_adj_2422)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20497_3_lut.init = 16'hcaca;
    LUT4 i20499_3_lut (.A(n21484), .B(n25278), .C(index_i[4]), .Z(n21486)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20499_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_3_i924_3_lut (.A(n908_adj_2638), .B(index_i[0]), .C(index_i[4]), 
         .Z(n924_adj_2419)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_3_i924_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_3_i891_3_lut (.A(n541_adj_2661), .B(n890_adj_2706), 
         .C(index_i[4]), .Z(n891_adj_2418)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_3_i891_3_lut.init = 16'hcaca;
    LUT4 i11272_2_lut_3_lut_4_lut (.A(n25058), .B(index_i[2]), .C(index_i[5]), 
         .D(n25053), .Z(n764_adj_2285)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11272_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 mux_192_Mux_3_i797_3_lut (.A(n412_adj_2636), .B(n796_adj_2760), 
         .C(index_i[4]), .Z(n797)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_3_i797_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_4_i270_3_lut (.A(n25066), .B(n25077), .C(index_i[3]), 
         .Z(n270)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_4_i270_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_3_i796_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n796_adj_2588)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C))+!A (B (C+!(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_3_i796_3_lut_4_lut_4_lut_4_lut.init = 16'hf07c;
    LUT4 mux_192_Mux_4_i348_3_lut (.A(n25047), .B(n25076), .C(index_i[3]), 
         .Z(n348_adj_2761)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_4_i348_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_3_i669_3_lut (.A(n653_adj_2366), .B(n668_adj_2740), 
         .C(index_i[4]), .Z(n669)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_3_i669_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_0_i397_3_lut (.A(n27521), .B(n27525), .C(index_q[3]), 
         .Z(n397_adj_2410)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i397_3_lut.init = 16'hcaca;
    PFUMX i18042 (.BLUT(n860_adj_2547), .ALUT(n891_adj_2545), .C0(index_i[5]), 
          .Z(n20372));
    LUT4 mux_192_Mux_4_i684_3_lut (.A(n85), .B(n108_adj_2732), .C(index_i[3]), 
         .Z(n684_adj_2474)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_4_i684_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_0_i1002_3_lut_3_lut_4_lut (.A(n25058), .B(index_i[2]), 
         .C(n38), .D(index_i[3]), .Z(n1002_adj_2271)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_0_i1002_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 i20509_3_lut (.A(n21472), .B(n21473), .C(index_i[4]), .Z(n21474)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20509_3_lut.init = 16'hcaca;
    LUT4 i18146_3_lut (.A(n20468), .B(n20469), .C(index_q[7]), .Z(n20476)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18146_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_8_i475_3_lut_3_lut_4_lut (.A(n25058), .B(index_i[2]), 
         .C(n24969), .D(index_i[3]), .Z(n475_adj_2695)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_8_i475_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 mux_192_Mux_3_i476_3_lut (.A(n460_adj_2553), .B(n285_adj_2549), 
         .C(index_i[4]), .Z(n476_adj_2406)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_3_i476_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_3_i413_3_lut (.A(n397_adj_2762), .B(n25035), .C(index_i[4]), 
         .Z(n413_adj_2405)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_3_i413_3_lut.init = 16'hcaca;
    LUT4 i18139_3_lut (.A(n20454), .B(n24248), .C(index_q[6]), .Z(n20469)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18139_3_lut.init = 16'hcaca;
    LUT4 i18148_3_lut (.A(n20472), .B(n20473), .C(index_q[7]), .Z(n20478)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18148_3_lut.init = 16'hcaca;
    LUT4 i18142_3_lut (.A(n20460), .B(n20461), .C(index_q[6]), .Z(n20472)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18142_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_0_i285_3_lut (.A(n25189), .B(n27522), .C(index_q[3]), 
         .Z(n285_adj_2665)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i285_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_3_i286_4_lut (.A(n93), .B(index_i[2]), .C(index_i[4]), 
         .D(n14096), .Z(n286)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_3_i286_4_lut.init = 16'h3aca;
    L6MUX21 i22454 (.D0(n24077), .D1(n24074), .SD(index_q[5]), .Z(n24078));
    LUT4 mux_193_Mux_0_i188_3_lut (.A(n25195), .B(n101_adj_2557), .C(index_q[3]), 
         .Z(n188_adj_2402)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i188_3_lut.init = 16'hcaca;
    LUT4 i18239_3_lut (.A(n20561), .B(n20562), .C(index_i[7]), .Z(n20569)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18239_3_lut.init = 16'hcaca;
    LUT4 i18232_3_lut (.A(n20547), .B(n23650), .C(index_i[6]), .Z(n20562)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18232_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_7_i890_3_lut_3_lut_4_lut (.A(n25058), .B(index_i[2]), 
         .C(n24970), .D(index_i[3]), .Z(n890_adj_2389)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_7_i890_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 i20156_3_lut (.A(n23611), .B(n124_adj_2376), .C(index_q[4]), 
         .Z(n21057)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20156_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_9_i124_3_lut_3_lut_4_lut (.A(n25058), .B(index_i[2]), 
         .C(n24969), .D(index_i[3]), .Z(n124_adj_2642)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_9_i124_3_lut_3_lut_4_lut.init = 16'h11f0;
    LUT4 i18241_3_lut (.A(n20565), .B(n20566), .C(index_i[7]), .Z(n20571)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18241_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_3_i747_3_lut (.A(n25178), .B(n404), .C(index_q[3]), 
         .Z(n747_adj_2396)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_3_i747_3_lut.init = 16'hcaca;
    LUT4 i18235_3_lut (.A(n23656), .B(n20554), .C(index_i[6]), .Z(n20565)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18235_3_lut.init = 16'hcaca;
    PFUMX i21552 (.BLUT(n23094), .ALUT(n23093), .C0(index_i[5]), .Z(n23095));
    PFUMX i22452 (.BLUT(n24076), .ALUT(n475_adj_2375), .C0(index_q[4]), 
          .Z(n24077));
    LUT4 mux_193_Mux_1_i986_3_lut (.A(n25194), .B(n25199), .C(index_q[3]), 
         .Z(n986_adj_2763)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_1_i986_3_lut.init = 16'hcaca;
    LUT4 i18608_3_lut (.A(n20931), .B(n20932), .C(index_q[7]), .Z(n20938)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18608_3_lut.init = 16'hcaca;
    LUT4 i18601_3_lut (.A(n20869), .B(n20872), .C(index_q[6]), .Z(n20931)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18601_3_lut.init = 16'hcaca;
    PFUMX i22449 (.BLUT(n24073), .ALUT(n24072), .C0(index_q[4]), .Z(n24074));
    LUT4 n25453_bdd_3_lut_23482 (.A(n25453), .B(n25452), .C(index_i[6]), 
         .Z(n25454)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n25453_bdd_3_lut_23482.init = 16'hcaca;
    LUT4 i18610_3_lut (.A(n22878), .B(n20936), .C(index_q[7]), .Z(n20940)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18610_3_lut.init = 16'hcaca;
    PFUMX i18215 (.BLUT(n12127), .ALUT(n62_adj_2764), .C0(index_i[5]), 
          .Z(n20545));
    LUT4 i17954_3_lut (.A(n20967), .B(n20970), .C(index_i[6]), .Z(n20284)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17954_3_lut.init = 16'hcaca;
    LUT4 i18179_3_lut (.A(n20503), .B(n20504), .C(index_i[7]), .Z(n20509)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18179_3_lut.init = 16'hcaca;
    LUT4 i18174_3_lut (.A(n20493), .B(n20494), .C(index_i[6]), .Z(n20504)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18174_3_lut.init = 16'hcaca;
    LUT4 i18208_3_lut (.A(n22938), .B(n20531), .C(index_i[7]), .Z(n20538)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18208_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_3_i158_3_lut (.A(n142_adj_2411), .B(n157_adj_2408), 
         .C(index_i[4]), .Z(n158)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_3_i158_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_3_i125_3_lut (.A(n46), .B(n30_adj_2480), .C(index_i[4]), 
         .Z(n125_adj_2393)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_3_i125_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_5_i924_4_lut_3_lut (.A(index_i[2]), .B(n14064), .C(index_i[4]), 
         .Z(n924)) /* synthesis lut_function=(!(A (B+(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_5_i924_4_lut_3_lut.init = 16'h5656;
    LUT4 i17914_3_lut (.A(n23068), .B(n26707), .C(index_i[7]), .Z(n20244)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17914_3_lut.init = 16'hcaca;
    LUT4 i18846_3_lut (.A(n21169), .B(n21170), .C(index_i[7]), .Z(n21176)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18846_3_lut.init = 16'hcaca;
    LUT4 i18839_3_lut (.A(n23811), .B(n20919), .C(index_i[6]), .Z(n21169)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18839_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_2_i700_3_lut_4_lut (.A(index_q[1]), .B(n25091), .C(index_q[4]), 
         .D(n684_adj_2518), .Z(n700_adj_2765)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_2_i700_3_lut_4_lut.init = 16'hefe0;
    LUT4 mux_193_Mux_3_i1018_3_lut_4_lut (.A(index_q[1]), .B(n25091), .C(index_q[4]), 
         .D(n19655), .Z(n1018_adj_2748)) /* synthesis lut_function=(A (C+!(D))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_3_i1018_3_lut_4_lut.init = 16'he0ef;
    LUT4 i18024_3_lut (.A(n20348), .B(n20349), .C(index_q[7]), .Z(n20354)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18024_3_lut.init = 16'hcaca;
    PFUMX i18153 (.BLUT(n31_adj_2540), .ALUT(n62), .C0(index_i[5]), .Z(n20483));
    LUT4 i18019_3_lut (.A(n20338), .B(n20339), .C(index_q[6]), .Z(n20349)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18019_3_lut.init = 16'hcaca;
    LUT4 n23436_bdd_3_lut (.A(n25216), .B(n444_adj_2766), .C(index_i[5]), 
         .Z(n23437)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n23436_bdd_3_lut.init = 16'hcaca;
    LUT4 i18978_3_lut (.A(n21301), .B(n21302), .C(index_q[7]), .Z(n21308)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18978_3_lut.init = 16'hcaca;
    LUT4 i18971_3_lut (.A(n23787), .B(n20833), .C(index_q[6]), .Z(n21301)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18971_3_lut.init = 16'hcaca;
    LUT4 i18084_3_lut (.A(n23400), .B(n20407), .C(index_q[7]), .Z(n20414)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18084_3_lut.init = 16'hcaca;
    LUT4 index_q_4__bdd_4_lut_21677 (.A(index_q[4]), .B(n24948), .C(index_q[7]), 
         .D(n24949), .Z(n22813)) /* synthesis lut_function=(A (C+!(D))+!A (B+!(C))) */ ;
    defparam index_q_4__bdd_4_lut_21677.init = 16'he5ef;
    PFUMX i18122 (.BLUT(n12110), .ALUT(n62_adj_2767), .C0(index_q[5]), 
          .Z(n20452));
    LUT4 n25041_bdd_4_lut (.A(n141), .B(index_i[5]), .C(index_i[4]), .D(n24941), 
         .Z(n25453)) /* synthesis lut_function=(A (B (D)+!B ((D)+!C))+!A (B (D)+!B (C (D)))) */ ;
    defparam n25041_bdd_4_lut.init = 16'hfe02;
    LUT4 mux_193_Mux_1_i732_3_lut (.A(n716_adj_2341), .B(n491_adj_2490), 
         .C(index_q[4]), .Z(n732_adj_2390)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_1_i732_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_6_i732_3_lut_4_lut (.A(n25193), .B(index_q[3]), .C(index_q[4]), 
         .D(n731_adj_2587), .Z(n732_adj_2747)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_6_i732_3_lut_4_lut.init = 16'hf909;
    LUT4 mux_193_Mux_6_i700_3_lut_4_lut (.A(n25193), .B(index_q[3]), .C(index_q[4]), 
         .D(n684_adj_2724), .Z(n700_adj_2745)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_6_i700_3_lut_4_lut.init = 16'h9f90;
    LUT4 i20526_3_lut (.A(n26765), .B(n23790), .C(index_i[5]), .Z(n20435)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20526_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_0_i526_3_lut (.A(n25076), .B(n25083), .C(index_i[3]), 
         .Z(n526)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_0_i526_3_lut.init = 16'hcaca;
    LUT4 i20530_3_lut (.A(n542_adj_2481), .B(n573_adj_2634), .C(index_i[5]), 
         .Z(n20429)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20530_3_lut.init = 16'hcaca;
    PFUMX i18091 (.BLUT(n31_adj_2538), .ALUT(n62_adj_2537), .C0(index_i[5]), 
          .Z(n20421));
    PFUMX i18029 (.BLUT(n31_adj_2534), .ALUT(n21250), .C0(index_i[5]), 
          .Z(n20359));
    LUT4 n23278_bdd_3_lut (.A(n25232), .B(n444_adj_2510), .C(index_q[5]), 
         .Z(n23279)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n23278_bdd_3_lut.init = 16'hcaca;
    LUT4 i20777_3_lut (.A(n20404), .B(n24174), .C(index_q[6]), .Z(n20413)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20777_3_lut.init = 16'hcaca;
    PFUMX i17998 (.BLUT(n31_adj_2530), .ALUT(n62_adj_2768), .C0(index_q[5]), 
          .Z(n20328));
    L6MUX21 i22434 (.D0(n24057), .D1(n24055), .SD(index_q[5]), .Z(n24058));
    LUT4 i20922_3_lut (.A(n20385), .B(n20386), .C(index_i[8]), .Z(n20388)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20922_3_lut.init = 16'hcaca;
    PFUMX i17967 (.BLUT(n31), .ALUT(n62_adj_2524), .C0(index_q[5]), .Z(n20297));
    LUT4 mux_192_Mux_0_i397_3_lut (.A(n27520), .B(n25088), .C(index_i[3]), 
         .Z(n397_adj_2374)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_0_i397_3_lut.init = 16'hcaca;
    LUT4 i11237_3_lut_4_lut (.A(index_q[4]), .B(n25096), .C(index_q[5]), 
         .D(n25188), .Z(n892_adj_2769)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11237_3_lut_4_lut.init = 16'hf8f0;
    LUT4 n25041_bdd_3_lut (.A(n25041), .B(n141), .C(index_i[4]), .Z(n25451)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n25041_bdd_3_lut.init = 16'hcaca;
    PFUMX i22432 (.BLUT(n24056), .ALUT(n285_adj_2608), .C0(index_q[4]), 
          .Z(n24057));
    LUT4 mux_193_Mux_10_i893_3_lut_4_lut (.A(n25095), .B(index_q[5]), .C(index_q[6]), 
         .D(n892_adj_2769), .Z(n893_adj_2420)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_10_i893_3_lut_4_lut.init = 16'hf101;
    LUT4 i18888_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[2]), .C(index_q[1]), 
         .D(index_q[3]), .Z(n21218)) /* synthesis lut_function=(A ((C (D))+!B)+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18888_3_lut_4_lut_4_lut.init = 16'he666;
    PFUMX i18062 (.BLUT(n158_adj_2521), .ALUT(n189_adj_2578), .C0(index_q[5]), 
          .Z(n20392));
    PFUMX i18063 (.BLUT(n221_adj_2770), .ALUT(n21363), .C0(index_q[5]), 
          .Z(n20393));
    LUT4 i18687_3_lut (.A(n21010), .B(n21011), .C(index_i[6]), .Z(n21017)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18687_3_lut.init = 16'hcaca;
    LUT4 i18688_3_lut (.A(n23862), .B(n21013), .C(index_i[6]), .Z(n21018)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18688_3_lut.init = 16'hcaca;
    LUT4 n612_bdd_3_lut (.A(n25205), .B(n25196), .C(index_q[3]), .Z(n24715)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n612_bdd_3_lut.init = 16'hcaca;
    PFUMX i18064 (.BLUT(n286_adj_2517), .ALUT(n317_adj_2515), .C0(index_q[5]), 
          .Z(n20394));
    LUT4 n612_bdd_3_lut_22946 (.A(n25194), .B(n141_adj_2357), .C(index_q[3]), 
         .Z(n24714)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n612_bdd_3_lut_22946.init = 16'hcaca;
    PFUMX i18065 (.BLUT(n349_adj_2771), .ALUT(n21366), .C0(index_q[5]), 
          .Z(n20395));
    LUT4 mux_193_Mux_12_i254_4_lut (.A(n24825), .B(n24853), .C(index_q[6]), 
         .D(n6_adj_2570), .Z(n254_adj_2371)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_12_i254_4_lut.init = 16'hca0a;
    LUT4 mux_192_Mux_12_i254_4_lut (.A(n24824), .B(n24854), .C(index_i[6]), 
         .D(n6), .Z(n254_adj_2370)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_12_i254_4_lut.init = 16'hca0a;
    LUT4 mux_193_Mux_9_i364_3_lut_3_lut_4_lut (.A(index_q[0]), .B(n25097), 
         .C(index_q[3]), .D(n24959), .Z(n364_adj_2353)) /* synthesis lut_function=(!(A (C (D))+!A (B (C (D))+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_9_i364_3_lut_3_lut_4_lut.init = 16'h0efe;
    LUT4 mux_192_Mux_0_i188_3_lut (.A(n25168), .B(n101), .C(index_i[3]), 
         .Z(n188)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_0_i188_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_0_i572_3_lut_4_lut (.A(index_q[0]), .B(n25097), .C(index_q[3]), 
         .D(n27523), .Z(n572_adj_2772)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i572_3_lut_4_lut.init = 16'hefe0;
    LUT4 i20192_3_lut (.A(n25226), .B(n124_adj_2773), .C(index_i[4]), 
         .Z(n20995)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20192_3_lut.init = 16'hcaca;
    LUT4 i9440_3_lut_4_lut (.A(index_q[0]), .B(n25097), .C(index_q[3]), 
         .D(index_q[4]), .Z(n12006)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9440_3_lut_4_lut.init = 16'h0e1e;
    LUT4 i20560_3_lut (.A(n286_adj_2774), .B(n317), .C(index_q[5]), .Z(n21317)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20560_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_5_i731_3_lut (.A(n27498), .B(n25088), .C(index_i[3]), 
         .Z(n731_adj_2358)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_5_i731_3_lut.init = 16'hcaca;
    PFUMX i22430 (.BLUT(n24054), .ALUT(n24053), .C0(index_q[4]), .Z(n24055));
    LUT4 mux_193_Mux_9_i124_3_lut_3_lut_4_lut (.A(index_q[0]), .B(n25097), 
         .C(index_q[3]), .D(n24980), .Z(n124_adj_2597)) /* synthesis lut_function=(!(A (C (D))+!A (B (C (D))+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_9_i124_3_lut_3_lut_4_lut.init = 16'h0efe;
    LUT4 n10509_bdd_3_lut_22969 (.A(n23092), .B(n23095), .C(index_i[4]), 
         .Z(n24732)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n10509_bdd_3_lut_22969.init = 16'hacac;
    LUT4 n46_bdd_3_lut_21512_3_lut_4_lut (.A(index_q[0]), .B(n25097), .C(index_q[4]), 
         .D(index_q[3]), .Z(n23054)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n46_bdd_3_lut_21512_3_lut_4_lut.init = 16'hf10f;
    LUT4 n24739_bdd_3_lut_24285 (.A(n24739), .B(n24732), .C(index_i[7]), 
         .Z(n24740)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n24739_bdd_3_lut_24285.init = 16'hcaca;
    LUT4 mux_193_Mux_3_i251_3_lut_4_lut (.A(index_q[0]), .B(n25097), .C(index_q[3]), 
         .D(n24959), .Z(n14996)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_3_i251_3_lut_4_lut.init = 16'hfe0e;
    LUT4 i11205_2_lut_rep_268_3_lut_4_lut (.A(index_q[0]), .B(n25097), .C(index_q[4]), 
         .D(index_q[3]), .Z(n24828)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11205_2_lut_rep_268_3_lut_4_lut.init = 16'hfef0;
    LUT4 i18510_4_lut_4_lut_3_lut_4_lut (.A(index_q[0]), .B(n25097), .C(index_q[4]), 
         .D(index_q[3]), .Z(n20840)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18510_4_lut_4_lut_3_lut_4_lut.init = 16'h11ef;
    L6MUX21 i21527 (.D0(n23067), .D1(n23065), .SD(index_i[6]), .Z(n23068));
    PFUMX i18066 (.BLUT(n413_adj_2509), .ALUT(n21369), .C0(index_q[5]), 
          .Z(n20396));
    LUT4 mux_193_Mux_8_i475_3_lut_3_lut_4_lut (.A(index_q[0]), .B(n25097), 
         .C(index_q[3]), .D(n24980), .Z(n475_adj_2705)) /* synthesis lut_function=(A (C+!(D))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_8_i475_3_lut_3_lut_4_lut.init = 16'he0ef;
    LUT4 mux_193_Mux_8_i653_3_lut_rep_257_3_lut_4_lut (.A(index_q[0]), .B(n25211), 
         .C(n24959), .D(index_q[3]), .Z(n24817)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(C+(D)))) */ ;
    defparam mux_193_Mux_8_i653_3_lut_rep_257_3_lut_4_lut.init = 16'h77f0;
    LUT4 index_i_0__bdd_4_lut_23047 (.A(index_i[0]), .B(index_i[3]), .C(index_i[1]), 
         .D(index_i[2]), .Z(n25278)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C))+!A (B (C (D)+!C !(D))+!B !(C+!(D))))) */ ;
    defparam index_i_0__bdd_4_lut_23047.init = 16'h16d3;
    LUT4 i20202_3_lut (.A(n620_adj_2775), .B(n14014), .C(index_i[4]), 
         .Z(n20981)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20202_3_lut.init = 16'hcaca;
    PFUMX i18067 (.BLUT(n21372), .ALUT(n507_adj_2776), .C0(index_q[5]), 
          .Z(n20397));
    PFUMX i18068 (.BLUT(n21375), .ALUT(n573_adj_2586), .C0(index_q[5]), 
          .Z(n20398));
    LUT4 i11208_3_lut_4_lut (.A(index_q[0]), .B(n25211), .C(n25090), .D(index_q[5]), 
         .Z(n318_adj_2367)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (C (D))) */ ;
    defparam i11208_3_lut_4_lut.init = 16'hf800;
    LUT4 n1018_bdd_4_lut_4_lut_4_lut_adj_79 (.A(index_q[0]), .B(n25211), 
         .C(index_q[4]), .D(index_q[3]), .Z(n23221)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (D))+!A (B (C (D)+!C !(D))+!B (D)))) */ ;
    defparam n1018_bdd_4_lut_4_lut_4_lut_adj_79.init = 16'h0c73;
    PFUMX i21525 (.BLUT(n23066), .ALUT(n62_adj_2348), .C0(index_i[5]), 
          .Z(n23067));
    LUT4 index_i_0__bdd_4_lut_23527 (.A(index_i[0]), .B(index_i[3]), .C(index_i[1]), 
         .D(index_i[2]), .Z(n25280)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C (D)))+!A !(B (C+!(D))+!B !(C+(D))))) */ ;
    defparam index_i_0__bdd_4_lut_23527.init = 16'h4ae7;
    LUT4 i18749_3_lut (.A(n21072), .B(n21073), .C(index_q[6]), .Z(n21079)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18749_3_lut.init = 16'hcaca;
    LUT4 i18750_3_lut (.A(n23963), .B(n21075), .C(index_q[6]), .Z(n21080)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18750_3_lut.init = 16'hcaca;
    LUT4 i17942_3_lut (.A(n20261), .B(n20262), .C(index_q[6]), .Z(n20272)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17942_3_lut.init = 16'hcaca;
    LUT4 i20205_3_lut (.A(n491_adj_2777), .B(n506), .C(index_i[4]), .Z(n20975)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20205_3_lut.init = 16'hcaca;
    PFUMX i23008 (.BLUT(n25217), .ALUT(n25218), .C0(index_i[0]), .Z(n25219));
    PFUMX i18069 (.BLUT(n605_adj_2502), .ALUT(n21378), .C0(index_q[5]), 
          .Z(n20399));
    LUT4 index_i_1__bdd_4_lut_23469 (.A(index_i[1]), .B(index_i[0]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n25282)) /* synthesis lut_function=(!(A (B (D)+!B (C+!(D)))+!A !(B (C (D)+!C !(D))+!B !((D)+!C)))) */ ;
    defparam index_i_1__bdd_4_lut_23469.init = 16'h429c;
    PFUMX i18070 (.BLUT(n669_adj_2498), .ALUT(n700_adj_2765), .C0(index_q[5]), 
          .Z(n20400));
    LUT4 i20583_3_lut (.A(n286_adj_2778), .B(n317_adj_2387), .C(index_i[5]), 
         .Z(n21285)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20583_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_9_i62_3_lut_4_lut_then_4_lut (.A(index_i[4]), .B(index_i[2]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n25285)) /* synthesis lut_function=(!(A (B (C+(D)))+!A (B+(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_9_i62_3_lut_4_lut_then_4_lut.init = 16'h222b;
    LUT4 index_q_6__bdd_4_lut_21761_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(n25091), .D(index_q[6]), .Z(n23059)) /* synthesis lut_function=(!(A (B (D)+!B (C (D)+!C !(D)))+!A (B (C (D))+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam index_q_6__bdd_4_lut_21761_4_lut.init = 16'h07fc;
    LUT4 mux_192_Mux_9_i62_3_lut_4_lut_else_4_lut (.A(index_i[4]), .B(index_i[2]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n25284)) /* synthesis lut_function=((B+(C (D)))+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_9_i62_3_lut_4_lut_else_4_lut.init = 16'hfddd;
    PFUMX i18071 (.BLUT(n732_adj_2496), .ALUT(n763_adj_2779), .C0(index_q[5]), 
          .Z(n20401));
    LUT4 n25458_bdd_3_lut (.A(n25458), .B(n25455), .C(index_i[5]), .Z(n25459)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n25458_bdd_3_lut.init = 16'hcaca;
    LUT4 i20585_3_lut (.A(n924_adj_2780), .B(n955), .C(index_q[5]), .Z(n21265)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20585_3_lut.init = 16'hcaca;
    LUT4 i18634_3_lut (.A(n141), .B(n25038), .C(index_i[3]), .Z(n20964)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18634_3_lut.init = 16'hcaca;
    LUT4 i18633_3_lut (.A(n85), .B(n25165), .C(index_i[3]), .Z(n20963)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18633_3_lut.init = 16'hcaca;
    LUT4 i18632_3_lut (.A(n27499), .B(n25166), .C(index_i[3]), .Z(n20962)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18632_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_6_i781_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), 
         .B(index_q[1]), .C(index_q[3]), .D(index_q[2]), .Z(n781_adj_2528)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A (B (C (D)+!C !(D))+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_6_i781_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hc837;
    LUT4 mux_193_Mux_8_i172_3_lut_rep_495 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n25055)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_8_i172_3_lut_rep_495.init = 16'h7c7c;
    PFUMX i24157 (.BLUT(n26779), .ALUT(n26778), .C0(index_q[3]), .Z(n26780));
    PFUMX i24154 (.BLUT(n26775), .ALUT(n26774), .C0(index_q[2]), .Z(n26776));
    LUT4 mux_193_Mux_0_i270_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n270_adj_2664)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C))+!A (B (C (D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i270_3_lut_3_lut_4_lut.init = 16'h0fc7;
    LUT4 mux_193_Mux_8_i205_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n205_adj_2711)) /* synthesis lut_function=(!(A (B (C)+!B !(C (D)+!C !(D)))+!A !(B ((D)+!C)+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_8_i205_3_lut_3_lut_4_lut.init = 16'h7c0f;
    LUT4 i11248_2_lut_rep_497 (.A(index_i[2]), .B(index_i[3]), .Z(n25057)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11248_2_lut_rep_497.init = 16'heeee;
    PFUMX i22421 (.BLUT(n24044), .ALUT(n24043), .C0(index_q[5]), .Z(n24045));
    L6MUX21 i18073 (.D0(n860_adj_2311), .D1(n891_adj_2305), .SD(index_q[5]), 
            .Z(n20403));
    PFUMX i21522 (.BLUT(n23064), .ALUT(n23063), .C0(index_i[5]), .Z(n23065));
    LUT4 mux_192_Mux_2_i908_3_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .D(index_i[3]), .Z(n908_adj_2289)) /* synthesis lut_function=(!(A (B+!(D))+!A !(B+!(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_2_i908_3_lut_4_lut_4_lut.init = 16'h6645;
    LUT4 mux_193_Mux_0_i443_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[0]), .D(index_q[3]), .Z(n443_adj_2413)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C (D))+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i443_3_lut_4_lut_4_lut_4_lut.init = 16'h0ed5;
    LUT4 i11552_2_lut_rep_386_3_lut (.A(index_i[2]), .B(index_i[3]), .C(index_i[1]), 
         .Z(n24946)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11552_2_lut_rep_386_3_lut.init = 16'hfefe;
    LUT4 i11374_2_lut_rep_498 (.A(index_i[0]), .B(index_i[1]), .Z(n25058)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11374_2_lut_rep_498.init = 16'h8888;
    LUT4 i11318_2_lut_rep_312_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[4]), .D(n25113), .Z(n24872)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11318_2_lut_rep_312_3_lut_4_lut.init = 16'hf8f0;
    LUT4 i11339_3_lut_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n14014)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (D))+!A (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11339_3_lut_3_lut_3_lut_4_lut.init = 16'h00f7;
    PFUMX i18092 (.BLUT(n94_adj_2487), .ALUT(n21384), .C0(index_i[5]), 
          .Z(n20422));
    LUT4 i11291_2_lut_rep_299_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n24859)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11291_2_lut_rep_299_3_lut_4_lut.init = 16'hf080;
    LUT4 i18631_3_lut (.A(n25038), .B(n27520), .C(index_i[3]), .Z(n20961)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18631_3_lut.init = 16'hcaca;
    LUT4 i11544_2_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(n25114), 
         .D(index_i[2]), .Z(n125_adj_2548)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11544_2_lut_3_lut_4_lut.init = 16'hf080;
    LUT4 mux_192_Mux_8_i635_3_lut_4_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n635_adj_2445)) /* synthesis lut_function=(!(A (B (C (D))+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_8_i635_3_lut_4_lut_3_lut_4_lut.init = 16'h0ff8;
    LUT4 i21405_then_3_lut (.A(index_i[0]), .B(index_i[4]), .C(index_i[3]), 
         .Z(n25291)) /* synthesis lut_function=(A (B)+!A (B (C)+!B !(C))) */ ;
    defparam i21405_then_3_lut.init = 16'hc9c9;
    LUT4 i11378_2_lut_2_lut_3_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .Z(n14053)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11378_2_lut_2_lut_3_lut.init = 16'h0808;
    LUT4 i1_2_lut_rep_294_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[4]), 
         .D(index_i[2]), .Z(n24854)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i1_2_lut_rep_294_3_lut_4_lut.init = 16'hf080;
    LUT4 mux_192_Mux_1_i348_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n348_adj_2751)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A (B ((D)+!C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_1_i348_3_lut_4_lut_4_lut_4_lut.init = 16'h38f0;
    LUT4 i21405_else_3_lut (.A(index_i[2]), .B(index_i[0]), .C(index_i[4]), 
         .D(index_i[3]), .Z(n25290)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)+!C !(D)))+!A (B (C+!(D))+!B !(C)))) */ ;
    defparam i21405_else_3_lut.init = 16'h1e38;
    LUT4 mux_193_Mux_8_i173_3_lut_3_lut_4_lut (.A(n25188), .B(index_q[2]), 
         .C(n25055), .D(index_q[3]), .Z(n173_adj_2738)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_8_i173_3_lut_3_lut_4_lut.init = 16'hf077;
    LUT4 mux_192_Mux_3_i796_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n796_adj_2760)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C))+!A (B (C+!(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_3_i796_3_lut_4_lut_4_lut_4_lut.init = 16'hf07c;
    LUT4 i18627_3_lut (.A(n25037), .B(n27520), .C(index_i[3]), .Z(n20957)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18627_3_lut.init = 16'hcaca;
    LUT4 i18626_3_lut (.A(n27499), .B(n108_adj_2732), .C(index_i[3]), 
         .Z(n20956)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18626_3_lut.init = 16'hcaca;
    LUT4 i18625_3_lut (.A(n85), .B(n25166), .C(index_i[3]), .Z(n20955)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18625_3_lut.init = 16'hcaca;
    LUT4 index_i_6__bdd_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(n25113), 
         .D(index_i[6]), .Z(n23094)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam index_i_6__bdd_3_lut_4_lut.init = 16'hf07f;
    PFUMX i24112 (.BLUT(n26705), .ALUT(n26704), .C0(index_i[3]), .Z(n26706));
    LUT4 mux_192_Mux_8_i526_3_lut_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n526_adj_2444)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_8_i526_3_lut_3_lut_3_lut_4_lut.init = 16'h0f70;
    PFUMX i24109 (.BLUT(n26701), .ALUT(n26700), .C0(index_i[2]), .Z(n26702));
    LUT4 index_i_6__bdd_4_lut_21700_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(n25057), .D(index_i[6]), .Z(n23093)) /* synthesis lut_function=(!(A (B (D)+!B (C (D)+!C !(D)))+!A (B (C (D))+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam index_i_6__bdd_4_lut_21700_4_lut.init = 16'h07fc;
    LUT4 i9579_3_lut_4_lut (.A(n25054), .B(index_q[2]), .C(index_q[5]), 
         .D(n25055), .Z(n12147)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9579_3_lut_4_lut.init = 16'hfe0e;
    LUT4 i2_2_lut_rep_482 (.A(index_q[1]), .B(index_q[3]), .Z(n25042)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i2_2_lut_rep_482.init = 16'heeee;
    LUT4 i20600_3_lut (.A(n26638), .B(n25295), .C(index_q[5]), .Z(n20311)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20600_3_lut.init = 16'hcaca;
    LUT4 i18624_3_lut (.A(n24941), .B(n25072), .C(index_i[3]), .Z(n20954)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18624_3_lut.init = 16'hcaca;
    LUT4 i11289_2_lut_rep_387_3_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .Z(n24947)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11289_2_lut_rep_387_3_lut.init = 16'hf8f8;
    LUT4 i20604_3_lut (.A(n542_adj_2637), .B(n573_adj_2592), .C(index_q[5]), 
         .Z(n20305)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20604_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_3_i1002_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n19673)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (D))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_3_i1002_3_lut_3_lut_4_lut.init = 16'hf708;
    LUT4 i19118_3_lut_3_lut_4_lut (.A(n25188), .B(index_q[2]), .C(n1001), 
         .D(index_q[3]), .Z(n21448)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19118_3_lut_3_lut_4_lut.init = 16'hf077;
    LUT4 mux_193_Mux_3_i93_3_lut_4_lut (.A(n25054), .B(index_q[2]), .C(index_q[3]), 
         .D(n25055), .Z(n93_adj_2621)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_3_i93_3_lut_4_lut.init = 16'hefe0;
    LUT4 i18620_3_lut (.A(n27520), .B(n25168), .C(index_i[3]), .Z(n20950)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18620_3_lut.init = 16'hcaca;
    LUT4 i11235_2_lut_3_lut_4_lut (.A(n25054), .B(index_q[2]), .C(index_q[5]), 
         .D(n25090), .Z(n764)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11235_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 mux_193_Mux_0_i1002_3_lut_3_lut_4_lut (.A(n25054), .B(index_q[2]), 
         .C(n1001), .D(index_q[3]), .Z(n1002)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i1002_3_lut_3_lut_4_lut.init = 16'hf011;
    PFUMX i18094 (.BLUT(n221_adj_2781), .ALUT(n252_adj_2782), .C0(index_i[5]), 
          .Z(n20424));
    LUT4 i22129_then_4_lut (.A(index_q[0]), .B(index_q[4]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n25294)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)+!C !(D))+!B (C (D)))) */ ;
    defparam i22129_then_4_lut.init = 16'hda0e;
    LUT4 mux_192_Mux_6_i812_3_lut_4_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n812_adj_2288)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(D))+!A !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_6_i812_3_lut_4_lut_3_lut_4_lut.init = 16'h7780;
    LUT4 i18619_3_lut (.A(n38), .B(n25037), .C(index_i[3]), .Z(n20949)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18619_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_7_i526_3_lut_3_lut_4_lut_4_lut_3_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n526_adj_2688)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(D))+!A !(D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_7_i526_3_lut_3_lut_4_lut_4_lut_3_lut_4_lut.init = 16'h887f;
    LUT4 i18583_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n20913)) /* synthesis lut_function=(A (B (C)+!B !(C (D)+!C !(D)))+!A !(B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18583_3_lut_4_lut_4_lut_4_lut.init = 16'h83f0;
    LUT4 i22129_else_4_lut (.A(index_q[0]), .B(index_q[4]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n25293)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C))+!A (B (C)+!B (C+(D)))) */ ;
    defparam i22129_else_4_lut.init = 16'hf178;
    LUT4 n123_bdd_3_lut_22962_3_lut_4_lut_4_lut_3_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n23646)) /* synthesis lut_function=(A (B (C)+!B !(D))+!A !(D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n123_bdd_3_lut_22962_3_lut_4_lut_4_lut_3_lut_4_lut.init = 16'h80f7;
    LUT4 i19214_3_lut_3_lut_4_lut (.A(n25163), .B(index_i[2]), .C(n38), 
         .D(index_i[3]), .Z(n21544)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19214_3_lut_3_lut_4_lut.init = 16'hf077;
    LUT4 i20619_3_lut (.A(n924_adj_2783), .B(n955_adj_2377), .C(index_i[5]), 
         .Z(n21141)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20619_3_lut.init = 16'hcaca;
    LUT4 i18617_3_lut (.A(n25168), .B(n24941), .C(index_i[3]), .Z(n20947)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18617_3_lut.init = 16'hcaca;
    PFUMX i18095 (.BLUT(n286_adj_2484), .ALUT(n21387), .C0(index_i[5]), 
          .Z(n20425));
    LUT4 i19200_3_lut_4_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n21530)) /* synthesis lut_function=(!(A (B (D)+!B !((D)+!C))+!A (B (C+(D))+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19200_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'h338f;
    LUT4 mux_192_Mux_8_i78_3_lut_4_lut (.A(n25163), .B(index_i[2]), .C(index_i[3]), 
         .D(n25059), .Z(n78)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_8_i78_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_192_Mux_8_i173_3_lut_3_lut_4_lut (.A(n25163), .B(index_i[2]), 
         .C(n25059), .D(index_i[3]), .Z(n173_adj_2784)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_8_i173_3_lut_3_lut_4_lut.init = 16'hf077;
    PFUMX i21519 (.BLUT(n23060), .ALUT(n23059), .C0(index_q[5]), .Z(n23061));
    LUT4 i11828_1_lut_2_lut (.A(index_q[1]), .B(index_q[3]), .Z(n541_adj_2262)) /* synthesis lut_function=(!(A+(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11828_1_lut_2_lut.init = 16'h1111;
    LUT4 i21130_2_lut_rep_301_2_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n24861)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i21130_2_lut_rep_301_2_lut_3_lut_4_lut.init = 16'h0007;
    LUT4 mux_192_Mux_6_i781_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n781_adj_2477)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A (B (C (D)+!C !(D))+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_6_i781_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hc837;
    LUT4 mux_193_Mux_9_i62_3_lut_4_lut_then_4_lut (.A(index_q[4]), .B(index_q[2]), 
         .C(index_q[1]), .D(index_q[0]), .Z(n25297)) /* synthesis lut_function=(!(A (B (C+(D)))+!A (B+(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_9_i62_3_lut_4_lut_then_4_lut.init = 16'h222b;
    LUT4 mux_193_Mux_9_i62_3_lut_4_lut_else_4_lut (.A(index_q[4]), .B(index_q[2]), 
         .C(index_q[1]), .D(index_q[0]), .Z(n25296)) /* synthesis lut_function=((B+(C (D)))+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_9_i62_3_lut_4_lut_else_4_lut.init = 16'hfddd;
    LUT4 i19205_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n21535)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A (B (C)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19205_3_lut_4_lut_4_lut.init = 16'h3c8c;
    L6MUX21 i21515 (.D0(n23056), .D1(n24798), .SD(index_q[6]), .Z(n23057));
    LUT4 mux_192_Mux_7_i315_3_lut_rep_478_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n25038)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_7_i315_3_lut_rep_478_3_lut.init = 16'h3838;
    PFUMX i18096 (.BLUT(n349_adj_2785), .ALUT(n21390), .C0(index_i[5]), 
          .Z(n20426));
    LUT4 mux_192_Mux_4_i1002_3_lut_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n1002_adj_2468)) /* synthesis lut_function=(A (B (C (D))+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_4_i1002_3_lut_3_lut_3_lut_4_lut.init = 16'hf007;
    LUT4 mux_192_Mux_7_i620_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n620_adj_2775)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A !(B (C+!(D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_7_i620_3_lut_4_lut_4_lut_4_lut.init = 16'h8c33;
    LUT4 mux_192_Mux_8_i93_3_lut_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n93_adj_2685)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (D))+!A (B ((D)+!C)+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_8_i93_3_lut_3_lut_4_lut_4_lut.init = 16'h08f3;
    LUT4 i19082_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n21412)) /* synthesis lut_function=(!(A (B (D)+!B !(D))+!A (B ((D)+!C)+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19082_3_lut_4_lut_4_lut_4_lut.init = 16'h33c8;
    LUT4 mux_192_Mux_7_i491_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n491_adj_2777)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(D))+!A (B (C+!(D))+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_7_i491_3_lut_4_lut_4_lut_4_lut.init = 16'h3780;
    LUT4 i11439_2_lut_rep_287_4_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n24847)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A (B+((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11439_2_lut_rep_287_4_lut_4_lut_4_lut_4_lut.init = 16'h0038;
    LUT4 mux_192_Mux_8_i70_3_lut_rep_499 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n25059)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_8_i70_3_lut_rep_499.init = 16'h7c7c;
    LUT4 n269_bdd_3_lut_22808_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n23860)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C))+!A (B (C (D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n269_bdd_3_lut_22808_3_lut_4_lut.init = 16'h0fc7;
    LUT4 mux_192_Mux_8_i205_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n205_adj_2696)) /* synthesis lut_function=(!(A (B (C)+!B !(C (D)+!C !(D)))+!A !(B ((D)+!C)+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_8_i205_3_lut_3_lut_4_lut.init = 16'h7c0f;
    PFUMX i21513 (.BLUT(n23055), .ALUT(n23054), .C0(index_q[5]), .Z(n23056));
    L6MUX21 i22399 (.D0(n24020), .D1(n24017), .SD(index_i[5]), .Z(n24021));
    PFUMX i22397 (.BLUT(n24019), .ALUT(n475_adj_2756), .C0(index_i[4]), 
          .Z(n24020));
    LUT4 i9578_3_lut_3_lut_4_lut (.A(n25163), .B(index_i[2]), .C(n157_adj_2313), 
         .D(index_i[4]), .Z(n12146)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9578_3_lut_3_lut_4_lut.init = 16'hf077;
    PFUMX i22394 (.BLUT(n24016), .ALUT(n24015), .C0(index_i[4]), .Z(n24017));
    LUT4 i21113_2_lut_rep_264_3_lut_4_lut (.A(n25163), .B(index_i[2]), .C(index_i[5]), 
         .D(n25053), .Z(n24824)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i21113_2_lut_rep_264_3_lut_4_lut.init = 16'h0f7f;
    L6MUX21 i22390 (.D0(n24013), .D1(n24011), .SD(index_i[5]), .Z(n24014));
    PFUMX i18101 (.BLUT(n669_adj_2478), .ALUT(n700_adj_2475), .C0(index_i[5]), 
          .Z(n20431));
    PFUMX i22388 (.BLUT(n21185), .ALUT(n24012), .C0(index_i[4]), .Z(n24013));
    PFUMX i18102 (.BLUT(n21402), .ALUT(n763_adj_2742), .C0(index_i[5]), 
          .Z(n20432));
    LUT4 i2_2_lut_rep_503 (.A(index_i[1]), .B(index_i[3]), .Z(n25063)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i2_2_lut_rep_503.init = 16'heeee;
    LUT4 i12128_1_lut_2_lut (.A(index_i[1]), .B(index_i[3]), .Z(n541_adj_2254)) /* synthesis lut_function=(!(A+(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i12128_1_lut_2_lut.init = 16'h1111;
    LUT4 mux_193_Mux_0_i316_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[3]), 
         .C(index_q[2]), .D(index_q[0]), .Z(n316_adj_2457)) /* synthesis lut_function=(!(A (B+(C))+!A !(B+(C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i316_3_lut_4_lut_4_lut_4_lut.init = 16'h5647;
    LUT4 i21000_2_lut_rep_504 (.A(index_i[0]), .B(index_i[1]), .Z(n25064)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i21000_2_lut_rep_504.init = 16'h9999;
    LUT4 i11471_2_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n668_adj_2260)) /* synthesis lut_function=(!(A ((D)+!B)+!A (B ((D)+!C)+!B (C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11471_2_lut_4_lut_4_lut_4_lut.init = 16'h00c9;
    LUT4 i9540_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(n25113), .D(index_i[4]), .Z(n189_adj_2596)) /* synthesis lut_function=(A (B (C (D)))+!A !(B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9540_3_lut_4_lut_4_lut_4_lut.init = 16'h9555;
    PFUMX i18103 (.BLUT(n21405), .ALUT(n828_adj_2710), .C0(index_i[5]), 
          .Z(n20433));
    PFUMX i22386 (.BLUT(n24010), .ALUT(n12177), .C0(n25113), .Z(n24011));
    L6MUX21 i22375 (.D0(n23997), .D1(n23995), .SD(index_i[5]), .Z(n23998));
    PFUMX i22373 (.BLUT(n23996), .ALUT(n285_adj_2549), .C0(index_i[4]), 
          .Z(n23997));
    PFUMX i22371 (.BLUT(n23994), .ALUT(n23993), .C0(index_i[4]), .Z(n23995));
    LUT4 i8416_2_lut_rep_568 (.A(index_i[4]), .B(index_i[5]), .Z(n25128)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i8416_2_lut_rep_568.init = 16'h8888;
    LUT4 i11575_3_lut_4_lut (.A(index_i[4]), .B(index_i[5]), .C(index_i[6]), 
         .D(index_i[3]), .Z(n509_adj_2252)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11575_3_lut_4_lut.init = 16'hf8f0;
    PFUMX i18104 (.BLUT(n860_adj_2472), .ALUT(n21408), .C0(index_i[5]), 
          .Z(n20434));
    PFUMX i22365 (.BLUT(n23988), .ALUT(n23987), .C0(index_i[5]), .Z(n23989));
    LUT4 mux_193_Mux_8_i301_3_lut_4_lut (.A(n25188), .B(index_q[2]), .C(index_q[3]), 
         .D(n25055), .Z(n301_adj_2571)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_8_i301_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_192_Mux_7_i45_3_lut_3_lut_rep_477_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n25037)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_7_i45_3_lut_3_lut_rep_477_3_lut.init = 16'h3939;
    LUT4 mux_192_Mux_5_i572_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n572_adj_2786)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A !(B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_5_i572_3_lut_4_lut_4_lut.init = 16'ha9a5;
    LUT4 i19202_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n21532)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !(B (C+!(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19202_3_lut_4_lut_4_lut.init = 16'ha5a9;
    LUT4 mux_192_Mux_5_i109_3_lut_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .Z(n109_adj_2565)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_5_i109_3_lut_3_lut_3_lut.init = 16'h3939;
    L6MUX21 i22360 (.D0(n23984), .D1(n23982), .SD(index_i[4]), .Z(n23985));
    LUT4 i11473_2_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n844_adj_2704)) /* synthesis lut_function=(A (B+!(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11473_2_lut_3_lut_4_lut.init = 16'h9ff9;
    PFUMX i22358 (.BLUT(n23983), .ALUT(n21158), .C0(index_i[5]), .Z(n23984));
    LUT4 mux_192_Mux_2_i604_3_lut_4_lut_4_lut_4_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n604_adj_2757)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)+!C !(D)))+!A (B (C)+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_2_i604_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'h3c9f;
    LUT4 mux_192_Mux_6_i573_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[4]), .D(n572_adj_2787), .Z(n573_adj_2712)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_6_i573_3_lut_4_lut.init = 16'hf909;
    L6MUX21 i23958 (.D0(n26502), .D1(n26498), .SD(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2126[7]));
    LUT4 i9604_3_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[4]), 
         .Z(n12174)) /* synthesis lut_function=(A (B)+!A !(B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9604_3_lut_4_lut_3_lut.init = 16'h9898;
    PFUMX i23956 (.BLUT(n26501), .ALUT(n26499), .C0(index_i[8]), .Z(n26502));
    PFUMX i22356 (.BLUT(n23981), .ALUT(n23980), .C0(index_i[3]), .Z(n23982));
    LUT4 mux_192_Mux_5_i251_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .Z(n251_adj_2551)) /* synthesis lut_function=(A (B)+!A (B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_5_i251_3_lut_3_lut.init = 16'hc9c9;
    PFUMX i23953 (.BLUT(n26497), .ALUT(n26496), .C0(index_i[8]), .Z(n26498));
    LUT4 mux_192_Mux_6_i498_3_lut_4_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n498)) /* synthesis lut_function=(A (B+!(C))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_6_i498_3_lut_4_lut_4_lut_3_lut.init = 16'h9b9b;
    PFUMX i22341 (.BLUT(n21062), .ALUT(n23962), .C0(index_q[5]), .Z(n23963));
    PFUMX i18123 (.BLUT(n94_adj_2464), .ALUT(n21417), .C0(index_q[5]), 
          .Z(n20453));
    PFUMX i22339 (.BLUT(n23960), .ALUT(n25017), .C0(index_q[3]), .Z(n23961));
    LUT4 mux_192_Mux_3_i347_3_lut_rep_505 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n25065)) /* synthesis lut_function=(A (B)+!A (B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_3_i347_3_lut_rep_505.init = 16'hc9c9;
    LUT4 mux_192_Mux_3_i396_3_lut_3_lut_rep_506 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n25066)) /* synthesis lut_function=(A (B+(C))+!A !(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_3_i396_3_lut_3_lut_rep_506.init = 16'ha9a9;
    LUT4 mux_192_Mux_6_i564_3_lut_4_lut_3_lut_rep_508 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n25068)) /* synthesis lut_function=(A (B)+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_6_i564_3_lut_4_lut_3_lut_rep_508.init = 16'hd9d9;
    LUT4 mux_192_Mux_5_i564_3_lut_rep_509 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n25069)) /* synthesis lut_function=(A (B (C))+!A !(B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_5_i564_3_lut_rep_509.init = 16'h9595;
    LUT4 mux_192_Mux_3_i676_3_lut_4_lut_3_lut_rep_510 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n25070)) /* synthesis lut_function=(A (B (C))+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_3_i676_3_lut_4_lut_3_lut_rep_510.init = 16'h9494;
    LUT4 mux_192_Mux_6_i356_3_lut_4_lut_3_lut_rep_511 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n25071)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_6_i356_3_lut_4_lut_3_lut_rep_511.init = 16'h4949;
    L6MUX21 i18124 (.D0(n21420), .D1(n21423), .SD(index_q[5]), .Z(n20454));
    LUT4 mux_192_Mux_7_i165_3_lut_3_lut_rep_512 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n25072)) /* synthesis lut_function=(A (B)+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_7_i165_3_lut_3_lut_rep_512.init = 16'h9c9c;
    LUT4 mux_192_Mux_3_i859_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n859_adj_2542)) /* synthesis lut_function=(!(A (B (D)+!B !(D))+!A (B (C+(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_3_i859_3_lut_3_lut_4_lut.init = 16'h339c;
    LUT4 i19193_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21523)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (D))+!A !(B (C (D))+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19193_3_lut_3_lut_4_lut.init = 16'h4933;
    PFUMX i18126 (.BLUT(n21426), .ALUT(n317_adj_2703), .C0(index_q[5]), 
          .Z(n20456));
    LUT4 n572_bdd_3_lut_22956_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n23651)) /* synthesis lut_function=(A (B (C+(D)))+!A (B ((D)+!C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n572_bdd_3_lut_22956_4_lut.init = 16'hcc94;
    LUT4 mux_192_Mux_2_i653_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n653_adj_2755)) /* synthesis lut_function=(A (B (C+!(D))+!B !(D))+!A !(B (C+!(D))+!B !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_2_i653_3_lut_4_lut.init = 16'h94aa;
    LUT4 mux_192_Mux_1_i93_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n93_adj_2753)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C+(D)))+!A !(B (C (D)+!C !(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_1_i93_3_lut_4_lut_4_lut.init = 16'h955a;
    PFUMX i18127 (.BLUT(n349_adj_2462), .ALUT(n21429), .C0(index_q[5]), 
          .Z(n20457));
    PFUMX i18152 (.BLUT(n20480), .ALUT(n20481), .C0(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_2141[1]));
    L6MUX21 i21501 (.D0(n23042), .D1(n23040), .SD(index_q[6]), .Z(n23043));
    L6MUX21 i18128 (.D0(n21432), .D1(n21435), .SD(index_q[5]), .Z(n20458));
    L6MUX21 i18129 (.D0(n21438), .D1(n21441), .SD(index_q[5]), .Z(n20459));
    PFUMX i18130 (.BLUT(n21444), .ALUT(n573_adj_2788), .C0(index_q[5]), 
          .Z(n20460));
    PFUMX i18245 (.BLUT(n20573), .ALUT(n20574), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2126[1]));
    LUT4 mux_192_Mux_6_i572_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n572_adj_2787)) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_6_i572_3_lut_4_lut.init = 16'hccd9;
    L6MUX21 i18131 (.D0(n21447), .D1(n636_adj_2295), .SD(index_q[5]), 
            .Z(n20461));
    PFUMX i18132 (.BLUT(n21450), .ALUT(n700_adj_2446), .C0(index_q[5]), 
          .Z(n20462));
    LUT4 i11398_3_lut_3_lut (.A(index_i[2]), .B(index_i[0]), .C(index_i[1]), 
         .Z(n38)) /* synthesis lut_function=(A (C)+!A (B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11398_3_lut_3_lut.init = 16'hf4f4;
    LUT4 i19217_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21547)) /* synthesis lut_function=(A (B (C)+!B (C (D)+!C !(D)))+!A !(B (C+!(D))+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19217_3_lut_4_lut_4_lut.init = 16'ha593;
    LUT4 mux_192_Mux_3_i397_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n397_adj_2762)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !(B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_3_i397_3_lut_4_lut_4_lut.init = 16'ha95a;
    LUT4 i19148_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21478)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A !(B (D)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19148_3_lut_3_lut_4_lut.init = 16'ha955;
    LUT4 i19227_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21557)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C+(D)))+!A (B (C)+!B !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19227_3_lut_4_lut_4_lut.init = 16'hc95a;
    LUT4 i20232_3_lut (.A(n109_adj_2327), .B(n124_adj_2612), .C(index_i[4]), 
         .Z(n20905)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20232_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_4_i349_3_lut_4_lut (.A(index_q[0]), .B(index_q[2]), 
         .C(index_q[4]), .D(n348_adj_2736), .Z(n349_adj_2719)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_4_i349_3_lut_4_lut.init = 16'hf606;
    L6MUX21 i18134 (.D0(n21453), .D1(n21456), .SD(index_q[5]), .Z(n20464));
    PFUMX i21499 (.BLUT(n23041), .ALUT(n62_adj_2319), .C0(index_q[5]), 
          .Z(n23042));
    LUT4 i11373_2_lut_rep_513 (.A(index_i[0]), .B(index_i[1]), .Z(n25073)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11373_2_lut_rep_513.init = 16'h2222;
    PFUMX i18136 (.BLUT(n924_adj_2458), .ALUT(n21462), .C0(index_q[5]), 
          .Z(n20466));
    LUT4 i15269_3_lut_3_lut (.A(index_q[0]), .B(index_q[2]), .C(index_q[3]), 
         .Z(n17532)) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i15269_3_lut_3_lut.init = 16'h6a6a;
    PFUMX i18137 (.BLUT(n987_adj_2789), .ALUT(n21465), .C0(index_q[5]), 
          .Z(n20467));
    LUT4 i20254_3_lut (.A(n620_adj_2273), .B(n13921), .C(index_q[4]), 
         .Z(n20883)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20254_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_0_i985_3_lut_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n985_adj_2790)) /* synthesis lut_function=(!(A (B+!(C))+!A (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_0_i985_3_lut_3_lut_3_lut.init = 16'h2525;
    LUT4 mux_192_Mux_4_i205_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n205_adj_2791)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_4_i205_3_lut_4_lut_4_lut.init = 16'h5a2a;
    PFUMX i21497 (.BLUT(n23039), .ALUT(n23038), .C0(index_q[5]), .Z(n23040));
    LUT4 mux_192_Mux_4_i723_3_lut_4_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n723)) /* synthesis lut_function=(A ((C)+!B)+!A !(B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_4_i723_3_lut_4_lut_4_lut_3_lut.init = 16'hb2b2;
    PFUMX i18613 (.BLUT(n20941), .ALUT(n20942), .C0(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_2141[7]));
    LUT4 i20257_3_lut (.A(n491_adj_2743), .B(n506_adj_2569), .C(index_q[4]), 
         .Z(n20877)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20257_3_lut.init = 16'hcaca;
    LUT4 i9580_3_lut_3_lut_4_lut (.A(n25188), .B(index_q[2]), .C(n15), 
         .D(index_q[4]), .Z(n12148)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9580_3_lut_3_lut_4_lut.init = 16'hf077;
    LUT4 mux_192_Mux_6_i157_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n157_adj_2792)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (D))+!A !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_6_i157_3_lut_4_lut_4_lut_4_lut.init = 16'h5d22;
    PFUMX i23006 (.BLUT(n25214), .ALUT(n25215), .C0(index_i[2]), .Z(n25216));
    LUT4 mux_192_Mux_6_i347_3_lut_4_lut_3_lut_rep_514 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n25074)) /* synthesis lut_function=(!(A (B+!(C))+!A ((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_6_i347_3_lut_4_lut_3_lut_rep_514.init = 16'h2424;
    LUT4 mux_192_Mux_4_i371_3_lut_4_lut_3_lut_rep_516 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n25076)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_4_i371_3_lut_4_lut_3_lut_rep_516.init = 16'h9292;
    LUT4 mux_192_Mux_6_i70_3_lut_rep_517 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n25077)) /* synthesis lut_function=(!(A (B+(C))+!A !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_6_i70_3_lut_rep_517.init = 16'h5252;
    LUT4 n908_bdd_3_lut_22805_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n23857)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A !(B ((D)+!C)+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n908_bdd_3_lut_22805_3_lut_4_lut.init = 16'h552c;
    LUT4 n21158_bdd_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n23983)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C))+!A !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n21158_bdd_3_lut_4_lut_4_lut.init = 16'h5a52;
    PFUMX i18183 (.BLUT(n20511), .ALUT(n20512), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2126[3]));
    LUT4 mux_192_Mux_2_i348_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n348_adj_2793)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_2_i348_3_lut_4_lut_4_lut.init = 16'h52a5;
    LUT4 mux_192_Mux_0_i812_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n812)) /* synthesis lut_function=(A (B (C+(D))+!B !(C))+!A (B (D)+!B !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_0_i812_3_lut_4_lut_4_lut_4_lut.init = 16'hcf92;
    LUT4 i19163_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21493)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C))+!A !(B ((D)+!C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19163_3_lut_4_lut_4_lut.init = 16'h925a;
    LUT4 i19055_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21385)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A !(B (C+!(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19055_3_lut_4_lut_4_lut.init = 16'ha52b;
    LUT4 mux_192_Mux_0_i491_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n491_adj_2386)) /* synthesis lut_function=(!(A (B (D)+!B !(C+!(D)))+!A ((C+!(D))+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_0_i491_3_lut_4_lut.init = 16'h24aa;
    LUT4 mux_192_Mux_5_i828_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[4]), .D(n25057), .Z(n828_adj_2759)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_5_i828_4_lut_4_lut.init = 16'hc66c;
    LUT4 mux_192_Mux_6_i732_3_lut_4_lut (.A(n25166), .B(index_i[3]), .C(index_i[4]), 
         .D(n412_adj_2636), .Z(n732_adj_2715)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_6_i732_3_lut_4_lut.init = 16'hf909;
    LUT4 i18536_3_lut (.A(n141_adj_2357), .B(n25160), .C(index_q[3]), 
         .Z(n20866)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18536_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_4_i14_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n978)) /* synthesis lut_function=(!(A (B+(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_4_i14_3_lut_3_lut.init = 16'h5656;
    LUT4 n526_bdd_3_lut_22966_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n23648)) /* synthesis lut_function=(!(A (B)+!A !(B (C+(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n526_bdd_3_lut_22966_3_lut_4_lut_4_lut.init = 16'h6663;
    PFUMX i18214 (.BLUT(n20542), .ALUT(n20543), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2126[2]));
    LUT4 i9491_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n526_adj_2283)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+(D)))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9491_3_lut_4_lut_4_lut.init = 16'h666c;
    LUT4 i18535_3_lut (.A(n85_adj_2600), .B(n25194), .C(index_q[3]), .Z(n20865)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18535_3_lut.init = 16'hcaca;
    LUT4 i9607_3_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[4]), 
         .Z(n12177)) /* synthesis lut_function=(!(A (B)+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9607_3_lut_4_lut_3_lut.init = 16'h6262;
    PFUMX i18248 (.BLUT(n20576), .ALUT(n20577), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2126[11]));
    LUT4 i18534_3_lut (.A(n27495), .B(n25193), .C(index_q[3]), .Z(n20864)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18534_3_lut.init = 16'hcaca;
    LUT4 i18533_3_lut (.A(n25160), .B(n27521), .C(index_q[3]), .Z(n20863)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18533_3_lut.init = 16'hcaca;
    LUT4 i18529_3_lut (.A(n25161), .B(n27521), .C(index_q[3]), .Z(n20859)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18529_3_lut.init = 16'hcaca;
    LUT4 i18528_3_lut (.A(n27495), .B(n108), .C(index_q[3]), .Z(n20858)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18528_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_6_i325_3_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n325_adj_2282)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_6_i325_3_lut_4_lut_3_lut.init = 16'h6d6d;
    PFUMX mux_192_Mux_14_i1023 (.BLUT(n511_adj_2606), .ALUT(n17770), .C0(index_i[9]), 
          .Z(quarter_wave_sample_register_i_15__N_2126[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 mux_192_Mux_7_i70_3_lut_rep_381_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n24941)) /* synthesis lut_function=(!(A (B)+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_7_i70_3_lut_rep_381_3_lut.init = 16'h6363;
    LUT4 mux_192_Mux_1_i746_3_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n746_adj_2794)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_1_i746_3_lut_4_lut_3_lut.init = 16'h8686;
    LUT4 i17333_4_lut (.A(n25095), .B(n892_adj_2769), .C(index_q[6]), 
         .D(index_q[5]), .Z(n19638)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D))))) */ ;
    defparam i17333_4_lut.init = 16'h3a35;
    LUT4 i18527_3_lut (.A(n85_adj_2600), .B(n25193), .C(index_q[3]), .Z(n20857)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18527_3_lut.init = 16'hcaca;
    LUT4 i20893_3_lut (.A(n19638), .B(n17788), .C(index_q[7]), .Z(n20891)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20893_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_1_i882_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n882)) /* synthesis lut_function=(A ((C)+!B)+!A !((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_1_i882_3_lut_3_lut.init = 16'ha6a6;
    LUT4 mux_192_Mux_7_i108_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n108_adj_2732)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_7_i108_3_lut_3_lut.init = 16'hc6c6;
    LUT4 mux_192_Mux_3_i507_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[4]), .D(n491_adj_2725), .Z(n507)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_3_i507_3_lut_4_lut.init = 16'h6f60;
    LUT4 i21077_2_lut_rep_265_3_lut_4_lut (.A(n25188), .B(index_q[2]), .C(index_q[5]), 
         .D(n25090), .Z(n24825)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21077_2_lut_rep_265_3_lut_4_lut.init = 16'h0f7f;
    LUT4 mux_192_Mux_0_i747_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n747)) /* synthesis lut_function=(!(A (B+!(C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_0_i747_3_lut_4_lut_4_lut_4_lut.init = 16'h6556;
    LUT4 mux_192_Mux_2_i731_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n731_adj_2754)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_2_i731_3_lut_4_lut_4_lut.init = 16'h6cc6;
    LUT4 i9515_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(n25113), .D(index_i[4]), .Z(n221_adj_2511)) /* synthesis lut_function=(!(A (B)+!A (B (C+(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9515_3_lut_4_lut_4_lut_4_lut.init = 16'h3336;
    LUT4 i21724_then_4_lut (.A(index_q[0]), .B(index_q[4]), .C(index_q[1]), 
         .D(index_q[3]), .Z(n25231)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam i21724_then_4_lut.init = 16'h3c69;
    LUT4 i18526_3_lut (.A(n25156), .B(n25205), .C(index_q[3]), .Z(n20856)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18526_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_1_i62_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[2]), 
         .C(index_q[4]), .D(index_q[3]), .Z(n62_adj_2767)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))+!A !(B (C)+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_1_i62_3_lut_4_lut_4_lut.init = 16'ha5a6;
    LUT4 i9605_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n12175)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B ((D)+!C)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9605_3_lut_4_lut_4_lut.init = 16'h6c3c;
    LUT4 n547_bdd_3_lut_4_lut (.A(index_q[0]), .B(index_q[2]), .C(n251_adj_2653), 
         .D(index_q[5]), .Z(n24042)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n547_bdd_3_lut_4_lut.init = 16'hf066;
    LUT4 mux_192_Mux_6_i442_3_lut_4_lut_3_lut_rep_519 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n25079)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_6_i442_3_lut_4_lut_3_lut_rep_519.init = 16'h6464;
    LUT4 mux_192_Mux_6_i7_3_lut_4_lut_3_lut_rep_520 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n25080)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_6_i7_3_lut_4_lut_3_lut_rep_520.init = 16'hd6d6;
    LUT4 mux_192_Mux_6_i483_3_lut_3_lut_rep_521 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n25081)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_6_i483_3_lut_3_lut_rep_521.init = 16'h6c6c;
    LUT4 mux_192_Mux_6_i29_3_lut_4_lut_3_lut_rep_522 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n25082)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_6_i29_3_lut_4_lut_3_lut_rep_522.init = 16'h6969;
    LUT4 mux_192_Mux_5_i652_3_lut_3_lut_rep_523 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n25083)) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_5_i652_3_lut_3_lut_rep_523.init = 16'h6a6a;
    LUT4 mux_192_Mux_6_i134_3_lut_4_lut_3_lut_rep_524 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n25084)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_6_i134_3_lut_4_lut_3_lut_rep_524.init = 16'h9696;
    LUT4 i18522_3_lut (.A(n27521), .B(n25195), .C(index_q[3]), .Z(n20852)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18522_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_5_i459_3_lut_4_lut_4_lut_3_lut_rep_525 (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[2]), .Z(n25085)) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_5_i459_3_lut_4_lut_4_lut_3_lut_rep_525.init = 16'h6b6b;
    LUT4 mux_192_Mux_5_i754_3_lut_4_lut_3_lut_rep_526 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n25086)) /* synthesis lut_function=(!(A (B)+!A ((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_5_i754_3_lut_4_lut_3_lut_rep_526.init = 16'h2626;
    LUT4 mux_192_Mux_5_i204_3_lut_3_lut_rep_527 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n25087)) /* synthesis lut_function=(!(A (B)+!A (B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_5_i204_3_lut_3_lut_rep_527.init = 16'h3636;
    LUT4 mux_192_Mux_5_i347_3_lut_4_lut_4_lut_3_lut_rep_528 (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[2]), .Z(n25088)) /* synthesis lut_function=(A ((C)+!B)+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_5_i347_3_lut_4_lut_4_lut_3_lut_rep_528.init = 16'hb6b6;
    PFUMX i18481 (.BLUT(n20809), .ALUT(n20810), .C0(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_2141[11]));
    LUT4 i18521_3_lut (.A(n1001), .B(n25161), .C(index_q[3]), .Z(n20851)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18521_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_5_i30_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n30_adj_2533)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A (B+!(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_5_i30_3_lut_4_lut.init = 16'hcc67;
    LUT4 n781_bdd_3_lut_4_lut_4_lut (.A(index_i[3]), .B(n781_adj_2302), 
         .C(index_i[4]), .D(n24969), .Z(n22893)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B ((D)+!C)+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n781_bdd_3_lut_4_lut_4_lut.init = 16'h5c0c;
    LUT4 i9523_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n12089)) /* synthesis lut_function=(!(A (B (D)+!B (C+!(D)))+!A !(B (D)+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9523_3_lut_4_lut_4_lut.init = 16'h4699;
    LUT4 mux_192_Mux_1_i301_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n301_adj_2415)) /* synthesis lut_function=(A (B (C+(D))+!B !(D))+!A !(B (C+(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_1_i301_3_lut_4_lut_4_lut.init = 16'h99b6;
    L6MUX21 i22312 (.D0(n23918), .D1(n23915), .SD(index_i[5]), .Z(n23919));
    LUT4 i8826_4_lut_4_lut (.A(index_i[3]), .B(index_i[0]), .C(index_i[1]), 
         .D(index_i[2]), .Z(n11355)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (D)+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i8826_4_lut_4_lut.init = 16'h0bf4;
    LUT4 mux_192_Mux_6_i475_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n475_adj_2756)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A !(B (C+(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_6_i475_3_lut_4_lut_4_lut.init = 16'h9936;
    LUT4 n173_bdd_3_lut (.A(n173_adj_2784), .B(n954_adj_2758), .C(index_i[4]), 
         .Z(n23387)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n173_bdd_3_lut.init = 16'hcaca;
    PFUMX i22310 (.BLUT(n23917), .ALUT(n23916), .C0(index_i[4]), .Z(n23918));
    LUT4 i19154_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21484)) /* synthesis lut_function=(!(A (B)+!A (B (C+(D))+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19154_3_lut_3_lut_4_lut.init = 16'h3326;
    LUT4 mux_192_Mux_5_i460_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n460_adj_2559)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A !(B (C)+!B !(C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_5_i460_3_lut_4_lut_4_lut.init = 16'h6b5a;
    LUT4 n604_bdd_3_lut_22972_3_lut_4_lut (.A(index_i[0]), .B(n25116), .C(index_i[4]), 
         .D(index_i[3]), .Z(n24736)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n604_bdd_3_lut_22972_3_lut_4_lut.init = 16'hf10f;
    LUT4 n396_bdd_3_lut_22051_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n23653)) /* synthesis lut_function=(A (B (C+(D))+!B ((D)+!C))+!A !(B (C+(D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n396_bdd_3_lut_22051_4_lut.init = 16'haa96;
    LUT4 mux_192_Mux_2_i491_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n491_adj_2795)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A !(B (C)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_2_i491_3_lut_4_lut_4_lut.init = 16'h6a5a;
    LUT4 mux_192_Mux_0_i142_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n142)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C))+!A !(B (C (D)+!C !(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_0_i142_3_lut_4_lut_4_lut.init = 16'ha569;
    LUT4 mux_192_Mux_0_i124_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n124_adj_2773)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A !(B (D)+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_0_i124_3_lut_4_lut_4_lut.init = 16'h6c99;
    LUT4 i19023_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21353)) /* synthesis lut_function=(A (B (C)+!B !(C (D)+!C !(D)))+!A (B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19023_3_lut_4_lut_4_lut.init = 16'hd6a5;
    LUT4 n483_bdd_3_lut_22787_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n23917)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C))+!A !(B (C+!(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n483_bdd_3_lut_22787_4_lut_4_lut.init = 16'h5ad6;
    LUT4 i19070_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21400)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19070_3_lut_4_lut.init = 16'h64cc;
    LUT4 i18660_4_lut_3_lut (.A(index_i[3]), .B(index_i[4]), .C(n24970), 
         .Z(n20990)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18660_4_lut_3_lut.init = 16'h6565;
    LUT4 i7177_2_lut_rep_530 (.A(index_q[3]), .B(index_q[4]), .Z(n25090)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i7177_2_lut_rep_530.init = 16'heeee;
    LUT4 mux_192_Mux_6_i924_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[4]), .D(n762_adj_2349), .Z(n924_adj_2783)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_6_i924_3_lut_4_lut.init = 16'h6f60;
    LUT4 i9471_3_lut_3_lut_4_lut (.A(index_q[3]), .B(index_q[4]), .C(n25180), 
         .D(index_q[0]), .Z(n605_adj_2686)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9471_3_lut_3_lut_4_lut.init = 16'h10fe;
    LUT4 i18881_then_4_lut (.A(index_q[2]), .B(index_q[1]), .C(index_q[4]), 
         .D(index_q[3]), .Z(n25238)) /* synthesis lut_function=(A (B (C+(D))+!B !(C))+!A !(B (C+(D))+!B !(C+!(D)))) */ ;
    defparam i18881_then_4_lut.init = 16'h9a97;
    LUT4 i9455_3_lut_4_lut (.A(index_q[3]), .B(index_q[4]), .C(n25197), 
         .D(n27522), .Z(n605_adj_2744)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9455_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i2_3_lut_4_lut_adj_80 (.A(index_q[3]), .B(index_q[4]), .C(index_q[5]), 
         .D(n25211), .Z(n17673)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i2_3_lut_4_lut_adj_80.init = 16'hfffe;
    LUT4 i11219_2_lut_rep_531 (.A(index_q[2]), .B(index_q[3]), .Z(n25091)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11219_2_lut_rep_531.init = 16'heeee;
    LUT4 i18519_3_lut (.A(n25195), .B(n25156), .C(index_q[3]), .Z(n20849)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18519_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_4_i221_3_lut_3_lut (.A(index_i[0]), .B(index_i[4]), 
         .C(n205_adj_2791), .Z(n221_adj_2781)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_4_i221_3_lut_3_lut.init = 16'h7474;
    LUT4 i21724_else_4_lut (.A(index_q[0]), .B(index_q[4]), .C(index_q[1]), 
         .D(index_q[3]), .Z(n25230)) /* synthesis lut_function=(!(A (B (C)+!B !(C (D)+!C !(D)))+!A (B ((D)+!C)+!B !((D)+!C)))) */ ;
    defparam i21724_else_4_lut.init = 16'h394b;
    LUT4 i11576_2_lut_rep_389_3_lut (.A(index_q[2]), .B(index_q[3]), .C(index_q[1]), 
         .Z(n24949)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11576_2_lut_rep_389_3_lut.init = 16'hfefe;
    LUT4 mux_192_Mux_2_i349_3_lut_3_lut (.A(index_i[0]), .B(index_i[4]), 
         .C(n348_adj_2793), .Z(n349_adj_2427)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_2_i349_3_lut_3_lut.init = 16'hd1d1;
    PFUMX i23024 (.BLUT(n25243), .ALUT(n25244), .C0(index_i[1]), .Z(n25245));
    LUT4 i21148_2_lut_rep_302_2_lut_3_lut_4_lut (.A(index_q[2]), .B(index_q[3]), 
         .C(index_q[1]), .D(index_q[0]), .Z(n24862)) /* synthesis lut_function=(!(A+(B+(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21148_2_lut_rep_302_2_lut_3_lut_4_lut.init = 16'h0111;
    LUT4 i21139_3_lut_3_lut (.A(index_q[3]), .B(index_q[2]), .C(index_q[5]), 
         .Z(n19828)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21139_3_lut_3_lut.init = 16'hfbfb;
    LUT4 i8828_4_lut_4_lut (.A(index_q[3]), .B(index_q[0]), .C(index_q[1]), 
         .D(index_q[2]), .Z(n11358)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (D)+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i8828_4_lut_4_lut.init = 16'h0bf4;
    LUT4 mux_192_Mux_5_i573_3_lut_3_lut (.A(index_i[0]), .B(index_i[4]), 
         .C(n572_adj_2786), .Z(n573_adj_2752)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_5_i573_3_lut_3_lut.init = 16'hd1d1;
    LUT4 i11281_2_lut_3_lut_3_lut (.A(index_q[3]), .B(index_q[1]), .C(index_q[0]), 
         .Z(n13956)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11281_2_lut_3_lut_3_lut.init = 16'h4040;
    LUT4 i18881_else_4_lut (.A(index_q[2]), .B(index_q[1]), .C(index_q[4]), 
         .D(index_q[3]), .Z(n25237)) /* synthesis lut_function=(!(A (B (C)+!B (C+(D)))+!A !(B (C (D)+!C !(D))+!B (C+!(D))))) */ ;
    defparam i18881_else_4_lut.init = 16'h581f;
    LUT4 n781_bdd_3_lut_4_lut_4_lut_adj_81 (.A(index_q[3]), .B(n781_adj_2307), 
         .C(index_q[4]), .D(n24956), .Z(n22876)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B ((D)+!C)+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n781_bdd_3_lut_4_lut_4_lut_adj_81.init = 16'h5c0c;
    LUT4 i10980_4_lut_4_lut (.A(index_q[3]), .B(index_q[2]), .C(index_q[0]), 
         .D(index_q[1]), .Z(n875)) /* synthesis lut_function=((B (C)+!B (D))+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i10980_4_lut_4_lut.init = 16'hf7d5;
    PFUMX i17920 (.BLUT(n20248), .ALUT(n20249), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2126[9]));
    LUT4 mux_193_Mux_1_i573_3_lut_4_lut_4_lut (.A(index_q[3]), .B(n557_adj_2647), 
         .C(index_q[4]), .D(n25160), .Z(n573_adj_2788)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B ((D)+!C)+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_1_i573_3_lut_4_lut_4_lut.init = 16'h5c0c;
    LUT4 i18360_3_lut_4_lut_3_lut (.A(index_q[3]), .B(index_q[4]), .C(n24980), 
         .Z(n20690)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18360_3_lut_4_lut_3_lut.init = 16'h6464;
    LUT4 mux_193_Mux_1_i987_3_lut_4_lut_4_lut (.A(index_q[3]), .B(n986_adj_2763), 
         .C(index_q[4]), .D(n25160), .Z(n987_adj_2789)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_1_i987_3_lut_4_lut_4_lut.init = 16'hc5c0;
    PFUMX i22307 (.BLUT(n23914), .ALUT(n23913), .C0(index_i[4]), .Z(n23915));
    LUT4 mux_193_Mux_2_i221_4_lut_4_lut (.A(index_q[3]), .B(index_q[4]), 
         .C(n24957), .D(n24857), .Z(n221_adj_2770)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (B+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_2_i221_4_lut_4_lut.init = 16'hf7c4;
    LUT4 i18569_4_lut_3_lut (.A(index_q[3]), .B(index_q[4]), .C(n24957), 
         .Z(n20899)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18569_4_lut_3_lut.init = 16'h6565;
    LUT4 mux_192_Mux_2_i763_4_lut_4_lut (.A(index_i[0]), .B(n12118), .C(index_i[4]), 
         .D(n157_adj_2792), .Z(n763_adj_2435)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_2_i763_4_lut_4_lut.init = 16'hdfd0;
    LUT4 mux_193_Mux_1_i890_4_lut_4_lut_4_lut_4_lut (.A(index_q[3]), .B(index_q[4]), 
         .C(n25156), .D(index_q[0]), .Z(n890_adj_2631)) /* synthesis lut_function=(!(A (B (D)+!B !(C))+!A (B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_1_i890_4_lut_4_lut_4_lut_4_lut.init = 16'h31fd;
    L6MUX21 i12810362_i1 (.D0(n21084), .D1(n21706), .SD(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_2141[0]));
    LUT4 mux_192_Mux_3_i700_3_lut_3_lut (.A(index_i[0]), .B(index_i[4]), 
         .C(n684_adj_2635), .Z(n700)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_3_i700_3_lut_3_lut.init = 16'h7474;
    LUT4 i9442_3_lut_3_lut (.A(index_q[3]), .B(index_q[4]), .C(n12007), 
         .Z(n12008)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9442_3_lut_3_lut.init = 16'h7474;
    LUT4 i11474_4_lut_4_lut (.A(index_i[3]), .B(index_i[2]), .C(index_i[0]), 
         .D(index_i[1]), .Z(n875_adj_2263)) /* synthesis lut_function=((B (C)+!B (D))+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11474_4_lut_4_lut.init = 16'hf7d5;
    LUT4 mux_192_Mux_1_i987_3_lut_4_lut_4_lut (.A(index_i[3]), .B(n986_adj_2683), 
         .C(index_i[4]), .D(n25038), .Z(n987)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_1_i987_3_lut_4_lut_4_lut.init = 16'hc5c0;
    LUT4 i18390_3_lut_4_lut_3_lut (.A(index_i[3]), .B(index_i[4]), .C(n24947), 
         .Z(n20720)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18390_3_lut_4_lut_3_lut.init = 16'h6464;
    L6MUX21 i12798356_i1 (.D0(n21022), .D1(n21786), .SD(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2126[0]));
    PFUMX i17951 (.BLUT(n20279), .ALUT(n20280), .C0(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_2141[5]));
    L6MUX21 i18825 (.D0(n21151), .D1(n21152), .SD(index_i[8]), .Z(n21155));
    PFUMX i18851 (.BLUT(n21179), .ALUT(n21180), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2126[8]));
    LUT4 i7171_2_lut_rep_535 (.A(index_q[3]), .B(index_q[4]), .Z(n25095)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i7171_2_lut_rep_535.init = 16'h8888;
    LUT4 i18989_3_lut_3_lut_4_lut (.A(index_q[3]), .B(index_q[4]), .C(n413), 
         .D(index_q[5]), .Z(n21319)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18989_3_lut_3_lut_4_lut.init = 16'h77f0;
    PFUMX mux_193_Mux_14_i1023 (.BLUT(n511), .ALUT(n19498), .C0(index_q[9]), 
          .Z(quarter_wave_sample_register_q_15__N_2141[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 mux_192_Mux_1_i890_4_lut_4_lut_4_lut_4_lut (.A(index_i[3]), .B(index_i[4]), 
         .C(n24941), .D(index_i[0]), .Z(n890_adj_2485)) /* synthesis lut_function=(!(A (B (D)+!B !(C))+!A (B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_1_i890_4_lut_4_lut_4_lut_4_lut.init = 16'h31fd;
    LUT4 i1_2_lut_rep_395_3_lut (.A(index_q[3]), .B(index_q[4]), .C(index_q[5]), 
         .Z(n24955)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_2_lut_rep_395_3_lut.init = 16'hf8f8;
    LUT4 i11247_2_lut_rep_536 (.A(index_q[2]), .B(index_q[3]), .Z(n25096)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11247_2_lut_rep_536.init = 16'h8888;
    LUT4 i20295_3_lut (.A(n109), .B(n124_adj_2536), .C(index_q[4]), .Z(n20819)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20295_3_lut.init = 16'hcaca;
    LUT4 i11577_2_lut_rep_344_3_lut (.A(index_q[2]), .B(index_q[3]), .C(index_q[1]), 
         .Z(n24904)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11577_2_lut_rep_344_3_lut.init = 16'h8080;
    LUT4 i2_2_lut_rep_388_3_lut_4_lut (.A(index_q[2]), .B(index_q[3]), .C(index_q[1]), 
         .D(index_q[0]), .Z(n24948)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i2_2_lut_rep_388_3_lut_4_lut.init = 16'h8000;
    LUT4 mux_193_Mux_7_i924_3_lut_3_lut_4_lut (.A(index_q[2]), .B(index_q[3]), 
         .C(index_q[4]), .D(n25188), .Z(n924_adj_2343)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_7_i924_3_lut_3_lut_4_lut.init = 16'h878f;
    LUT4 i18362_3_lut_3_lut_3_lut_4_lut (.A(index_q[2]), .B(index_q[3]), 
         .C(index_q[4]), .D(index_q[1]), .Z(n20692)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18362_3_lut_3_lut_3_lut_4_lut.init = 16'h878f;
    PFUMX i18028 (.BLUT(n20356), .ALUT(n20357), .C0(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_2141[3]));
    LUT4 mux_192_Mux_4_i142_3_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[3]), 
         .C(index_i[2]), .Z(n142_adj_2716)) /* synthesis lut_function=(A (B (C))+!A !(B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_4_i142_3_lut_4_lut_3_lut.init = 16'h9595;
    LUT4 i11226_2_lut_rep_310_3_lut_4_lut (.A(index_q[2]), .B(index_q[3]), 
         .C(index_q[4]), .D(n25188), .Z(n24870)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11226_2_lut_rep_310_3_lut_4_lut.init = 16'hf8f0;
    L6MUX21 i18949 (.D0(n21275), .D1(n21276), .SD(index_q[8]), .Z(n21279));
    LUT4 i17528_1_lut_2_lut (.A(index_q[2]), .B(index_q[3]), .Z(n19858)) /* synthesis lut_function=(!(A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i17528_1_lut_2_lut.init = 16'h7777;
    LUT4 mux_192_Mux_0_i572_3_lut_4_lut (.A(index_i[0]), .B(n25116), .C(index_i[3]), 
         .D(n25087), .Z(n572)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_0_i572_3_lut_4_lut.init = 16'hefe0;
    PFUMX i18983 (.BLUT(n21311), .ALUT(n21312), .C0(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_2141[8]));
    PFUMX i18059 (.BLUT(n20387), .ALUT(n20388), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2126[5]));
    LUT4 i11655_2_lut_2_lut_3_lut (.A(index_q[2]), .B(index_q[3]), .C(index_q[0]), 
         .Z(n14330)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11655_2_lut_2_lut_3_lut.init = 16'h0808;
    LUT4 i11418_2_lut_rep_537 (.A(index_q[1]), .B(index_q[2]), .Z(n25097)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11418_2_lut_rep_537.init = 16'heeee;
    PFUMX i18090 (.BLUT(n20418), .ALUT(n20419), .C0(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_2141[2]));
    PFUMX i19186 (.BLUT(n21514), .ALUT(n21515), .C0(index_i[4]), .Z(n21516));
    LUT4 mux_193_Mux_3_i1002_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n19655)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (D))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_3_i1002_3_lut_3_lut_4_lut.init = 16'hf708;
    LUT4 mux_192_Mux_3_i251_3_lut_4_lut (.A(index_i[0]), .B(n25116), .C(index_i[3]), 
         .D(n24985), .Z(n14998)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_3_i251_3_lut_4_lut.init = 16'hfe0e;
    PFUMX i19189 (.BLUT(n21517), .ALUT(n21518), .C0(index_i[4]), .Z(n21519));
    LUT4 mux_193_Mux_9_i93_3_lut_3_lut_3_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .Z(n93_adj_2354)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_9_i93_3_lut_3_lut_3_lut.init = 16'hc1c1;
    LUT4 mux_193_Mux_4_i236_3_lut_4_lut_4_lut_3_lut_rep_463_4_lut (.A(index_q[1]), 
         .B(index_q[2]), .C(index_q[3]), .D(index_q[0]), .Z(n25023)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_4_i236_3_lut_4_lut_4_lut_3_lut_rep_463_4_lut.init = 16'hf01f;
    LUT4 i11567_2_lut_rep_279_2_lut_3_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[0]), .Z(n24839)) /* synthesis lut_function=(A (C)+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11567_2_lut_rep_279_2_lut_3_lut.init = 16'hf1f1;
    PFUMX i18121 (.BLUT(n20449), .ALUT(n20450), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2126[4]));
    LUT4 mux_192_Mux_3_i747_3_lut (.A(n25079), .B(n498), .C(index_i[3]), 
         .Z(n747_adj_2290)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_3_i747_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_0_i46_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[0]), .D(index_q[3]), .Z(n46_adj_2730)) /* synthesis lut_function=(A ((D)+!B)+!A (B (D)+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i46_3_lut_4_lut_4_lut_4_lut.init = 16'hfe33;
    LUT4 n21359_bdd_3_lut_3_lut (.A(index_q[1]), .B(n526_adj_2499), .C(index_q[4]), 
         .Z(n23396)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n21359_bdd_3_lut_3_lut.init = 16'h5c5c;
    LUT4 quarter_wave_sample_register_i_11__I_0_3_lut (.A(quarter_wave_sample_register_i[11]), 
         .B(o_val_pipeline_i_0__15__N_2157[11]), .C(phase_negation_i[1]), 
         .Z(o_val_pipeline_i_0__15__N_2164)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[14] 77[8])
    defparam quarter_wave_sample_register_i_11__I_0_3_lut.init = 16'hcaca;
    LUT4 i18864_3_lut_4_lut_3_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .D(index_q[0]), .Z(n21194)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18864_3_lut_4_lut_3_lut_4_lut.init = 16'h0fe0;
    LUT4 i11213_2_lut_rep_361_3_lut (.A(index_q[1]), .B(index_q[2]), .C(index_q[3]), 
         .Z(n24921)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11213_2_lut_rep_361_3_lut.init = 16'he0e0;
    LUT4 i11214_2_lut_rep_296_3_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[4]), .D(index_q[3]), .Z(n24856)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11214_2_lut_rep_296_3_lut_4_lut.init = 16'hfef0;
    LUT4 i10967_2_lut_rep_396_3_lut (.A(index_q[1]), .B(index_q[2]), .C(index_q[0]), 
         .Z(n24956)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i10967_2_lut_rep_396_3_lut.init = 16'hfefe;
    LUT4 mux_193_Mux_9_i285_3_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .D(index_q[0]), .Z(n285_adj_2591)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_9_i285_3_lut_4_lut_4_lut.init = 16'hc0c1;
    LUT4 mux_193_Mux_2_i173_3_lut_3_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .D(index_q[0]), .Z(n173_adj_2577)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_2_i173_3_lut_3_lut_4_lut.init = 16'h0e1e;
    LUT4 i11204_2_lut_rep_315_3_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .D(index_q[0]), .Z(n24875)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11204_2_lut_rep_315_3_lut_4_lut.init = 16'hf0e0;
    LUT4 mux_193_Mux_5_i954_3_lut_3_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .D(index_q[0]), .Z(n954_adj_2508)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B (C)+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_5_i954_3_lut_3_lut_4_lut_4_lut.init = 16'h0c1c;
    L6MUX21 i18149 (.D0(n20474), .D1(n20475), .SD(index_q[7]), .Z(n20479));
    LUT4 n46_bdd_3_lut_21511_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[4]), .D(index_q[3]), .Z(n23051)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C+(D)))+!A (B (C (D)+!C !(D))+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n46_bdd_3_lut_21511_4_lut_4_lut_4_lut.init = 16'hc10f;
    L6MUX21 i22257 (.D0(n23861), .D1(n23858), .SD(index_i[5]), .Z(n23862));
    LUT4 mux_193_Mux_8_i716_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[0]), .D(index_q[3]), .Z(n716_adj_2734)) /* synthesis lut_function=(!(A (B (D))+!A (B (D)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_8_i716_3_lut_4_lut_4_lut_4_lut.init = 16'h33fe;
    PFUMX i22255 (.BLUT(n23860), .ALUT(n23859), .C0(index_i[4]), .Z(n23861));
    LUT4 mux_192_Mux_2_i221_4_lut_4_lut (.A(index_i[3]), .B(index_i[4]), 
         .C(n24970), .D(n24859), .Z(n221_adj_2424)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (B+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_2_i221_4_lut_4_lut.init = 16'hf7c4;
    LUT4 i9482_3_lut_3_lut (.A(index_i[3]), .B(index_i[4]), .C(n12047), 
         .Z(n12048)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9482_3_lut_3_lut.init = 16'h7474;
    LUT4 mux_192_Mux_2_i507_3_lut_3_lut (.A(index_i[0]), .B(index_i[4]), 
         .C(n491_adj_2795), .Z(n507_adj_2429)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_2_i507_3_lut_3_lut.init = 16'h7474;
    LUT4 mux_193_Mux_5_i781_3_lut_4_lut_4_lut (.A(index_q[1]), .B(n25178), 
         .C(index_q[3]), .D(n25011), .Z(n781_adj_2676)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_5_i781_3_lut_4_lut_4_lut.init = 16'hfc5c;
    PFUMX i22252 (.BLUT(n23857), .ALUT(n908_adj_2750), .C0(index_i[4]), 
          .Z(n23858));
    LUT4 mux_192_Mux_1_i62_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[4]), .D(index_i[3]), .Z(n62_adj_2764)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))+!A !(B (C)+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_1_i62_3_lut_4_lut_4_lut.init = 16'ha5a6;
    LUT4 n543_bdd_3_lut_4_lut (.A(index_i[0]), .B(index_i[2]), .C(n251_adj_2562), 
         .D(index_i[5]), .Z(n23986)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n543_bdd_3_lut_4_lut.init = 16'hf066;
    LUT4 i19022_3_lut_4_lut_4_lut (.A(index_i[0]), .B(n25083), .C(index_i[3]), 
         .D(n25122), .Z(n21352)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19022_3_lut_4_lut_4_lut.init = 16'hcfc5;
    LUT4 mux_192_Mux_4_i349_3_lut_4_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[4]), .D(n348_adj_2761), .Z(n349_adj_2785)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_4_i349_3_lut_4_lut.init = 16'hf606;
    L6MUX21 i22234 (.D0(n23840), .D1(n23837), .SD(index_q[5]), .Z(n23841));
    PFUMX i22232 (.BLUT(n15_adj_2531), .ALUT(n23838), .C0(index_q[4]), 
          .Z(n23840));
    LUT4 mux_192_Mux_4_i252_4_lut_4_lut (.A(index_i[0]), .B(index_i[3]), 
         .C(n25116), .D(index_i[4]), .Z(n252_adj_2782)) /* synthesis lut_function=(!(A (B (D)+!B !(D))+!A !(B ((D)+!C)+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_4_i252_4_lut_4_lut.init = 16'h669d;
    LUT4 mux_192_Mux_3_i444_3_lut_4_lut (.A(index_i[0]), .B(index_i[3]), 
         .C(n25122), .D(index_i[4]), .Z(n444)) /* synthesis lut_function=(!(A (B (D)+!B (C (D)))+!A !(B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_3_i444_3_lut_4_lut.init = 16'h46aa;
    PFUMX i22229 (.BLUT(n23836), .ALUT(n23835), .C0(index_q[4]), .Z(n23837));
    LUT4 i15276_3_lut_3_lut (.A(index_i[0]), .B(index_i[2]), .C(index_i[3]), 
         .Z(n17539)) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i15276_3_lut_3_lut.init = 16'h6a6a;
    LUT4 i11342_2_lut_rep_485 (.A(index_i[0]), .B(index_i[1]), .Z(n25045)) /* synthesis lut_function=((B)+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11342_2_lut_rep_485.init = 16'hdddd;
    LUT4 i18828_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n21158)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (D))+!A !(D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18828_3_lut_4_lut_4_lut_4_lut.init = 16'ha25d;
    LUT4 mux_192_Mux_1_i908_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n908_adj_2750)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+(D)))+!A (B (C+(D))+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_1_i908_3_lut_4_lut_4_lut_4_lut.init = 16'h332d;
    LUT4 i1_2_lut_rep_445 (.A(index_q[6]), .B(index_q[7]), .Z(n25005)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_2_lut_rep_445.init = 16'heeee;
    LUT4 mux_192_Mux_6_i540_3_lut_3_lut_3_lut_rep_678 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27518)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_6_i540_3_lut_3_lut_3_lut_rep_678.init = 16'h9393;
    L6MUX21 i18242 (.D0(n20567), .D1(n20568), .SD(index_i[7]), .Z(n20572));
    PFUMX i19198 (.BLUT(n21526), .ALUT(n21527), .C0(index_i[4]), .Z(n21528));
    LUT4 i11325_3_lut_3_lut_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[0]), 
         .Z(n85)) /* synthesis lut_function=(!(A ((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11325_3_lut_3_lut_3_lut.init = 16'h5d5d;
    PFUMX i19201 (.BLUT(n21529), .ALUT(n21530), .C0(index_i[4]), .Z(n21531));
    LUT4 mux_192_Mux_0_i635_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n635)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_0_i635_3_lut_4_lut_4_lut.init = 16'hfd0a;
    LUT4 i11280_3_lut_3_lut (.A(index_q[1]), .B(index_q[0]), .C(index_q[2]), 
         .Z(n85_adj_2600)) /* synthesis lut_function=(!(A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11280_3_lut_3_lut.init = 16'h7575;
    LUT4 i9480_3_lut_4_lut (.A(index_i[0]), .B(n25116), .C(index_i[3]), 
         .D(index_i[4]), .Z(n12046)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9480_3_lut_4_lut.init = 16'h0e1e;
    LUT4 n476_bdd_3_lut_21855_3_lut (.A(index_i[1]), .B(index_i[4]), .C(n124_adj_2459), 
         .Z(n22932)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n476_bdd_3_lut_21855_3_lut.init = 16'hd1d1;
    LUT4 mux_192_Mux_6_i300_3_lut_rep_487 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n25047)) /* synthesis lut_function=(A (B+!(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_6_i300_3_lut_rep_487.init = 16'hdada;
    LUT4 quarter_wave_sample_register_i_10__I_0_3_lut (.A(quarter_wave_sample_register_i[10]), 
         .B(o_val_pipeline_i_0__15__N_2157[10]), .C(phase_negation_i[1]), 
         .Z(o_val_pipeline_i_0__15__N_2166)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[14] 77[8])
    defparam quarter_wave_sample_register_i_10__I_0_3_lut.init = 16'hcaca;
    LUT4 i19190_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21520)) /* synthesis lut_function=(!(A (B (C (D))+!B (C (D)+!C !(D)))+!A !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19190_3_lut_4_lut_4_lut.init = 16'h5aad;
    LUT4 n277_bdd_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n23914)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n277_bdd_3_lut_4_lut_4_lut.init = 16'ha5ad;
    LUT4 i19076_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21406)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19076_3_lut_4_lut_4_lut.init = 16'hda5a;
    L6MUX21 i18254 (.D0(n20582), .D1(n20583), .SD(index_q[8]), .Z(n20584));
    LUT4 i18596_4_lut_4_lut_3_lut_4_lut (.A(index_i[0]), .B(n25116), .C(index_i[4]), 
         .D(index_i[3]), .Z(n20926)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18596_4_lut_4_lut_3_lut_4_lut.init = 16'h11ef;
    PFUMX i19204 (.BLUT(n21532), .ALUT(n21533), .C0(index_i[4]), .Z(n21534));
    L6MUX21 i18257 (.D0(n20585), .D1(n20586), .SD(index_i[8]), .Z(n20587));
    L6MUX21 i22206 (.D0(n23810), .D1(n23808), .SD(index_i[5]), .Z(n23811));
    PFUMX i19207 (.BLUT(n21535), .ALUT(n21536), .C0(index_i[4]), .Z(n21537));
    PFUMX i22204 (.BLUT(n23809), .ALUT(n285), .C0(index_i[4]), .Z(n23810));
    LUT4 i21090_2_lut_rep_450 (.A(index_q[4]), .B(index_q[3]), .Z(n25010)) /* synthesis lut_function=(A+!(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21090_2_lut_rep_450.init = 16'hbbbb;
    LUT4 i20522_3_lut_4_lut (.A(index_q[4]), .B(index_q[3]), .C(n25259), 
         .D(n746), .Z(n763_adj_2391)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20522_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i11269_2_lut_rep_272_3_lut_4_lut (.A(index_i[0]), .B(n25116), .C(index_i[4]), 
         .D(index_i[3]), .Z(n24832)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11269_2_lut_rep_272_3_lut_4_lut.init = 16'hfef0;
    LUT4 i17500_2_lut_rep_544 (.A(index_q[5]), .B(index_q[4]), .Z(n25104)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i17500_2_lut_rep_544.init = 16'h8888;
    LUT4 i11971_2_lut_rep_451 (.A(index_q[2]), .B(index_q[0]), .Z(n25011)) /* synthesis lut_function=(A (B)) */ ;
    defparam i11971_2_lut_rep_451.init = 16'h8888;
    LUT4 i11197_3_lut_4_lut (.A(index_q[5]), .B(index_q[4]), .C(index_q[6]), 
         .D(index_q[3]), .Z(n509)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11197_3_lut_4_lut.init = 16'hf8f0;
    LUT4 mux_193_Mux_0_i236_3_lut_3_lut (.A(index_q[0]), .B(index_q[2]), 
         .C(index_q[3]), .Z(n236_adj_2666)) /* synthesis lut_function=(A (B+(C))+!A !(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i236_3_lut_3_lut.init = 16'ha9a9;
    LUT4 mux_192_Mux_0_i364_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n364_adj_2373)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A ((C+!(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_0_i364_3_lut_3_lut_4_lut.init = 16'hdb55;
    LUT4 i19173_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21503)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D))+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19173_3_lut_4_lut.init = 16'hccdb;
    LUT4 i19212_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21542)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C))+!A !(B (C)+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19212_3_lut_4_lut_4_lut.init = 16'h5ad3;
    PFUMX i22202 (.BLUT(n78), .ALUT(n23807), .C0(index_i[4]), .Z(n23808));
    PFUMX i22184 (.BLUT(n23789), .ALUT(n23788), .C0(index_i[4]), .Z(n23790));
    LUT4 n23394_bdd_3_lut (.A(n23394), .B(n476_adj_2470), .C(index_q[5]), 
         .Z(n23395)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n23394_bdd_3_lut.init = 16'hcaca;
    L6MUX21 i22181 (.D0(n23786), .D1(n23783), .SD(index_q[5]), .Z(n23787));
    PFUMX i22179 (.BLUT(n23785), .ALUT(n23784), .C0(index_q[4]), .Z(n23786));
    LUT4 i19176_3_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[3]), .C(index_i[2]), 
         .D(index_i[0]), .Z(n21506)) /* synthesis lut_function=(A (B (D)+!B (C (D)+!C !(D)))+!A (B (D)+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19176_3_lut_4_lut_4_lut.init = 16'hfc13;
    PFUMX i19213 (.BLUT(n21541), .ALUT(n21542), .C0(index_i[4]), .Z(n21543));
    LUT4 mux_193_Mux_6_i332_3_lut_4_lut_3_lut_3_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[0]), .Z(n332)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_6_i332_3_lut_4_lut_3_lut_3_lut.init = 16'h3d3d;
    LUT4 i10957_2_lut_rep_420_3_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .Z(n24980)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i10957_2_lut_rep_420_3_lut.init = 16'hf8f8;
    PFUMX i19376 (.BLUT(n21704), .ALUT(n21705), .C0(index_q[8]), .Z(n21706));
    LUT4 i18074_4_lut_4_lut (.A(index_q[4]), .B(index_q[5]), .C(n25225), 
         .D(n908_adj_2702), .Z(n20404)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam i18074_4_lut_4_lut.init = 16'hd1c0;
    LUT4 i20992_2_lut_rep_456 (.A(index_i[1]), .B(index_i[2]), .Z(n25016)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20992_2_lut_rep_456.init = 16'h9999;
    LUT4 n22_bdd_2_lut_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[3]), 
         .Z(n23632)) /* synthesis lut_function=(A (B+(C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n22_bdd_2_lut_3_lut.init = 16'hf9f9;
    LUT4 i11275_3_lut_rep_321_4_lut (.A(n25113), .B(index_i[4]), .C(index_i[5]), 
         .D(n25163), .Z(n24881)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11275_3_lut_rep_321_4_lut.init = 16'hf8f0;
    LUT4 mux_192_Mux_0_i93_3_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .Z(n93_adj_2737)) /* synthesis lut_function=(A (B)+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_0_i93_3_lut_3_lut.init = 16'h9c9c;
    PFUMX i22176 (.BLUT(n301_adj_2571), .ALUT(n23782), .C0(index_q[4]), 
          .Z(n23783));
    LUT4 n23398_bdd_3_lut_21892 (.A(n25222), .B(n23396), .C(index_q[5]), 
         .Z(n23399)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n23398_bdd_3_lut_21892.init = 16'hcaca;
    LUT4 mux_192_Mux_5_i781_3_lut_4_lut_4_lut (.A(index_i[1]), .B(n25079), 
         .C(index_i[3]), .D(n25033), .Z(n781_adj_2550)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_5_i781_3_lut_4_lut_4_lut.init = 16'hfc5c;
    LUT4 i18937_3_lut (.A(n23841), .B(n21252), .C(index_q[6]), .Z(n21267)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18937_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_6_i924_3_lut_4_lut (.A(index_q[2]), .B(index_q[3]), 
         .C(index_q[4]), .D(n762_adj_2337), .Z(n924_adj_2780)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_6_i924_3_lut_4_lut.init = 16'h6f60;
    PFUMX i19219 (.BLUT(n21547), .ALUT(n21548), .C0(index_i[4]), .Z(n21549));
    PFUMX i19222 (.BLUT(n21550), .ALUT(n21551), .C0(index_i[4]), .Z(n21552));
    PFUMX i21407 (.BLUT(n22937), .ALUT(n22933), .C0(index_i[6]), .Z(n22938));
    LUT4 mux_193_Mux_3_i94_3_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[4]), .D(n93_adj_2621), .Z(n94_adj_2723)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_3_i94_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_193_Mux_3_i62_3_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[4]), .D(n812_adj_2296), .Z(n62_adj_2768)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_3_i62_3_lut_4_lut.init = 16'h6f60;
    PFUMX i9449 (.BLUT(n12171), .ALUT(n12172), .C0(n19858), .Z(n12015));
    LUT4 i5507_1_lut_rep_457 (.A(index_q[0]), .Z(n25017)) /* synthesis lut_function=(!(A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i5507_1_lut_rep_457.init = 16'h5555;
    PFUMX i19225 (.BLUT(n21553), .ALUT(n21554), .C0(index_i[4]), .Z(n21555));
    LUT4 mux_192_Mux_6_i700_3_lut_4_lut (.A(n25166), .B(index_i[3]), .C(index_i[4]), 
         .D(n684_adj_2733), .Z(n700_adj_2714)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_6_i700_3_lut_4_lut.init = 16'h9f90;
    LUT4 mux_192_Mux_9_i364_3_lut_3_lut_4_lut (.A(index_i[0]), .B(n25116), 
         .C(index_i[3]), .D(n24985), .Z(n364_adj_2380)) /* synthesis lut_function=(!(A (C (D))+!A (B (C (D))+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_9_i364_3_lut_3_lut_4_lut.init = 16'h0efe;
    PFUMX i19456 (.BLUT(n21784), .ALUT(n21785), .C0(index_i[8]), .Z(n21786));
    LUT4 mux_193_Mux_2_i349_3_lut_3_lut (.A(index_q[0]), .B(index_q[4]), 
         .C(n348_adj_2539), .Z(n349_adj_2771)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_2_i349_3_lut_3_lut.init = 16'hd1d1;
    LUT4 mux_193_Mux_5_i573_3_lut_3_lut (.A(index_q[0]), .B(index_q[4]), 
         .C(n572_adj_2624), .Z(n573_adj_2684)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_5_i573_3_lut_3_lut.init = 16'hd1d1;
    LUT4 mux_193_Mux_2_i763_4_lut_4_lut (.A(index_q[0]), .B(n12093), .C(index_q[4]), 
         .D(n157_adj_2535), .Z(n763_adj_2779)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_2_i763_4_lut_4_lut.init = 16'hdfd0;
    LUT4 i11340_2_lut_rep_553 (.A(index_i[2]), .B(index_i[3]), .Z(n25113)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11340_2_lut_rep_553.init = 16'h8888;
    LUT4 i8007_3_lut_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), .C(index_i[1]), 
         .D(index_i[0]), .Z(n157_adj_2554)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(D))+!A !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i8007_3_lut_3_lut_4_lut.init = 16'h7780;
    LUT4 i15286_3_lut_3_lut_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n17549)) /* synthesis lut_function=(!(A (B (C)+!B !(C (D)+!C !(D)))+!A !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i15286_3_lut_3_lut_3_lut_4_lut.init = 16'h780f;
    LUT4 mux_192_Mux_7_i924_3_lut_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[4]), .D(n25163), .Z(n924_adj_2321)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_7_i924_3_lut_3_lut_4_lut.init = 16'h878f;
    LUT4 i11536_2_lut_rep_362_3_lut (.A(index_i[2]), .B(index_i[3]), .C(index_i[1]), 
         .Z(n24922)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11536_2_lut_rep_362_3_lut.init = 16'h8080;
    LUT4 mux_193_Mux_3_i700_3_lut_3_lut (.A(index_q[0]), .B(index_q[4]), 
         .C(n684_adj_2278), .Z(n700_adj_2739)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_3_i700_3_lut_3_lut.init = 16'h7474;
    LUT4 i18392_3_lut_3_lut_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[4]), .D(index_i[1]), .Z(n20722)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i18392_3_lut_3_lut_3_lut_4_lut.init = 16'h878f;
    LUT4 i15285_3_lut_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), .C(index_i[1]), 
         .D(index_i[0]), .Z(n17548)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i15285_3_lut_3_lut_4_lut.init = 16'hf078;
    LUT4 i9493_3_lut_3_lut_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n541_adj_2661)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9493_3_lut_3_lut_3_lut_4_lut.init = 16'h870f;
    LUT4 i11261_2_lut_rep_311_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[4]), .D(n25163), .Z(n24871)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11261_2_lut_rep_311_3_lut_4_lut.init = 16'hf8f0;
    LUT4 i9557_3_lut_4_lut_3_lut_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[0]), .D(index_i[1]), .Z(n875_adj_2279)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9557_3_lut_4_lut_3_lut_3_lut_4_lut.init = 16'h878f;
    LUT4 mux_192_Mux_6_i636_4_lut_4_lut (.A(index_i[1]), .B(index_i[4]), 
         .C(n635_adj_2476), .D(n14321), .Z(n636_adj_2713)) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_6_i636_4_lut_4_lut.init = 16'hf3d1;
    LUT4 i2_2_lut_rep_385_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), .C(index_i[1]), 
         .D(index_i[0]), .Z(n24945)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i2_2_lut_rep_385_3_lut_4_lut.init = 16'h8000;
    LUT4 i9543_3_lut_4_lut_4_lut (.A(index_q[0]), .B(n588), .C(index_q[4]), 
         .D(n25097), .Z(n12109)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B ((D)+!C)+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9543_3_lut_4_lut_4_lut.init = 16'h5c0c;
    LUT4 i18912_3_lut_4_lut_4_lut (.A(index_q[0]), .B(n25177), .C(index_q[3]), 
         .D(n25097), .Z(n21242)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18912_3_lut_4_lut_4_lut.init = 16'hc5c0;
    LUT4 i9539_2_lut_rep_405_3_lut (.A(index_i[2]), .B(index_i[3]), .C(index_i[4]), 
         .Z(n24965)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9539_2_lut_rep_405_3_lut.init = 16'h8080;
    PFUMX i15267 (.BLUT(n17528), .ALUT(n17529), .C0(index_q[4]), .Z(n17530));
    LUT4 i11646_2_lut_2_lut_3_lut (.A(index_i[2]), .B(index_i[3]), .C(index_i[0]), 
         .Z(n14321)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11646_2_lut_2_lut_3_lut.init = 16'h0808;
    LUT4 mux_193_Mux_2_i859_3_lut_4_lut_4_lut (.A(index_q[0]), .B(n25173), 
         .C(index_q[3]), .D(n25097), .Z(n859_adj_2310)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B ((D)+!C)+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_2_i859_3_lut_4_lut_4_lut.init = 16'h5c0c;
    LUT4 i12094_2_lut_rep_554 (.A(index_i[3]), .B(index_i[4]), .Z(n25114)) /* synthesis lut_function=(A (B)) */ ;
    defparam i12094_2_lut_rep_554.init = 16'h8888;
    LUT4 mux_192_Mux_1_i732_3_lut (.A(n716_adj_2332), .B(n491), .C(index_i[4]), 
         .Z(n732)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_1_i732_3_lut.init = 16'hcaca;
    LUT4 i18957_3_lut_3_lut_4_lut (.A(index_i[3]), .B(index_i[4]), .C(n413_adj_2407), 
         .D(index_i[5]), .Z(n21287)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(C+(D)))) */ ;
    defparam i18957_3_lut_3_lut_4_lut.init = 16'h77f0;
    LUT4 i9542_3_lut_3_lut_3_lut_4_lut (.A(index_i[3]), .B(index_i[4]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n444_adj_2766)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C))+!A (C))) */ ;
    defparam i9542_3_lut_3_lut_3_lut_4_lut.init = 16'h0f87;
    LUT4 mux_193_Mux_2_i507_3_lut_3_lut (.A(index_q[0]), .B(index_q[4]), 
         .C(n491_adj_2522), .Z(n507_adj_2776)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_2_i507_3_lut_3_lut.init = 16'h7474;
    LUT4 mux_193_Mux_4_i221_3_lut_3_lut (.A(index_q[0]), .B(index_q[4]), 
         .C(n205), .Z(n221_adj_2717)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_4_i221_3_lut_3_lut.init = 16'h7474;
    LUT4 quarter_wave_sample_register_i_13__I_0_3_lut (.A(quarter_wave_sample_register_i[13]), 
         .B(o_val_pipeline_i_0__15__N_2157[13]), .C(phase_negation_i[1]), 
         .Z(o_val_pipeline_i_0__15__N_2160)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[14] 77[8])
    defparam quarter_wave_sample_register_i_13__I_0_3_lut.init = 16'hcaca;
    LUT4 i20859_3_lut (.A(n20528), .B(n23637), .C(index_i[6]), .Z(n20537)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20859_3_lut.init = 16'hcaca;
    LUT4 i18779_3_lut_4_lut_4_lut (.A(index_q[0]), .B(n25180), .C(index_q[3]), 
         .D(n25211), .Z(n21109)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18779_3_lut_4_lut_4_lut.init = 16'hcfc5;
    LUT4 mux_193_Mux_4_i142_3_lut_4_lut_3_lut (.A(index_q[0]), .B(index_q[3]), 
         .C(index_q[2]), .Z(n142_adj_2749)) /* synthesis lut_function=(A (B (C))+!A !(B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_4_i142_3_lut_4_lut_3_lut.init = 16'h9595;
    LUT4 mux_192_Mux_0_i986_3_lut (.A(n25081), .B(n985_adj_2790), .C(index_i[3]), 
         .Z(n986_adj_2270)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_0_i986_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_0_i333_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n333)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B (D))) */ ;
    defparam mux_192_Mux_0_i333_3_lut_3_lut_4_lut.init = 16'hf10e;
    LUT4 mux_192_Mux_0_i971_3_lut (.A(n25087), .B(n25164), .C(index_i[3]), 
         .Z(n971_adj_2269)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_0_i971_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_0_i939_4_lut (.A(n978), .B(n25073), .C(index_i[3]), 
         .D(index_i[2]), .Z(n939_adj_2267)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_0_i939_4_lut.init = 16'hfaca;
    LUT4 mux_192_Mux_0_i923_3_lut (.A(n25041), .B(n27520), .C(index_i[3]), 
         .Z(n923_adj_2266)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_0_i923_3_lut.init = 16'hcaca;
    LUT4 i10954_2_lut_rep_462 (.A(index_q[0]), .B(index_q[1]), .Z(n25022)) /* synthesis lut_function=((B)+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i10954_2_lut_rep_462.init = 16'hdddd;
    LUT4 mux_193_Mux_4_i252_4_lut_4_lut (.A(index_q[0]), .B(index_q[3]), 
         .C(n25097), .D(index_q[4]), .Z(n252_adj_2718)) /* synthesis lut_function=(!(A (B (D)+!B !(D))+!A !(B ((D)+!C)+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_4_i252_4_lut_4_lut.init = 16'h669d;
    LUT4 mux_193_Mux_0_i635_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n635_adj_2796)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i635_3_lut_4_lut_4_lut.init = 16'hfd0a;
    LUT4 i9535_2_lut_rep_556 (.A(index_i[1]), .B(index_i[2]), .Z(n25116)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9535_2_lut_rep_556.init = 16'heeee;
    LUT4 i19330_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n21660)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (D))+!A !(D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19330_3_lut_4_lut_4_lut_4_lut.init = 16'ha25d;
    LUT4 mux_192_Mux_0_i46_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .D(index_i[3]), .Z(n46_adj_2741)) /* synthesis lut_function=(A ((D)+!B)+!A (B (D)+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_0_i46_3_lut_4_lut_4_lut_4_lut.init = 16'hfe33;
    LUT4 mux_193_Mux_3_i444_3_lut_4_lut (.A(index_q[0]), .B(index_q[3]), 
         .C(n25211), .D(index_q[4]), .Z(n444_adj_2735)) /* synthesis lut_function=(!(A (B (D)+!B (C (D)))+!A !(B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_3_i444_3_lut_4_lut.init = 16'h46aa;
    LUT4 n851_bdd_3_lut_22831_4_lut_4_lut (.A(index_q[0]), .B(index_q[2]), 
         .C(index_q[1]), .D(index_q[3]), .Z(n23836)) /* synthesis lut_function=(A (B+!((D)+!C))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n851_bdd_3_lut_22831_4_lut_4_lut.init = 16'h99b9;
    LUT4 i2_3_lut_4_lut_adj_82 (.A(index_i[5]), .B(index_i[6]), .C(index_i[7]), 
         .D(n25114), .Z(n19504)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i2_3_lut_4_lut_adj_82.init = 16'hfffe;
    LUT4 i11555_2_lut_rep_338_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[0]), 
         .Z(n24898)) /* synthesis lut_function=(A (C)+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11555_2_lut_rep_338_3_lut.init = 16'hf1f1;
    LUT4 i11284_2_lut_rep_360_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[3]), 
         .Z(n24920)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11284_2_lut_rep_360_3_lut.init = 16'he0e0;
    LUT4 mux_192_Mux_4_i236_3_lut_4_lut_3_lut_rep_475_4_lut (.A(index_i[1]), 
         .B(index_i[2]), .C(index_i[3]), .D(index_i[0]), .Z(n25035)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_4_i236_3_lut_4_lut_3_lut_rep_475_4_lut.init = 16'hf01f;
    LUT4 i18082_3_lut (.A(n24165), .B(n20403), .C(index_q[6]), .Z(n20412)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18082_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_9_i93_3_lut_3_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .Z(n93_adj_2388)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_9_i93_3_lut_3_lut_3_lut.init = 16'hc1c1;
    LUT4 mux_192_Mux_0_i716_3_lut (.A(n25086), .B(n25069), .C(index_i[3]), 
         .Z(n716)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_0_i716_3_lut.init = 16'hcaca;
    LUT4 i11419_2_lut_rep_409_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[0]), 
         .Z(n24969)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11419_2_lut_rep_409_3_lut.init = 16'hfefe;
    LUT4 i12289_2_lut_rep_298_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[4]), .D(index_i[3]), .Z(n24858)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i12289_2_lut_rep_298_3_lut_4_lut.init = 16'hfef0;
    LUT4 i19052_3_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[3]), 
         .D(index_i[0]), .Z(n21382)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19052_3_lut_3_lut_4_lut.init = 16'h0fe0;
    LUT4 i20785_3_lut (.A(n12008), .B(n892), .C(index_q[6]), .Z(n21305)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20785_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_4_i491_3_lut_4_lut_4_lut (.A(index_q[2]), .B(n25194), 
         .C(index_q[3]), .D(n25054), .Z(n491_adj_2617)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_4_i491_3_lut_4_lut_4_lut.init = 16'hfc5c;
    LUT4 mux_192_Mux_2_i173_3_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n173_adj_2707)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_2_i173_3_lut_3_lut_4_lut.init = 16'h0e1e;
    LUT4 mux_192_Mux_5_i954_3_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n954_adj_2758)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B (C)+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_5_i954_3_lut_4_lut_4_lut.init = 16'h0c1c;
    LUT4 mux_193_Mux_0_i923_3_lut (.A(n25196), .B(n27521), .C(index_q[3]), 
         .Z(n923)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i923_3_lut.init = 16'hcaca;
    LUT4 i18940_3_lut (.A(n21257), .B(n24078), .C(index_q[6]), .Z(n21270)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18940_3_lut.init = 16'hcaca;
    LUT4 i18939_3_lut (.A(n24058), .B(n21256), .C(index_q[6]), .Z(n21269)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18939_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_0_i526_3_lut (.A(n25204), .B(n25180), .C(index_q[3]), 
         .Z(n526_adj_2261)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i526_3_lut.init = 16'hcaca;
    LUT4 n10509_bdd_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[4]), .D(index_i[3]), .Z(n24733)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C+(D)))+!A (B (C (D)+!C !(D))+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n10509_bdd_3_lut_4_lut_4_lut_4_lut.init = 16'hc10f;
    LUT4 mux_192_Mux_0_i653_3_lut (.A(n24941), .B(n25077), .C(index_i[3]), 
         .Z(n653)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_0_i653_3_lut.init = 16'hcaca;
    LUT4 i20876_3_lut (.A(n27397), .B(n24046), .C(index_q[6]), .Z(n21268)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20876_3_lut.init = 16'hcaca;
    LUT4 i11294_2_lut_rep_323_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n24883)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11294_2_lut_rep_323_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i20799_3_lut (.A(n12048), .B(n892_adj_2663), .C(index_i[6]), 
         .Z(n21173)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20799_3_lut.init = 16'hcaca;
    LUT4 mux_192_Mux_9_i285_3_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n285_adj_2639)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_9_i285_3_lut_4_lut_4_lut.init = 16'hc0c1;
    LUT4 mux_192_Mux_8_i716_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .D(index_i[3]), .Z(n716_adj_2720)) /* synthesis lut_function=(!(A (B (D))+!A (B (D)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_8_i716_3_lut_4_lut_4_lut_4_lut.init = 16'h33fe;
    LUT4 i19230_3_lut_3_lut_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[3]), 
         .Z(n21560)) /* synthesis lut_function=(A (C)+!A (B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19230_3_lut_3_lut_3_lut.init = 16'he5e5;
    LUT4 mux_193_Mux_5_i924_4_lut_3_lut (.A(index_q[2]), .B(n14799), .C(index_q[4]), 
         .Z(n924_adj_2466)) /* synthesis lut_function=(!(A (B+(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_5_i924_4_lut_3_lut.init = 16'h5656;
    PFUMX i19329 (.BLUT(n21657), .ALUT(n21658), .C0(index_q[4]), .Z(n21659));
    LUT4 i18816_3_lut (.A(n24014), .B(n24021), .C(index_i[6]), .Z(n21146)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18816_3_lut.init = 16'hcaca;
    L6MUX21 i18607 (.D0(n20929), .D1(n20930), .SD(index_q[7]), .Z(n20937));
    LUT4 i21004_2_lut_rep_465 (.A(index_q[1]), .B(index_q[2]), .Z(n25025)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i21004_2_lut_rep_465.init = 16'h9999;
    LUT4 mux_192_Mux_0_i620_3_lut (.A(n25165), .B(n25066), .C(index_i[3]), 
         .Z(n620)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_192_Mux_0_i620_3_lut.init = 16'hcaca;
    LUT4 i18815_3_lut (.A(n23998), .B(n21132), .C(index_i[6]), .Z(n21145)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18815_3_lut.init = 16'hcaca;
    LUT4 n262_bdd_2_lut_22539_3_lut (.A(index_q[1]), .B(index_q[2]), .C(index_q[3]), 
         .Z(n24169)) /* synthesis lut_function=(A (B+(C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n262_bdd_2_lut_22539_3_lut.init = 16'hf9f9;
    LUT4 i20883_3_lut (.A(n27412), .B(n23990), .C(index_i[6]), .Z(n21144)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20883_3_lut.init = 16'hcaca;
    LUT4 mux_193_Mux_0_i93_3_lut_3_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .Z(n93_adj_2731)) /* synthesis lut_function=(A (B)+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_193_Mux_0_i93_3_lut_3_lut.init = 16'h9c9c;
    LUT4 i12242_2_lut_rep_466 (.A(index_q[2]), .B(index_q[0]), .Z(n25026)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i12242_2_lut_rep_466.init = 16'heeee;
    LUT4 i15298_3_lut_4_lut (.A(index_q[2]), .B(index_q[0]), .C(n25042), 
         .D(index_q[4]), .Z(n286_adj_2774)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;
    defparam i15298_3_lut_4_lut.init = 16'hfe00;
    LUT4 mux_192_Mux_8_i653_3_lut_rep_255_3_lut_4_lut (.A(index_i[0]), .B(n25122), 
         .C(n24985), .D(index_i[3]), .Z(n24815)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(C+(D)))) */ ;
    defparam mux_192_Mux_8_i653_3_lut_rep_255_3_lut_4_lut.init = 16'h77f0;
    L6MUX21 i22054 (.D0(n23655), .D1(n23652), .SD(index_i[5]), .Z(n23656));
    PFUMX i22052 (.BLUT(n23654), .ALUT(n23653), .C0(index_i[4]), .Z(n23655));
    PFUMX i22049 (.BLUT(n23651), .ALUT(n24847), .C0(index_i[4]), .Z(n23652));
    PFUMX i19332 (.BLUT(n21660), .ALUT(n21661), .C0(index_q[4]), .Z(n21662));
    L6MUX21 i22047 (.D0(n23649), .D1(n23647), .SD(index_i[4]), .Z(n23650));
    PFUMX i22045 (.BLUT(n24859), .ALUT(n23648), .C0(index_i[5]), .Z(n23649));
    LUT4 i17994_3_lut (.A(n20319), .B(n20320), .C(index_q[7]), .Z(n20324)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i17994_3_lut.init = 16'hcaca;
    PFUMX i22043 (.BLUT(n23646), .ALUT(n23645), .C0(index_i[5]), .Z(n23647));
    PFUMX i18692 (.BLUT(n21020), .ALUT(n21021), .C0(index_i[8]), .Z(n21022));
    LUT4 i12121_2_lut_rep_471 (.A(index_i[2]), .B(index_i[0]), .Z(n25031)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i12121_2_lut_rep_471.init = 16'heeee;
    LUT4 i15296_3_lut_4_lut (.A(index_i[2]), .B(index_i[0]), .C(n25063), 
         .D(index_i[4]), .Z(n286_adj_2778)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;
    defparam i15296_3_lut_4_lut.init = 16'hfe00;
    L6MUX21 i22035 (.D0(n23636), .D1(n23634), .SD(index_i[5]), .Z(n23637));
    PFUMX i22033 (.BLUT(n572_adj_2786), .ALUT(n23635), .C0(index_i[4]), 
          .Z(n23636));
    PFUMX i22031 (.BLUT(n23633), .ALUT(n23632), .C0(index_i[4]), .Z(n23634));
    L6MUX21 i22029 (.D0(n24802), .D1(n23627), .SD(index_i[4]), .Z(n23631));
    LUT4 i21092_2_lut_rep_472 (.A(index_i[4]), .B(index_i[3]), .Z(n25032)) /* synthesis lut_function=(A+!(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i21092_2_lut_rep_472.init = 16'hbbbb;
    LUT4 i20753_3_lut_4_lut (.A(index_i[4]), .B(index_i[3]), .C(n25245), 
         .D(n746_adj_2794), .Z(n763)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20753_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i11292_2_lut_rep_425_3_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .Z(n24985)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i11292_2_lut_rep_425_3_lut.init = 16'he0e0;
    LUT4 i11386_2_lut_rep_473 (.A(index_i[2]), .B(index_i[0]), .Z(n25033)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11386_2_lut_rep_473.init = 16'h8888;
    LUT4 i1_2_lut_rep_293_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[4]), 
         .D(index_q[2]), .Z(n24853)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_2_lut_rep_293_3_lut_4_lut.init = 16'hf080;
    LUT4 n250_bdd_3_lut_3_lut_4_lut_4_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n24244)) /* synthesis lut_function=(A (B (C)+!B !(D))+!A !(D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n250_bdd_3_lut_3_lut_4_lut_4_lut_3_lut_4_lut.init = 16'h80f7;
    L6MUX21 i21378 (.D0(n22894), .D1(n22892), .SD(index_i[6]), .Z(n22895));
    PFUMX i21374 (.BLUT(n62_adj_2348), .ALUT(n22891), .C0(index_i[5]), 
          .Z(n22892));
    LUT4 mux_192_Mux_7_i141_3_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n141)) /* synthesis lut_function=(A ((C)+!B)+!A (B+!(C))) */ ;
    defparam mux_192_Mux_7_i141_3_lut_4_lut_3_lut.init = 16'he7e7;
    PFUMX i19345 (.BLUT(n21673), .ALUT(n21674), .C0(index_q[4]), .Z(n21675));
    PFUMX i19347 (.BLUT(n557_adj_2603), .ALUT(n572_adj_2772), .C0(index_q[4]), 
          .Z(n21677));
    PFUMX i22025 (.BLUT(n23626), .ALUT(n23625), .C0(index_i[5]), .Z(n23627));
    PFUMX i19348 (.BLUT(n589_adj_2324), .ALUT(n604_adj_2335), .C0(index_q[4]), 
          .Z(n21678));
    PFUMX i19349 (.BLUT(n620_adj_2322), .ALUT(n635_adj_2796), .C0(index_q[4]), 
          .Z(n21679));
    PFUMX i19350 (.BLUT(n653_adj_2320), .ALUT(n668_adj_2610), .C0(index_q[4]), 
          .Z(n21680));
    CCU2D add_358_13 (.A0(quarter_wave_sample_register_q[12]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_q[13]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17304), .COUT(n17305), 
          .S0(o_val_pipeline_q_0__15__N_2189[12]), .S1(o_val_pipeline_q_0__15__N_2189[13]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(80[29:60])
    defparam add_358_13.INIT0 = 16'hf555;
    defparam add_358_13.INIT1 = 16'hf555;
    defparam add_358_13.INJECT1_0 = "NO";
    defparam add_358_13.INJECT1_1 = "NO";
    PFUMX i19351 (.BLUT(n684_adj_2488), .ALUT(n699_adj_2598), .C0(index_q[4]), 
          .Z(n21681));
    PFUMX i19352 (.BLUT(n716_adj_2318), .ALUT(n731_adj_2746), .C0(index_q[4]), 
          .Z(n21682));
    PFUMX i18754 (.BLUT(n21082), .ALUT(n21083), .C0(index_q[8]), .Z(n21084));
    PFUMX i21376 (.BLUT(n22893), .ALUT(n20990), .C0(index_i[5]), .Z(n22894));
    L6MUX21 i21369 (.D0(n22877), .D1(n22875), .SD(index_q[6]), .Z(n22878));
    PFUMX i21367 (.BLUT(n22876), .ALUT(n20899), .C0(index_q[5]), .Z(n22877));
    PFUMX i19353 (.BLUT(n747_adj_2503), .ALUT(n762_adj_2640), .C0(index_q[4]), 
          .Z(n21683));
    PFUMX i21365 (.BLUT(n62_adj_2319), .ALUT(n22874), .C0(index_q[5]), 
          .Z(n22875));
    PFUMX i19354 (.BLUT(n781_adj_2492), .ALUT(n796_adj_2286), .C0(index_q[4]), 
          .Z(n21684));
    PFUMX i19355 (.BLUT(n812_adj_2645), .ALUT(n11927), .C0(index_q[4]), 
          .Z(n21685));
    PFUMX i22013 (.BLUT(n23610), .ALUT(n27522), .C0(index_q[3]), .Z(n23611));
    PFUMX i18821 (.BLUT(n21143), .ALUT(n21144), .C0(index_i[7]), .Z(n21151));
    L6MUX21 i21350 (.D0(n22855), .D1(n24785), .SD(index_i[6]), .Z(n22856));
    
endmodule
//
// Verilog Description of module \nco(OW=12)_U1 
//

module \nco(OW=12)_U1  (increment, o_phase, GND_net, i_ref_clk_c, i_resetb_N_301) /* synthesis syn_module_defined=1 */ ;
    input [30:0]increment;
    output [11:0]o_phase;
    input GND_net;
    input i_ref_clk_c;
    input i_resetb_N_301;
    
    wire i_ref_clk_c /* synthesis SET_AS_NETWORK=i_ref_clk_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(22[12:21])
    
    wire n17448;
    wire [31:0]n133;
    
    wire n17449, n17447;
    wire [31:0]n233;
    
    wire n17446, n17445, n17444, n17443, n17442, n17441, n17440, 
        n17439, n17453, n17452, n17451, n17450;
    
    CCU2D phase_register_505_add_4_22 (.A0(increment[20]), .B0(o_phase[0]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[21]), .B1(o_phase[1]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17448), .COUT(n17449), .S0(n133[20]), 
          .S1(n133[21]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_505_add_4_22.INIT0 = 16'h5666;
    defparam phase_register_505_add_4_22.INIT1 = 16'h5666;
    defparam phase_register_505_add_4_22.INJECT1_0 = "NO";
    defparam phase_register_505_add_4_22.INJECT1_1 = "NO";
    CCU2D phase_register_505_add_4_20 (.A0(increment[18]), .B0(n233[18]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[19]), .B1(n233[19]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17447), .COUT(n17448), .S0(n133[18]), 
          .S1(n133[19]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_505_add_4_20.INIT0 = 16'h5666;
    defparam phase_register_505_add_4_20.INIT1 = 16'h5666;
    defparam phase_register_505_add_4_20.INJECT1_0 = "NO";
    defparam phase_register_505_add_4_20.INJECT1_1 = "NO";
    CCU2D phase_register_505_add_4_18 (.A0(increment[16]), .B0(n233[16]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[17]), .B1(n233[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17446), .COUT(n17447), .S0(n133[16]), 
          .S1(n133[17]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_505_add_4_18.INIT0 = 16'h5666;
    defparam phase_register_505_add_4_18.INIT1 = 16'h5666;
    defparam phase_register_505_add_4_18.INJECT1_0 = "NO";
    defparam phase_register_505_add_4_18.INJECT1_1 = "NO";
    CCU2D phase_register_505_add_4_16 (.A0(increment[14]), .B0(n233[14]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[15]), .B1(n233[15]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17445), .COUT(n17446), .S0(n133[14]), 
          .S1(n133[15]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_505_add_4_16.INIT0 = 16'h5666;
    defparam phase_register_505_add_4_16.INIT1 = 16'h5666;
    defparam phase_register_505_add_4_16.INJECT1_0 = "NO";
    defparam phase_register_505_add_4_16.INJECT1_1 = "NO";
    CCU2D phase_register_505_add_4_14 (.A0(increment[12]), .B0(n233[12]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[13]), .B1(n233[13]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17444), .COUT(n17445), .S0(n133[12]), 
          .S1(n133[13]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_505_add_4_14.INIT0 = 16'h5666;
    defparam phase_register_505_add_4_14.INIT1 = 16'h5666;
    defparam phase_register_505_add_4_14.INJECT1_0 = "NO";
    defparam phase_register_505_add_4_14.INJECT1_1 = "NO";
    CCU2D phase_register_505_add_4_12 (.A0(increment[10]), .B0(n233[10]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[11]), .B1(n233[11]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17443), .COUT(n17444), .S0(n133[10]), 
          .S1(n133[11]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_505_add_4_12.INIT0 = 16'h5666;
    defparam phase_register_505_add_4_12.INIT1 = 16'h5666;
    defparam phase_register_505_add_4_12.INJECT1_0 = "NO";
    defparam phase_register_505_add_4_12.INJECT1_1 = "NO";
    CCU2D phase_register_505_add_4_10 (.A0(increment[8]), .B0(n233[8]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[9]), .B1(n233[9]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17442), .COUT(n17443), .S0(n133[8]), 
          .S1(n133[9]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_505_add_4_10.INIT0 = 16'h5666;
    defparam phase_register_505_add_4_10.INIT1 = 16'h5666;
    defparam phase_register_505_add_4_10.INJECT1_0 = "NO";
    defparam phase_register_505_add_4_10.INJECT1_1 = "NO";
    CCU2D phase_register_505_add_4_8 (.A0(increment[6]), .B0(n233[6]), .C0(GND_net), 
          .D0(GND_net), .A1(increment[7]), .B1(n233[7]), .C1(GND_net), 
          .D1(GND_net), .CIN(n17441), .COUT(n17442), .S0(n133[6]), .S1(n133[7]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_505_add_4_8.INIT0 = 16'h5666;
    defparam phase_register_505_add_4_8.INIT1 = 16'h5666;
    defparam phase_register_505_add_4_8.INJECT1_0 = "NO";
    defparam phase_register_505_add_4_8.INJECT1_1 = "NO";
    CCU2D phase_register_505_add_4_6 (.A0(increment[4]), .B0(n233[4]), .C0(GND_net), 
          .D0(GND_net), .A1(increment[5]), .B1(n233[5]), .C1(GND_net), 
          .D1(GND_net), .CIN(n17440), .COUT(n17441), .S0(n133[4]), .S1(n133[5]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_505_add_4_6.INIT0 = 16'h5666;
    defparam phase_register_505_add_4_6.INIT1 = 16'h5666;
    defparam phase_register_505_add_4_6.INJECT1_0 = "NO";
    defparam phase_register_505_add_4_6.INJECT1_1 = "NO";
    CCU2D phase_register_505_add_4_4 (.A0(increment[2]), .B0(n233[2]), .C0(GND_net), 
          .D0(GND_net), .A1(increment[3]), .B1(n233[3]), .C1(GND_net), 
          .D1(GND_net), .CIN(n17439), .COUT(n17440), .S0(n133[2]), .S1(n133[3]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_505_add_4_4.INIT0 = 16'h5666;
    defparam phase_register_505_add_4_4.INIT1 = 16'h5666;
    defparam phase_register_505_add_4_4.INJECT1_0 = "NO";
    defparam phase_register_505_add_4_4.INJECT1_1 = "NO";
    CCU2D phase_register_505_add_4_2 (.A0(increment[0]), .B0(n233[0]), .C0(GND_net), 
          .D0(GND_net), .A1(increment[1]), .B1(n233[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n17439), .S1(n133[1]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_505_add_4_2.INIT0 = 16'h7000;
    defparam phase_register_505_add_4_2.INIT1 = 16'h5666;
    defparam phase_register_505_add_4_2.INJECT1_0 = "NO";
    defparam phase_register_505_add_4_2.INJECT1_1 = "NO";
    FD1S3DX phase_register_505__i0 (.D(n133[0]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(n233[0])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_505__i0.GSR = "DISABLED";
    LUT4 i15209_2_lut (.A(increment[0]), .B(n233[0]), .Z(n133[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i15209_2_lut.init = 16'h6666;
    CCU2D phase_register_505_add_4_32 (.A0(increment[30]), .B0(o_phase[10]), 
          .C0(GND_net), .D0(GND_net), .A1(o_phase[11]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n17453), .S0(n133[30]), .S1(n133[31]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_505_add_4_32.INIT0 = 16'h5666;
    defparam phase_register_505_add_4_32.INIT1 = 16'hfaaa;
    defparam phase_register_505_add_4_32.INJECT1_0 = "NO";
    defparam phase_register_505_add_4_32.INJECT1_1 = "NO";
    FD1S3DX phase_register_505__i31 (.D(n133[31]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(o_phase[11])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_505__i31.GSR = "DISABLED";
    FD1S3DX phase_register_505__i30 (.D(n133[30]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(o_phase[10])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_505__i30.GSR = "DISABLED";
    FD1S3DX phase_register_505__i29 (.D(n133[29]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(o_phase[9])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_505__i29.GSR = "DISABLED";
    FD1S3DX phase_register_505__i28 (.D(n133[28]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(o_phase[8])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_505__i28.GSR = "DISABLED";
    FD1S3DX phase_register_505__i27 (.D(n133[27]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(o_phase[7])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_505__i27.GSR = "DISABLED";
    FD1S3DX phase_register_505__i26 (.D(n133[26]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(o_phase[6])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_505__i26.GSR = "DISABLED";
    FD1S3DX phase_register_505__i25 (.D(n133[25]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(o_phase[5])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_505__i25.GSR = "DISABLED";
    FD1S3DX phase_register_505__i24 (.D(n133[24]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(o_phase[4])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_505__i24.GSR = "DISABLED";
    FD1S3DX phase_register_505__i23 (.D(n133[23]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(o_phase[3])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_505__i23.GSR = "DISABLED";
    FD1S3DX phase_register_505__i22 (.D(n133[22]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(o_phase[2])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_505__i22.GSR = "DISABLED";
    FD1S3DX phase_register_505__i21 (.D(n133[21]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(o_phase[1])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_505__i21.GSR = "DISABLED";
    FD1S3DX phase_register_505__i20 (.D(n133[20]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(o_phase[0])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_505__i20.GSR = "DISABLED";
    FD1S3DX phase_register_505__i19 (.D(n133[19]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(n233[19])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_505__i19.GSR = "DISABLED";
    FD1S3DX phase_register_505__i18 (.D(n133[18]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(n233[18])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_505__i18.GSR = "DISABLED";
    FD1S3DX phase_register_505__i17 (.D(n133[17]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(n233[17])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_505__i17.GSR = "DISABLED";
    FD1S3DX phase_register_505__i16 (.D(n133[16]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(n233[16])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_505__i16.GSR = "DISABLED";
    FD1S3DX phase_register_505__i15 (.D(n133[15]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(n233[15])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_505__i15.GSR = "DISABLED";
    FD1S3DX phase_register_505__i14 (.D(n133[14]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(n233[14])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_505__i14.GSR = "DISABLED";
    FD1S3DX phase_register_505__i13 (.D(n133[13]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(n233[13])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_505__i13.GSR = "DISABLED";
    FD1S3DX phase_register_505__i12 (.D(n133[12]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(n233[12])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_505__i12.GSR = "DISABLED";
    FD1S3DX phase_register_505__i11 (.D(n133[11]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(n233[11])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_505__i11.GSR = "DISABLED";
    FD1S3DX phase_register_505__i10 (.D(n133[10]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(n233[10])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_505__i10.GSR = "DISABLED";
    FD1S3DX phase_register_505__i9 (.D(n133[9]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(n233[9])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_505__i9.GSR = "DISABLED";
    FD1S3DX phase_register_505__i8 (.D(n133[8]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(n233[8])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_505__i8.GSR = "DISABLED";
    FD1S3DX phase_register_505__i7 (.D(n133[7]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(n233[7])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_505__i7.GSR = "DISABLED";
    FD1S3DX phase_register_505__i6 (.D(n133[6]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(n233[6])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_505__i6.GSR = "DISABLED";
    FD1S3DX phase_register_505__i5 (.D(n133[5]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(n233[5])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_505__i5.GSR = "DISABLED";
    FD1S3DX phase_register_505__i4 (.D(n133[4]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(n233[4])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_505__i4.GSR = "DISABLED";
    FD1S3DX phase_register_505__i3 (.D(n133[3]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(n233[3])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_505__i3.GSR = "DISABLED";
    FD1S3DX phase_register_505__i2 (.D(n133[2]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(n233[2])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_505__i2.GSR = "DISABLED";
    FD1S3DX phase_register_505__i1 (.D(n133[1]), .CK(i_ref_clk_c), .CD(i_resetb_N_301), 
            .Q(n233[1])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_505__i1.GSR = "DISABLED";
    CCU2D phase_register_505_add_4_30 (.A0(increment[28]), .B0(o_phase[8]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[29]), .B1(o_phase[9]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17452), .COUT(n17453), .S0(n133[28]), 
          .S1(n133[29]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_505_add_4_30.INIT0 = 16'h5666;
    defparam phase_register_505_add_4_30.INIT1 = 16'h5666;
    defparam phase_register_505_add_4_30.INJECT1_0 = "NO";
    defparam phase_register_505_add_4_30.INJECT1_1 = "NO";
    CCU2D phase_register_505_add_4_28 (.A0(increment[26]), .B0(o_phase[6]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[27]), .B1(o_phase[7]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17451), .COUT(n17452), .S0(n133[26]), 
          .S1(n133[27]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_505_add_4_28.INIT0 = 16'h5666;
    defparam phase_register_505_add_4_28.INIT1 = 16'h5666;
    defparam phase_register_505_add_4_28.INJECT1_0 = "NO";
    defparam phase_register_505_add_4_28.INJECT1_1 = "NO";
    CCU2D phase_register_505_add_4_26 (.A0(increment[24]), .B0(o_phase[4]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[25]), .B1(o_phase[5]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17450), .COUT(n17451), .S0(n133[24]), 
          .S1(n133[25]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_505_add_4_26.INIT0 = 16'h5666;
    defparam phase_register_505_add_4_26.INIT1 = 16'h5666;
    defparam phase_register_505_add_4_26.INJECT1_0 = "NO";
    defparam phase_register_505_add_4_26.INJECT1_1 = "NO";
    CCU2D phase_register_505_add_4_24 (.A0(increment[22]), .B0(o_phase[2]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[23]), .B1(o_phase[3]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17449), .COUT(n17450), .S0(n133[22]), 
          .S1(n133[23]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_505_add_4_24.INIT0 = 16'h5666;
    defparam phase_register_505_add_4_24.INIT1 = 16'h5666;
    defparam phase_register_505_add_4_24.INJECT1_0 = "NO";
    defparam phase_register_505_add_4_24.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module efb_inst
//

module efb_inst (i_ref_clk_c, i_resetb_N_301, n27585, wb_lo_data_7__N_96, 
            wb_we, \wb_addr[7] , \wb_addr[6] , \wb_addr[5] , \wb_addr[4] , 
            \wb_addr[3] , \wb_addr[2] , \wb_addr[1] , \wb_addr[0] , 
            \wb_odata[7] , \wb_odata[6] , \wb_odata[5] , \wb_odata[4] , 
            \wb_odata[3] , \wb_odata[2] , \wb_odata[1] , \wb_odata[0] , 
            pll_data_o, pll_ack, wb_lo_data, wb_lo_ack, pll_clk, pll_rst, 
            pll_stb, pll_we, pll_addr, pll_data_i, GND_net, VCC_net) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;
    input i_ref_clk_c;
    input i_resetb_N_301;
    input n27585;
    input wb_lo_data_7__N_96;
    input wb_we;
    input \wb_addr[7] ;
    input \wb_addr[6] ;
    input \wb_addr[5] ;
    input \wb_addr[4] ;
    input \wb_addr[3] ;
    input \wb_addr[2] ;
    input \wb_addr[1] ;
    input \wb_addr[0] ;
    input \wb_odata[7] ;
    input \wb_odata[6] ;
    input \wb_odata[5] ;
    input \wb_odata[4] ;
    input \wb_odata[3] ;
    input \wb_odata[2] ;
    input \wb_odata[1] ;
    input \wb_odata[0] ;
    input [7:0]pll_data_o;
    input pll_ack;
    output [7:0]wb_lo_data;
    output wb_lo_ack;
    output pll_clk;
    output pll_rst;
    output pll_stb;
    output pll_we;
    output [4:0]pll_addr;
    output [7:0]pll_data_i;
    input GND_net;
    input VCC_net;
    
    wire i_ref_clk_c /* synthesis SET_AS_NETWORK=i_ref_clk_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(22[12:21])
    
    EFB EFBInst_0 (.WBCLKI(i_ref_clk_c), .WBRSTI(i_resetb_N_301), .WBCYCI(n27585), 
        .WBSTBI(wb_lo_data_7__N_96), .WBWEI(wb_we), .WBADRI0(\wb_addr[0] ), 
        .WBADRI1(\wb_addr[1] ), .WBADRI2(\wb_addr[2] ), .WBADRI3(\wb_addr[3] ), 
        .WBADRI4(\wb_addr[4] ), .WBADRI5(\wb_addr[5] ), .WBADRI6(\wb_addr[6] ), 
        .WBADRI7(\wb_addr[7] ), .WBDATI0(\wb_odata[0] ), .WBDATI1(\wb_odata[1] ), 
        .WBDATI2(\wb_odata[2] ), .WBDATI3(\wb_odata[3] ), .WBDATI4(\wb_odata[4] ), 
        .WBDATI5(\wb_odata[5] ), .WBDATI6(\wb_odata[6] ), .WBDATI7(\wb_odata[7] ), 
        .I2C1SCLI(GND_net), .I2C1SDAI(GND_net), .I2C2SCLI(GND_net), .I2C2SDAI(GND_net), 
        .SPISCKI(GND_net), .SPIMISOI(GND_net), .SPIMOSII(GND_net), .SPISCSN(GND_net), 
        .TCCLKI(GND_net), .TCRSTN(GND_net), .TCIC(GND_net), .UFMSN(VCC_net), 
        .PLL0DATI0(pll_data_o[0]), .PLL0DATI1(pll_data_o[1]), .PLL0DATI2(pll_data_o[2]), 
        .PLL0DATI3(pll_data_o[3]), .PLL0DATI4(pll_data_o[4]), .PLL0DATI5(pll_data_o[5]), 
        .PLL0DATI6(pll_data_o[6]), .PLL0DATI7(pll_data_o[7]), .PLL0ACKI(pll_ack), 
        .PLL1DATI0(GND_net), .PLL1DATI1(GND_net), .PLL1DATI2(GND_net), 
        .PLL1DATI3(GND_net), .PLL1DATI4(GND_net), .PLL1DATI5(GND_net), 
        .PLL1DATI6(GND_net), .PLL1DATI7(GND_net), .PLL1ACKI(GND_net), 
        .WBDATO0(wb_lo_data[0]), .WBDATO1(wb_lo_data[1]), .WBDATO2(wb_lo_data[2]), 
        .WBDATO3(wb_lo_data[3]), .WBDATO4(wb_lo_data[4]), .WBDATO5(wb_lo_data[5]), 
        .WBDATO6(wb_lo_data[6]), .WBDATO7(wb_lo_data[7]), .WBACKO(wb_lo_ack), 
        .PLLCLKO(pll_clk), .PLLRSTO(pll_rst), .PLL0STBO(pll_stb), .PLLWEO(pll_we), 
        .PLLADRO0(pll_addr[0]), .PLLADRO1(pll_addr[1]), .PLLADRO2(pll_addr[2]), 
        .PLLADRO3(pll_addr[3]), .PLLADRO4(pll_addr[4]), .PLLDATO0(pll_data_i[0]), 
        .PLLDATO1(pll_data_i[1]), .PLLDATO2(pll_data_i[2]), .PLLDATO3(pll_data_i[3]), 
        .PLLDATO4(pll_data_i[4]), .PLLDATO5(pll_data_i[5]), .PLLDATO6(pll_data_i[6]), 
        .PLLDATO7(pll_data_i[7])) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=8, LSE_LCOL=10, LSE_RCOL=3, LSE_LLINE=179, LSE_RLINE=191 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(179[10] 191[3])
    defparam EFBInst_0.EFB_I2C1 = "DISABLED";
    defparam EFBInst_0.EFB_I2C2 = "DISABLED";
    defparam EFBInst_0.EFB_SPI = "DISABLED";
    defparam EFBInst_0.EFB_TC = "DISABLED";
    defparam EFBInst_0.EFB_TC_PORTMODE = "WB";
    defparam EFBInst_0.EFB_UFM = "DISABLED";
    defparam EFBInst_0.EFB_WB_CLK_FREQ = "50.0";
    defparam EFBInst_0.DEV_DENSITY = "6900L";
    defparam EFBInst_0.UFM_INIT_PAGES = 0;
    defparam EFBInst_0.UFM_INIT_START_PAGE = 0;
    defparam EFBInst_0.UFM_INIT_ALL_ZEROS = "ENABLED";
    defparam EFBInst_0.UFM_INIT_FILE_NAME = "NONE";
    defparam EFBInst_0.UFM_INIT_FILE_FORMAT = "HEX";
    defparam EFBInst_0.I2C1_ADDRESSING = "7BIT";
    defparam EFBInst_0.I2C2_ADDRESSING = "7BIT";
    defparam EFBInst_0.I2C1_SLAVE_ADDR = "0b1000001";
    defparam EFBInst_0.I2C2_SLAVE_ADDR = "0b1000010";
    defparam EFBInst_0.I2C1_BUS_PERF = "100kHz";
    defparam EFBInst_0.I2C2_BUS_PERF = "100kHz";
    defparam EFBInst_0.I2C1_CLK_DIVIDER = 1;
    defparam EFBInst_0.I2C2_CLK_DIVIDER = 1;
    defparam EFBInst_0.I2C1_GEN_CALL = "DISABLED";
    defparam EFBInst_0.I2C2_GEN_CALL = "DISABLED";
    defparam EFBInst_0.I2C1_WAKEUP = "DISABLED";
    defparam EFBInst_0.I2C2_WAKEUP = "DISABLED";
    defparam EFBInst_0.SPI_MODE = "MASTER";
    defparam EFBInst_0.SPI_CLK_DIVIDER = 1;
    defparam EFBInst_0.SPI_LSB_FIRST = "DISABLED";
    defparam EFBInst_0.SPI_CLK_INV = "DISABLED";
    defparam EFBInst_0.SPI_PHASE_ADJ = "DISABLED";
    defparam EFBInst_0.SPI_SLAVE_HANDSHAKE = "DISABLED";
    defparam EFBInst_0.SPI_INTR_TXRDY = "DISABLED";
    defparam EFBInst_0.SPI_INTR_RXRDY = "DISABLED";
    defparam EFBInst_0.SPI_INTR_TXOVR = "DISABLED";
    defparam EFBInst_0.SPI_INTR_RXOVR = "DISABLED";
    defparam EFBInst_0.SPI_WAKEUP = "DISABLED";
    defparam EFBInst_0.TC_MODE = "CTCM";
    defparam EFBInst_0.TC_SCLK_SEL = "PCLOCK";
    defparam EFBInst_0.TC_CCLK_SEL = 1;
    defparam EFBInst_0.GSR = "ENABLED";
    defparam EFBInst_0.TC_TOP_SET = 65535;
    defparam EFBInst_0.TC_OCR_SET = 32767;
    defparam EFBInst_0.TC_OC_MODE = "TOGGLE";
    defparam EFBInst_0.TC_RESETN = "ENABLED";
    defparam EFBInst_0.TC_TOP_SEL = "OFF";
    defparam EFBInst_0.TC_OV_INT = "OFF";
    defparam EFBInst_0.TC_OCR_INT = "OFF";
    defparam EFBInst_0.TC_ICR_INT = "OFF";
    defparam EFBInst_0.TC_OVERFLOW = "DISABLED";
    defparam EFBInst_0.TC_ICAPTURE = "DISABLED";
    
endmodule
//
// Verilog Description of module clock_phase_shifter
//

module clock_phase_shifter (q_clk_p_c, i_clk_2f_N_2249, q_clk_n_c, i_clk_p_c, 
            lo_pll_out, i_clk_n_c) /* synthesis syn_module_defined=1 */ ;
    output q_clk_p_c;
    input i_clk_2f_N_2249;
    input q_clk_n_c;
    output i_clk_p_c;
    input lo_pll_out;
    input i_clk_n_c;
    
    wire i_clk_2f_N_2249 /* synthesis is_inv_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/clock_phase_shifter.v(11[21:28])
    wire lo_pll_out /* synthesis is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(159[6:16])
    
    FD1S3AX o_clk_q_10 (.D(q_clk_n_c), .CK(i_clk_2f_N_2249), .Q(q_clk_p_c)) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=21, LSE_RCOL=2, LSE_LLINE=160, LSE_RLINE=164 */ ;   // d:/documents/git_local/fm_modulator/rtl/clock_phase_shifter.v(17[8] 19[4])
    defparam o_clk_q_10.GSR = "DISABLED";
    FD1S3AX o_clk_i_9 (.D(i_clk_n_c), .CK(lo_pll_out), .Q(i_clk_p_c)) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=21, LSE_RCOL=2, LSE_LLINE=160, LSE_RLINE=164 */ ;   // d:/documents/git_local/fm_modulator/rtl/clock_phase_shifter.v(13[8] 15[4])
    defparam o_clk_i_9.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module TSALL
// module not written out since it is a black-box. 
//

//
// Verilog Description of module \rxuartlite(CLOCKS_PER_BAUD=20) 
//

module \rxuartlite(CLOCKS_PER_BAUD=20)  (i_ref_clk_c, \rx_data[0] , rx_stb, 
            i_wbu_uart_rx_c, chg_counter, i_ref_clk_c_enable_180, chg_counter_23__N_406, 
            GND_net, \rx_data[6] , \rx_data[5] , \rx_data[4] , \rx_data[3] , 
            \rx_data[2] , \rx_data[1] ) /* synthesis syn_module_defined=1 */ ;
    input i_ref_clk_c;
    output \rx_data[0] ;
    output rx_stb;
    input i_wbu_uart_rx_c;
    output [23:0]chg_counter;
    input i_ref_clk_c_enable_180;
    output chg_counter_23__N_406;
    input GND_net;
    output \rx_data[6] ;
    output \rx_data[5] ;
    output \rx_data[4] ;
    output \rx_data[3] ;
    output \rx_data[2] ;
    output \rx_data[1] ;
    
    wire i_ref_clk_c /* synthesis SET_AS_NETWORK=i_ref_clk_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(22[12:21])
    
    wire qq_uart, q_uart, ck_uart, o_data_7__N_418;
    wire [7:0]data_reg;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(142[12:20])
    wire [3:0]state;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(75[13:18])
    
    wire i_ref_clk_c_enable_355;
    wire [3:0]state_3__N_322;
    
    wire half_baud_time, half_baud_time_N_457;
    wire [23:0]baud_counter;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(78[17:29])
    
    wire i_ref_clk_c_enable_416, n24981;
    wire [23:0]baud_counter_23__N_421;
    
    wire n25240, n25241;
    wire [23:0]n534;
    
    wire zero_baud_counter, i_ref_clk_c_enable_147, n14854, n24903, 
        n24886, n17337, half_baud_time_N_458, n17336, n17335, n17334, 
        n17333, n17332, n17331, n17330, n17329, n17328, n17327, 
        n17394;
    wire [23:0]n290;
    
    wire n17393, n17392, zero_baud_counter_N_454, n17391, n17390, 
        n17389, n17388, n17387, n17386, n17318, n17385, n17384, 
        n17383, n25014, n23729, n23728, n19721, n11693, n46, n19719, 
        n25, n19737, n19727, n19683, n19723, n19675, n17317, n17316, 
        state_3__N_415, n17315, n25013, n24845, n17314, n17313, 
        n17312, data_reg_7__N_416, n17311, n17310, n17309, n172, 
        n17705, i_ref_clk_c_enable_351, n17308, n17307;
    wire [3:0]n560;
    
    FD1S3AY qq_uart_70 (.D(q_uart), .CK(i_ref_clk_c), .Q(qq_uart)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(90[9] 91[66])
    defparam qq_uart_70.GSR = "DISABLED";
    FD1S3AY ck_uart_71 (.D(qq_uart), .CK(i_ref_clk_c), .Q(ck_uart)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(90[9] 91[66])
    defparam ck_uart_71.GSR = "DISABLED";
    FD1P3AX o_data__i1 (.D(data_reg[0]), .SP(o_data_7__N_418), .CK(i_ref_clk_c), 
            .Q(\rx_data[0] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(155[9] 161[18])
    defparam o_data__i1.GSR = "DISABLED";
    FD1P3AY state_i0 (.D(state_3__N_322[0]), .SP(i_ref_clk_c_enable_355), 
            .CK(i_ref_clk_c), .Q(state[0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(116[9] 134[5])
    defparam state_i0.GSR = "DISABLED";
    FD1S3AX half_baud_time_73 (.D(half_baud_time_N_457), .CK(i_ref_clk_c), 
            .Q(half_baud_time)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(111[9] 112[70])
    defparam half_baud_time_73.GSR = "DISABLED";
    FD1S3AX o_wr_76 (.D(o_data_7__N_418), .CK(i_ref_clk_c), .Q(rx_stb)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(155[9] 161[18])
    defparam o_wr_76.GSR = "DISABLED";
    FD1S3AY q_uart_69 (.D(i_wbu_uart_rx_c), .CK(i_ref_clk_c), .Q(q_uart)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(90[9] 91[66])
    defparam q_uart_69.GSR = "DISABLED";
    FD1P3JX baud_counter_i1 (.D(baud_counter_23__N_421[1]), .SP(i_ref_clk_c_enable_416), 
            .PD(n24981), .CK(i_ref_clk_c), .Q(baud_counter[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i1.GSR = "DISABLED";
    FD1P3JX baud_counter_i4 (.D(baud_counter_23__N_421[4]), .SP(i_ref_clk_c_enable_416), 
            .PD(n24981), .CK(i_ref_clk_c), .Q(baud_counter[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i4.GSR = "DISABLED";
    PFUMX i23022 (.BLUT(n25240), .ALUT(n25241), .C0(state[3]), .Z(state_3__N_322[3]));
    FD1P3IX chg_counter__i0 (.D(n534[0]), .SP(i_ref_clk_c_enable_180), .CD(chg_counter_23__N_406), 
            .CK(i_ref_clk_c), .Q(chg_counter[0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[34])
    defparam chg_counter__i0.GSR = "DISABLED";
    FD1P3AY zero_baud_counter_79 (.D(n14854), .SP(i_ref_clk_c_enable_147), 
            .CK(i_ref_clk_c), .Q(zero_baud_counter)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(187[9] 195[29])
    defparam zero_baud_counter_79.GSR = "DISABLED";
    LUT4 i2_3_lut_4_lut (.A(state[0]), .B(n24903), .C(zero_baud_counter), 
         .D(ck_uart), .Z(o_data_7__N_418)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(144[27:48])
    defparam i2_3_lut_4_lut.init = 16'h1000;
    LUT4 i2_3_lut_4_lut_adj_74 (.A(n24981), .B(n24886), .C(state[3]), 
         .D(zero_baud_counter), .Z(i_ref_clk_c_enable_416)) /* synthesis lut_function=(A+!(B (C (D)))) */ ;
    defparam i2_3_lut_4_lut_adj_74.init = 16'hbfff;
    FD1P3IX chg_counter__i23 (.D(n534[23]), .SP(i_ref_clk_c_enable_180), 
            .CD(chg_counter_23__N_406), .CK(i_ref_clk_c), .Q(chg_counter[23])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[34])
    defparam chg_counter__i23.GSR = "DISABLED";
    FD1P3IX chg_counter__i22 (.D(n534[22]), .SP(i_ref_clk_c_enable_180), 
            .CD(chg_counter_23__N_406), .CK(i_ref_clk_c), .Q(chg_counter[22])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[34])
    defparam chg_counter__i22.GSR = "DISABLED";
    FD1P3IX chg_counter__i21 (.D(n534[21]), .SP(i_ref_clk_c_enable_180), 
            .CD(chg_counter_23__N_406), .CK(i_ref_clk_c), .Q(chg_counter[21])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[34])
    defparam chg_counter__i21.GSR = "DISABLED";
    FD1P3IX chg_counter__i20 (.D(n534[20]), .SP(i_ref_clk_c_enable_180), 
            .CD(chg_counter_23__N_406), .CK(i_ref_clk_c), .Q(chg_counter[20])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[34])
    defparam chg_counter__i20.GSR = "DISABLED";
    FD1P3IX chg_counter__i19 (.D(n534[19]), .SP(i_ref_clk_c_enable_180), 
            .CD(chg_counter_23__N_406), .CK(i_ref_clk_c), .Q(chg_counter[19])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[34])
    defparam chg_counter__i19.GSR = "DISABLED";
    FD1P3IX chg_counter__i18 (.D(n534[18]), .SP(i_ref_clk_c_enable_180), 
            .CD(chg_counter_23__N_406), .CK(i_ref_clk_c), .Q(chg_counter[18])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[34])
    defparam chg_counter__i18.GSR = "DISABLED";
    FD1P3IX chg_counter__i17 (.D(n534[17]), .SP(i_ref_clk_c_enable_180), 
            .CD(chg_counter_23__N_406), .CK(i_ref_clk_c), .Q(chg_counter[17])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[34])
    defparam chg_counter__i17.GSR = "DISABLED";
    FD1P3IX chg_counter__i16 (.D(n534[16]), .SP(i_ref_clk_c_enable_180), 
            .CD(chg_counter_23__N_406), .CK(i_ref_clk_c), .Q(chg_counter[16])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[34])
    defparam chg_counter__i16.GSR = "DISABLED";
    FD1P3IX chg_counter__i15 (.D(n534[15]), .SP(i_ref_clk_c_enable_180), 
            .CD(chg_counter_23__N_406), .CK(i_ref_clk_c), .Q(chg_counter[15])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[34])
    defparam chg_counter__i15.GSR = "DISABLED";
    FD1P3IX chg_counter__i14 (.D(n534[14]), .SP(i_ref_clk_c_enable_180), 
            .CD(chg_counter_23__N_406), .CK(i_ref_clk_c), .Q(chg_counter[14])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[34])
    defparam chg_counter__i14.GSR = "DISABLED";
    FD1P3IX chg_counter__i13 (.D(n534[13]), .SP(i_ref_clk_c_enable_180), 
            .CD(chg_counter_23__N_406), .CK(i_ref_clk_c), .Q(chg_counter[13])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[34])
    defparam chg_counter__i13.GSR = "DISABLED";
    FD1P3IX chg_counter__i12 (.D(n534[12]), .SP(i_ref_clk_c_enable_180), 
            .CD(chg_counter_23__N_406), .CK(i_ref_clk_c), .Q(chg_counter[12])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[34])
    defparam chg_counter__i12.GSR = "DISABLED";
    FD1P3IX chg_counter__i11 (.D(n534[11]), .SP(i_ref_clk_c_enable_180), 
            .CD(chg_counter_23__N_406), .CK(i_ref_clk_c), .Q(chg_counter[11])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[34])
    defparam chg_counter__i11.GSR = "DISABLED";
    FD1P3IX chg_counter__i10 (.D(n534[10]), .SP(i_ref_clk_c_enable_180), 
            .CD(chg_counter_23__N_406), .CK(i_ref_clk_c), .Q(chg_counter[10])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[34])
    defparam chg_counter__i10.GSR = "DISABLED";
    FD1P3IX chg_counter__i9 (.D(n534[9]), .SP(i_ref_clk_c_enable_180), .CD(chg_counter_23__N_406), 
            .CK(i_ref_clk_c), .Q(chg_counter[9])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[34])
    defparam chg_counter__i9.GSR = "DISABLED";
    FD1P3IX chg_counter__i8 (.D(n534[8]), .SP(i_ref_clk_c_enable_180), .CD(chg_counter_23__N_406), 
            .CK(i_ref_clk_c), .Q(chg_counter[8])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[34])
    defparam chg_counter__i8.GSR = "DISABLED";
    FD1P3IX chg_counter__i7 (.D(n534[7]), .SP(i_ref_clk_c_enable_180), .CD(chg_counter_23__N_406), 
            .CK(i_ref_clk_c), .Q(chg_counter[7])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[34])
    defparam chg_counter__i7.GSR = "DISABLED";
    FD1P3IX chg_counter__i6 (.D(n534[6]), .SP(i_ref_clk_c_enable_180), .CD(chg_counter_23__N_406), 
            .CK(i_ref_clk_c), .Q(chg_counter[6])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[34])
    defparam chg_counter__i6.GSR = "DISABLED";
    FD1P3IX chg_counter__i5 (.D(n534[5]), .SP(i_ref_clk_c_enable_180), .CD(chg_counter_23__N_406), 
            .CK(i_ref_clk_c), .Q(chg_counter[5])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[34])
    defparam chg_counter__i5.GSR = "DISABLED";
    FD1P3IX chg_counter__i4 (.D(n534[4]), .SP(i_ref_clk_c_enable_180), .CD(chg_counter_23__N_406), 
            .CK(i_ref_clk_c), .Q(chg_counter[4])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[34])
    defparam chg_counter__i4.GSR = "DISABLED";
    FD1P3IX chg_counter__i3 (.D(n534[3]), .SP(i_ref_clk_c_enable_180), .CD(chg_counter_23__N_406), 
            .CK(i_ref_clk_c), .Q(chg_counter[3])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[34])
    defparam chg_counter__i3.GSR = "DISABLED";
    FD1P3IX chg_counter__i2 (.D(n534[2]), .SP(i_ref_clk_c_enable_180), .CD(chg_counter_23__N_406), 
            .CK(i_ref_clk_c), .Q(chg_counter[2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[34])
    defparam chg_counter__i2.GSR = "DISABLED";
    FD1P3IX chg_counter__i1 (.D(n534[1]), .SP(i_ref_clk_c_enable_180), .CD(chg_counter_23__N_406), 
            .CK(i_ref_clk_c), .Q(chg_counter[1])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[34])
    defparam chg_counter__i1.GSR = "DISABLED";
    CCU2D sub_375_add_2_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n17337), .S0(half_baud_time_N_458));
    defparam sub_375_add_2_cout.INIT0 = 16'h0000;
    defparam sub_375_add_2_cout.INIT1 = 16'h0000;
    defparam sub_375_add_2_cout.INJECT1_0 = "NO";
    defparam sub_375_add_2_cout.INJECT1_1 = "NO";
    CCU2D sub_375_add_2_22 (.A0(chg_counter[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17336), .COUT(n17337));
    defparam sub_375_add_2_22.INIT0 = 16'h5555;
    defparam sub_375_add_2_22.INIT1 = 16'h5555;
    defparam sub_375_add_2_22.INJECT1_0 = "NO";
    defparam sub_375_add_2_22.INJECT1_1 = "NO";
    CCU2D sub_375_add_2_20 (.A0(chg_counter[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17335), .COUT(n17336));
    defparam sub_375_add_2_20.INIT0 = 16'h5555;
    defparam sub_375_add_2_20.INIT1 = 16'h5555;
    defparam sub_375_add_2_20.INJECT1_0 = "NO";
    defparam sub_375_add_2_20.INJECT1_1 = "NO";
    CCU2D sub_375_add_2_18 (.A0(chg_counter[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17334), .COUT(n17335));
    defparam sub_375_add_2_18.INIT0 = 16'h5555;
    defparam sub_375_add_2_18.INIT1 = 16'h5555;
    defparam sub_375_add_2_18.INJECT1_0 = "NO";
    defparam sub_375_add_2_18.INJECT1_1 = "NO";
    CCU2D sub_375_add_2_16 (.A0(chg_counter[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17333), .COUT(n17334));
    defparam sub_375_add_2_16.INIT0 = 16'h5555;
    defparam sub_375_add_2_16.INIT1 = 16'h5555;
    defparam sub_375_add_2_16.INJECT1_0 = "NO";
    defparam sub_375_add_2_16.INJECT1_1 = "NO";
    CCU2D sub_375_add_2_14 (.A0(chg_counter[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17332), .COUT(n17333));
    defparam sub_375_add_2_14.INIT0 = 16'h5555;
    defparam sub_375_add_2_14.INIT1 = 16'h5555;
    defparam sub_375_add_2_14.INJECT1_0 = "NO";
    defparam sub_375_add_2_14.INJECT1_1 = "NO";
    CCU2D sub_375_add_2_12 (.A0(chg_counter[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17331), .COUT(n17332));
    defparam sub_375_add_2_12.INIT0 = 16'h5555;
    defparam sub_375_add_2_12.INIT1 = 16'h5555;
    defparam sub_375_add_2_12.INJECT1_0 = "NO";
    defparam sub_375_add_2_12.INJECT1_1 = "NO";
    CCU2D sub_375_add_2_10 (.A0(chg_counter[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17330), .COUT(n17331));
    defparam sub_375_add_2_10.INIT0 = 16'h5555;
    defparam sub_375_add_2_10.INIT1 = 16'h5555;
    defparam sub_375_add_2_10.INJECT1_0 = "NO";
    defparam sub_375_add_2_10.INJECT1_1 = "NO";
    CCU2D sub_375_add_2_8 (.A0(chg_counter[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17329), .COUT(n17330));
    defparam sub_375_add_2_8.INIT0 = 16'h5555;
    defparam sub_375_add_2_8.INIT1 = 16'h5555;
    defparam sub_375_add_2_8.INJECT1_0 = "NO";
    defparam sub_375_add_2_8.INJECT1_1 = "NO";
    CCU2D sub_375_add_2_6 (.A0(chg_counter[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17328), .COUT(n17329));
    defparam sub_375_add_2_6.INIT0 = 16'h5555;
    defparam sub_375_add_2_6.INIT1 = 16'h5555;
    defparam sub_375_add_2_6.INJECT1_0 = "NO";
    defparam sub_375_add_2_6.INJECT1_1 = "NO";
    CCU2D sub_375_add_2_4 (.A0(chg_counter[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17327), .COUT(n17328));
    defparam sub_375_add_2_4.INIT0 = 16'h5555;
    defparam sub_375_add_2_4.INIT1 = 16'h5555;
    defparam sub_375_add_2_4.INJECT1_0 = "NO";
    defparam sub_375_add_2_4.INJECT1_1 = "NO";
    CCU2D sub_375_add_2_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(chg_counter[3]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n17327));
    defparam sub_375_add_2_2.INIT0 = 16'h0000;
    defparam sub_375_add_2_2.INIT1 = 16'h5aaa;
    defparam sub_375_add_2_2.INJECT1_0 = "NO";
    defparam sub_375_add_2_2.INJECT1_1 = "NO";
    CCU2D sub_49_add_2_25 (.A0(baud_counter[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n17394), .S0(n290[23]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_25.INIT0 = 16'h5555;
    defparam sub_49_add_2_25.INIT1 = 16'h0000;
    defparam sub_49_add_2_25.INJECT1_0 = "NO";
    defparam sub_49_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_49_add_2_23 (.A0(baud_counter[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17393), .COUT(n17394), .S0(n290[21]), 
          .S1(n290[22]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_23.INIT0 = 16'h5555;
    defparam sub_49_add_2_23.INIT1 = 16'h5555;
    defparam sub_49_add_2_23.INJECT1_0 = "NO";
    defparam sub_49_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_49_add_2_21 (.A0(baud_counter[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17392), .COUT(n17393), .S0(n290[19]), 
          .S1(n290[20]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_21.INIT0 = 16'h5555;
    defparam sub_49_add_2_21.INIT1 = 16'h5555;
    defparam sub_49_add_2_21.INJECT1_0 = "NO";
    defparam sub_49_add_2_21.INJECT1_1 = "NO";
    LUT4 zero_baud_counter_I_0_2_lut (.A(zero_baud_counter), .B(state[3]), 
         .Z(zero_baud_counter_N_454)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(175[11:52])
    defparam zero_baud_counter_I_0_2_lut.init = 16'h2222;
    CCU2D sub_49_add_2_19 (.A0(baud_counter[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17391), .COUT(n17392), .S0(n290[17]), 
          .S1(n290[18]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_19.INIT0 = 16'h5555;
    defparam sub_49_add_2_19.INIT1 = 16'h5555;
    defparam sub_49_add_2_19.INJECT1_0 = "NO";
    defparam sub_49_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_49_add_2_17 (.A0(baud_counter[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17390), .COUT(n17391), .S0(n290[15]), 
          .S1(n290[16]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_17.INIT0 = 16'h5555;
    defparam sub_49_add_2_17.INIT1 = 16'h5555;
    defparam sub_49_add_2_17.INJECT1_0 = "NO";
    defparam sub_49_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_49_add_2_15 (.A0(baud_counter[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17389), .COUT(n17390), .S0(n290[13]), 
          .S1(n290[14]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_15.INIT0 = 16'h5555;
    defparam sub_49_add_2_15.INIT1 = 16'h5555;
    defparam sub_49_add_2_15.INJECT1_0 = "NO";
    defparam sub_49_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_49_add_2_13 (.A0(baud_counter[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17388), .COUT(n17389), .S0(n290[11]), 
          .S1(n290[12]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_13.INIT0 = 16'h5555;
    defparam sub_49_add_2_13.INIT1 = 16'h5555;
    defparam sub_49_add_2_13.INJECT1_0 = "NO";
    defparam sub_49_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_49_add_2_11 (.A0(baud_counter[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17387), .COUT(n17388), .S0(n290[9]), .S1(n290[10]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_11.INIT0 = 16'h5555;
    defparam sub_49_add_2_11.INIT1 = 16'h5555;
    defparam sub_49_add_2_11.INJECT1_0 = "NO";
    defparam sub_49_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_49_add_2_9 (.A0(baud_counter[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17386), .COUT(n17387), .S0(n290[7]), .S1(n290[8]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_9.INIT0 = 16'h5555;
    defparam sub_49_add_2_9.INIT1 = 16'h5555;
    defparam sub_49_add_2_9.INJECT1_0 = "NO";
    defparam sub_49_add_2_9.INJECT1_1 = "NO";
    CCU2D add_90_25 (.A0(chg_counter[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n17318), .S0(n534[23]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:33])
    defparam add_90_25.INIT0 = 16'h5aaa;
    defparam add_90_25.INIT1 = 16'h0000;
    defparam add_90_25.INJECT1_0 = "NO";
    defparam add_90_25.INJECT1_1 = "NO";
    CCU2D sub_49_add_2_7 (.A0(baud_counter[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17385), .COUT(n17386), .S0(n290[5]), .S1(n290[6]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_7.INIT0 = 16'h5555;
    defparam sub_49_add_2_7.INIT1 = 16'h5555;
    defparam sub_49_add_2_7.INJECT1_0 = "NO";
    defparam sub_49_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_49_add_2_5 (.A0(baud_counter[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17384), .COUT(n17385), .S0(n290[3]), .S1(n290[4]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_5.INIT0 = 16'h5555;
    defparam sub_49_add_2_5.INIT1 = 16'h5555;
    defparam sub_49_add_2_5.INJECT1_0 = "NO";
    defparam sub_49_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_49_add_2_3 (.A0(baud_counter[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17383), .COUT(n17384), .S0(n290[1]), .S1(n290[2]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_3.INIT0 = 16'h5555;
    defparam sub_49_add_2_3.INIT1 = 16'h5555;
    defparam sub_49_add_2_3.INJECT1_0 = "NO";
    defparam sub_49_add_2_3.INJECT1_1 = "NO";
    LUT4 n4_bdd_4_lut (.A(n25014), .B(state[0]), .C(state[1]), .D(ck_uart), 
         .Z(n23729)) /* synthesis lut_function=(A (C+(D))+!A !(B (C)+!B !(C))) */ ;
    defparam n4_bdd_4_lut.init = 16'hbeb4;
    LUT4 n4_bdd_2_lut_22407 (.A(ck_uart), .B(half_baud_time), .Z(n23728)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam n4_bdd_2_lut_22407.init = 16'hbbbb;
    LUT4 qq_uart_I_0_2_lut (.A(qq_uart), .B(ck_uart), .Z(chg_counter_23__N_406)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(100[6:24])
    defparam qq_uart_I_0_2_lut.init = 16'h6666;
    CCU2D sub_49_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(baud_counter[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n17383), .S1(n290[0]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_1.INIT0 = 16'hF000;
    defparam sub_49_add_2_1.INIT1 = 16'h5555;
    defparam sub_49_add_2_1.INJECT1_0 = "NO";
    defparam sub_49_add_2_1.INJECT1_1 = "NO";
    LUT4 i1_4_lut (.A(n19721), .B(n11693), .C(n46), .D(n19719), .Z(i_ref_clk_c_enable_147)) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;
    defparam i1_4_lut.init = 16'hccdc;
    LUT4 i17409_4_lut (.A(baud_counter[18]), .B(baud_counter[23]), .C(baud_counter[3]), 
         .D(baud_counter[16]), .Z(n19721)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17409_4_lut.init = 16'hfffe;
    LUT4 i22_4_lut (.A(n25), .B(n19737), .C(n19727), .D(n19683), .Z(n46)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i22_4_lut.init = 16'h0002;
    LUT4 i17407_4_lut (.A(baud_counter[19]), .B(baud_counter[13]), .C(baud_counter[2]), 
         .D(baud_counter[14]), .Z(n19719)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17407_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut (.A(baud_counter[10]), .B(baud_counter[0]), .Z(n25)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut.init = 16'h4444;
    LUT4 i17425_4_lut (.A(baud_counter[12]), .B(n19723), .C(n19675), .D(baud_counter[11]), 
         .Z(n19737)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17425_4_lut.init = 16'hfffe;
    LUT4 i17415_4_lut (.A(baud_counter[8]), .B(baud_counter[1]), .C(baud_counter[9]), 
         .D(baud_counter[6]), .Z(n19727)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17415_4_lut.init = 16'hfffe;
    LUT4 i17372_2_lut (.A(baud_counter[20]), .B(baud_counter[5]), .Z(n19683)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i17372_2_lut.init = 16'heeee;
    LUT4 i17411_4_lut (.A(baud_counter[21]), .B(baud_counter[7]), .C(baud_counter[4]), 
         .D(baud_counter[15]), .Z(n19723)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i17411_4_lut.init = 16'hfffe;
    LUT4 i17364_2_lut (.A(baud_counter[17]), .B(baud_counter[22]), .Z(n19675)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i17364_2_lut.init = 16'heeee;
    LUT4 i11426_3_lut_4_lut (.A(state[0]), .B(n24903), .C(zero_baud_counter_N_454), 
         .D(n290[1]), .Z(baud_counter_23__N_421[1])) /* synthesis lut_function=(A (B (C+(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(144[27:48])
    defparam i11426_3_lut_4_lut.init = 16'hddd0;
    LUT4 i21137_3_lut_3_lut_4_lut (.A(state[0]), .B(n24903), .C(zero_baud_counter_N_454), 
         .D(n24981), .Z(n14854)) /* synthesis lut_function=(!(A (B (C+(D))+!B (D))+!A (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(144[27:48])
    defparam i21137_3_lut_3_lut_4_lut.init = 16'h002f;
    LUT4 i11425_3_lut_4_lut (.A(state[0]), .B(n24903), .C(zero_baud_counter_N_454), 
         .D(n290[4]), .Z(baud_counter_23__N_421[4])) /* synthesis lut_function=(A (B (C+(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(144[27:48])
    defparam i11425_3_lut_4_lut.init = 16'hddd0;
    LUT4 i10916_3_lut_4_lut (.A(state[0]), .B(n24903), .C(zero_baud_counter_N_454), 
         .D(n290[0]), .Z(baud_counter_23__N_421[0])) /* synthesis lut_function=(A (B (C+(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(144[27:48])
    defparam i10916_3_lut_4_lut.init = 16'hddd0;
    LUT4 i1_2_lut_3_lut_4_lut (.A(state[0]), .B(n24903), .C(zero_baud_counter_N_454), 
         .D(n24981), .Z(n11693)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(144[27:48])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfff2;
    CCU2D add_90_23 (.A0(chg_counter[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17317), .COUT(n17318), .S0(n534[21]), 
          .S1(n534[22]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:33])
    defparam add_90_23.INIT0 = 16'h5aaa;
    defparam add_90_23.INIT1 = 16'h5aaa;
    defparam add_90_23.INJECT1_0 = "NO";
    defparam add_90_23.INJECT1_1 = "NO";
    CCU2D add_90_21 (.A0(chg_counter[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17316), .COUT(n17317), .S0(n534[19]), 
          .S1(n534[20]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:33])
    defparam add_90_21.INIT0 = 16'h5aaa;
    defparam add_90_21.INIT1 = 16'h5aaa;
    defparam add_90_21.INJECT1_0 = "NO";
    defparam add_90_21.INJECT1_1 = "NO";
    LUT4 i2_3_lut_4_lut_adj_75 (.A(ck_uart), .B(n25014), .C(zero_baud_counter), 
         .D(state_3__N_415), .Z(i_ref_clk_c_enable_355)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(125[15:47])
    defparam i2_3_lut_4_lut_adj_75.init = 16'hfff8;
    CCU2D add_90_19 (.A0(chg_counter[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17315), .COUT(n17316), .S0(n534[17]), 
          .S1(n534[18]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:33])
    defparam add_90_19.INIT0 = 16'h5aaa;
    defparam add_90_19.INIT1 = 16'h5aaa;
    defparam add_90_19.INJECT1_0 = "NO";
    defparam add_90_19.INJECT1_1 = "NO";
    LUT4 i2_2_lut_rep_285_4_lut (.A(state[3]), .B(state[0]), .C(n25013), 
         .D(ck_uart), .Z(n24845)) /* synthesis lut_function=(A (B (D)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(125[15:47])
    defparam i2_2_lut_rep_285_4_lut.init = 16'ha800;
    CCU2D add_90_17 (.A0(chg_counter[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17314), .COUT(n17315), .S0(n534[15]), 
          .S1(n534[16]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:33])
    defparam add_90_17.INIT0 = 16'h5aaa;
    defparam add_90_17.INIT1 = 16'h5aaa;
    defparam add_90_17.INJECT1_0 = "NO";
    defparam add_90_17.INJECT1_1 = "NO";
    CCU2D add_90_15 (.A0(chg_counter[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17313), .COUT(n17314), .S0(n534[13]), 
          .S1(n534[14]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:33])
    defparam add_90_15.INIT0 = 16'h5aaa;
    defparam add_90_15.INIT1 = 16'h5aaa;
    defparam add_90_15.INJECT1_0 = "NO";
    defparam add_90_15.INJECT1_1 = "NO";
    CCU2D add_90_13 (.A0(chg_counter[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17312), .COUT(n17313), .S0(n534[11]), 
          .S1(n534[12]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:33])
    defparam add_90_13.INIT0 = 16'h5aaa;
    defparam add_90_13.INIT1 = 16'h5aaa;
    defparam add_90_13.INJECT1_0 = "NO";
    defparam add_90_13.INJECT1_1 = "NO";
    LUT4 zero_baud_counter_I_0_82_2_lut_3_lut_4_lut (.A(state[3]), .B(n25013), 
         .C(zero_baud_counter), .D(state[0]), .Z(data_reg_7__N_416)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(144[27:48])
    defparam zero_baud_counter_I_0_82_2_lut_3_lut_4_lut.init = 16'hf0d0;
    CCU2D add_90_11 (.A0(chg_counter[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17311), .COUT(n17312), .S0(n534[9]), .S1(n534[10]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:33])
    defparam add_90_11.INIT0 = 16'h5aaa;
    defparam add_90_11.INIT1 = 16'h5aaa;
    defparam add_90_11.INJECT1_0 = "NO";
    defparam add_90_11.INJECT1_1 = "NO";
    CCU2D add_90_9 (.A0(chg_counter[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(chg_counter[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n17310), .COUT(n17311), .S0(n534[7]), .S1(n534[8]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:33])
    defparam add_90_9.INIT0 = 16'h5aaa;
    defparam add_90_9.INIT1 = 16'h5aaa;
    defparam add_90_9.INJECT1_0 = "NO";
    defparam add_90_9.INJECT1_1 = "NO";
    CCU2D add_90_7 (.A0(chg_counter[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(chg_counter[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n17309), .COUT(n17310), .S0(n534[5]), .S1(n534[6]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:33])
    defparam add_90_7.INIT0 = 16'h5aaa;
    defparam add_90_7.INIT1 = 16'h5aaa;
    defparam add_90_7.INJECT1_0 = "NO";
    defparam add_90_7.INJECT1_1 = "NO";
    LUT4 state_3__I_0_80_i1_4_lut (.A(n172), .B(n17705), .C(state_3__N_415), 
         .D(n24845), .Z(state_3__N_322[0])) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C))+!A !((C+(D))+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(125[11] 134[5])
    defparam state_3__I_0_80_i1_4_lut.init = 16'h5f53;
    FD1P3IX baud_counter_i23 (.D(n290[23]), .SP(i_ref_clk_c_enable_351), 
            .CD(n11693), .CK(i_ref_clk_c), .Q(baud_counter[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i23.GSR = "DISABLED";
    LUT4 i21_2_lut (.A(ck_uart), .B(half_baud_time), .Z(n172)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(121[7:35])
    defparam i21_2_lut.init = 16'h4444;
    LUT4 i3_4_lut (.A(state[0]), .B(state[2]), .C(state[1]), .D(state[3]), 
         .Z(state_3__N_415)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i3_4_lut.init = 16'h8000;
    CCU2D add_90_5 (.A0(chg_counter[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(chg_counter[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n17308), .COUT(n17309), .S0(n534[3]), .S1(n534[4]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:33])
    defparam add_90_5.INIT0 = 16'h5aaa;
    defparam add_90_5.INIT1 = 16'h5aaa;
    defparam add_90_5.INJECT1_0 = "NO";
    defparam add_90_5.INJECT1_1 = "NO";
    CCU2D add_90_3 (.A0(chg_counter[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(chg_counter[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n17307), .COUT(n17308), .S0(n534[1]), .S1(n534[2]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:33])
    defparam add_90_3.INIT0 = 16'h5aaa;
    defparam add_90_3.INIT1 = 16'h5aaa;
    defparam add_90_3.INJECT1_0 = "NO";
    defparam add_90_3.INJECT1_1 = "NO";
    LUT4 ck_uart_N_448_I_0_2_lut (.A(ck_uart), .B(half_baud_time_N_458), 
         .Z(half_baud_time_N_457)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(112[21:69])
    defparam ck_uart_N_448_I_0_2_lut.init = 16'h4444;
    CCU2D add_90_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(chg_counter[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n17307), .S1(n534[0]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:33])
    defparam add_90_1.INIT0 = 16'hF000;
    defparam add_90_1.INIT1 = 16'h5555;
    defparam add_90_1.INJECT1_0 = "NO";
    defparam add_90_1.INJECT1_1 = "NO";
    FD1P3IX baud_counter_i22 (.D(n290[22]), .SP(i_ref_clk_c_enable_351), 
            .CD(n11693), .CK(i_ref_clk_c), .Q(baud_counter[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i22.GSR = "DISABLED";
    FD1P3IX baud_counter_i21 (.D(n290[21]), .SP(i_ref_clk_c_enable_351), 
            .CD(n11693), .CK(i_ref_clk_c), .Q(baud_counter[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i21.GSR = "DISABLED";
    FD1P3IX baud_counter_i20 (.D(n290[20]), .SP(i_ref_clk_c_enable_351), 
            .CD(n11693), .CK(i_ref_clk_c), .Q(baud_counter[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i20.GSR = "DISABLED";
    FD1P3IX baud_counter_i19 (.D(n290[19]), .SP(i_ref_clk_c_enable_351), 
            .CD(n11693), .CK(i_ref_clk_c), .Q(baud_counter[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i19.GSR = "DISABLED";
    FD1P3IX baud_counter_i18 (.D(n290[18]), .SP(i_ref_clk_c_enable_351), 
            .CD(n11693), .CK(i_ref_clk_c), .Q(baud_counter[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i18.GSR = "DISABLED";
    FD1P3IX baud_counter_i17 (.D(n290[17]), .SP(i_ref_clk_c_enable_351), 
            .CD(n11693), .CK(i_ref_clk_c), .Q(baud_counter[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i17.GSR = "DISABLED";
    FD1P3IX baud_counter_i16 (.D(n290[16]), .SP(i_ref_clk_c_enable_351), 
            .CD(n11693), .CK(i_ref_clk_c), .Q(baud_counter[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i16.GSR = "DISABLED";
    FD1P3IX baud_counter_i15 (.D(n290[15]), .SP(i_ref_clk_c_enable_351), 
            .CD(n11693), .CK(i_ref_clk_c), .Q(baud_counter[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i15.GSR = "DISABLED";
    FD1P3IX baud_counter_i14 (.D(n290[14]), .SP(i_ref_clk_c_enable_351), 
            .CD(n11693), .CK(i_ref_clk_c), .Q(baud_counter[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i14.GSR = "DISABLED";
    FD1P3IX baud_counter_i13 (.D(n290[13]), .SP(i_ref_clk_c_enable_351), 
            .CD(n11693), .CK(i_ref_clk_c), .Q(baud_counter[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i13.GSR = "DISABLED";
    FD1P3IX baud_counter_i12 (.D(n290[12]), .SP(i_ref_clk_c_enable_351), 
            .CD(n11693), .CK(i_ref_clk_c), .Q(baud_counter[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i12.GSR = "DISABLED";
    FD1P3IX baud_counter_i11 (.D(n290[11]), .SP(i_ref_clk_c_enable_351), 
            .CD(n11693), .CK(i_ref_clk_c), .Q(baud_counter[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i11.GSR = "DISABLED";
    FD1P3IX baud_counter_i10 (.D(n290[10]), .SP(i_ref_clk_c_enable_351), 
            .CD(n11693), .CK(i_ref_clk_c), .Q(baud_counter[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i10.GSR = "DISABLED";
    FD1P3IX baud_counter_i9 (.D(n290[9]), .SP(i_ref_clk_c_enable_351), .CD(n11693), 
            .CK(i_ref_clk_c), .Q(baud_counter[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i9.GSR = "DISABLED";
    FD1P3IX baud_counter_i8 (.D(n290[8]), .SP(i_ref_clk_c_enable_351), .CD(n11693), 
            .CK(i_ref_clk_c), .Q(baud_counter[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i8.GSR = "DISABLED";
    FD1P3IX baud_counter_i7 (.D(n290[7]), .SP(i_ref_clk_c_enable_351), .CD(n11693), 
            .CK(i_ref_clk_c), .Q(baud_counter[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i7.GSR = "DISABLED";
    FD1P3IX baud_counter_i6 (.D(n290[6]), .SP(i_ref_clk_c_enable_351), .CD(n11693), 
            .CK(i_ref_clk_c), .Q(baud_counter[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i6.GSR = "DISABLED";
    FD1P3IX baud_counter_i5 (.D(n290[5]), .SP(i_ref_clk_c_enable_351), .CD(n11693), 
            .CK(i_ref_clk_c), .Q(baud_counter[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i5.GSR = "DISABLED";
    LUT4 i9653_1_lut (.A(zero_baud_counter), .Z(i_ref_clk_c_enable_351)) /* synthesis lut_function=(!(A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(187[9] 195[29])
    defparam i9653_1_lut.init = 16'h5555;
    FD1P3IX baud_counter_i3 (.D(n290[3]), .SP(i_ref_clk_c_enable_351), .CD(n11693), 
            .CK(i_ref_clk_c), .Q(baud_counter[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i3.GSR = "DISABLED";
    FD1P3IX baud_counter_i2 (.D(n290[2]), .SP(i_ref_clk_c_enable_351), .CD(n11693), 
            .CK(i_ref_clk_c), .Q(baud_counter[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i2.GSR = "DISABLED";
    FD1P3AY state_i3 (.D(state_3__N_322[3]), .SP(i_ref_clk_c_enable_355), 
            .CK(i_ref_clk_c), .Q(state[3])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(116[9] 134[5])
    defparam state_i3.GSR = "DISABLED";
    FD1P3AY state_i2 (.D(state_3__N_322[2]), .SP(i_ref_clk_c_enable_355), 
            .CK(i_ref_clk_c), .Q(state[2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(116[9] 134[5])
    defparam state_i2.GSR = "DISABLED";
    FD1P3AY state_i1 (.D(state_3__N_322[1]), .SP(i_ref_clk_c_enable_355), 
            .CK(i_ref_clk_c), .Q(state[1])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(116[9] 134[5])
    defparam state_i1.GSR = "DISABLED";
    FD1P3AX o_data__i7 (.D(data_reg[6]), .SP(o_data_7__N_418), .CK(i_ref_clk_c), 
            .Q(\rx_data[6] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(155[9] 161[18])
    defparam o_data__i7.GSR = "DISABLED";
    FD1P3AX o_data__i6 (.D(data_reg[5]), .SP(o_data_7__N_418), .CK(i_ref_clk_c), 
            .Q(\rx_data[5] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(155[9] 161[18])
    defparam o_data__i6.GSR = "DISABLED";
    FD1P3AX o_data__i5 (.D(data_reg[4]), .SP(o_data_7__N_418), .CK(i_ref_clk_c), 
            .Q(\rx_data[4] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(155[9] 161[18])
    defparam o_data__i5.GSR = "DISABLED";
    FD1P3AX o_data__i4 (.D(data_reg[3]), .SP(o_data_7__N_418), .CK(i_ref_clk_c), 
            .Q(\rx_data[3] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(155[9] 161[18])
    defparam o_data__i4.GSR = "DISABLED";
    FD1P3AX o_data__i3 (.D(data_reg[2]), .SP(o_data_7__N_418), .CK(i_ref_clk_c), 
            .Q(\rx_data[2] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(155[9] 161[18])
    defparam o_data__i3.GSR = "DISABLED";
    FD1P3AX o_data__i2 (.D(data_reg[1]), .SP(o_data_7__N_418), .CK(i_ref_clk_c), 
            .Q(\rx_data[1] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(155[9] 161[18])
    defparam o_data__i2.GSR = "DISABLED";
    LUT4 state_3__I_0_80_i3_4_lut (.A(n172), .B(n560[2]), .C(state_3__N_415), 
         .D(n24845), .Z(state_3__N_322[2])) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A !(B+(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(125[11] 134[5])
    defparam state_3__I_0_80_i3_4_lut.init = 16'h5f5c;
    LUT4 i2_3_lut_rep_421 (.A(half_baud_time), .B(ck_uart), .C(state_3__N_415), 
         .Z(n24981)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(171[6:57])
    defparam i2_3_lut_rep_421.init = 16'h2020;
    LUT4 i1_2_lut_rep_453 (.A(state[2]), .B(state[1]), .Z(n25013)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(144[27:48])
    defparam i1_2_lut_rep_453.init = 16'heeee;
    LUT4 i1_2_lut_3_lut_4_lut_adj_76 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(state[3]), .Z(n17705)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(144[27:48])
    defparam i1_2_lut_3_lut_4_lut_adj_76.init = 16'h0ef0;
    LUT4 state_3__I_0_80_i4_4_lut_else_4_lut (.A(state[0]), .B(n24845), 
         .C(state[2]), .D(state[1]), .Z(n25240)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(125[11] 134[5])
    defparam state_3__I_0_80_i4_4_lut_else_4_lut.init = 16'heccc;
    LUT4 i1_2_lut_rep_343_3_lut (.A(state[2]), .B(state[1]), .C(state[3]), 
         .Z(n24903)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(144[27:48])
    defparam i1_2_lut_rep_343_3_lut.init = 16'hefef;
    LUT4 i1_2_lut_rep_326_3_lut_4_lut (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(state[3]), .Z(n24886)) /* synthesis lut_function=(A+(B+!(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(144[27:48])
    defparam i1_2_lut_rep_326_3_lut_4_lut.init = 16'hefff;
    LUT4 i1_3_lut_rep_454 (.A(state[2]), .B(state[1]), .C(state[0]), .D(state[3]), 
         .Z(n25014)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(144[27:48])
    defparam i1_3_lut_rep_454.init = 16'hfe00;
    LUT4 i735_2_lut_3_lut_4_lut_4_lut (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(state[3]), .Z(n560[2])) /* synthesis lut_function=(A (((D)+!C)+!B)+!A !(((D)+!C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(144[27:48])
    defparam i735_2_lut_3_lut_4_lut_4_lut.init = 16'haa6a;
    LUT4 state_3__I_0_80_i4_4_lut_then_4_lut (.A(n172), .B(state[0]), .C(state[2]), 
         .D(state[1]), .Z(n25241)) /* synthesis lut_function=(!(A (B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(125[11] 134[5])
    defparam state_3__I_0_80_i4_4_lut_then_4_lut.init = 16'h7fff;
    PFUMX i22126 (.BLUT(n23729), .ALUT(n23728), .C0(state_3__N_415), .Z(state_3__N_322[1]));
    FD1P3JX baud_counter_i0 (.D(baud_counter_23__N_421[0]), .SP(i_ref_clk_c_enable_416), 
            .PD(n24981), .CK(i_ref_clk_c), .Q(baud_counter[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i0.GSR = "DISABLED";
    FD1P3AX data_reg_i0_i0 (.D(data_reg[1]), .SP(data_reg_7__N_416), .CK(i_ref_clk_c), 
            .Q(data_reg[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(143[9] 145[42])
    defparam data_reg_i0_i0.GSR = "DISABLED";
    FD1P3AX data_reg_i0_i7 (.D(qq_uart), .SP(data_reg_7__N_416), .CK(i_ref_clk_c), 
            .Q(data_reg[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(143[9] 145[42])
    defparam data_reg_i0_i7.GSR = "DISABLED";
    FD1P3AX data_reg_i0_i6 (.D(data_reg[7]), .SP(data_reg_7__N_416), .CK(i_ref_clk_c), 
            .Q(data_reg[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(143[9] 145[42])
    defparam data_reg_i0_i6.GSR = "DISABLED";
    FD1P3AX data_reg_i0_i5 (.D(data_reg[6]), .SP(data_reg_7__N_416), .CK(i_ref_clk_c), 
            .Q(data_reg[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(143[9] 145[42])
    defparam data_reg_i0_i5.GSR = "DISABLED";
    FD1P3AX data_reg_i0_i4 (.D(data_reg[5]), .SP(data_reg_7__N_416), .CK(i_ref_clk_c), 
            .Q(data_reg[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(143[9] 145[42])
    defparam data_reg_i0_i4.GSR = "DISABLED";
    FD1P3AX data_reg_i0_i3 (.D(data_reg[4]), .SP(data_reg_7__N_416), .CK(i_ref_clk_c), 
            .Q(data_reg[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(143[9] 145[42])
    defparam data_reg_i0_i3.GSR = "DISABLED";
    FD1P3AX data_reg_i0_i2 (.D(data_reg[3]), .SP(data_reg_7__N_416), .CK(i_ref_clk_c), 
            .Q(data_reg[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(143[9] 145[42])
    defparam data_reg_i0_i2.GSR = "DISABLED";
    FD1P3AX data_reg_i0_i1 (.D(data_reg[2]), .SP(data_reg_7__N_416), .CK(i_ref_clk_c), 
            .Q(data_reg[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=54, LSE_RCOL=102, LSE_LLINE=54, LSE_RLINE=54 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(143[9] 145[42])
    defparam data_reg_i0_i1.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module dynamic_pll
//

module dynamic_pll (i_clk_2f_N_2249, lo_pll_out, i_ref_clk_c, pll_clk, 
            pll_rst, pll_stb, pll_we, pll_data_i, pll_addr, pll_data_o, 
            pll_ack, GND_net) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;
    output i_clk_2f_N_2249;
    output lo_pll_out;
    input i_ref_clk_c;
    input pll_clk;
    input pll_rst;
    input pll_stb;
    input pll_we;
    input [7:0]pll_data_i;
    input [4:0]pll_addr;
    output [7:0]pll_data_o;
    output pll_ack;
    input GND_net;
    
    wire i_clk_2f_N_2249 /* synthesis is_inv_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/clock_phase_shifter.v(11[21:28])
    wire lo_pll_out /* synthesis is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(159[6:16])
    wire i_ref_clk_c /* synthesis SET_AS_NETWORK=i_ref_clk_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(22[12:21])
    
    INV i24691 (.A(lo_pll_out), .Z(i_clk_2f_N_2249));
    EHXPLLJ PLLInst_0 (.CLKI(i_ref_clk_c), .CLKFB(lo_pll_out), .PHASESEL0(GND_net), 
            .PHASESEL1(GND_net), .PHASEDIR(GND_net), .PHASESTEP(GND_net), 
            .LOADREG(GND_net), .STDBY(GND_net), .PLLWAKESYNC(GND_net), 
            .RST(GND_net), .RESETC(GND_net), .RESETD(GND_net), .RESETM(GND_net), 
            .ENCLKOP(GND_net), .ENCLKOS(GND_net), .ENCLKOS2(GND_net), 
            .ENCLKOS3(GND_net), .PLLCLK(pll_clk), .PLLRST(pll_rst), .PLLSTB(pll_stb), 
            .PLLWE(pll_we), .PLLDATI0(pll_data_i[0]), .PLLDATI1(pll_data_i[1]), 
            .PLLDATI2(pll_data_i[2]), .PLLDATI3(pll_data_i[3]), .PLLDATI4(pll_data_i[4]), 
            .PLLDATI5(pll_data_i[5]), .PLLDATI6(pll_data_i[6]), .PLLDATI7(pll_data_i[7]), 
            .PLLADDR0(pll_addr[0]), .PLLADDR1(pll_addr[1]), .PLLADDR2(pll_addr[2]), 
            .PLLADDR3(pll_addr[3]), .PLLADDR4(pll_addr[4]), .CLKOP(lo_pll_out), 
            .PLLDATO0(pll_data_o[0]), .PLLDATO1(pll_data_o[1]), .PLLDATO2(pll_data_o[2]), 
            .PLLDATO3(pll_data_o[3]), .PLLDATO4(pll_data_o[4]), .PLLDATO5(pll_data_o[5]), 
            .PLLDATO6(pll_data_o[6]), .PLLDATO7(pll_data_o[7]), .PLLACK(pll_ack)) /* synthesis FREQUENCY_PIN_CLKOP="96.000000", FREQUENCY_PIN_CLKI="12.000000", ICP_CURRENT="7", LPF_RESISTOR="8", syn_instantiated=1, LSE_LINE_FILE_ID=8, LSE_LCOL=13, LSE_RCOL=5, LSE_LLINE=166, LSE_RLINE=177 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(166[13] 177[5])
    defparam PLLInst_0.CLKI_DIV = 1;
    defparam PLLInst_0.CLKFB_DIV = 8;
    defparam PLLInst_0.CLKOP_DIV = 5;
    defparam PLLInst_0.CLKOS_DIV = 1;
    defparam PLLInst_0.CLKOS2_DIV = 1;
    defparam PLLInst_0.CLKOS3_DIV = 1;
    defparam PLLInst_0.CLKOP_ENABLE = "ENABLED";
    defparam PLLInst_0.CLKOS_ENABLE = "DISABLED";
    defparam PLLInst_0.CLKOS2_ENABLE = "DISABLED";
    defparam PLLInst_0.CLKOS3_ENABLE = "DISABLED";
    defparam PLLInst_0.VCO_BYPASS_A0 = "DISABLED";
    defparam PLLInst_0.VCO_BYPASS_B0 = "DISABLED";
    defparam PLLInst_0.VCO_BYPASS_C0 = "DISABLED";
    defparam PLLInst_0.VCO_BYPASS_D0 = "DISABLED";
    defparam PLLInst_0.CLKOP_CPHASE = 4;
    defparam PLLInst_0.CLKOS_CPHASE = 0;
    defparam PLLInst_0.CLKOS2_CPHASE = 0;
    defparam PLLInst_0.CLKOS3_CPHASE = 0;
    defparam PLLInst_0.CLKOP_FPHASE = 0;
    defparam PLLInst_0.CLKOS_FPHASE = 0;
    defparam PLLInst_0.CLKOS2_FPHASE = 0;
    defparam PLLInst_0.CLKOS3_FPHASE = 0;
    defparam PLLInst_0.FEEDBK_PATH = "CLKOP";
    defparam PLLInst_0.FRACN_ENABLE = "ENABLED";
    defparam PLLInst_0.FRACN_DIV = 2731;
    defparam PLLInst_0.CLKOP_TRIM_POL = "RISING";
    defparam PLLInst_0.CLKOP_TRIM_DELAY = 0;
    defparam PLLInst_0.CLKOS_TRIM_POL = "FALLING";
    defparam PLLInst_0.CLKOS_TRIM_DELAY = 0;
    defparam PLLInst_0.PLL_USE_WB = "ENABLED";
    defparam PLLInst_0.PREDIVIDER_MUXA1 = 0;
    defparam PLLInst_0.PREDIVIDER_MUXB1 = 0;
    defparam PLLInst_0.PREDIVIDER_MUXC1 = 0;
    defparam PLLInst_0.PREDIVIDER_MUXD1 = 0;
    defparam PLLInst_0.OUTDIVIDER_MUXA2 = "DIVA";
    defparam PLLInst_0.OUTDIVIDER_MUXB2 = "DIVB";
    defparam PLLInst_0.OUTDIVIDER_MUXC2 = "DIVC";
    defparam PLLInst_0.OUTDIVIDER_MUXD2 = "DIVD";
    defparam PLLInst_0.PLL_LOCK_MODE = 0;
    defparam PLLInst_0.STDBY_ENABLE = "DISABLED";
    defparam PLLInst_0.DPHASE_SOURCE = "DISABLED";
    defparam PLLInst_0.PLLRST_ENA = "DISABLED";
    defparam PLLInst_0.MRST_ENA = "DISABLED";
    defparam PLLInst_0.DCRST_ENA = "DISABLED";
    defparam PLLInst_0.DDRST_ENA = "DISABLED";
    defparam PLLInst_0.INTFB_WAKE = "DISABLED";
    
endmodule
//
// Verilog Description of module \txuartlite(TIMING_BITS=24,CLOCKS_PER_BAUD=20) 
//

module \txuartlite(TIMING_BITS=24,CLOCKS_PER_BAUD=20)  (i_ref_clk_c, i_ref_clk_c_enable_329, 
            \lcl_data_7__N_511[0] , zero_baud_counter_N_526, zero_baud_counter, 
            zero_baud_counter_N_525, o_wbu_uart_tx_c, n24992, GND_net, 
            \lcl_data[7] , n27530, \lcl_data[6] , \lcl_data_7__N_511[6] , 
            \lcl_data[5] , \lcl_data_7__N_511[5] , \lcl_data[4] , \lcl_data_7__N_511[4] , 
            \lcl_data[3] , \lcl_data_7__N_511[3] , \lcl_data[2] , \lcl_data_7__N_511[2] , 
            \lcl_data[1] , \lcl_data_7__N_511[1] , n24890, \state[0] , 
            o_busy_N_536, tx_busy, n17568) /* synthesis syn_module_defined=1 */ ;
    input i_ref_clk_c;
    input i_ref_clk_c_enable_329;
    input \lcl_data_7__N_511[0] ;
    output zero_baud_counter_N_526;
    output zero_baud_counter;
    input zero_baud_counter_N_525;
    output o_wbu_uart_tx_c;
    input n24992;
    input GND_net;
    output \lcl_data[7] ;
    input n27530;
    output \lcl_data[6] ;
    input \lcl_data_7__N_511[6] ;
    output \lcl_data[5] ;
    input \lcl_data_7__N_511[5] ;
    output \lcl_data[4] ;
    input \lcl_data_7__N_511[4] ;
    output \lcl_data[3] ;
    input \lcl_data_7__N_511[3] ;
    output \lcl_data[2] ;
    input \lcl_data_7__N_511[2] ;
    output \lcl_data[1] ;
    input \lcl_data_7__N_511[1] ;
    output n24890;
    output \state[0] ;
    output o_busy_N_536;
    output tx_busy;
    input n17568;
    
    wire i_ref_clk_c /* synthesis SET_AS_NETWORK=i_ref_clk_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(22[12:21])
    wire [7:0]lcl_data;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(84[12:20])
    
    wire n41, zero_baud_counter_N_528, n46, n42;
    wire [23:0]baud_counter;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(82[17:29])
    wire [23:0]baud_counter_23__N_483;
    
    wire n40, n25234, n25235;
    wire [3:0]state;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(83[12:17])
    
    wire n25236, n30, n25227, n25228, n25229, n17382;
    wire [23:0]n108;
    
    wire n25000, n11539, n17381, n17380, n17379, n17378, n17377, 
        n17376, n17375, n17374, n17373, n17372, n17371;
    wire [23:0]n133;
    
    wire n8934;
    wire [3:0]n27;
    
    wire n25, n44, n38, n26;
    
    FD1P3AY lcl_data_i0 (.D(\lcl_data_7__N_511[0] ), .SP(i_ref_clk_c_enable_329), 
            .CK(i_ref_clk_c), .Q(lcl_data[0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=55, LSE_RCOL=112, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(139[9] 143[40])
    defparam lcl_data_i0.GSR = "DISABLED";
    LUT4 i10921_4_lut (.A(n41), .B(zero_baud_counter_N_528), .C(n46), 
         .D(n42), .Z(zero_baud_counter_N_526)) /* synthesis lut_function=(A (B)+!A (B+!(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(221[12] 224[43])
    defparam i10921_4_lut.init = 16'hcccd;
    FD1S3AY zero_baud_counter_49 (.D(zero_baud_counter_N_525), .CK(i_ref_clk_c), 
            .Q(zero_baud_counter)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=55, LSE_RCOL=112, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam zero_baud_counter_49.GSR = "DISABLED";
    FD1S3AX baud_counter_i0 (.D(baud_counter_23__N_483[0]), .CK(i_ref_clk_c), 
            .Q(baud_counter[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=55, LSE_RCOL=112, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i0.GSR = "DISABLED";
    FD1P3IX o_uart_tx_48 (.D(lcl_data[0]), .SP(i_ref_clk_c_enable_329), 
            .CD(n24992), .CK(i_ref_clk_c), .Q(o_wbu_uart_tx_c)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=55, LSE_RCOL=112, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(154[9] 158[29])
    defparam o_uart_tx_48.GSR = "DISABLED";
    LUT4 i16_4_lut (.A(baud_counter[21]), .B(baud_counter[7]), .C(baud_counter[4]), 
         .D(baud_counter[15]), .Z(n40)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(207[24:43])
    defparam i16_4_lut.init = 16'hfffe;
    PFUMX i23018 (.BLUT(n25234), .ALUT(n25235), .C0(state[3]), .Z(n25236));
    LUT4 i6_2_lut (.A(baud_counter[17]), .B(baud_counter[22]), .Z(n30)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(207[24:43])
    defparam i6_2_lut.init = 16'heeee;
    PFUMX i23014 (.BLUT(n25227), .ALUT(n25228), .C0(state[2]), .Z(n25229));
    CCU2D sub_36_add_2_25 (.A0(baud_counter[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n17382), .S0(n108[23]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_25.INIT0 = 16'h5555;
    defparam sub_36_add_2_25.INIT1 = 16'h0000;
    defparam sub_36_add_2_25.INJECT1_0 = "NO";
    defparam sub_36_add_2_25.INJECT1_1 = "NO";
    LUT4 i1_2_lut_4_lut (.A(n25000), .B(state[2]), .C(state[1]), .D(zero_baud_counter), 
         .Z(n11539)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;
    defparam i1_2_lut_4_lut.init = 16'hff80;
    CCU2D sub_36_add_2_23 (.A0(baud_counter[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17381), .COUT(n17382), .S0(n108[21]), 
          .S1(n108[22]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_23.INIT0 = 16'h5555;
    defparam sub_36_add_2_23.INIT1 = 16'h5555;
    defparam sub_36_add_2_23.INJECT1_0 = "NO";
    defparam sub_36_add_2_23.INJECT1_1 = "NO";
    FD1S3IX baud_counter_i23 (.D(n108[23]), .CK(i_ref_clk_c), .CD(n11539), 
            .Q(baud_counter[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=55, LSE_RCOL=112, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i23.GSR = "DISABLED";
    CCU2D sub_36_add_2_21 (.A0(baud_counter[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17380), .COUT(n17381), .S0(n108[19]), 
          .S1(n108[20]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_21.INIT0 = 16'h5555;
    defparam sub_36_add_2_21.INIT1 = 16'h5555;
    defparam sub_36_add_2_21.INJECT1_0 = "NO";
    defparam sub_36_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_36_add_2_19 (.A0(baud_counter[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17379), .COUT(n17380), .S0(n108[17]), 
          .S1(n108[18]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_19.INIT0 = 16'h5555;
    defparam sub_36_add_2_19.INIT1 = 16'h5555;
    defparam sub_36_add_2_19.INJECT1_0 = "NO";
    defparam sub_36_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_36_add_2_17 (.A0(baud_counter[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17378), .COUT(n17379), .S0(n108[15]), 
          .S1(n108[16]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_17.INIT0 = 16'h5555;
    defparam sub_36_add_2_17.INIT1 = 16'h5555;
    defparam sub_36_add_2_17.INJECT1_0 = "NO";
    defparam sub_36_add_2_17.INJECT1_1 = "NO";
    LUT4 i2_4_lut (.A(n25000), .B(zero_baud_counter), .C(state[2]), .D(state[1]), 
         .Z(zero_baud_counter_N_528)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i2_4_lut.init = 16'h0008;
    CCU2D sub_36_add_2_15 (.A0(baud_counter[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17377), .COUT(n17378), .S0(n108[13]), 
          .S1(n108[14]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_15.INIT0 = 16'h5555;
    defparam sub_36_add_2_15.INIT1 = 16'h5555;
    defparam sub_36_add_2_15.INJECT1_0 = "NO";
    defparam sub_36_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_36_add_2_13 (.A0(baud_counter[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17376), .COUT(n17377), .S0(n108[11]), 
          .S1(n108[12]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_13.INIT0 = 16'h5555;
    defparam sub_36_add_2_13.INIT1 = 16'h5555;
    defparam sub_36_add_2_13.INJECT1_0 = "NO";
    defparam sub_36_add_2_13.INJECT1_1 = "NO";
    FD1S3IX baud_counter_i22 (.D(n108[22]), .CK(i_ref_clk_c), .CD(n11539), 
            .Q(baud_counter[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=55, LSE_RCOL=112, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i22.GSR = "DISABLED";
    FD1S3IX baud_counter_i21 (.D(n108[21]), .CK(i_ref_clk_c), .CD(n11539), 
            .Q(baud_counter[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=55, LSE_RCOL=112, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i21.GSR = "DISABLED";
    FD1S3IX baud_counter_i20 (.D(n108[20]), .CK(i_ref_clk_c), .CD(n11539), 
            .Q(baud_counter[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=55, LSE_RCOL=112, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i20.GSR = "DISABLED";
    FD1S3IX baud_counter_i19 (.D(n108[19]), .CK(i_ref_clk_c), .CD(n11539), 
            .Q(baud_counter[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=55, LSE_RCOL=112, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i19.GSR = "DISABLED";
    FD1S3IX baud_counter_i18 (.D(n108[18]), .CK(i_ref_clk_c), .CD(n11539), 
            .Q(baud_counter[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=55, LSE_RCOL=112, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i18.GSR = "DISABLED";
    FD1S3IX baud_counter_i17 (.D(n108[17]), .CK(i_ref_clk_c), .CD(n11539), 
            .Q(baud_counter[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=55, LSE_RCOL=112, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i17.GSR = "DISABLED";
    FD1S3IX baud_counter_i16 (.D(n108[16]), .CK(i_ref_clk_c), .CD(n11539), 
            .Q(baud_counter[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=55, LSE_RCOL=112, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i16.GSR = "DISABLED";
    FD1S3IX baud_counter_i15 (.D(n108[15]), .CK(i_ref_clk_c), .CD(n11539), 
            .Q(baud_counter[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=55, LSE_RCOL=112, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i15.GSR = "DISABLED";
    FD1S3IX baud_counter_i14 (.D(n108[14]), .CK(i_ref_clk_c), .CD(n11539), 
            .Q(baud_counter[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=55, LSE_RCOL=112, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i14.GSR = "DISABLED";
    FD1S3IX baud_counter_i13 (.D(n108[13]), .CK(i_ref_clk_c), .CD(n11539), 
            .Q(baud_counter[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=55, LSE_RCOL=112, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i13.GSR = "DISABLED";
    FD1S3IX baud_counter_i12 (.D(n108[12]), .CK(i_ref_clk_c), .CD(n11539), 
            .Q(baud_counter[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=55, LSE_RCOL=112, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i12.GSR = "DISABLED";
    FD1S3IX baud_counter_i11 (.D(n108[11]), .CK(i_ref_clk_c), .CD(n11539), 
            .Q(baud_counter[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=55, LSE_RCOL=112, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i11.GSR = "DISABLED";
    FD1S3IX baud_counter_i10 (.D(n108[10]), .CK(i_ref_clk_c), .CD(n11539), 
            .Q(baud_counter[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=55, LSE_RCOL=112, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i10.GSR = "DISABLED";
    FD1S3IX baud_counter_i9 (.D(n108[9]), .CK(i_ref_clk_c), .CD(n11539), 
            .Q(baud_counter[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=55, LSE_RCOL=112, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i9.GSR = "DISABLED";
    FD1S3IX baud_counter_i8 (.D(n108[8]), .CK(i_ref_clk_c), .CD(n11539), 
            .Q(baud_counter[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=55, LSE_RCOL=112, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i8.GSR = "DISABLED";
    FD1S3IX baud_counter_i7 (.D(n108[7]), .CK(i_ref_clk_c), .CD(n11539), 
            .Q(baud_counter[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=55, LSE_RCOL=112, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i7.GSR = "DISABLED";
    FD1S3IX baud_counter_i6 (.D(n108[6]), .CK(i_ref_clk_c), .CD(n11539), 
            .Q(baud_counter[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=55, LSE_RCOL=112, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i6.GSR = "DISABLED";
    FD1S3IX baud_counter_i5 (.D(n108[5]), .CK(i_ref_clk_c), .CD(n11539), 
            .Q(baud_counter[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=55, LSE_RCOL=112, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i5.GSR = "DISABLED";
    FD1S3AX baud_counter_i4 (.D(baud_counter_23__N_483[4]), .CK(i_ref_clk_c), 
            .Q(baud_counter[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=55, LSE_RCOL=112, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i4.GSR = "DISABLED";
    FD1S3IX baud_counter_i3 (.D(n108[3]), .CK(i_ref_clk_c), .CD(n11539), 
            .Q(baud_counter[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=55, LSE_RCOL=112, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i3.GSR = "DISABLED";
    FD1S3IX baud_counter_i2 (.D(n108[2]), .CK(i_ref_clk_c), .CD(n11539), 
            .Q(baud_counter[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=55, LSE_RCOL=112, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i2.GSR = "DISABLED";
    FD1S3AX baud_counter_i1 (.D(baud_counter_23__N_483[1]), .CK(i_ref_clk_c), 
            .Q(baud_counter[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=55, LSE_RCOL=112, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i1.GSR = "DISABLED";
    FD1P3IX lcl_data_i7 (.D(n27530), .SP(zero_baud_counter), .CD(n24992), 
            .CK(i_ref_clk_c), .Q(\lcl_data[7] )) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=55, LSE_RCOL=112, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(139[9] 143[40])
    defparam lcl_data_i7.GSR = "DISABLED";
    CCU2D sub_36_add_2_11 (.A0(baud_counter[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17375), .COUT(n17376), .S0(n108[9]), .S1(n108[10]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_11.INIT0 = 16'h5555;
    defparam sub_36_add_2_11.INIT1 = 16'h5555;
    defparam sub_36_add_2_11.INJECT1_0 = "NO";
    defparam sub_36_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_36_add_2_9 (.A0(baud_counter[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17374), .COUT(n17375), .S0(n108[7]), .S1(n108[8]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_9.INIT0 = 16'h5555;
    defparam sub_36_add_2_9.INIT1 = 16'h5555;
    defparam sub_36_add_2_9.INJECT1_0 = "NO";
    defparam sub_36_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_36_add_2_7 (.A0(baud_counter[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17373), .COUT(n17374), .S0(n108[5]), .S1(n108[6]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_7.INIT0 = 16'h5555;
    defparam sub_36_add_2_7.INIT1 = 16'h5555;
    defparam sub_36_add_2_7.INJECT1_0 = "NO";
    defparam sub_36_add_2_7.INJECT1_1 = "NO";
    FD1P3AY lcl_data_i6 (.D(\lcl_data_7__N_511[6] ), .SP(i_ref_clk_c_enable_329), 
            .CK(i_ref_clk_c), .Q(\lcl_data[6] )) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=55, LSE_RCOL=112, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(139[9] 143[40])
    defparam lcl_data_i6.GSR = "DISABLED";
    CCU2D sub_36_add_2_5 (.A0(baud_counter[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17372), .COUT(n17373), .S0(n108[3]), .S1(n108[4]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_5.INIT0 = 16'h5555;
    defparam sub_36_add_2_5.INIT1 = 16'h5555;
    defparam sub_36_add_2_5.INJECT1_0 = "NO";
    defparam sub_36_add_2_5.INJECT1_1 = "NO";
    FD1P3AY lcl_data_i5 (.D(\lcl_data_7__N_511[5] ), .SP(i_ref_clk_c_enable_329), 
            .CK(i_ref_clk_c), .Q(\lcl_data[5] )) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=55, LSE_RCOL=112, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(139[9] 143[40])
    defparam lcl_data_i5.GSR = "DISABLED";
    FD1P3AY lcl_data_i4 (.D(\lcl_data_7__N_511[4] ), .SP(i_ref_clk_c_enable_329), 
            .CK(i_ref_clk_c), .Q(\lcl_data[4] )) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=55, LSE_RCOL=112, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(139[9] 143[40])
    defparam lcl_data_i4.GSR = "DISABLED";
    FD1P3AY lcl_data_i3 (.D(\lcl_data_7__N_511[3] ), .SP(i_ref_clk_c_enable_329), 
            .CK(i_ref_clk_c), .Q(\lcl_data[3] )) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=55, LSE_RCOL=112, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(139[9] 143[40])
    defparam lcl_data_i3.GSR = "DISABLED";
    FD1P3AY lcl_data_i2 (.D(\lcl_data_7__N_511[2] ), .SP(i_ref_clk_c_enable_329), 
            .CK(i_ref_clk_c), .Q(\lcl_data[2] )) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=55, LSE_RCOL=112, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(139[9] 143[40])
    defparam lcl_data_i2.GSR = "DISABLED";
    FD1P3AY lcl_data_i1 (.D(\lcl_data_7__N_511[1] ), .SP(i_ref_clk_c_enable_329), 
            .CK(i_ref_clk_c), .Q(\lcl_data[1] )) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=55, LSE_RCOL=112, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(139[9] 143[40])
    defparam lcl_data_i1.GSR = "DISABLED";
    CCU2D sub_36_add_2_3 (.A0(baud_counter[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17371), .COUT(n17372), .S0(n108[1]), .S1(n108[2]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_3.INIT0 = 16'h5555;
    defparam sub_36_add_2_3.INIT1 = 16'h5555;
    defparam sub_36_add_2_3.INJECT1_0 = "NO";
    defparam sub_36_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_36_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(baud_counter[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n17371), .S1(n108[0]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_1.INIT0 = 16'hF000;
    defparam sub_36_add_2_1.INIT1 = 16'h5555;
    defparam sub_36_add_2_1.INJECT1_0 = "NO";
    defparam sub_36_add_2_1.INJECT1_1 = "NO";
    LUT4 baud_counter_23__I_10_i5_4_lut (.A(n24992), .B(n133[4]), .C(n24890), 
         .D(zero_baud_counter_N_528), .Z(baud_counter_23__N_483[4])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((C+(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(217[12] 224[43])
    defparam baud_counter_23__I_10_i5_4_lut.init = 16'ha0ac;
    LUT4 i11405_2_lut (.A(n108[4]), .B(zero_baud_counter), .Z(n133[4])) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(224[4:43])
    defparam i11405_2_lut.init = 16'heeee;
    LUT4 baud_counter_23__I_10_i2_4_lut (.A(n24992), .B(n133[1]), .C(n24890), 
         .D(zero_baud_counter_N_528), .Z(baud_counter_23__N_483[1])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((C+(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(217[12] 224[43])
    defparam baud_counter_23__I_10_i2_4_lut.init = 16'ha0ac;
    LUT4 i11406_2_lut (.A(n108[1]), .B(zero_baud_counter), .Z(n133[1])) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(224[4:43])
    defparam i11406_2_lut.init = 16'heeee;
    LUT4 i17_4_lut (.A(baud_counter[18]), .B(baud_counter[23]), .C(baud_counter[3]), 
         .D(baud_counter[16]), .Z(n41)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(207[24:43])
    defparam i17_4_lut.init = 16'hfffe;
    LUT4 i688_4_lut (.A(state[2]), .B(state[3]), .C(state[1]), .D(\state[0] ), 
         .Z(o_busy_N_536)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;
    defparam i688_4_lut.init = 16'hccc8;
    LUT4 i21048_2_lut (.A(o_busy_N_536), .B(zero_baud_counter), .Z(n8934)) /* synthesis lut_function=(!(A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(97[8] 113[6])
    defparam i21048_2_lut.init = 16'h7777;
    LUT4 state_504_mux_6_i2_4_lut (.A(state[1]), .B(n24992), .C(o_busy_N_536), 
         .D(\state[0] ), .Z(n27[1])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(110[14:26])
    defparam state_504_mux_6_i2_4_lut.init = 16'h353a;
    FD1P3AX state_504__i3 (.D(n25236), .SP(zero_baud_counter), .CK(i_ref_clk_c), 
            .Q(state[3]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(110[14:26])
    defparam state_504__i3.GSR = "DISABLED";
    LUT4 state_504_mux_6_i3_4_lut_then_4_lut (.A(n24992), .B(\state[0] ), 
         .C(state[1]), .D(state[3]), .Z(n25228)) /* synthesis lut_function=(!(A (B (C+(D))+!B (D))+!A !(((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(110[14:26])
    defparam state_504_mux_6_i3_4_lut_then_4_lut.init = 16'h553f;
    LUT4 state_504_mux_6_i3_4_lut_else_4_lut (.A(n24992), .B(\state[0] ), 
         .C(state[1]), .D(state[3]), .Z(n25227)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A !(B (C+(D))+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(110[14:26])
    defparam state_504_mux_6_i3_4_lut_else_4_lut.init = 16'h54c0;
    LUT4 baud_counter_23__I_10_i1_4_lut (.A(n24992), .B(n133[0]), .C(n24890), 
         .D(zero_baud_counter_N_528), .Z(baud_counter_23__N_483[0])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((C+(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(217[12] 224[43])
    defparam baud_counter_23__I_10_i1_4_lut.init = 16'ha0ac;
    LUT4 i10918_2_lut (.A(n108[0]), .B(zero_baud_counter), .Z(n133[0])) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(224[4:43])
    defparam i10918_2_lut.init = 16'heeee;
    LUT4 i1_2_lut_rep_440 (.A(\state[0] ), .B(state[3]), .Z(n25000)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_440.init = 16'h8888;
    LUT4 i2_3_lut_rep_330_4_lut (.A(\state[0] ), .B(state[3]), .C(state[1]), 
         .D(state[2]), .Z(n24890)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i2_3_lut_rep_330_4_lut.init = 16'h8000;
    FD1S3JX r_busy_45 (.D(n8934), .CK(i_ref_clk_c), .PD(n24992), .Q(tx_busy)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=55, LSE_RCOL=112, LSE_LLINE=63, LSE_RLINE=63 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(92[9] 114[5])
    defparam r_busy_45.GSR = "DISABLED";
    LUT4 state_504_mux_6_i4_4_lut_then_4_lut (.A(n24992), .B(state[2]), 
         .C(\state[0] ), .D(state[1]), .Z(n25235)) /* synthesis lut_function=(!(A (B+(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(110[14:26])
    defparam state_504_mux_6_i4_4_lut_then_4_lut.init = 16'h5557;
    FD1P3AX state_504__i2 (.D(n25229), .SP(zero_baud_counter), .CK(i_ref_clk_c), 
            .Q(state[2]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(110[14:26])
    defparam state_504__i2.GSR = "DISABLED";
    FD1P3AX state_504__i1 (.D(n27[1]), .SP(zero_baud_counter), .CK(i_ref_clk_c), 
            .Q(state[1]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(110[14:26])
    defparam state_504__i1.GSR = "DISABLED";
    FD1P3AX state_504__i0 (.D(n17568), .SP(zero_baud_counter), .CK(i_ref_clk_c), 
            .Q(\state[0] ));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(110[14:26])
    defparam state_504__i0.GSR = "DISABLED";
    LUT4 i22_4_lut (.A(n25), .B(n44), .C(n38), .D(n26), .Z(n46)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(207[24:43])
    defparam i22_4_lut.init = 16'hfffe;
    LUT4 i18_4_lut (.A(baud_counter[19]), .B(baud_counter[13]), .C(baud_counter[2]), 
         .D(baud_counter[14]), .Z(n42)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(207[24:43])
    defparam i18_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut (.A(baud_counter[10]), .B(baud_counter[0]), .Z(n25)) /* synthesis lut_function=(A+!(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(207[24:43])
    defparam i1_2_lut.init = 16'hbbbb;
    LUT4 i20_4_lut (.A(baud_counter[12]), .B(n40), .C(n30), .D(baud_counter[11]), 
         .Z(n44)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(207[24:43])
    defparam i20_4_lut.init = 16'hfffe;
    LUT4 i14_4_lut (.A(baud_counter[8]), .B(baud_counter[1]), .C(baud_counter[9]), 
         .D(baud_counter[6]), .Z(n38)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(207[24:43])
    defparam i14_4_lut.init = 16'hfffe;
    LUT4 i2_2_lut (.A(baud_counter[20]), .B(baud_counter[5]), .Z(n26)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(207[24:43])
    defparam i2_2_lut.init = 16'heeee;
    LUT4 state_504_mux_6_i4_4_lut_else_4_lut (.A(state[2]), .B(\state[0] ), 
         .C(state[1]), .Z(n25234)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(110[14:26])
    defparam state_504_mux_6_i4_4_lut_else_4_lut.init = 16'h8080;
    
endmodule
