// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.11.3.469
// Netlist written on Wed Jan 13 21:49:59 2021
//
// Verilog Description of module top
//

module top (i_ref_clk, i_resetb, i_wbu_uart_rx, o_wbu_uart_tx, o_baseband_i, 
            o_baseband_q, dac_clk_p, dac_clk_n, i_clk_p, i_clk_n, 
            q_clk_p, q_clk_n) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(4[8:11])
    input i_ref_clk;   // d:/documents/git_local/fm_modulator/rtl/top.v(22[12:21])
    input i_resetb;   // d:/documents/git_local/fm_modulator/rtl/top.v(22[23:31])
    input i_wbu_uart_rx;   // d:/documents/git_local/fm_modulator/rtl/top.v(24[12:25])
    output o_wbu_uart_tx;   // d:/documents/git_local/fm_modulator/rtl/top.v(25[13:26])
    output [9:0]o_baseband_i;   // d:/documents/git_local/fm_modulator/rtl/top.v(27[38:50])
    output [9:0]o_baseband_q;   // d:/documents/git_local/fm_modulator/rtl/top.v(27[52:64])
    output dac_clk_p;   // d:/documents/git_local/fm_modulator/rtl/top.v(28[49:58])
    output dac_clk_n;   // d:/documents/git_local/fm_modulator/rtl/top.v(28[60:69])
    output i_clk_p;   // d:/documents/git_local/fm_modulator/rtl/top.v(28[13:20])
    output i_clk_n;   // d:/documents/git_local/fm_modulator/rtl/top.v(28[22:29])
    output q_clk_p;   // d:/documents/git_local/fm_modulator/rtl/top.v(28[31:38])
    output q_clk_n;   // d:/documents/git_local/fm_modulator/rtl/top.v(28[40:47])
    
    wire i_ref_clk_c /* synthesis is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(22[12:21])
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(28[49:58])
    wire o_baseband_i_c_15 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[37:47])
    wire o_baseband_i_c_14 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[37:47])
    wire o_baseband_i_c_13 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[37:47])
    wire o_baseband_i_c_12 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[37:47])
    wire o_baseband_i_c_11 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[37:47])
    wire o_baseband_i_c_10 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[37:47])
    wire n3655 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[37:47])
    wire o_baseband_i_c_8 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[37:47])
    wire o_baseband_i_c_7 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[37:47])
    wire o_baseband_q_c_15 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[49:59])
    wire o_baseband_q_c_14 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[49:59])
    wire o_baseband_q_c_13 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[49:59])
    wire o_baseband_q_c_12 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[49:59])
    wire o_baseband_q_c_11 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[49:59])
    wire o_baseband_q_c_10 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[49:59])
    wire n3656 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[49:59])
    wire o_baseband_q_c_8 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[49:59])
    wire o_baseband_q_c_7 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[49:59])
    wire lo_pll_out /* synthesis is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(160[6:16])
    wire i_clk_2f_N_2249 /* synthesis is_inv_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/clock_phase_shifter.v(11[21:28])
    
    wire GND_net, VCC_net, i_resetb_c, i_wbu_uart_rx_c, o_wbu_uart_tx_c, 
        o_baseband_i_c_9, o_baseband_q_c_9, i_clk_p_c, q_clk_p_c, dac_clk_n_c, 
        i_resetb_N_301, rx_stb;
    wire [7:0]rx_data;   // d:/documents/git_local/fm_modulator/rtl/top.v(51[12:19])
    
    wire tx_busy, wb_cyc, wb_stb, wb_we;
    wire [29:0]wb_addr;   // d:/documents/git_local/fm_modulator/rtl/top.v(68[13:20])
    wire [31:0]wb_odata;   // d:/documents/git_local/fm_modulator/rtl/top.v(69[13:21])
    
    wire wb_ack, wb_err;
    wire [31:0]wb_idata;   // d:/documents/git_local/fm_modulator/rtl/top.v(74[12:20])
    wire [29:0]bus_err_address;   // d:/documents/git_local/fm_modulator/rtl/top.v(98[12:27])
    
    wire wb_fm_ack;
    wire [31:0]wb_fm_data;   // d:/documents/git_local/fm_modulator/rtl/top.v(102[13:23])
    wire [31:0]wb_smpl_data;   // d:/documents/git_local/fm_modulator/rtl/top.v(105[12:24])
    
    wire wb_smpl_ack;
    wire [23:0]chg_counter;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(97[17:28])
    wire [7:0]wb_lo_data;   // d:/documents/git_local/fm_modulator/rtl/top.v(138[12:22])
    
    wire wb_lo_ack, pll_clk, pll_rst, pll_stb, pll_we, pll_ack;
    wire [7:0]pll_data_i;   // d:/documents/git_local/fm_modulator/rtl/top.v(144[12:22])
    wire [7:0]pll_data_o;   // d:/documents/git_local/fm_modulator/rtl/top.v(144[24:34])
    wire [4:0]pll_addr;   // d:/documents/git_local/fm_modulator/rtl/top.v(145[12:20])
    wire [31:0]smpl_register;   // d:/documents/git_local/fm_modulator/rtl/top.v(198[13:26])
    wire [31:0]power_counter;   // d:/documents/git_local/fm_modulator/rtl/top.v(198[28:41])
    
    wire smpl_interrupt, none_sel, wb_fm_data_31__N_63, wb_lo_data_7__N_96, 
        n20801, n20799, n20695;
    wire [31:0]wb_smpl_data_31__N_64;
    wire [31:0]power_counter_31__N_232;
    wire [30:0]power_counter_31__N_201;
    wire [31:0]power_counter_31__N_129;
    
    wire wb_smpl_sel_N_311;
    wire [31:0]wb_idata_31__N_266;
    wire [31:0]wb_idata_31__N_1;
    
    wire chg_counter_23__N_406, n26701, n26730, n20749;
    wire [3:0]state_adj_3085;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(83[12:17])
    wire [7:0]lcl_data;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(84[12:20])
    
    wire zero_baud_counter, o_busy_N_536, n20797;
    wire [7:0]lcl_data_7__N_511;
    
    wire n20745, i_clk_n_c, q_clk_n_c, dac_clk_p_c_enable_273, n20787, 
        n20739, n12737, n21212, n2161, n2160, n2159, n2158, n26695, 
        n2156, n2155, n2154, n26696, n2151, n2150, n2149, n2148, 
        n2147, n26702, n20733, n26703, n26704, n2143, n2141, n2140, 
        n2139, n2138, n2137, n2136, n2135, n2134, n2132, n2131, 
        n2, n7, dac_clk_p_c_enable_175, n26784, n17552, n17551, 
        n17557, n17539, n17569, n17550, n17568, n17549, n17567, 
        n9474, n17548, n17566, n21184, n20755, n20719, n17547, 
        n38, n34, n17565, n21043, n21039, n17545, n17564, n17543, 
        n26699, n9898, n20701, n26762, n26947, n26946, n17563, 
        n17542, n20977, n17562, n20971, n26924, n17561, n17540, 
        n26910, n17560, n17541, n17559, n26897, n17844, dac_clk_p_c_enable_403, 
        n20377, n17546, n17558, n17555, n17554, n17553, n17544, 
        n26694, n17556, dac_clk_p_c_enable_322, n2_adj_3033, n1, n2_adj_3034, 
        n1_adj_3035, n2_adj_3036, n2_adj_3037, n1_adj_3038, n2_adj_3039, 
        n1_adj_3040, n2_adj_3041, n4, n1_adj_3042, n2_adj_3043, n1_adj_3044, 
        n2_adj_3045, n1_adj_3046, n2_adj_3047, n1_adj_3048, n2_adj_3049, 
        n1_adj_3050, n2_adj_3051, n1_adj_3052, n21228, n26805, n2_adj_3053, 
        n2_adj_3054, n1_adj_3055, n2_adj_3056, n2_adj_3057, n21281, 
        n21277, n21226, n2_adj_3058, n2_adj_3059, n1_adj_3060, n2_adj_3061, 
        n1_adj_3062, n2_adj_3063, n1_adj_3064, n2_adj_3065, n1_adj_3066, 
        n2_adj_3067, n1_adj_3068, n2_adj_3069, n2_adj_3070, n2_adj_3071, 
        n1_adj_3072, n2_adj_3073, n1_adj_3074, n2_adj_3075, n1_adj_3076, 
        n2_adj_3077, n2_adj_3078, n1_adj_3079, n2_adj_3080, n1_adj_3081, 
        n2_adj_3082, n1_adj_3083, n21271, n21267, n21265, n29502, 
        n29501, n21261, n21259;
    
    VHI i2 (.Z(VCC_net));
    GSR GSR_INST (.GSR(i_resetb_N_301)) /* synthesis syn_instantiated=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(33[5:28])
    \rxuartlite(CLOCKS_PER_BAUD=10000)  rxtransport (.dac_clk_p_c(dac_clk_p_c), 
            .\rx_data[0] (rx_data[0]), .rx_stb(rx_stb), .i_wbu_uart_rx_c(i_wbu_uart_rx_c), 
            .chg_counter({chg_counter}), .dac_clk_p_c_enable_175(dac_clk_p_c_enable_175), 
            .chg_counter_23__N_406(chg_counter_23__N_406), .GND_net(GND_net), 
            .\rx_data[6] (rx_data[6]), .\rx_data[5] (rx_data[5]), .\rx_data[4] (rx_data[4]), 
            .\rx_data[3] (rx_data[3]), .\rx_data[2] (rx_data[2]), .\rx_data[1] (rx_data[1])) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(53[57:105])
    hbbus genbus (.dac_clk_p_c(dac_clk_p_c), .wb_we(wb_we), .wb_odata({wb_odata}), 
          .wb_stb(wb_stb), .wb_cyc(wb_cyc), .wb_err(wb_err), .wb_ack(wb_ack), 
          .\wb_idata[0] (wb_idata[0]), .wb_addr({wb_addr}), .\wb_idata[2] (wb_idata[2]), 
          .\wb_idata[3] (wb_idata[3]), .\wb_idata[4] (wb_idata[4]), .\wb_idata[5] (wb_idata[5]), 
          .\wb_idata[6] (wb_idata[6]), .\wb_idata[7] (wb_idata[7]), .\wb_idata[8] (wb_idata[8]), 
          .\wb_idata[9] (wb_idata[9]), .\wb_idata[10] (wb_idata[10]), .\wb_idata[11] (wb_idata[11]), 
          .\wb_idata[12] (wb_idata[12]), .\wb_idata[13] (wb_idata[13]), 
          .\wb_idata[14] (wb_idata[14]), .\wb_idata[15] (wb_idata[15]), 
          .\wb_idata[16] (wb_idata[16]), .\wb_idata[17] (wb_idata[17]), 
          .\wb_idata[18] (wb_idata[18]), .\wb_idata[19] (wb_idata[19]), 
          .\wb_idata[20] (wb_idata[20]), .\wb_idata[21] (wb_idata[21]), 
          .\wb_idata[22] (wb_idata[22]), .\wb_idata[23] (wb_idata[23]), 
          .\wb_idata[24] (wb_idata[24]), .\wb_idata[25] (wb_idata[25]), 
          .\wb_idata[26] (wb_idata[26]), .\wb_idata[27] (wb_idata[27]), 
          .\wb_idata[28] (wb_idata[28]), .\wb_idata[29] (wb_idata[29]), 
          .\wb_idata[30] (wb_idata[30]), .\wb_idata[31] (wb_idata[31]), 
          .n2(n2), .GND_net(GND_net), .n12737(n12737), .n29502(n29502), 
          .VCC_net(VCC_net), .rx_stb(rx_stb), .\rx_data[4] (rx_data[4]), 
          .\rx_data[3] (rx_data[3]), .\rx_data[1] (rx_data[1]), .\rx_data[0] (rx_data[0]), 
          .\rx_data[5] (rx_data[5]), .\rx_data[2] (rx_data[2]), .\rx_data[6] (rx_data[6]), 
          .tx_busy(tx_busy), .n26910(n26910), .\lcl_data[1] (lcl_data[1]), 
          .\lcl_data_7__N_511[0] (lcl_data_7__N_511[0]), .\lcl_data[4] (lcl_data[4]), 
          .\lcl_data_7__N_511[3] (lcl_data_7__N_511[3]), .\lcl_data[5] (lcl_data[5]), 
          .\lcl_data_7__N_511[4] (lcl_data_7__N_511[4]), .\lcl_data[6] (lcl_data[6]), 
          .\lcl_data_7__N_511[5] (lcl_data_7__N_511[5]), .zero_baud_counter(zero_baud_counter), 
          .dac_clk_p_c_enable_322(dac_clk_p_c_enable_322), .\lcl_data[7] (lcl_data[7]), 
          .\lcl_data_7__N_511[6] (lcl_data_7__N_511[6]), .\lcl_data[3] (lcl_data[3]), 
          .\lcl_data_7__N_511[2] (lcl_data_7__N_511[2]), .\lcl_data[2] (lcl_data[2]), 
          .\lcl_data_7__N_511[1] (lcl_data_7__N_511[1]), .o_busy_N_536(o_busy_N_536), 
          .\state[0] (state_adj_3085[0]), .n17844(n17844)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(77[7] 93[22])
    FD1S3AX wb_smpl_data_i0 (.D(wb_smpl_data_31__N_64[0]), .CK(dac_clk_p_c), 
            .Q(wb_smpl_data[0]));   // d:/documents/git_local/fm_modulator/rtl/top.v(215[9] 223[10])
    defparam wb_smpl_data_i0.GSR = "DISABLED";
    FD1S3AX power_counter_i0 (.D(power_counter_31__N_129[0]), .CK(dac_clk_p_c), 
            .Q(power_counter[0])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 232[54])
    defparam power_counter_i0.GSR = "DISABLED";
    FD1S3AX wb_idata_i0 (.D(wb_idata_31__N_1[0]), .CK(dac_clk_p_c), .Q(wb_idata[0]));   // d:/documents/git_local/fm_modulator/rtl/top.v(268[9] 276[22])
    defparam wb_idata_i0.GSR = "DISABLED";
    FD1S3JX wb_ack_70 (.D(n4), .CK(dac_clk_p_c), .PD(wb_smpl_ack), .Q(wb_ack)) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(265[9] 266[57])
    defparam wb_ack_70.GSR = "DISABLED";
    PUR PUR_INST (.PUR(i_resetb_N_301)) /* synthesis syn_instantiated=1 */ ;
    defparam PUR_INST.RST_PULSE = 1;
    FD1S3IX wb_smpl_ack_63 (.D(wb_stb), .CK(dac_clk_p_c), .CD(wb_smpl_sel_N_311), 
            .Q(wb_smpl_ack)) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(201[9] 202[44])
    defparam wb_smpl_ack_63.GSR = "DISABLED";
    fm_generator_wb_slave wb_fm_data_31__I_0 (.dac_clk_p_c(dac_clk_p_c), .wb_odata({wb_odata}), 
            .i_resetb_N_301(i_resetb_N_301), .wb_fm_data({wb_fm_data}), 
            .wb_fm_ack(wb_fm_ack), .wb_fm_data_31__N_63(wb_fm_data_31__N_63), 
            .GND_net(GND_net), .\wb_addr[0] (wb_addr[0]), .\wb_addr[1] (wb_addr[1]), 
            .\power_counter[1] (power_counter[1]), .\smpl_register[1] (smpl_register[1]), 
            .n2161(n2161), .n26946(n26946), .n38(n38), .n34(n34), .\wb_addr[8] (wb_addr[8]), 
            .\wb_addr[12] (wb_addr[12]), .n26947(n26947), .\wb_addr[15] (wb_addr[15]), 
            .\wb_addr[9] (wb_addr[9]), .i_resetb_c(i_resetb_c), .n20739(n20739), 
            .n2(n2_adj_3077), .\smpl_register[5] (smpl_register[5]), .n26694(n26694), 
            .n2_adj_1(n2_adj_3053), .\smpl_register[20] (smpl_register[20]), 
            .n26704(n26704), .n2_adj_2(n2_adj_3056), .\smpl_register[18] (smpl_register[18]), 
            .n26703(n26703), .n2_adj_3(n2_adj_3057), .\smpl_register[17] (smpl_register[17]), 
            .n26702(n26702), .n2_adj_4(n2_adj_3058), .\smpl_register[16] (smpl_register[16]), 
            .n26701(n26701), .n2_adj_5(n2_adj_3036), .\smpl_register[29] (smpl_register[29]), 
            .n26699(n26699), .n2_adj_6(n2_adj_3069), .\smpl_register[10] (smpl_register[10]), 
            .n26696(n26696), .n2_adj_7(n2_adj_3070), .\smpl_register[9] (smpl_register[9]), 
            .n26695(n26695), .n20755(n20755), .n21184(n21184), .n20749(n20749), 
            .n20719(n20719), .o_baseband_q_c_7(o_baseband_q_c_7), .o_baseband_i_c_7(o_baseband_i_c_7), 
            .o_baseband_i_c_15(o_baseband_i_c_15), .o_baseband_i_c_14(o_baseband_i_c_14), 
            .o_baseband_i_c_13(o_baseband_i_c_13), .o_baseband_i_c_12(o_baseband_i_c_12), 
            .o_baseband_i_c_11(o_baseband_i_c_11), .o_baseband_i_c_10(o_baseband_i_c_10), 
            .n3655(n3655), .o_baseband_i_c_8(o_baseband_i_c_8), .n29501(n29501), 
            .o_baseband_q_c_15(o_baseband_q_c_15), .o_baseband_q_c_14(o_baseband_q_c_14), 
            .o_baseband_q_c_13(o_baseband_q_c_13), .o_baseband_q_c_12(o_baseband_q_c_12), 
            .o_baseband_q_c_11(o_baseband_q_c_11), .o_baseband_q_c_10(o_baseband_q_c_10), 
            .n3656(n3656), .o_baseband_q_c_8(o_baseband_q_c_8)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(124[2] 135[2])
    FD1P3AX smpl_register_i0_i0 (.D(wb_odata[0]), .SP(dac_clk_p_c_enable_273), 
            .CK(dac_clk_p_c), .Q(smpl_register[0]));   // d:/documents/git_local/fm_modulator/rtl/top.v(205[9] 213[6])
    defparam smpl_register_i0_i0.GSR = "DISABLED";
    FD1S3IX wb_err_68 (.D(none_sel), .CK(dac_clk_p_c), .CD(n2), .Q(wb_err));   // d:/documents/git_local/fm_modulator/rtl/top.v(254[9] 255[34])
    defparam wb_err_68.GSR = "DISABLED";
    LUT4 i1_2_lut (.A(n34), .B(wb_addr[9]), .Z(n20749)) /* synthesis lut_function=(A+!(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[23:49])
    defparam i1_2_lut.init = 16'hbbbb;
    OB o_baseband_i_pad_7 (.I(o_baseband_i_c_14), .O(o_baseband_i[7]));   // d:/documents/git_local/fm_modulator/rtl/top.v(27[38:50])
    OB o_baseband_i_pad_8 (.I(o_baseband_i_c_15), .O(o_baseband_i[8]));   // d:/documents/git_local/fm_modulator/rtl/top.v(27[38:50])
    FD1P3AX bus_err_address_i0_i0 (.D(wb_addr[0]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[0])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(258[9] 260[31])
    defparam bus_err_address_i0_i0.GSR = "DISABLED";
    PFUMX mux_393_Mux_3_i3 (.BLUT(n1_adj_3081), .ALUT(n2_adj_3080), .C0(wb_addr[1]), 
          .Z(n2159));
    OB o_baseband_i_pad_9 (.I(o_baseband_i_c_9), .O(o_baseband_i[9]));   // d:/documents/git_local/fm_modulator/rtl/top.v(27[38:50])
    OB o_wbu_uart_tx_pad (.I(o_wbu_uart_tx_c), .O(o_wbu_uart_tx));   // d:/documents/git_local/fm_modulator/rtl/top.v(25[13:26])
    LUT4 mux_393_Mux_25_i2_3_lut (.A(bus_err_address[23]), .B(power_counter[25]), 
         .C(wb_addr[0]), .Z(n2_adj_3043)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(216[3] 223[10])
    defparam mux_393_Mux_25_i2_3_lut.init = 16'hcaca;
    PFUMX mux_393_Mux_2_i3 (.BLUT(n1_adj_3083), .ALUT(n2_adj_3082), .C0(wb_addr[1]), 
          .Z(n2160));
    CCU2D add_34_27 (.A0(power_counter[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17551), .COUT(n17552), .S0(power_counter_31__N_232[25]), 
          .S1(power_counter_31__N_232[26]));   // d:/documents/git_local/fm_modulator/rtl/top.v(230[21:41])
    defparam add_34_27.INIT0 = 16'h5aaa;
    defparam add_34_27.INIT1 = 16'h5aaa;
    defparam add_34_27.INJECT1_0 = "NO";
    defparam add_34_27.INJECT1_1 = "NO";
    PFUMX mux_393_Mux_23_i3 (.BLUT(n1_adj_3048), .ALUT(n2_adj_3047), .C0(wb_addr[1]), 
          .Z(n2139));
    PFUMX mux_393_Mux_24_i3 (.BLUT(n1_adj_3046), .ALUT(n2_adj_3045), .C0(wb_addr[1]), 
          .Z(n2138));
    PFUMX mux_393_Mux_4_i3 (.BLUT(n1_adj_3079), .ALUT(n2_adj_3078), .C0(wb_addr[1]), 
          .Z(n2158));
    PFUMX mux_393_Mux_6_i3 (.BLUT(n1_adj_3076), .ALUT(n2_adj_3075), .C0(wb_addr[1]), 
          .Z(n2156));
    PFUMX mux_393_Mux_7_i3 (.BLUT(n1_adj_3074), .ALUT(n2_adj_3073), .C0(wb_addr[1]), 
          .Z(n2155));
    PFUMX mux_393_Mux_25_i3 (.BLUT(n1_adj_3044), .ALUT(n2_adj_3043), .C0(wb_addr[1]), 
          .Z(n2137));
    LUT4 i1_4_lut (.A(n21271), .B(n38), .C(n26946), .D(n20701), .Z(dac_clk_p_c_enable_273)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut.init = 16'h0100;
    LUT4 i1_4_lut_adj_139 (.A(n20695), .B(wb_addr[1]), .C(wb_addr[12]), 
         .D(n26947), .Z(n20701)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_4_lut_adj_139.init = 16'h0200;
    LUT4 i1_2_lut_adj_140 (.A(wb_addr[0]), .B(wb_addr[15]), .Z(n20695)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_140.init = 16'h8888;
    PFUMX mux_393_Mux_8_i3 (.BLUT(n1_adj_3072), .ALUT(n2_adj_3071), .C0(wb_addr[1]), 
          .Z(n2154));
    LUT4 i17650_2_lut (.A(wb_addr[2]), .B(wb_addr[3]), .Z(n9474)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i17650_2_lut.init = 16'heeee;
    FD1P3AX smpl_register_i0_i31 (.D(wb_odata[31]), .SP(dac_clk_p_c_enable_273), 
            .CK(dac_clk_p_c), .Q(smpl_register[31]));   // d:/documents/git_local/fm_modulator/rtl/top.v(205[9] 213[6])
    defparam smpl_register_i0_i31.GSR = "DISABLED";
    LUT4 i1_3_lut_4_lut (.A(wb_addr[1]), .B(n26897), .C(wb_addr[15]), 
         .D(n26946), .Z(n20719)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[23:49])
    defparam i1_3_lut_4_lut.init = 16'hffef;
    FD1P3AX smpl_register_i0_i30 (.D(wb_odata[30]), .SP(dac_clk_p_c_enable_273), 
            .CK(dac_clk_p_c), .Q(smpl_register[30]));   // d:/documents/git_local/fm_modulator/rtl/top.v(205[9] 213[6])
    defparam smpl_register_i0_i30.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i29 (.D(wb_odata[29]), .SP(dac_clk_p_c_enable_273), 
            .CK(dac_clk_p_c), .Q(smpl_register[29]));   // d:/documents/git_local/fm_modulator/rtl/top.v(205[9] 213[6])
    defparam smpl_register_i0_i29.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i28 (.D(wb_odata[28]), .SP(dac_clk_p_c_enable_273), 
            .CK(dac_clk_p_c), .Q(smpl_register[28]));   // d:/documents/git_local/fm_modulator/rtl/top.v(205[9] 213[6])
    defparam smpl_register_i0_i28.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i27 (.D(wb_odata[27]), .SP(dac_clk_p_c_enable_273), 
            .CK(dac_clk_p_c), .Q(smpl_register[27]));   // d:/documents/git_local/fm_modulator/rtl/top.v(205[9] 213[6])
    defparam smpl_register_i0_i27.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i26 (.D(wb_odata[26]), .SP(dac_clk_p_c_enable_273), 
            .CK(dac_clk_p_c), .Q(smpl_register[26]));   // d:/documents/git_local/fm_modulator/rtl/top.v(205[9] 213[6])
    defparam smpl_register_i0_i26.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i25 (.D(wb_odata[25]), .SP(dac_clk_p_c_enable_273), 
            .CK(dac_clk_p_c), .Q(smpl_register[25]));   // d:/documents/git_local/fm_modulator/rtl/top.v(205[9] 213[6])
    defparam smpl_register_i0_i25.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i24 (.D(wb_odata[24]), .SP(dac_clk_p_c_enable_273), 
            .CK(dac_clk_p_c), .Q(smpl_register[24]));   // d:/documents/git_local/fm_modulator/rtl/top.v(205[9] 213[6])
    defparam smpl_register_i0_i24.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i23 (.D(wb_odata[23]), .SP(dac_clk_p_c_enable_273), 
            .CK(dac_clk_p_c), .Q(smpl_register[23]));   // d:/documents/git_local/fm_modulator/rtl/top.v(205[9] 213[6])
    defparam smpl_register_i0_i23.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i22 (.D(wb_odata[22]), .SP(dac_clk_p_c_enable_273), 
            .CK(dac_clk_p_c), .Q(smpl_register[22]));   // d:/documents/git_local/fm_modulator/rtl/top.v(205[9] 213[6])
    defparam smpl_register_i0_i22.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i21 (.D(wb_odata[21]), .SP(dac_clk_p_c_enable_273), 
            .CK(dac_clk_p_c), .Q(smpl_register[21]));   // d:/documents/git_local/fm_modulator/rtl/top.v(205[9] 213[6])
    defparam smpl_register_i0_i21.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i20 (.D(wb_odata[20]), .SP(dac_clk_p_c_enable_273), 
            .CK(dac_clk_p_c), .Q(smpl_register[20]));   // d:/documents/git_local/fm_modulator/rtl/top.v(205[9] 213[6])
    defparam smpl_register_i0_i20.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i19 (.D(wb_odata[19]), .SP(dac_clk_p_c_enable_273), 
            .CK(dac_clk_p_c), .Q(smpl_register[19]));   // d:/documents/git_local/fm_modulator/rtl/top.v(205[9] 213[6])
    defparam smpl_register_i0_i19.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i18 (.D(wb_odata[18]), .SP(dac_clk_p_c_enable_273), 
            .CK(dac_clk_p_c), .Q(smpl_register[18]));   // d:/documents/git_local/fm_modulator/rtl/top.v(205[9] 213[6])
    defparam smpl_register_i0_i18.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i17 (.D(wb_odata[17]), .SP(dac_clk_p_c_enable_273), 
            .CK(dac_clk_p_c), .Q(smpl_register[17]));   // d:/documents/git_local/fm_modulator/rtl/top.v(205[9] 213[6])
    defparam smpl_register_i0_i17.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i16 (.D(wb_odata[16]), .SP(dac_clk_p_c_enable_273), 
            .CK(dac_clk_p_c), .Q(smpl_register[16]));   // d:/documents/git_local/fm_modulator/rtl/top.v(205[9] 213[6])
    defparam smpl_register_i0_i16.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i15 (.D(wb_odata[15]), .SP(dac_clk_p_c_enable_273), 
            .CK(dac_clk_p_c), .Q(smpl_register[15]));   // d:/documents/git_local/fm_modulator/rtl/top.v(205[9] 213[6])
    defparam smpl_register_i0_i15.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i14 (.D(wb_odata[14]), .SP(dac_clk_p_c_enable_273), 
            .CK(dac_clk_p_c), .Q(smpl_register[14]));   // d:/documents/git_local/fm_modulator/rtl/top.v(205[9] 213[6])
    defparam smpl_register_i0_i14.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i13 (.D(wb_odata[13]), .SP(dac_clk_p_c_enable_273), 
            .CK(dac_clk_p_c), .Q(smpl_register[13]));   // d:/documents/git_local/fm_modulator/rtl/top.v(205[9] 213[6])
    defparam smpl_register_i0_i13.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i12 (.D(wb_odata[12]), .SP(dac_clk_p_c_enable_273), 
            .CK(dac_clk_p_c), .Q(smpl_register[12]));   // d:/documents/git_local/fm_modulator/rtl/top.v(205[9] 213[6])
    defparam smpl_register_i0_i12.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i11 (.D(wb_odata[11]), .SP(dac_clk_p_c_enable_273), 
            .CK(dac_clk_p_c), .Q(smpl_register[11]));   // d:/documents/git_local/fm_modulator/rtl/top.v(205[9] 213[6])
    defparam smpl_register_i0_i11.GSR = "DISABLED";
    LUT4 wb_idata_31__I_0_i32_4_lut (.A(wb_smpl_data[31]), .B(wb_fm_data[31]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_1[31])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(271[8] 276[22])
    defparam wb_idata_31__I_0_i32_4_lut.init = 16'hcac0;
    FD1P3AX smpl_register_i0_i10 (.D(wb_odata[10]), .SP(dac_clk_p_c_enable_273), 
            .CK(dac_clk_p_c), .Q(smpl_register[10]));   // d:/documents/git_local/fm_modulator/rtl/top.v(205[9] 213[6])
    defparam smpl_register_i0_i10.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i9 (.D(wb_odata[9]), .SP(dac_clk_p_c_enable_273), 
            .CK(dac_clk_p_c), .Q(smpl_register[9]));   // d:/documents/git_local/fm_modulator/rtl/top.v(205[9] 213[6])
    defparam smpl_register_i0_i9.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i8 (.D(wb_odata[8]), .SP(dac_clk_p_c_enable_273), 
            .CK(dac_clk_p_c), .Q(smpl_register[8]));   // d:/documents/git_local/fm_modulator/rtl/top.v(205[9] 213[6])
    defparam smpl_register_i0_i8.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i7 (.D(wb_odata[7]), .SP(dac_clk_p_c_enable_273), 
            .CK(dac_clk_p_c), .Q(smpl_register[7]));   // d:/documents/git_local/fm_modulator/rtl/top.v(205[9] 213[6])
    defparam smpl_register_i0_i7.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i6 (.D(wb_odata[6]), .SP(dac_clk_p_c_enable_273), 
            .CK(dac_clk_p_c), .Q(smpl_register[6]));   // d:/documents/git_local/fm_modulator/rtl/top.v(205[9] 213[6])
    defparam smpl_register_i0_i6.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i5 (.D(wb_odata[5]), .SP(dac_clk_p_c_enable_273), 
            .CK(dac_clk_p_c), .Q(smpl_register[5]));   // d:/documents/git_local/fm_modulator/rtl/top.v(205[9] 213[6])
    defparam smpl_register_i0_i5.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i4 (.D(wb_odata[4]), .SP(dac_clk_p_c_enable_273), 
            .CK(dac_clk_p_c), .Q(smpl_register[4]));   // d:/documents/git_local/fm_modulator/rtl/top.v(205[9] 213[6])
    defparam smpl_register_i0_i4.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i3 (.D(wb_odata[3]), .SP(dac_clk_p_c_enable_273), 
            .CK(dac_clk_p_c), .Q(smpl_register[3]));   // d:/documents/git_local/fm_modulator/rtl/top.v(205[9] 213[6])
    defparam smpl_register_i0_i3.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i2 (.D(wb_odata[2]), .SP(dac_clk_p_c_enable_273), 
            .CK(dac_clk_p_c), .Q(smpl_register[2]));   // d:/documents/git_local/fm_modulator/rtl/top.v(205[9] 213[6])
    defparam smpl_register_i0_i2.GSR = "DISABLED";
    FD1P3AX smpl_register_i0_i1 (.D(wb_odata[1]), .SP(dac_clk_p_c_enable_273), 
            .CK(dac_clk_p_c), .Q(smpl_register[1]));   // d:/documents/git_local/fm_modulator/rtl/top.v(205[9] 213[6])
    defparam smpl_register_i0_i1.GSR = "DISABLED";
    PFUMX mux_393_Mux_11_i3 (.BLUT(n1_adj_3068), .ALUT(n2_adj_3067), .C0(wb_addr[1]), 
          .Z(n2151));
    LUT4 i1_4_lut_adj_141 (.A(n21261), .B(n21281), .C(n21277), .D(chg_counter_23__N_406), 
         .Z(dac_clk_p_c_enable_175)) /* synthesis lut_function=((((D)+!C)+!B)+!A) */ ;
    defparam i1_4_lut_adj_141.init = 16'hff7f;
    LUT4 i18899_4_lut (.A(chg_counter[2]), .B(chg_counter[7]), .C(chg_counter[10]), 
         .D(chg_counter[11]), .Z(n21261)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i18899_4_lut.init = 16'h8000;
    LUT4 i18919_4_lut (.A(n21226), .B(n21267), .C(n21265), .D(n21228), 
         .Z(n21281)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i18919_4_lut.init = 16'h8000;
    LUT4 i18915_4_lut (.A(chg_counter[18]), .B(n21259), .C(n21212), .D(chg_counter[3]), 
         .Z(n21277)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i18915_4_lut.init = 16'h8000;
    LUT4 i18865_2_lut (.A(chg_counter[9]), .B(chg_counter[5]), .Z(n21226)) /* synthesis lut_function=(A (B)) */ ;
    defparam i18865_2_lut.init = 16'h8888;
    LUT4 i18905_4_lut (.A(chg_counter[1]), .B(chg_counter[15]), .C(chg_counter[16]), 
         .D(chg_counter[14]), .Z(n21267)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i18905_4_lut.init = 16'h8000;
    LUT4 i18903_4_lut (.A(chg_counter[23]), .B(chg_counter[8]), .C(chg_counter[17]), 
         .D(chg_counter[13]), .Z(n21265)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i18903_4_lut.init = 16'h8000;
    LUT4 i18867_2_lut (.A(chg_counter[12]), .B(chg_counter[19]), .Z(n21228)) /* synthesis lut_function=(A (B)) */ ;
    defparam i18867_2_lut.init = 16'h8888;
    LUT4 i18897_4_lut (.A(chg_counter[20]), .B(chg_counter[6]), .C(chg_counter[21]), 
         .D(chg_counter[0]), .Z(n21259)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i18897_4_lut.init = 16'h8000;
    LUT4 i18851_2_lut (.A(chg_counter[22]), .B(chg_counter[4]), .Z(n21212)) /* synthesis lut_function=(A (B)) */ ;
    defparam i18851_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_142 (.A(wb_addr[8]), .B(n26762), .C(n21043), .D(wb_addr[9]), 
         .Z(none_sel)) /* synthesis lut_function=(A (B+(C))+!A (B+(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[23:49])
    defparam i1_4_lut_adj_142.init = 16'hfcfd;
    LUT4 i_resetb_I_0_1_lut (.A(i_resetb_c), .Z(i_resetb_N_301)) /* synthesis lut_function=(!(A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(31[16:25])
    defparam i_resetb_I_0_1_lut.init = 16'h5555;
    LUT4 i1_4_lut_adj_143 (.A(n26946), .B(n38), .C(n34), .D(n20977), 
         .Z(wb_fm_data_31__N_63)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut_adj_143.init = 16'h0100;
    LUT4 i1_4_lut_adj_144 (.A(wb_addr[8]), .B(wb_addr[12]), .C(n20971), 
         .D(wb_addr[9]), .Z(n20977)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_4_lut_adj_144.init = 16'h1000;
    LUT4 i1_2_lut_adj_145 (.A(wb_addr[15]), .B(wb_stb), .Z(n20971)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_145.init = 16'h8888;
    LUT4 i763_1_lut (.A(o_baseband_i_c_15), .Z(o_baseband_i_c_9)) /* synthesis lut_function=(!(A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(113[31:66])
    defparam i763_1_lut.init = 16'h5555;
    LUT4 i1_2_lut_rep_407_3_lut_4_lut (.A(n26946), .B(wb_addr[12]), .C(n21043), 
         .D(n38), .Z(n26730)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[23:49])
    defparam i1_2_lut_rep_407_3_lut_4_lut.init = 16'hfffe;
    LUT4 i11133_2_lut (.A(smpl_register[22]), .B(wb_addr[0]), .Z(n1_adj_3050)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(216[3] 223[10])
    defparam i11133_2_lut.init = 16'h8888;
    LUT4 mux_392_i1_4_lut (.A(smpl_interrupt), .B(n21039), .C(n7), .D(n9898), 
         .Z(wb_smpl_data_31__N_64[0])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(216[3] 223[10])
    defparam mux_392_i1_4_lut.init = 16'hca0a;
    LUT4 mux_393_Mux_21_i2_3_lut (.A(bus_err_address[19]), .B(power_counter[21]), 
         .C(wb_addr[0]), .Z(n2_adj_3051)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(216[3] 223[10])
    defparam mux_393_Mux_21_i2_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut (.A(wb_addr[3]), .B(wb_addr[2]), .C(wb_addr[0]), .Z(n21039)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_3_lut.init = 16'h1010;
    LUT4 i7402_3_lut (.A(smpl_register[0]), .B(power_counter[0]), .C(wb_addr[1]), 
         .Z(n9898)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(216[3] 223[10])
    defparam i7402_3_lut.init = 16'hcaca;
    LUT4 i11132_2_lut (.A(smpl_register[21]), .B(wb_addr[0]), .Z(n1_adj_3052)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(216[3] 223[10])
    defparam i11132_2_lut.init = 16'h8888;
    LUT4 mux_393_Mux_20_i2_3_lut (.A(bus_err_address[18]), .B(power_counter[20]), 
         .C(wb_addr[0]), .Z(n2_adj_3053)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(216[3] 223[10])
    defparam mux_393_Mux_20_i2_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_146 (.A(wb_addr[1]), .B(wb_addr[2]), .C(wb_addr[0]), 
         .D(wb_addr[3]), .Z(n7)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(210[4:8])
    defparam i1_4_lut_adj_146.init = 16'hfffb;
    LUT4 mux_393_Mux_19_i2_3_lut (.A(bus_err_address[17]), .B(power_counter[19]), 
         .C(wb_addr[0]), .Z(n2_adj_3054)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(216[3] 223[10])
    defparam mux_393_Mux_19_i2_3_lut.init = 16'hcaca;
    LUT4 i11130_2_lut (.A(smpl_register[19]), .B(wb_addr[0]), .Z(n1_adj_3055)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(216[3] 223[10])
    defparam i11130_2_lut.init = 16'h8888;
    LUT4 mux_393_Mux_18_i2_3_lut (.A(bus_err_address[16]), .B(power_counter[18]), 
         .C(wb_addr[0]), .Z(n2_adj_3056)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(216[3] 223[10])
    defparam mux_393_Mux_18_i2_3_lut.init = 16'hcaca;
    LUT4 mux_393_Mux_17_i2_3_lut (.A(bus_err_address[15]), .B(power_counter[17]), 
         .C(wb_addr[0]), .Z(n2_adj_3057)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(216[3] 223[10])
    defparam mux_393_Mux_17_i2_3_lut.init = 16'hcaca;
    LUT4 mux_393_Mux_16_i2_3_lut (.A(bus_err_address[14]), .B(power_counter[16]), 
         .C(wb_addr[0]), .Z(n2_adj_3058)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(216[3] 223[10])
    defparam mux_393_Mux_16_i2_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_147 (.A(n20797), .B(n20799), .C(n20801), .D(n20787), 
         .Z(n38)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[23:49])
    defparam i1_4_lut_adj_147.init = 16'hfffe;
    LUT4 i1_2_lut_adj_148 (.A(wb_addr[11]), .B(wb_addr[16]), .Z(n20797)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[23:49])
    defparam i1_2_lut_adj_148.init = 16'heeee;
    LUT4 i1_4_lut_adj_149 (.A(wb_addr[17]), .B(wb_addr[14]), .C(wb_addr[23]), 
         .D(wb_addr[20]), .Z(n20799)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[23:49])
    defparam i1_4_lut_adj_149.init = 16'hfffe;
    LUT4 i1_4_lut_adj_150 (.A(wb_addr[25]), .B(wb_addr[10]), .C(wb_addr[26]), 
         .D(wb_addr[21]), .Z(n20801)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[23:49])
    defparam i1_4_lut_adj_150.init = 16'hfffe;
    LUT4 i1_2_lut_adj_151 (.A(wb_addr[27]), .B(wb_addr[18]), .Z(n20787)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[23:49])
    defparam i1_2_lut_adj_151.init = 16'heeee;
    LUT4 i1_4_lut_adj_152 (.A(wb_addr[28]), .B(wb_addr[19]), .C(wb_addr[13]), 
         .D(wb_addr[29]), .Z(n34)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[23:49])
    defparam i1_4_lut_adj_152.init = 16'hfffe;
    LUT4 mux_393_Mux_15_i2_3_lut (.A(bus_err_address[13]), .B(power_counter[15]), 
         .C(wb_addr[0]), .Z(n2_adj_3059)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(216[3] 223[10])
    defparam mux_393_Mux_15_i2_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_77_i1_3_lut (.A(power_counter_31__N_232[0]), 
         .B(power_counter_31__N_201[0]), .C(power_counter[31]), .Z(power_counter_31__N_129[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(232[4:54])
    defparam power_counter_31__I_0_77_i1_3_lut.init = 16'hcaca;
    LUT4 wb_idata_31__I_0_i1_3_lut (.A(wb_idata_31__N_266[0]), .B(wb_fm_data[0]), 
         .C(wb_fm_ack), .Z(wb_idata_31__N_1[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(271[8] 276[22])
    defparam wb_idata_31__I_0_i1_3_lut.init = 16'hcaca;
    LUT4 mux_59_i1_4_lut (.A(wb_lo_data[0]), .B(wb_smpl_data[0]), .C(wb_smpl_ack), 
         .D(wb_lo_ack), .Z(wb_idata_31__N_266[0])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(273[8] 276[22])
    defparam mux_59_i1_4_lut.init = 16'hcac0;
    LUT4 i1_2_lut_adj_153 (.A(wb_fm_ack), .B(wb_lo_ack), .Z(n4)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(266[13:56])
    defparam i1_2_lut_adj_153.init = 16'heeee;
    LUT4 i11126_2_lut (.A(smpl_register[15]), .B(wb_addr[0]), .Z(n1_adj_3060)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(216[3] 223[10])
    defparam i11126_2_lut.init = 16'h8888;
    PFUMX mux_393_Mux_26_i3 (.BLUT(n1_adj_3042), .ALUT(n2_adj_3041), .C0(wb_addr[1]), 
          .Z(n2136));
    LUT4 i1_2_lut_adj_154 (.A(wb_addr[15]), .B(n34), .Z(n21043)) /* synthesis lut_function=((B)+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[23:49])
    defparam i1_2_lut_adj_154.init = 16'hdddd;
    LUT4 i11113_2_lut (.A(smpl_register[2]), .B(wb_addr[0]), .Z(n1_adj_3083)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(216[3] 223[10])
    defparam i11113_2_lut.init = 16'h8888;
    PFUMX mux_393_Mux_12_i3 (.BLUT(n1_adj_3066), .ALUT(n2_adj_3065), .C0(wb_addr[1]), 
          .Z(n2150));
    PFUMX mux_393_Mux_27_i3 (.BLUT(n1_adj_3040), .ALUT(n2_adj_3039), .C0(wb_addr[1]), 
          .Z(n2135));
    LUT4 mux_393_Mux_14_i2_3_lut (.A(bus_err_address[12]), .B(power_counter[14]), 
         .C(wb_addr[0]), .Z(n2_adj_3061)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(216[3] 223[10])
    defparam mux_393_Mux_14_i2_3_lut.init = 16'hcaca;
    LUT4 i11125_2_lut (.A(smpl_register[14]), .B(wb_addr[0]), .Z(n1_adj_3062)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(216[3] 223[10])
    defparam i11125_2_lut.init = 16'h8888;
    LUT4 mux_393_Mux_31_i2_3_lut (.A(bus_err_address[29]), .B(power_counter[31]), 
         .C(wb_addr[0]), .Z(n2_adj_3033)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(216[3] 223[10])
    defparam mux_393_Mux_31_i2_3_lut.init = 16'hcaca;
    LUT4 i11142_2_lut (.A(smpl_register[31]), .B(wb_addr[0]), .Z(n1)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(216[3] 223[10])
    defparam i11142_2_lut.init = 16'h8888;
    LUT4 mux_393_Mux_30_i2_3_lut (.A(bus_err_address[28]), .B(power_counter[30]), 
         .C(wb_addr[0]), .Z(n2_adj_3034)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(216[3] 223[10])
    defparam mux_393_Mux_30_i2_3_lut.init = 16'hcaca;
    LUT4 i11141_2_lut (.A(smpl_register[30]), .B(wb_addr[0]), .Z(n1_adj_3035)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(216[3] 223[10])
    defparam i11141_2_lut.init = 16'h8888;
    LUT4 mux_393_Mux_13_i2_3_lut (.A(bus_err_address[11]), .B(power_counter[13]), 
         .C(wb_addr[0]), .Z(n2_adj_3063)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(216[3] 223[10])
    defparam mux_393_Mux_13_i2_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n38), .B(n26805), .C(n26924), .D(n21043), 
         .Z(wb_smpl_sel_N_311)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[23:49])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 mux_393_Mux_29_i2_3_lut (.A(bus_err_address[27]), .B(power_counter[29]), 
         .C(wb_addr[0]), .Z(n2_adj_3036)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(216[3] 223[10])
    defparam mux_393_Mux_29_i2_3_lut.init = 16'hcaca;
    LUT4 i11124_2_lut (.A(smpl_register[13]), .B(wb_addr[0]), .Z(n1_adj_3064)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(216[3] 223[10])
    defparam i11124_2_lut.init = 16'h8888;
    LUT4 mux_393_Mux_28_i2_3_lut (.A(bus_err_address[26]), .B(power_counter[28]), 
         .C(wb_addr[0]), .Z(n2_adj_3037)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(216[3] 223[10])
    defparam mux_393_Mux_28_i2_3_lut.init = 16'hcaca;
    LUT4 i11139_2_lut (.A(smpl_register[28]), .B(wb_addr[0]), .Z(n1_adj_3038)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(216[3] 223[10])
    defparam i11139_2_lut.init = 16'h8888;
    LUT4 mux_393_Mux_27_i2_3_lut (.A(bus_err_address[25]), .B(power_counter[27]), 
         .C(wb_addr[0]), .Z(n2_adj_3039)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(216[3] 223[10])
    defparam mux_393_Mux_27_i2_3_lut.init = 16'hcaca;
    LUT4 i11138_2_lut (.A(smpl_register[27]), .B(wb_addr[0]), .Z(n1_adj_3040)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(216[3] 223[10])
    defparam i11138_2_lut.init = 16'h8888;
    LUT4 mux_393_Mux_12_i2_3_lut (.A(bus_err_address[10]), .B(power_counter[12]), 
         .C(wb_addr[0]), .Z(n2_adj_3065)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(216[3] 223[10])
    defparam mux_393_Mux_12_i2_3_lut.init = 16'hcaca;
    PFUMX mux_393_Mux_28_i3 (.BLUT(n1_adj_3038), .ALUT(n2_adj_3037), .C0(wb_addr[1]), 
          .Z(n2134));
    PFUMX mux_393_Mux_13_i3 (.BLUT(n1_adj_3064), .ALUT(n2_adj_3063), .C0(wb_addr[1]), 
          .Z(n2149));
    CCU2D add_34_25 (.A0(power_counter[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17550), .COUT(n17551), .S0(power_counter_31__N_232[23]), 
          .S1(power_counter_31__N_232[24]));   // d:/documents/git_local/fm_modulator/rtl/top.v(230[21:41])
    defparam add_34_25.INIT0 = 16'h5aaa;
    defparam add_34_25.INIT1 = 16'h5aaa;
    defparam add_34_25.INJECT1_0 = "NO";
    defparam add_34_25.INJECT1_1 = "NO";
    CCU2D add_35_31 (.A0(power_counter[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17569), .S0(power_counter_31__N_201[29]), 
          .S1(power_counter_31__N_201[30]));   // d:/documents/git_local/fm_modulator/rtl/top.v(232[27:53])
    defparam add_35_31.INIT0 = 16'h5aaa;
    defparam add_35_31.INIT1 = 16'h5aaa;
    defparam add_35_31.INJECT1_0 = "NO";
    defparam add_35_31.INJECT1_1 = "NO";
    LUT4 i11123_2_lut (.A(smpl_register[12]), .B(wb_addr[0]), .Z(n1_adj_3066)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(216[3] 223[10])
    defparam i11123_2_lut.init = 16'h8888;
    PFUMX mux_393_Mux_30_i3 (.BLUT(n1_adj_3035), .ALUT(n2_adj_3034), .C0(wb_addr[1]), 
          .Z(n2132));
    LUT4 mux_393_Mux_26_i2_3_lut (.A(bus_err_address[24]), .B(power_counter[26]), 
         .C(wb_addr[0]), .Z(n2_adj_3041)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(216[3] 223[10])
    defparam mux_393_Mux_26_i2_3_lut.init = 16'hcaca;
    PFUMX mux_393_Mux_31_i3 (.BLUT(n1), .ALUT(n2_adj_3033), .C0(wb_addr[1]), 
          .Z(n2131));
    LUT4 i11137_2_lut (.A(smpl_register[26]), .B(wb_addr[0]), .Z(n1_adj_3042)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(216[3] 223[10])
    defparam i11137_2_lut.init = 16'h8888;
    PFUMX mux_393_Mux_14_i3 (.BLUT(n1_adj_3062), .ALUT(n2_adj_3061), .C0(wb_addr[1]), 
          .Z(n2148));
    CCU2D add_34_23 (.A0(power_counter[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17549), .COUT(n17550), .S0(power_counter_31__N_232[21]), 
          .S1(power_counter_31__N_232[22]));   // d:/documents/git_local/fm_modulator/rtl/top.v(230[21:41])
    defparam add_34_23.INIT0 = 16'h5aaa;
    defparam add_34_23.INIT1 = 16'h5aaa;
    defparam add_34_23.INJECT1_0 = "NO";
    defparam add_34_23.INJECT1_1 = "NO";
    FD1S3AX wb_idata_i31 (.D(wb_idata_31__N_1[31]), .CK(dac_clk_p_c), .Q(wb_idata[31]));   // d:/documents/git_local/fm_modulator/rtl/top.v(268[9] 276[22])
    defparam wb_idata_i31.GSR = "DISABLED";
    LUT4 wb_idata_31__I_0_i31_4_lut (.A(wb_smpl_data[30]), .B(wb_fm_data[30]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_1[30])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(271[8] 276[22])
    defparam wb_idata_31__I_0_i31_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i30_4_lut (.A(wb_smpl_data[29]), .B(wb_fm_data[29]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_1[29])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(271[8] 276[22])
    defparam wb_idata_31__I_0_i30_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i29_4_lut (.A(wb_smpl_data[28]), .B(wb_fm_data[28]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_1[28])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(271[8] 276[22])
    defparam wb_idata_31__I_0_i29_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i28_4_lut (.A(wb_smpl_data[27]), .B(wb_fm_data[27]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_1[27])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(271[8] 276[22])
    defparam wb_idata_31__I_0_i28_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i27_4_lut (.A(wb_smpl_data[26]), .B(wb_fm_data[26]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_1[26])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(271[8] 276[22])
    defparam wb_idata_31__I_0_i27_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i26_4_lut (.A(wb_smpl_data[25]), .B(wb_fm_data[25]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_1[25])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(271[8] 276[22])
    defparam wb_idata_31__I_0_i26_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i25_4_lut (.A(wb_smpl_data[24]), .B(wb_fm_data[24]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_1[24])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(271[8] 276[22])
    defparam wb_idata_31__I_0_i25_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i24_4_lut (.A(wb_smpl_data[23]), .B(wb_fm_data[23]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_1[23])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(271[8] 276[22])
    defparam wb_idata_31__I_0_i24_4_lut.init = 16'hcac0;
    LUT4 i22625_4_lut (.A(n26730), .B(n26924), .C(n26947), .D(n7), .Z(dac_clk_p_c_enable_403)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(205[9] 213[6])
    defparam i22625_4_lut.init = 16'h0010;
    LUT4 i10095_1_lut (.A(wb_idata[1]), .Z(n12737)) /* synthesis lut_function=(!(A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(268[9] 276[22])
    defparam i10095_1_lut.init = 16'h5555;
    LUT4 wb_idata_31__I_0_i23_4_lut (.A(wb_smpl_data[22]), .B(wb_fm_data[22]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_1[22])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(271[8] 276[22])
    defparam wb_idata_31__I_0_i23_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i22_4_lut (.A(wb_smpl_data[21]), .B(wb_fm_data[21]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_1[21])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(271[8] 276[22])
    defparam wb_idata_31__I_0_i22_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i21_4_lut (.A(wb_smpl_data[20]), .B(wb_fm_data[20]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_1[20])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(271[8] 276[22])
    defparam wb_idata_31__I_0_i21_4_lut.init = 16'hcac0;
    LUT4 i11136_2_lut (.A(smpl_register[25]), .B(wb_addr[0]), .Z(n1_adj_3044)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(216[3] 223[10])
    defparam i11136_2_lut.init = 16'h8888;
    LUT4 wb_idata_31__I_0_i20_4_lut (.A(wb_smpl_data[19]), .B(wb_fm_data[19]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_1[19])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(271[8] 276[22])
    defparam wb_idata_31__I_0_i20_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i19_4_lut (.A(wb_smpl_data[18]), .B(wb_fm_data[18]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_1[18])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(271[8] 276[22])
    defparam wb_idata_31__I_0_i19_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i18_4_lut (.A(wb_smpl_data[17]), .B(wb_fm_data[17]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_1[17])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(271[8] 276[22])
    defparam wb_idata_31__I_0_i18_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i17_4_lut (.A(wb_smpl_data[16]), .B(wb_fm_data[16]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_1[16])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(271[8] 276[22])
    defparam wb_idata_31__I_0_i17_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i16_4_lut (.A(wb_smpl_data[15]), .B(wb_fm_data[15]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_1[15])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(271[8] 276[22])
    defparam wb_idata_31__I_0_i16_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i15_4_lut (.A(wb_smpl_data[14]), .B(wb_fm_data[14]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_1[14])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(271[8] 276[22])
    defparam wb_idata_31__I_0_i15_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i14_4_lut (.A(wb_smpl_data[13]), .B(wb_fm_data[13]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_1[13])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(271[8] 276[22])
    defparam wb_idata_31__I_0_i14_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i13_4_lut (.A(wb_smpl_data[12]), .B(wb_fm_data[12]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_1[12])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(271[8] 276[22])
    defparam wb_idata_31__I_0_i13_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i12_4_lut (.A(wb_smpl_data[11]), .B(wb_fm_data[11]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_1[11])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(271[8] 276[22])
    defparam wb_idata_31__I_0_i12_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i11_4_lut (.A(wb_smpl_data[10]), .B(wb_fm_data[10]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_1[10])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(271[8] 276[22])
    defparam wb_idata_31__I_0_i11_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i10_4_lut (.A(wb_smpl_data[9]), .B(wb_fm_data[9]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_1[9])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(271[8] 276[22])
    defparam wb_idata_31__I_0_i10_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i9_4_lut (.A(wb_smpl_data[8]), .B(wb_fm_data[8]), 
         .C(wb_fm_ack), .D(wb_smpl_ack), .Z(wb_idata_31__N_1[8])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(271[8] 276[22])
    defparam wb_idata_31__I_0_i9_4_lut.init = 16'hcac0;
    LUT4 i1_2_lut_rep_601 (.A(wb_addr[9]), .B(wb_addr[8]), .Z(n26924)) /* synthesis lut_function=(A+!(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[23:49])
    defparam i1_2_lut_rep_601.init = 16'hbbbb;
    LUT4 i18909_3_lut_4_lut (.A(wb_addr[9]), .B(wb_addr[8]), .C(n34), 
         .D(n9474), .Z(n21271)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[23:49])
    defparam i18909_3_lut_4_lut.init = 16'hfffb;
    LUT4 wb_idata_31__I_0_i8_3_lut (.A(wb_idata_31__N_266[7]), .B(wb_fm_data[7]), 
         .C(wb_fm_ack), .Z(wb_idata_31__N_1[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(271[8] 276[22])
    defparam wb_idata_31__I_0_i8_3_lut.init = 16'hcaca;
    LUT4 mux_59_i8_4_lut (.A(wb_lo_data[7]), .B(wb_smpl_data[7]), .C(wb_smpl_ack), 
         .D(wb_lo_ack), .Z(wb_idata_31__N_266[7])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(273[8] 276[22])
    defparam mux_59_i8_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i7_3_lut (.A(wb_idata_31__N_266[6]), .B(wb_fm_data[6]), 
         .C(wb_fm_ack), .Z(wb_idata_31__N_1[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(271[8] 276[22])
    defparam wb_idata_31__I_0_i7_3_lut.init = 16'hcaca;
    LUT4 mux_59_i7_4_lut (.A(wb_lo_data[6]), .B(wb_smpl_data[6]), .C(wb_smpl_ack), 
         .D(wb_lo_ack), .Z(wb_idata_31__N_266[6])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(273[8] 276[22])
    defparam mux_59_i7_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i6_3_lut (.A(wb_idata_31__N_266[5]), .B(wb_fm_data[5]), 
         .C(wb_fm_ack), .Z(wb_idata_31__N_1[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(271[8] 276[22])
    defparam wb_idata_31__I_0_i6_3_lut.init = 16'hcaca;
    LUT4 mux_59_i6_4_lut (.A(wb_lo_data[5]), .B(wb_smpl_data[5]), .C(wb_smpl_ack), 
         .D(wb_lo_ack), .Z(wb_idata_31__N_266[5])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(273[8] 276[22])
    defparam mux_59_i6_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i5_3_lut (.A(wb_idata_31__N_266[4]), .B(wb_fm_data[4]), 
         .C(wb_fm_ack), .Z(wb_idata_31__N_1[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(271[8] 276[22])
    defparam wb_idata_31__I_0_i5_3_lut.init = 16'hcaca;
    LUT4 mux_59_i5_4_lut (.A(wb_lo_data[4]), .B(wb_smpl_data[4]), .C(wb_smpl_ack), 
         .D(wb_lo_ack), .Z(wb_idata_31__N_266[4])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(273[8] 276[22])
    defparam mux_59_i5_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i4_3_lut (.A(wb_idata_31__N_266[3]), .B(wb_fm_data[3]), 
         .C(wb_fm_ack), .Z(wb_idata_31__N_1[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(271[8] 276[22])
    defparam wb_idata_31__I_0_i4_3_lut.init = 16'hcaca;
    LUT4 mux_59_i4_4_lut (.A(wb_lo_data[3]), .B(wb_smpl_data[3]), .C(wb_smpl_ack), 
         .D(wb_lo_ack), .Z(wb_idata_31__N_266[3])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(273[8] 276[22])
    defparam mux_59_i4_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i3_3_lut (.A(wb_idata_31__N_266[2]), .B(wb_fm_data[2]), 
         .C(wb_fm_ack), .Z(wb_idata_31__N_1[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(271[8] 276[22])
    defparam wb_idata_31__I_0_i3_3_lut.init = 16'hcaca;
    LUT4 mux_59_i3_4_lut (.A(wb_lo_data[2]), .B(wb_smpl_data[2]), .C(wb_smpl_ack), 
         .D(wb_lo_ack), .Z(wb_idata_31__N_266[2])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(273[8] 276[22])
    defparam mux_59_i3_4_lut.init = 16'hcac0;
    LUT4 wb_idata_31__I_0_i2_3_lut (.A(wb_idata_31__N_266[1]), .B(wb_fm_data[1]), 
         .C(wb_fm_ack), .Z(wb_idata_31__N_1[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(271[8] 276[22])
    defparam wb_idata_31__I_0_i2_3_lut.init = 16'hcaca;
    LUT4 mux_59_i2_4_lut (.A(wb_lo_data[1]), .B(wb_smpl_data[1]), .C(wb_smpl_ack), 
         .D(wb_lo_ack), .Z(wb_idata_31__N_266[1])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(273[8] 276[22])
    defparam mux_59_i2_4_lut.init = 16'hcac0;
    LUT4 power_counter_31__I_0_77_i31_3_lut (.A(power_counter_31__N_232[30]), 
         .B(power_counter_31__N_201[30]), .C(power_counter[31]), .Z(power_counter_31__N_129[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(232[4:54])
    defparam power_counter_31__I_0_77_i31_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_77_i30_3_lut (.A(power_counter_31__N_232[29]), 
         .B(power_counter_31__N_201[29]), .C(power_counter[31]), .Z(power_counter_31__N_129[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(232[4:54])
    defparam power_counter_31__I_0_77_i30_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_77_i29_3_lut (.A(power_counter_31__N_232[28]), 
         .B(power_counter_31__N_201[28]), .C(power_counter[31]), .Z(power_counter_31__N_129[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(232[4:54])
    defparam power_counter_31__I_0_77_i29_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_77_i28_3_lut (.A(power_counter_31__N_232[27]), 
         .B(power_counter_31__N_201[27]), .C(power_counter[31]), .Z(power_counter_31__N_129[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(232[4:54])
    defparam power_counter_31__I_0_77_i28_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_77_i27_3_lut (.A(power_counter_31__N_232[26]), 
         .B(power_counter_31__N_201[26]), .C(power_counter[31]), .Z(power_counter_31__N_129[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(232[4:54])
    defparam power_counter_31__I_0_77_i27_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_77_i26_3_lut (.A(power_counter_31__N_232[25]), 
         .B(power_counter_31__N_201[25]), .C(power_counter[31]), .Z(power_counter_31__N_129[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(232[4:54])
    defparam power_counter_31__I_0_77_i26_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_77_i25_3_lut (.A(power_counter_31__N_232[24]), 
         .B(power_counter_31__N_201[24]), .C(power_counter[31]), .Z(power_counter_31__N_129[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(232[4:54])
    defparam power_counter_31__I_0_77_i25_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_77_i24_3_lut (.A(power_counter_31__N_232[23]), 
         .B(power_counter_31__N_201[23]), .C(power_counter[31]), .Z(power_counter_31__N_129[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(232[4:54])
    defparam power_counter_31__I_0_77_i24_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_77_i23_3_lut (.A(power_counter_31__N_232[22]), 
         .B(power_counter_31__N_201[22]), .C(power_counter[31]), .Z(power_counter_31__N_129[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(232[4:54])
    defparam power_counter_31__I_0_77_i23_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_77_i22_3_lut (.A(power_counter_31__N_232[21]), 
         .B(power_counter_31__N_201[21]), .C(power_counter[31]), .Z(power_counter_31__N_129[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(232[4:54])
    defparam power_counter_31__I_0_77_i22_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_77_i21_3_lut (.A(power_counter_31__N_232[20]), 
         .B(power_counter_31__N_201[20]), .C(power_counter[31]), .Z(power_counter_31__N_129[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(232[4:54])
    defparam power_counter_31__I_0_77_i21_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_77_i20_3_lut (.A(power_counter_31__N_232[19]), 
         .B(power_counter_31__N_201[19]), .C(power_counter[31]), .Z(power_counter_31__N_129[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(232[4:54])
    defparam power_counter_31__I_0_77_i20_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_77_i19_3_lut (.A(power_counter_31__N_232[18]), 
         .B(power_counter_31__N_201[18]), .C(power_counter[31]), .Z(power_counter_31__N_129[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(232[4:54])
    defparam power_counter_31__I_0_77_i19_3_lut.init = 16'hcaca;
    CCU2D add_35_29 (.A0(power_counter[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17568), .COUT(n17569), .S0(power_counter_31__N_201[27]), 
          .S1(power_counter_31__N_201[28]));   // d:/documents/git_local/fm_modulator/rtl/top.v(232[27:53])
    defparam add_35_29.INIT0 = 16'h5aaa;
    defparam add_35_29.INIT1 = 16'h5aaa;
    defparam add_35_29.INJECT1_0 = "NO";
    defparam add_35_29.INJECT1_1 = "NO";
    LUT4 power_counter_31__I_0_77_i18_3_lut (.A(power_counter_31__N_232[17]), 
         .B(power_counter_31__N_201[17]), .C(power_counter[31]), .Z(power_counter_31__N_129[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(232[4:54])
    defparam power_counter_31__I_0_77_i18_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_77_i17_3_lut (.A(power_counter_31__N_232[16]), 
         .B(power_counter_31__N_201[16]), .C(power_counter[31]), .Z(power_counter_31__N_129[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(232[4:54])
    defparam power_counter_31__I_0_77_i17_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_77_i16_3_lut (.A(power_counter_31__N_232[15]), 
         .B(power_counter_31__N_201[15]), .C(power_counter[31]), .Z(power_counter_31__N_129[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(232[4:54])
    defparam power_counter_31__I_0_77_i16_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_77_i15_3_lut (.A(power_counter_31__N_232[14]), 
         .B(power_counter_31__N_201[14]), .C(power_counter[31]), .Z(power_counter_31__N_129[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(232[4:54])
    defparam power_counter_31__I_0_77_i15_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_77_i14_3_lut (.A(power_counter_31__N_232[13]), 
         .B(power_counter_31__N_201[13]), .C(power_counter[31]), .Z(power_counter_31__N_129[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(232[4:54])
    defparam power_counter_31__I_0_77_i14_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_77_i13_3_lut (.A(power_counter_31__N_232[12]), 
         .B(power_counter_31__N_201[12]), .C(power_counter[31]), .Z(power_counter_31__N_129[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(232[4:54])
    defparam power_counter_31__I_0_77_i13_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_77_i12_3_lut (.A(power_counter_31__N_232[11]), 
         .B(power_counter_31__N_201[11]), .C(power_counter[31]), .Z(power_counter_31__N_129[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(232[4:54])
    defparam power_counter_31__I_0_77_i12_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_77_i11_3_lut (.A(power_counter_31__N_232[10]), 
         .B(power_counter_31__N_201[10]), .C(power_counter[31]), .Z(power_counter_31__N_129[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(232[4:54])
    defparam power_counter_31__I_0_77_i11_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_77_i10_3_lut (.A(power_counter_31__N_232[9]), 
         .B(power_counter_31__N_201[9]), .C(power_counter[31]), .Z(power_counter_31__N_129[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(232[4:54])
    defparam power_counter_31__I_0_77_i10_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_77_i9_3_lut (.A(power_counter_31__N_232[8]), 
         .B(power_counter_31__N_201[8]), .C(power_counter[31]), .Z(power_counter_31__N_129[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(232[4:54])
    defparam power_counter_31__I_0_77_i9_3_lut.init = 16'hcaca;
    LUT4 mux_393_Mux_11_i2_3_lut (.A(bus_err_address[9]), .B(power_counter[11]), 
         .C(wb_addr[0]), .Z(n2_adj_3067)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(216[3] 223[10])
    defparam mux_393_Mux_11_i2_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_77_i8_3_lut (.A(power_counter_31__N_232[7]), 
         .B(power_counter_31__N_201[7]), .C(power_counter[31]), .Z(power_counter_31__N_129[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(232[4:54])
    defparam power_counter_31__I_0_77_i8_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_77_i7_3_lut (.A(power_counter_31__N_232[6]), 
         .B(power_counter_31__N_201[6]), .C(power_counter[31]), .Z(power_counter_31__N_129[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(232[4:54])
    defparam power_counter_31__I_0_77_i7_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_77_i6_3_lut (.A(power_counter_31__N_232[5]), 
         .B(power_counter_31__N_201[5]), .C(power_counter[31]), .Z(power_counter_31__N_129[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(232[4:54])
    defparam power_counter_31__I_0_77_i6_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_77_i5_3_lut (.A(power_counter_31__N_232[4]), 
         .B(power_counter_31__N_201[4]), .C(power_counter[31]), .Z(power_counter_31__N_129[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(232[4:54])
    defparam power_counter_31__I_0_77_i5_3_lut.init = 16'hcaca;
    LUT4 i11122_2_lut (.A(smpl_register[11]), .B(wb_addr[0]), .Z(n1_adj_3068)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(216[3] 223[10])
    defparam i11122_2_lut.init = 16'h8888;
    LUT4 power_counter_31__I_0_77_i4_3_lut (.A(power_counter_31__N_232[3]), 
         .B(power_counter_31__N_201[3]), .C(power_counter[31]), .Z(power_counter_31__N_129[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(232[4:54])
    defparam power_counter_31__I_0_77_i4_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_77_i3_3_lut (.A(power_counter_31__N_232[2]), 
         .B(power_counter_31__N_201[2]), .C(power_counter[31]), .Z(power_counter_31__N_129[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(232[4:54])
    defparam power_counter_31__I_0_77_i3_3_lut.init = 16'hcaca;
    LUT4 power_counter_31__I_0_77_i2_3_lut (.A(power_counter_31__N_232[1]), 
         .B(power_counter_31__N_201[1]), .C(power_counter[31]), .Z(power_counter_31__N_129[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(232[4:54])
    defparam power_counter_31__I_0_77_i2_3_lut.init = 16'hcaca;
    LUT4 i847_1_lut (.A(o_baseband_q_c_15), .Z(o_baseband_q_c_9)) /* synthesis lut_function=(!(A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(114[31:66])
    defparam i847_1_lut.init = 16'h5555;
    LUT4 dac_clk_p_I_0_1_lut (.A(dac_clk_p_c), .Z(dac_clk_n_c)) /* synthesis lut_function=(!(A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(46[20:30])
    defparam dac_clk_p_I_0_1_lut.init = 16'h5555;
    LUT4 mux_393_Mux_10_i2_3_lut (.A(bus_err_address[8]), .B(power_counter[10]), 
         .C(wb_addr[0]), .Z(n2_adj_3069)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(216[3] 223[10])
    defparam mux_393_Mux_10_i2_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_574 (.A(wb_addr[12]), .B(wb_addr[8]), .Z(n26897)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[23:49])
    defparam i1_2_lut_rep_574.init = 16'heeee;
    PFUMX mux_393_Mux_15_i3 (.BLUT(n1_adj_3060), .ALUT(n2_adj_3059), .C0(wb_addr[1]), 
          .Z(n2147));
    LUT4 mux_393_Mux_2_i2_3_lut (.A(bus_err_address[0]), .B(power_counter[2]), 
         .C(wb_addr[0]), .Z(n2_adj_3082)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(216[3] 223[10])
    defparam mux_393_Mux_2_i2_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_rep_461_3_lut (.A(wb_addr[12]), .B(wb_addr[8]), .C(wb_addr[1]), 
         .Z(n26784)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[23:49])
    defparam i1_2_lut_rep_461_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_3_lut (.A(wb_addr[12]), .B(wb_addr[8]), .C(wb_addr[0]), 
         .Z(n20745)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[23:49])
    defparam i1_2_lut_3_lut.init = 16'hfefe;
    LUT4 i1_4_lut_adj_155 (.A(n26784), .B(n20733), .C(n34), .D(wb_addr[0]), 
         .Z(n20739)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[23:49])
    defparam i1_4_lut_adj_155.init = 16'hfffe;
    CCU2D add_34_21 (.A0(power_counter[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17548), .COUT(n17549), .S0(power_counter_31__N_232[19]), 
          .S1(power_counter_31__N_232[20]));   // d:/documents/git_local/fm_modulator/rtl/top.v(230[21:41])
    defparam add_34_21.INIT0 = 16'h5aaa;
    defparam add_34_21.INIT1 = 16'h5aaa;
    defparam add_34_21.INJECT1_0 = "NO";
    defparam add_34_21.INJECT1_1 = "NO";
    LUT4 mux_393_Mux_9_i2_3_lut (.A(bus_err_address[7]), .B(power_counter[9]), 
         .C(wb_addr[0]), .Z(n2_adj_3070)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(216[3] 223[10])
    defparam mux_393_Mux_9_i2_3_lut.init = 16'hcaca;
    LUT4 mux_393_Mux_8_i2_3_lut (.A(bus_err_address[6]), .B(power_counter[8]), 
         .C(wb_addr[0]), .Z(n2_adj_3071)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(216[3] 223[10])
    defparam mux_393_Mux_8_i2_3_lut.init = 16'hcaca;
    LUT4 i11119_2_lut (.A(smpl_register[8]), .B(wb_addr[0]), .Z(n1_adj_3072)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(216[3] 223[10])
    defparam i11119_2_lut.init = 16'h8888;
    LUT4 mux_393_Mux_7_i2_3_lut (.A(bus_err_address[5]), .B(power_counter[7]), 
         .C(wb_addr[0]), .Z(n2_adj_3073)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(216[3] 223[10])
    defparam mux_393_Mux_7_i2_3_lut.init = 16'hcaca;
    LUT4 i11118_2_lut (.A(smpl_register[7]), .B(wb_addr[0]), .Z(n1_adj_3074)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(216[3] 223[10])
    defparam i11118_2_lut.init = 16'h8888;
    LUT4 mux_393_Mux_24_i2_3_lut (.A(bus_err_address[22]), .B(power_counter[24]), 
         .C(wb_addr[0]), .Z(n2_adj_3045)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(216[3] 223[10])
    defparam mux_393_Mux_24_i2_3_lut.init = 16'hcaca;
    LUT4 o_clk_q_I_0_1_lut (.A(q_clk_p_c), .Z(q_clk_n_c)) /* synthesis lut_function=(!(A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/clock_phase_shifter.v(18[16:24])
    defparam o_clk_q_I_0_1_lut.init = 16'h5555;
    LUT4 mux_393_Mux_6_i2_3_lut (.A(bus_err_address[4]), .B(power_counter[6]), 
         .C(wb_addr[0]), .Z(n2_adj_3075)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(216[3] 223[10])
    defparam mux_393_Mux_6_i2_3_lut.init = 16'hcaca;
    LUT4 i11117_2_lut (.A(smpl_register[6]), .B(wb_addr[0]), .Z(n1_adj_3076)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(216[3] 223[10])
    defparam i11117_2_lut.init = 16'h8888;
    LUT4 mux_393_Mux_5_i2_3_lut (.A(bus_err_address[3]), .B(power_counter[5]), 
         .C(wb_addr[0]), .Z(n2_adj_3077)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(216[3] 223[10])
    defparam mux_393_Mux_5_i2_3_lut.init = 16'hcaca;
    LUT4 mux_393_Mux_4_i2_3_lut (.A(bus_err_address[2]), .B(power_counter[4]), 
         .C(wb_addr[0]), .Z(n2_adj_3078)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(216[3] 223[10])
    defparam mux_393_Mux_4_i2_3_lut.init = 16'hcaca;
    LUT4 i11115_2_lut (.A(smpl_register[4]), .B(wb_addr[0]), .Z(n1_adj_3079)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(216[3] 223[10])
    defparam i11115_2_lut.init = 16'h8888;
    LUT4 i6_2_lut_rep_623 (.A(wb_addr[22]), .B(wb_addr[24]), .Z(n26946)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[23:49])
    defparam i6_2_lut_rep_623.init = 16'heeee;
    LUT4 i1_2_lut_rep_482_3_lut (.A(wb_addr[22]), .B(wb_addr[24]), .C(wb_addr[12]), 
         .Z(n26805)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[23:49])
    defparam i1_2_lut_rep_482_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_rep_439_3_lut_4_lut (.A(wb_addr[22]), .B(wb_addr[24]), 
         .C(n38), .D(wb_addr[12]), .Z(n26762)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[23:49])
    defparam i1_2_lut_rep_439_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_3_lut_adj_156 (.A(wb_addr[22]), .B(wb_addr[24]), .C(wb_addr[9]), 
         .Z(n20733)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[23:49])
    defparam i1_2_lut_3_lut_adj_156.init = 16'hefef;
    LUT4 i1_2_lut_rep_624 (.A(wb_stb), .B(wb_we), .Z(n26947)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(126[39:58])
    defparam i1_2_lut_rep_624.init = 16'h8888;
    LUT4 i18823_2_lut_3_lut (.A(wb_stb), .B(wb_we), .C(wb_addr[0]), .Z(n21184)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(126[39:58])
    defparam i18823_2_lut_3_lut.init = 16'h8080;
    LUT4 i11135_2_lut (.A(smpl_register[24]), .B(wb_addr[0]), .Z(n1_adj_3046)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(216[3] 223[10])
    defparam i11135_2_lut.init = 16'h8888;
    LUT4 o_clk_i_I_0_1_lut (.A(i_clk_p_c), .Z(i_clk_n_c)) /* synthesis lut_function=(!(A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/clock_phase_shifter.v(14[16:24])
    defparam o_clk_i_I_0_1_lut.init = 16'h5555;
    PFUMX mux_393_Mux_19_i3 (.BLUT(n1_adj_3055), .ALUT(n2_adj_3054), .C0(wb_addr[1]), 
          .Z(n2143));
    LUT4 mux_393_Mux_3_i2_3_lut (.A(bus_err_address[1]), .B(power_counter[3]), 
         .C(wb_addr[0]), .Z(n2_adj_3080)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(216[3] 223[10])
    defparam mux_393_Mux_3_i2_3_lut.init = 16'hcaca;
    VLO i1 (.Z(GND_net));
    PFUMX mux_393_Mux_21_i3 (.BLUT(n1_adj_3052), .ALUT(n2_adj_3051), .C0(wb_addr[1]), 
          .Z(n2141));
    LUT4 i1_4_lut_adj_157 (.A(n26946), .B(n20749), .C(wb_addr[15]), .D(n20745), 
         .Z(n20755)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(244[23:49])
    defparam i1_4_lut_adj_157.init = 16'hffef;
    PFUMX mux_393_Mux_22_i3 (.BLUT(n1_adj_3050), .ALUT(n2_adj_3049), .C0(wb_addr[1]), 
          .Z(n2140));
    LUT4 i11114_2_lut (.A(smpl_register[3]), .B(wb_addr[0]), .Z(n1_adj_3081)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(216[3] 223[10])
    defparam i11114_2_lut.init = 16'h8888;
    LUT4 mux_393_Mux_23_i2_3_lut (.A(bus_err_address[21]), .B(power_counter[23]), 
         .C(wb_addr[0]), .Z(n2_adj_3047)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(216[3] 223[10])
    defparam mux_393_Mux_23_i2_3_lut.init = 16'hcaca;
    TSALL TSALL_INST (.TSALL(GND_net));
    LUT4 i11134_2_lut (.A(smpl_register[23]), .B(wb_addr[0]), .Z(n1_adj_3048)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(216[3] 223[10])
    defparam i11134_2_lut.init = 16'h8888;
    FD1S3AX wb_idata_i30 (.D(wb_idata_31__N_1[30]), .CK(dac_clk_p_c), .Q(wb_idata[30]));   // d:/documents/git_local/fm_modulator/rtl/top.v(268[9] 276[22])
    defparam wb_idata_i30.GSR = "DISABLED";
    FD1S3AX wb_idata_i29 (.D(wb_idata_31__N_1[29]), .CK(dac_clk_p_c), .Q(wb_idata[29]));   // d:/documents/git_local/fm_modulator/rtl/top.v(268[9] 276[22])
    defparam wb_idata_i29.GSR = "DISABLED";
    FD1S3AX wb_idata_i28 (.D(wb_idata_31__N_1[28]), .CK(dac_clk_p_c), .Q(wb_idata[28]));   // d:/documents/git_local/fm_modulator/rtl/top.v(268[9] 276[22])
    defparam wb_idata_i28.GSR = "DISABLED";
    FD1S3AX wb_idata_i27 (.D(wb_idata_31__N_1[27]), .CK(dac_clk_p_c), .Q(wb_idata[27]));   // d:/documents/git_local/fm_modulator/rtl/top.v(268[9] 276[22])
    defparam wb_idata_i27.GSR = "DISABLED";
    FD1S3AX wb_idata_i26 (.D(wb_idata_31__N_1[26]), .CK(dac_clk_p_c), .Q(wb_idata[26]));   // d:/documents/git_local/fm_modulator/rtl/top.v(268[9] 276[22])
    defparam wb_idata_i26.GSR = "DISABLED";
    FD1S3AX wb_idata_i25 (.D(wb_idata_31__N_1[25]), .CK(dac_clk_p_c), .Q(wb_idata[25]));   // d:/documents/git_local/fm_modulator/rtl/top.v(268[9] 276[22])
    defparam wb_idata_i25.GSR = "DISABLED";
    FD1S3AX wb_idata_i24 (.D(wb_idata_31__N_1[24]), .CK(dac_clk_p_c), .Q(wb_idata[24]));   // d:/documents/git_local/fm_modulator/rtl/top.v(268[9] 276[22])
    defparam wb_idata_i24.GSR = "DISABLED";
    FD1S3AX wb_idata_i23 (.D(wb_idata_31__N_1[23]), .CK(dac_clk_p_c), .Q(wb_idata[23]));   // d:/documents/git_local/fm_modulator/rtl/top.v(268[9] 276[22])
    defparam wb_idata_i23.GSR = "DISABLED";
    FD1P3AX smpl_interrupt_65 (.D(wb_odata[0]), .SP(dac_clk_p_c_enable_403), 
            .CK(dac_clk_p_c), .Q(smpl_interrupt)) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(205[9] 213[6])
    defparam smpl_interrupt_65.GSR = "DISABLED";
    LUT4 i3_4_lut (.A(wb_addr[9]), .B(wb_addr[8]), .C(wb_cyc), .D(n20377), 
         .Z(wb_lo_data_7__N_96)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i3_4_lut.init = 16'h8000;
    FD1S3AX wb_idata_i22 (.D(wb_idata_31__N_1[22]), .CK(dac_clk_p_c), .Q(wb_idata[22]));   // d:/documents/git_local/fm_modulator/rtl/top.v(268[9] 276[22])
    defparam wb_idata_i22.GSR = "DISABLED";
    LUT4 i2_4_lut (.A(n34), .B(wb_addr[15]), .C(n38), .D(n26805), .Z(n20377)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i2_4_lut.init = 16'h0004;
    CCU2D add_35_27 (.A0(power_counter[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17567), .COUT(n17568), .S0(power_counter_31__N_201[25]), 
          .S1(power_counter_31__N_201[26]));   // d:/documents/git_local/fm_modulator/rtl/top.v(232[27:53])
    defparam add_35_27.INIT0 = 16'h5aaa;
    defparam add_35_27.INIT1 = 16'h5aaa;
    defparam add_35_27.INJECT1_0 = "NO";
    defparam add_35_27.INJECT1_1 = "NO";
    LUT4 mux_393_Mux_22_i2_3_lut (.A(bus_err_address[20]), .B(power_counter[22]), 
         .C(wb_addr[0]), .Z(n2_adj_3049)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(216[3] 223[10])
    defparam mux_393_Mux_22_i2_3_lut.init = 16'hcaca;
    FD1S3AX wb_idata_i21 (.D(wb_idata_31__N_1[21]), .CK(dac_clk_p_c), .Q(wb_idata[21]));   // d:/documents/git_local/fm_modulator/rtl/top.v(268[9] 276[22])
    defparam wb_idata_i21.GSR = "DISABLED";
    efb_inst wb_lo_data_7__I_0 (.dac_clk_p_c(dac_clk_p_c), .i_resetb_N_301(i_resetb_N_301), 
            .wb_cyc(wb_cyc), .wb_lo_data_7__N_96(wb_lo_data_7__N_96), .wb_we(wb_we), 
            .\wb_addr[7] (wb_addr[7]), .\wb_addr[6] (wb_addr[6]), .\wb_addr[5] (wb_addr[5]), 
            .\wb_addr[4] (wb_addr[4]), .\wb_addr[3] (wb_addr[3]), .\wb_addr[2] (wb_addr[2]), 
            .\wb_addr[1] (wb_addr[1]), .\wb_addr[0] (wb_addr[0]), .\wb_odata[7] (wb_odata[7]), 
            .\wb_odata[6] (wb_odata[6]), .\wb_odata[5] (wb_odata[5]), .\wb_odata[4] (wb_odata[4]), 
            .\wb_odata[3] (wb_odata[3]), .\wb_odata[2] (wb_odata[2]), .\wb_odata[1] (wb_odata[1]), 
            .\wb_odata[0] (wb_odata[0]), .pll_data_o({pll_data_o}), .pll_ack(pll_ack), 
            .wb_lo_data({wb_lo_data}), .wb_lo_ack(wb_lo_ack), .pll_clk(pll_clk), 
            .pll_rst(pll_rst), .pll_stb(pll_stb), .pll_we(pll_we), .pll_addr({pll_addr}), 
            .pll_data_i({pll_data_i}), .GND_net(GND_net), .VCC_net(VCC_net)) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(180[10] 192[3])
    clock_phase_shifter clock_phase_shifter_inst (.q_clk_p_c(q_clk_p_c), .i_clk_2f_N_2249(i_clk_2f_N_2249), 
            .q_clk_n_c(q_clk_n_c), .i_clk_p_c(i_clk_p_c), .lo_pll_out(lo_pll_out), 
            .i_clk_n_c(i_clk_n_c)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(161[21] 165[2])
    FD1S3AX wb_idata_i20 (.D(wb_idata_31__N_1[20]), .CK(dac_clk_p_c), .Q(wb_idata[20]));   // d:/documents/git_local/fm_modulator/rtl/top.v(268[9] 276[22])
    defparam wb_idata_i20.GSR = "DISABLED";
    sys_clk sys_clk_inst (.i_ref_clk_c(i_ref_clk_c), .dac_clk_p_c(dac_clk_p_c), 
            .GND_net(GND_net)) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(37[10:54])
    CCU2D add_35_25 (.A0(power_counter[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17566), .COUT(n17567), .S0(power_counter_31__N_201[23]), 
          .S1(power_counter_31__N_201[24]));   // d:/documents/git_local/fm_modulator/rtl/top.v(232[27:53])
    defparam add_35_25.INIT0 = 16'h5aaa;
    defparam add_35_25.INIT1 = 16'h5aaa;
    defparam add_35_25.INJECT1_0 = "NO";
    defparam add_35_25.INJECT1_1 = "NO";
    CCU2D add_34_19 (.A0(power_counter[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17547), .COUT(n17548), .S0(power_counter_31__N_232[17]), 
          .S1(power_counter_31__N_232[18]));   // d:/documents/git_local/fm_modulator/rtl/top.v(230[21:41])
    defparam add_34_19.INIT0 = 16'h5aaa;
    defparam add_34_19.INIT1 = 16'h5aaa;
    defparam add_34_19.INJECT1_0 = "NO";
    defparam add_34_19.INJECT1_1 = "NO";
    CCU2D add_35_23 (.A0(power_counter[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17565), .COUT(n17566), .S0(power_counter_31__N_201[21]), 
          .S1(power_counter_31__N_201[22]));   // d:/documents/git_local/fm_modulator/rtl/top.v(232[27:53])
    defparam add_35_23.INIT0 = 16'h5aaa;
    defparam add_35_23.INIT1 = 16'h5aaa;
    defparam add_35_23.INJECT1_0 = "NO";
    defparam add_35_23.INJECT1_1 = "NO";
    CCU2D add_34_17 (.A0(power_counter[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17546), .COUT(n17547), .S0(power_counter_31__N_232[15]), 
          .S1(power_counter_31__N_232[16]));   // d:/documents/git_local/fm_modulator/rtl/top.v(230[21:41])
    defparam add_34_17.INIT0 = 16'h5aaa;
    defparam add_34_17.INIT1 = 16'h5aaa;
    defparam add_34_17.INJECT1_0 = "NO";
    defparam add_34_17.INJECT1_1 = "NO";
    CCU2D add_35_21 (.A0(power_counter[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17564), .COUT(n17565), .S0(power_counter_31__N_201[19]), 
          .S1(power_counter_31__N_201[20]));   // d:/documents/git_local/fm_modulator/rtl/top.v(232[27:53])
    defparam add_35_21.INIT0 = 16'h5aaa;
    defparam add_35_21.INIT1 = 16'h5aaa;
    defparam add_35_21.INJECT1_0 = "NO";
    defparam add_35_21.INJECT1_1 = "NO";
    OB o_baseband_i_pad_6 (.I(o_baseband_i_c_13), .O(o_baseband_i[6]));   // d:/documents/git_local/fm_modulator/rtl/top.v(27[38:50])
    FD1S3AX wb_idata_i19 (.D(wb_idata_31__N_1[19]), .CK(dac_clk_p_c), .Q(wb_idata[19]));   // d:/documents/git_local/fm_modulator/rtl/top.v(268[9] 276[22])
    defparam wb_idata_i19.GSR = "DISABLED";
    FD1S3AX wb_idata_i18 (.D(wb_idata_31__N_1[18]), .CK(dac_clk_p_c), .Q(wb_idata[18]));   // d:/documents/git_local/fm_modulator/rtl/top.v(268[9] 276[22])
    defparam wb_idata_i18.GSR = "DISABLED";
    FD1S3AX wb_idata_i17 (.D(wb_idata_31__N_1[17]), .CK(dac_clk_p_c), .Q(wb_idata[17]));   // d:/documents/git_local/fm_modulator/rtl/top.v(268[9] 276[22])
    defparam wb_idata_i17.GSR = "DISABLED";
    FD1S3AX wb_idata_i16 (.D(wb_idata_31__N_1[16]), .CK(dac_clk_p_c), .Q(wb_idata[16]));   // d:/documents/git_local/fm_modulator/rtl/top.v(268[9] 276[22])
    defparam wb_idata_i16.GSR = "DISABLED";
    FD1S3AX wb_idata_i15 (.D(wb_idata_31__N_1[15]), .CK(dac_clk_p_c), .Q(wb_idata[15]));   // d:/documents/git_local/fm_modulator/rtl/top.v(268[9] 276[22])
    defparam wb_idata_i15.GSR = "DISABLED";
    FD1S3AX wb_idata_i14 (.D(wb_idata_31__N_1[14]), .CK(dac_clk_p_c), .Q(wb_idata[14]));   // d:/documents/git_local/fm_modulator/rtl/top.v(268[9] 276[22])
    defparam wb_idata_i14.GSR = "DISABLED";
    FD1S3AX wb_idata_i13 (.D(wb_idata_31__N_1[13]), .CK(dac_clk_p_c), .Q(wb_idata[13]));   // d:/documents/git_local/fm_modulator/rtl/top.v(268[9] 276[22])
    defparam wb_idata_i13.GSR = "DISABLED";
    FD1S3AX wb_idata_i12 (.D(wb_idata_31__N_1[12]), .CK(dac_clk_p_c), .Q(wb_idata[12]));   // d:/documents/git_local/fm_modulator/rtl/top.v(268[9] 276[22])
    defparam wb_idata_i12.GSR = "DISABLED";
    FD1S3AX wb_idata_i11 (.D(wb_idata_31__N_1[11]), .CK(dac_clk_p_c), .Q(wb_idata[11]));   // d:/documents/git_local/fm_modulator/rtl/top.v(268[9] 276[22])
    defparam wb_idata_i11.GSR = "DISABLED";
    FD1S3AX wb_idata_i10 (.D(wb_idata_31__N_1[10]), .CK(dac_clk_p_c), .Q(wb_idata[10]));   // d:/documents/git_local/fm_modulator/rtl/top.v(268[9] 276[22])
    defparam wb_idata_i10.GSR = "DISABLED";
    FD1S3AX wb_idata_i9 (.D(wb_idata_31__N_1[9]), .CK(dac_clk_p_c), .Q(wb_idata[9]));   // d:/documents/git_local/fm_modulator/rtl/top.v(268[9] 276[22])
    defparam wb_idata_i9.GSR = "DISABLED";
    FD1S3AX wb_idata_i8 (.D(wb_idata_31__N_1[8]), .CK(dac_clk_p_c), .Q(wb_idata[8]));   // d:/documents/git_local/fm_modulator/rtl/top.v(268[9] 276[22])
    defparam wb_idata_i8.GSR = "DISABLED";
    FD1S3AX wb_idata_i7 (.D(wb_idata_31__N_1[7]), .CK(dac_clk_p_c), .Q(wb_idata[7]));   // d:/documents/git_local/fm_modulator/rtl/top.v(268[9] 276[22])
    defparam wb_idata_i7.GSR = "DISABLED";
    FD1S3AX wb_idata_i6 (.D(wb_idata_31__N_1[6]), .CK(dac_clk_p_c), .Q(wb_idata[6]));   // d:/documents/git_local/fm_modulator/rtl/top.v(268[9] 276[22])
    defparam wb_idata_i6.GSR = "DISABLED";
    FD1S3AX wb_idata_i5 (.D(wb_idata_31__N_1[5]), .CK(dac_clk_p_c), .Q(wb_idata[5]));   // d:/documents/git_local/fm_modulator/rtl/top.v(268[9] 276[22])
    defparam wb_idata_i5.GSR = "DISABLED";
    FD1S3AX wb_idata_i4 (.D(wb_idata_31__N_1[4]), .CK(dac_clk_p_c), .Q(wb_idata[4]));   // d:/documents/git_local/fm_modulator/rtl/top.v(268[9] 276[22])
    defparam wb_idata_i4.GSR = "DISABLED";
    FD1S3AX wb_idata_i3 (.D(wb_idata_31__N_1[3]), .CK(dac_clk_p_c), .Q(wb_idata[3]));   // d:/documents/git_local/fm_modulator/rtl/top.v(268[9] 276[22])
    defparam wb_idata_i3.GSR = "DISABLED";
    FD1S3AX wb_idata_i2 (.D(wb_idata_31__N_1[2]), .CK(dac_clk_p_c), .Q(wb_idata[2]));   // d:/documents/git_local/fm_modulator/rtl/top.v(268[9] 276[22])
    defparam wb_idata_i2.GSR = "DISABLED";
    FD1S3AX wb_idata_i1 (.D(wb_idata_31__N_1[1]), .CK(dac_clk_p_c), .Q(wb_idata[1]));   // d:/documents/git_local/fm_modulator/rtl/top.v(268[9] 276[22])
    defparam wb_idata_i1.GSR = "DISABLED";
    CCU2D add_34_15 (.A0(power_counter[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17545), .COUT(n17546), .S0(power_counter_31__N_232[13]), 
          .S1(power_counter_31__N_232[14]));   // d:/documents/git_local/fm_modulator/rtl/top.v(230[21:41])
    defparam add_34_15.INIT0 = 16'h5aaa;
    defparam add_34_15.INIT1 = 16'h5aaa;
    defparam add_34_15.INJECT1_0 = "NO";
    defparam add_34_15.INJECT1_1 = "NO";
    CCU2D add_35_19 (.A0(power_counter[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17563), .COUT(n17564), .S0(power_counter_31__N_201[17]), 
          .S1(power_counter_31__N_201[18]));   // d:/documents/git_local/fm_modulator/rtl/top.v(232[27:53])
    defparam add_35_19.INIT0 = 16'h5aaa;
    defparam add_35_19.INIT1 = 16'h5aaa;
    defparam add_35_19.INJECT1_0 = "NO";
    defparam add_35_19.INJECT1_1 = "NO";
    CCU2D add_34_5 (.A0(power_counter[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17540), .COUT(n17541), .S0(power_counter_31__N_232[3]), 
          .S1(power_counter_31__N_232[4]));   // d:/documents/git_local/fm_modulator/rtl/top.v(230[21:41])
    defparam add_34_5.INIT0 = 16'h5aaa;
    defparam add_34_5.INIT1 = 16'h5aaa;
    defparam add_34_5.INJECT1_0 = "NO";
    defparam add_34_5.INJECT1_1 = "NO";
    CCU2D add_35_17 (.A0(power_counter[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17562), .COUT(n17563), .S0(power_counter_31__N_201[15]), 
          .S1(power_counter_31__N_201[16]));   // d:/documents/git_local/fm_modulator/rtl/top.v(232[27:53])
    defparam add_35_17.INIT0 = 16'h5aaa;
    defparam add_35_17.INIT1 = 16'h5aaa;
    defparam add_35_17.INJECT1_0 = "NO";
    defparam add_35_17.INJECT1_1 = "NO";
    CCU2D add_35_15 (.A0(power_counter[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17561), .COUT(n17562), .S0(power_counter_31__N_201[13]), 
          .S1(power_counter_31__N_201[14]));   // d:/documents/git_local/fm_modulator/rtl/top.v(232[27:53])
    defparam add_35_15.INIT0 = 16'h5aaa;
    defparam add_35_15.INIT1 = 16'h5aaa;
    defparam add_35_15.INJECT1_0 = "NO";
    defparam add_35_15.INJECT1_1 = "NO";
    CCU2D add_35_13 (.A0(power_counter[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17560), .COUT(n17561), .S0(power_counter_31__N_201[11]), 
          .S1(power_counter_31__N_201[12]));   // d:/documents/git_local/fm_modulator/rtl/top.v(232[27:53])
    defparam add_35_13.INIT0 = 16'h5aaa;
    defparam add_35_13.INIT1 = 16'h5aaa;
    defparam add_35_13.INJECT1_0 = "NO";
    defparam add_35_13.INJECT1_1 = "NO";
    CCU2D add_35_11 (.A0(power_counter[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17559), .COUT(n17560), .S0(power_counter_31__N_201[9]), 
          .S1(power_counter_31__N_201[10]));   // d:/documents/git_local/fm_modulator/rtl/top.v(232[27:53])
    defparam add_35_11.INIT0 = 16'h5aaa;
    defparam add_35_11.INIT1 = 16'h5aaa;
    defparam add_35_11.INJECT1_0 = "NO";
    defparam add_35_11.INJECT1_1 = "NO";
    CCU2D add_34_9 (.A0(power_counter[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17542), .COUT(n17543), .S0(power_counter_31__N_232[7]), 
          .S1(power_counter_31__N_232[8]));   // d:/documents/git_local/fm_modulator/rtl/top.v(230[21:41])
    defparam add_34_9.INIT0 = 16'h5aaa;
    defparam add_34_9.INIT1 = 16'h5aaa;
    defparam add_34_9.INJECT1_0 = "NO";
    defparam add_34_9.INJECT1_1 = "NO";
    CCU2D add_35_9 (.A0(power_counter[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17558), .COUT(n17559), .S0(power_counter_31__N_201[7]), 
          .S1(power_counter_31__N_201[8]));   // d:/documents/git_local/fm_modulator/rtl/top.v(232[27:53])
    defparam add_35_9.INIT0 = 16'h5aaa;
    defparam add_35_9.INIT1 = 16'h5aaa;
    defparam add_35_9.INJECT1_0 = "NO";
    defparam add_35_9.INJECT1_1 = "NO";
    CCU2D add_35_7 (.A0(power_counter[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17557), .COUT(n17558), .S0(power_counter_31__N_201[5]), 
          .S1(power_counter_31__N_201[6]));   // d:/documents/git_local/fm_modulator/rtl/top.v(232[27:53])
    defparam add_35_7.INIT0 = 16'h5aaa;
    defparam add_35_7.INIT1 = 16'h5aaa;
    defparam add_35_7.INJECT1_0 = "NO";
    defparam add_35_7.INJECT1_1 = "NO";
    CCU2D add_34_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(power_counter[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n17539), .S1(power_counter_31__N_232[0]));   // d:/documents/git_local/fm_modulator/rtl/top.v(230[21:41])
    defparam add_34_1.INIT0 = 16'hF000;
    defparam add_34_1.INIT1 = 16'h5555;
    defparam add_34_1.INJECT1_0 = "NO";
    defparam add_34_1.INJECT1_1 = "NO";
    CCU2D add_35_5 (.A0(power_counter[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17556), .COUT(n17557), .S0(power_counter_31__N_201[3]), 
          .S1(power_counter_31__N_201[4]));   // d:/documents/git_local/fm_modulator/rtl/top.v(232[27:53])
    defparam add_35_5.INIT0 = 16'h5aaa;
    defparam add_35_5.INIT1 = 16'h5aaa;
    defparam add_35_5.INJECT1_0 = "NO";
    defparam add_35_5.INJECT1_1 = "NO";
    CCU2D add_35_3 (.A0(power_counter[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17555), .COUT(n17556), .S0(power_counter_31__N_201[1]), 
          .S1(power_counter_31__N_201[2]));   // d:/documents/git_local/fm_modulator/rtl/top.v(232[27:53])
    defparam add_35_3.INIT0 = 16'h5aaa;
    defparam add_35_3.INIT1 = 16'h5aaa;
    defparam add_35_3.INJECT1_0 = "NO";
    defparam add_35_3.INJECT1_1 = "NO";
    CCU2D add_34_3 (.A0(power_counter[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17539), .COUT(n17540), .S0(power_counter_31__N_232[1]), 
          .S1(power_counter_31__N_232[2]));   // d:/documents/git_local/fm_modulator/rtl/top.v(230[21:41])
    defparam add_34_3.INIT0 = 16'h5aaa;
    defparam add_34_3.INIT1 = 16'h5aaa;
    defparam add_34_3.INJECT1_0 = "NO";
    defparam add_34_3.INJECT1_1 = "NO";
    CCU2D add_35_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(power_counter[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n17555), .S1(power_counter_31__N_201[0]));   // d:/documents/git_local/fm_modulator/rtl/top.v(232[27:53])
    defparam add_35_1.INIT0 = 16'hF000;
    defparam add_35_1.INIT1 = 16'h5555;
    defparam add_35_1.INJECT1_0 = "NO";
    defparam add_35_1.INJECT1_1 = "NO";
    CCU2D add_34_13 (.A0(power_counter[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17544), .COUT(n17545), .S0(power_counter_31__N_232[11]), 
          .S1(power_counter_31__N_232[12]));   // d:/documents/git_local/fm_modulator/rtl/top.v(230[21:41])
    defparam add_34_13.INIT0 = 16'h5aaa;
    defparam add_34_13.INIT1 = 16'h5aaa;
    defparam add_34_13.INJECT1_0 = "NO";
    defparam add_34_13.INJECT1_1 = "NO";
    CCU2D add_34_33 (.A0(power_counter[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n17554), .S0(power_counter_31__N_232[31]));   // d:/documents/git_local/fm_modulator/rtl/top.v(230[21:41])
    defparam add_34_33.INIT0 = 16'h5aaa;
    defparam add_34_33.INIT1 = 16'h0000;
    defparam add_34_33.INJECT1_0 = "NO";
    defparam add_34_33.INJECT1_1 = "NO";
    CCU2D add_34_7 (.A0(power_counter[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17541), .COUT(n17542), .S0(power_counter_31__N_232[5]), 
          .S1(power_counter_31__N_232[6]));   // d:/documents/git_local/fm_modulator/rtl/top.v(230[21:41])
    defparam add_34_7.INIT0 = 16'h5aaa;
    defparam add_34_7.INIT1 = 16'h5aaa;
    defparam add_34_7.INJECT1_0 = "NO";
    defparam add_34_7.INJECT1_1 = "NO";
    CCU2D add_34_31 (.A0(power_counter[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17553), .COUT(n17554), .S0(power_counter_31__N_232[29]), 
          .S1(power_counter_31__N_232[30]));   // d:/documents/git_local/fm_modulator/rtl/top.v(230[21:41])
    defparam add_34_31.INIT0 = 16'h5aaa;
    defparam add_34_31.INIT1 = 16'h5aaa;
    defparam add_34_31.INJECT1_0 = "NO";
    defparam add_34_31.INJECT1_1 = "NO";
    FD1P3AX power_counter_i31 (.D(n29502), .SP(power_counter_31__N_232[31]), 
            .CK(dac_clk_p_c), .Q(power_counter[31])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 232[54])
    defparam power_counter_i31.GSR = "DISABLED";
    FD1S3AX power_counter_i30 (.D(power_counter_31__N_129[30]), .CK(dac_clk_p_c), 
            .Q(power_counter[30])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 232[54])
    defparam power_counter_i30.GSR = "DISABLED";
    FD1S3AX power_counter_i29 (.D(power_counter_31__N_129[29]), .CK(dac_clk_p_c), 
            .Q(power_counter[29])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 232[54])
    defparam power_counter_i29.GSR = "DISABLED";
    FD1S3AX power_counter_i28 (.D(power_counter_31__N_129[28]), .CK(dac_clk_p_c), 
            .Q(power_counter[28])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 232[54])
    defparam power_counter_i28.GSR = "DISABLED";
    FD1S3AX power_counter_i27 (.D(power_counter_31__N_129[27]), .CK(dac_clk_p_c), 
            .Q(power_counter[27])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 232[54])
    defparam power_counter_i27.GSR = "DISABLED";
    FD1S3AX power_counter_i26 (.D(power_counter_31__N_129[26]), .CK(dac_clk_p_c), 
            .Q(power_counter[26])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 232[54])
    defparam power_counter_i26.GSR = "DISABLED";
    FD1S3AX power_counter_i25 (.D(power_counter_31__N_129[25]), .CK(dac_clk_p_c), 
            .Q(power_counter[25])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 232[54])
    defparam power_counter_i25.GSR = "DISABLED";
    FD1S3AX power_counter_i24 (.D(power_counter_31__N_129[24]), .CK(dac_clk_p_c), 
            .Q(power_counter[24])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 232[54])
    defparam power_counter_i24.GSR = "DISABLED";
    FD1S3AX power_counter_i23 (.D(power_counter_31__N_129[23]), .CK(dac_clk_p_c), 
            .Q(power_counter[23])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 232[54])
    defparam power_counter_i23.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i29 (.D(wb_addr[29]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[29])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(258[9] 260[31])
    defparam bus_err_address_i0_i29.GSR = "DISABLED";
    CCU2D add_34_11 (.A0(power_counter[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17543), .COUT(n17544), .S0(power_counter_31__N_232[9]), 
          .S1(power_counter_31__N_232[10]));   // d:/documents/git_local/fm_modulator/rtl/top.v(230[21:41])
    defparam add_34_11.INIT0 = 16'h5aaa;
    defparam add_34_11.INIT1 = 16'h5aaa;
    defparam add_34_11.INJECT1_0 = "NO";
    defparam add_34_11.INJECT1_1 = "NO";
    CCU2D add_34_29 (.A0(power_counter[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(power_counter[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17552), .COUT(n17553), .S0(power_counter_31__N_232[27]), 
          .S1(power_counter_31__N_232[28]));   // d:/documents/git_local/fm_modulator/rtl/top.v(230[21:41])
    defparam add_34_29.INIT0 = 16'h5aaa;
    defparam add_34_29.INIT1 = 16'h5aaa;
    defparam add_34_29.INJECT1_0 = "NO";
    defparam add_34_29.INJECT1_1 = "NO";
    FD1P3AX bus_err_address_i0_i28 (.D(wb_addr[28]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[28])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(258[9] 260[31])
    defparam bus_err_address_i0_i28.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i27 (.D(wb_addr[27]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[27])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(258[9] 260[31])
    defparam bus_err_address_i0_i27.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i26 (.D(wb_addr[26]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[26])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(258[9] 260[31])
    defparam bus_err_address_i0_i26.GSR = "DISABLED";
    FD1S3AX power_counter_i22 (.D(power_counter_31__N_129[22]), .CK(dac_clk_p_c), 
            .Q(power_counter[22])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 232[54])
    defparam power_counter_i22.GSR = "DISABLED";
    FD1S3AX power_counter_i21 (.D(power_counter_31__N_129[21]), .CK(dac_clk_p_c), 
            .Q(power_counter[21])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 232[54])
    defparam power_counter_i21.GSR = "DISABLED";
    FD1S3AX power_counter_i20 (.D(power_counter_31__N_129[20]), .CK(dac_clk_p_c), 
            .Q(power_counter[20])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 232[54])
    defparam power_counter_i20.GSR = "DISABLED";
    FD1S3AX power_counter_i19 (.D(power_counter_31__N_129[19]), .CK(dac_clk_p_c), 
            .Q(power_counter[19])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 232[54])
    defparam power_counter_i19.GSR = "DISABLED";
    FD1S3AX power_counter_i18 (.D(power_counter_31__N_129[18]), .CK(dac_clk_p_c), 
            .Q(power_counter[18])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 232[54])
    defparam power_counter_i18.GSR = "DISABLED";
    FD1S3AX power_counter_i17 (.D(power_counter_31__N_129[17]), .CK(dac_clk_p_c), 
            .Q(power_counter[17])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 232[54])
    defparam power_counter_i17.GSR = "DISABLED";
    FD1S3AX power_counter_i16 (.D(power_counter_31__N_129[16]), .CK(dac_clk_p_c), 
            .Q(power_counter[16])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 232[54])
    defparam power_counter_i16.GSR = "DISABLED";
    FD1S3AX power_counter_i15 (.D(power_counter_31__N_129[15]), .CK(dac_clk_p_c), 
            .Q(power_counter[15])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 232[54])
    defparam power_counter_i15.GSR = "DISABLED";
    FD1S3AX power_counter_i14 (.D(power_counter_31__N_129[14]), .CK(dac_clk_p_c), 
            .Q(power_counter[14])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 232[54])
    defparam power_counter_i14.GSR = "DISABLED";
    FD1S3AX power_counter_i13 (.D(power_counter_31__N_129[13]), .CK(dac_clk_p_c), 
            .Q(power_counter[13])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 232[54])
    defparam power_counter_i13.GSR = "DISABLED";
    FD1S3AX power_counter_i12 (.D(power_counter_31__N_129[12]), .CK(dac_clk_p_c), 
            .Q(power_counter[12])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 232[54])
    defparam power_counter_i12.GSR = "DISABLED";
    FD1S3AX power_counter_i11 (.D(power_counter_31__N_129[11]), .CK(dac_clk_p_c), 
            .Q(power_counter[11])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 232[54])
    defparam power_counter_i11.GSR = "DISABLED";
    FD1S3AX power_counter_i10 (.D(power_counter_31__N_129[10]), .CK(dac_clk_p_c), 
            .Q(power_counter[10])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 232[54])
    defparam power_counter_i10.GSR = "DISABLED";
    FD1S3AX power_counter_i9 (.D(power_counter_31__N_129[9]), .CK(dac_clk_p_c), 
            .Q(power_counter[9])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 232[54])
    defparam power_counter_i9.GSR = "DISABLED";
    FD1S3AX power_counter_i8 (.D(power_counter_31__N_129[8]), .CK(dac_clk_p_c), 
            .Q(power_counter[8])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 232[54])
    defparam power_counter_i8.GSR = "DISABLED";
    FD1S3AX power_counter_i7 (.D(power_counter_31__N_129[7]), .CK(dac_clk_p_c), 
            .Q(power_counter[7])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 232[54])
    defparam power_counter_i7.GSR = "DISABLED";
    FD1S3AX power_counter_i6 (.D(power_counter_31__N_129[6]), .CK(dac_clk_p_c), 
            .Q(power_counter[6])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 232[54])
    defparam power_counter_i6.GSR = "DISABLED";
    FD1S3AX power_counter_i5 (.D(power_counter_31__N_129[5]), .CK(dac_clk_p_c), 
            .Q(power_counter[5])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 232[54])
    defparam power_counter_i5.GSR = "DISABLED";
    FD1S3AX power_counter_i4 (.D(power_counter_31__N_129[4]), .CK(dac_clk_p_c), 
            .Q(power_counter[4])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 232[54])
    defparam power_counter_i4.GSR = "DISABLED";
    FD1S3AX power_counter_i3 (.D(power_counter_31__N_129[3]), .CK(dac_clk_p_c), 
            .Q(power_counter[3])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 232[54])
    defparam power_counter_i3.GSR = "DISABLED";
    FD1S3AX power_counter_i2 (.D(power_counter_31__N_129[2]), .CK(dac_clk_p_c), 
            .Q(power_counter[2])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 232[54])
    defparam power_counter_i2.GSR = "DISABLED";
    FD1S3AX power_counter_i1 (.D(power_counter_31__N_129[1]), .CK(dac_clk_p_c), 
            .Q(power_counter[1])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(227[9] 232[54])
    defparam power_counter_i1.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i31 (.D(n2131), .CK(dac_clk_p_c), .CD(n9474), 
            .Q(wb_smpl_data[31]));   // d:/documents/git_local/fm_modulator/rtl/top.v(215[9] 223[10])
    defparam wb_smpl_data_i31.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i30 (.D(n2132), .CK(dac_clk_p_c), .CD(n9474), 
            .Q(wb_smpl_data[30]));   // d:/documents/git_local/fm_modulator/rtl/top.v(215[9] 223[10])
    defparam wb_smpl_data_i30.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i29 (.D(n26699), .CK(dac_clk_p_c), .CD(n9474), 
            .Q(wb_smpl_data[29]));   // d:/documents/git_local/fm_modulator/rtl/top.v(215[9] 223[10])
    defparam wb_smpl_data_i29.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i28 (.D(n2134), .CK(dac_clk_p_c), .CD(n9474), 
            .Q(wb_smpl_data[28]));   // d:/documents/git_local/fm_modulator/rtl/top.v(215[9] 223[10])
    defparam wb_smpl_data_i28.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i27 (.D(n2135), .CK(dac_clk_p_c), .CD(n9474), 
            .Q(wb_smpl_data[27]));   // d:/documents/git_local/fm_modulator/rtl/top.v(215[9] 223[10])
    defparam wb_smpl_data_i27.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i26 (.D(n2136), .CK(dac_clk_p_c), .CD(n9474), 
            .Q(wb_smpl_data[26]));   // d:/documents/git_local/fm_modulator/rtl/top.v(215[9] 223[10])
    defparam wb_smpl_data_i26.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i25 (.D(n2137), .CK(dac_clk_p_c), .CD(n9474), 
            .Q(wb_smpl_data[25]));   // d:/documents/git_local/fm_modulator/rtl/top.v(215[9] 223[10])
    defparam wb_smpl_data_i25.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i24 (.D(n2138), .CK(dac_clk_p_c), .CD(n9474), 
            .Q(wb_smpl_data[24]));   // d:/documents/git_local/fm_modulator/rtl/top.v(215[9] 223[10])
    defparam wb_smpl_data_i24.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i25 (.D(wb_addr[25]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[25])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(258[9] 260[31])
    defparam bus_err_address_i0_i25.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i24 (.D(wb_addr[24]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[24])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(258[9] 260[31])
    defparam bus_err_address_i0_i24.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i23 (.D(wb_addr[23]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[23])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(258[9] 260[31])
    defparam bus_err_address_i0_i23.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i22 (.D(wb_addr[22]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[22])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(258[9] 260[31])
    defparam bus_err_address_i0_i22.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i21 (.D(wb_addr[21]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[21])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(258[9] 260[31])
    defparam bus_err_address_i0_i21.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i20 (.D(wb_addr[20]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[20])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(258[9] 260[31])
    defparam bus_err_address_i0_i20.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i19 (.D(wb_addr[19]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[19])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(258[9] 260[31])
    defparam bus_err_address_i0_i19.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i18 (.D(wb_addr[18]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[18])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(258[9] 260[31])
    defparam bus_err_address_i0_i18.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i17 (.D(wb_addr[17]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[17])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(258[9] 260[31])
    defparam bus_err_address_i0_i17.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i16 (.D(wb_addr[16]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[16])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(258[9] 260[31])
    defparam bus_err_address_i0_i16.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i15 (.D(wb_addr[15]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[15])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(258[9] 260[31])
    defparam bus_err_address_i0_i15.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i14 (.D(wb_addr[14]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[14])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(258[9] 260[31])
    defparam bus_err_address_i0_i14.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i13 (.D(wb_addr[13]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[13])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(258[9] 260[31])
    defparam bus_err_address_i0_i13.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i12 (.D(wb_addr[12]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[12])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(258[9] 260[31])
    defparam bus_err_address_i0_i12.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i11 (.D(wb_addr[11]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[11])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(258[9] 260[31])
    defparam bus_err_address_i0_i11.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i10 (.D(wb_addr[10]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[10])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(258[9] 260[31])
    defparam bus_err_address_i0_i10.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i9 (.D(wb_addr[9]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[9])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(258[9] 260[31])
    defparam bus_err_address_i0_i9.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i8 (.D(wb_addr[8]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[8])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(258[9] 260[31])
    defparam bus_err_address_i0_i8.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i7 (.D(wb_addr[7]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[7])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(258[9] 260[31])
    defparam bus_err_address_i0_i7.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i6 (.D(wb_addr[6]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[6])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(258[9] 260[31])
    defparam bus_err_address_i0_i6.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i5 (.D(wb_addr[5]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[5])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(258[9] 260[31])
    defparam bus_err_address_i0_i5.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i4 (.D(wb_addr[4]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[4])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(258[9] 260[31])
    defparam bus_err_address_i0_i4.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i3 (.D(wb_addr[3]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[3])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(258[9] 260[31])
    defparam bus_err_address_i0_i3.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i2 (.D(wb_addr[2]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[2])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(258[9] 260[31])
    defparam bus_err_address_i0_i2.GSR = "DISABLED";
    FD1P3AX bus_err_address_i0_i1 (.D(wb_addr[1]), .SP(wb_err), .CK(dac_clk_p_c), 
            .Q(bus_err_address[1])) /* synthesis lse_init_val=0 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(258[9] 260[31])
    defparam bus_err_address_i0_i1.GSR = "DISABLED";
    LUT4 m1_lut (.Z(n29502)) /* synthesis lut_function=1, syn_instantiated=1 */ ;
    defparam m1_lut.init = 16'hffff;
    FD1S3IX wb_smpl_data_i23 (.D(n2139), .CK(dac_clk_p_c), .CD(n9474), 
            .Q(wb_smpl_data[23]));   // d:/documents/git_local/fm_modulator/rtl/top.v(215[9] 223[10])
    defparam wb_smpl_data_i23.GSR = "DISABLED";
    OB o_baseband_i_pad_5 (.I(o_baseband_i_c_12), .O(o_baseband_i[5]));   // d:/documents/git_local/fm_modulator/rtl/top.v(27[38:50])
    OB o_baseband_i_pad_4 (.I(o_baseband_i_c_11), .O(o_baseband_i[4]));   // d:/documents/git_local/fm_modulator/rtl/top.v(27[38:50])
    OB o_baseband_i_pad_3 (.I(o_baseband_i_c_10), .O(o_baseband_i[3]));   // d:/documents/git_local/fm_modulator/rtl/top.v(27[38:50])
    OB o_baseband_i_pad_2 (.I(n3655), .O(o_baseband_i[2]));   // d:/documents/git_local/fm_modulator/rtl/top.v(27[38:50])
    OB o_baseband_i_pad_1 (.I(o_baseband_i_c_8), .O(o_baseband_i[1]));   // d:/documents/git_local/fm_modulator/rtl/top.v(27[38:50])
    OB o_baseband_i_pad_0 (.I(o_baseband_i_c_7), .O(o_baseband_i[0]));   // d:/documents/git_local/fm_modulator/rtl/top.v(27[38:50])
    OB o_baseband_q_pad_9 (.I(o_baseband_q_c_9), .O(o_baseband_q[9]));   // d:/documents/git_local/fm_modulator/rtl/top.v(27[52:64])
    OB o_baseband_q_pad_8 (.I(o_baseband_q_c_15), .O(o_baseband_q[8]));   // d:/documents/git_local/fm_modulator/rtl/top.v(27[52:64])
    OB o_baseband_q_pad_7 (.I(o_baseband_q_c_14), .O(o_baseband_q[7]));   // d:/documents/git_local/fm_modulator/rtl/top.v(27[52:64])
    OB o_baseband_q_pad_6 (.I(o_baseband_q_c_13), .O(o_baseband_q[6]));   // d:/documents/git_local/fm_modulator/rtl/top.v(27[52:64])
    OB o_baseband_q_pad_5 (.I(o_baseband_q_c_12), .O(o_baseband_q[5]));   // d:/documents/git_local/fm_modulator/rtl/top.v(27[52:64])
    OB o_baseband_q_pad_4 (.I(o_baseband_q_c_11), .O(o_baseband_q[4]));   // d:/documents/git_local/fm_modulator/rtl/top.v(27[52:64])
    OB o_baseband_q_pad_3 (.I(o_baseband_q_c_10), .O(o_baseband_q[3]));   // d:/documents/git_local/fm_modulator/rtl/top.v(27[52:64])
    OB o_baseband_q_pad_2 (.I(n3656), .O(o_baseband_q[2]));   // d:/documents/git_local/fm_modulator/rtl/top.v(27[52:64])
    OB o_baseband_q_pad_1 (.I(o_baseband_q_c_8), .O(o_baseband_q[1]));   // d:/documents/git_local/fm_modulator/rtl/top.v(27[52:64])
    OB o_baseband_q_pad_0 (.I(o_baseband_q_c_7), .O(o_baseband_q[0]));   // d:/documents/git_local/fm_modulator/rtl/top.v(27[52:64])
    OB dac_clk_p_pad (.I(dac_clk_p_c), .O(dac_clk_p));   // d:/documents/git_local/fm_modulator/rtl/top.v(28[49:58])
    OB dac_clk_n_pad (.I(dac_clk_n_c), .O(dac_clk_n));   // d:/documents/git_local/fm_modulator/rtl/top.v(28[60:69])
    OB i_clk_p_pad (.I(i_clk_p_c), .O(i_clk_p));   // d:/documents/git_local/fm_modulator/rtl/top.v(28[13:20])
    OB i_clk_n_pad (.I(i_clk_n_c), .O(i_clk_n));   // d:/documents/git_local/fm_modulator/rtl/top.v(28[22:29])
    OB q_clk_p_pad (.I(q_clk_p_c), .O(q_clk_p));   // d:/documents/git_local/fm_modulator/rtl/top.v(28[31:38])
    OB q_clk_n_pad (.I(q_clk_n_c), .O(q_clk_n));   // d:/documents/git_local/fm_modulator/rtl/top.v(28[40:47])
    IB i_ref_clk_pad (.I(i_ref_clk), .O(i_ref_clk_c));   // d:/documents/git_local/fm_modulator/rtl/top.v(22[12:21])
    IB i_resetb_pad (.I(i_resetb), .O(i_resetb_c));   // d:/documents/git_local/fm_modulator/rtl/top.v(22[23:31])
    IB i_wbu_uart_rx_pad (.I(i_wbu_uart_rx), .O(i_wbu_uart_rx_c));   // d:/documents/git_local/fm_modulator/rtl/top.v(24[12:25])
    FD1S3IX wb_smpl_data_i4 (.D(n2158), .CK(dac_clk_p_c), .CD(n9474), 
            .Q(wb_smpl_data[4]));   // d:/documents/git_local/fm_modulator/rtl/top.v(215[9] 223[10])
    defparam wb_smpl_data_i4.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i22 (.D(n2140), .CK(dac_clk_p_c), .CD(n9474), 
            .Q(wb_smpl_data[22]));   // d:/documents/git_local/fm_modulator/rtl/top.v(215[9] 223[10])
    defparam wb_smpl_data_i22.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i3 (.D(n2159), .CK(dac_clk_p_c), .CD(n9474), 
            .Q(wb_smpl_data[3]));   // d:/documents/git_local/fm_modulator/rtl/top.v(215[9] 223[10])
    defparam wb_smpl_data_i3.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i21 (.D(n2141), .CK(dac_clk_p_c), .CD(n9474), 
            .Q(wb_smpl_data[21]));   // d:/documents/git_local/fm_modulator/rtl/top.v(215[9] 223[10])
    defparam wb_smpl_data_i21.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i2 (.D(n2160), .CK(dac_clk_p_c), .CD(n9474), 
            .Q(wb_smpl_data[2]));   // d:/documents/git_local/fm_modulator/rtl/top.v(215[9] 223[10])
    defparam wb_smpl_data_i2.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i20 (.D(n26704), .CK(dac_clk_p_c), .CD(n9474), 
            .Q(wb_smpl_data[20]));   // d:/documents/git_local/fm_modulator/rtl/top.v(215[9] 223[10])
    defparam wb_smpl_data_i20.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i1 (.D(n2161), .CK(dac_clk_p_c), .CD(n9474), 
            .Q(wb_smpl_data[1]));   // d:/documents/git_local/fm_modulator/rtl/top.v(215[9] 223[10])
    defparam wb_smpl_data_i1.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i19 (.D(n2143), .CK(dac_clk_p_c), .CD(n9474), 
            .Q(wb_smpl_data[19]));   // d:/documents/git_local/fm_modulator/rtl/top.v(215[9] 223[10])
    defparam wb_smpl_data_i19.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i18 (.D(n26703), .CK(dac_clk_p_c), .CD(n9474), 
            .Q(wb_smpl_data[18]));   // d:/documents/git_local/fm_modulator/rtl/top.v(215[9] 223[10])
    defparam wb_smpl_data_i18.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i17 (.D(n26702), .CK(dac_clk_p_c), .CD(n9474), 
            .Q(wb_smpl_data[17]));   // d:/documents/git_local/fm_modulator/rtl/top.v(215[9] 223[10])
    defparam wb_smpl_data_i17.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i16 (.D(n26701), .CK(dac_clk_p_c), .CD(n9474), 
            .Q(wb_smpl_data[16]));   // d:/documents/git_local/fm_modulator/rtl/top.v(215[9] 223[10])
    defparam wb_smpl_data_i16.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i15 (.D(n2147), .CK(dac_clk_p_c), .CD(n9474), 
            .Q(wb_smpl_data[15]));   // d:/documents/git_local/fm_modulator/rtl/top.v(215[9] 223[10])
    defparam wb_smpl_data_i15.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i14 (.D(n2148), .CK(dac_clk_p_c), .CD(n9474), 
            .Q(wb_smpl_data[14]));   // d:/documents/git_local/fm_modulator/rtl/top.v(215[9] 223[10])
    defparam wb_smpl_data_i14.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i13 (.D(n2149), .CK(dac_clk_p_c), .CD(n9474), 
            .Q(wb_smpl_data[13]));   // d:/documents/git_local/fm_modulator/rtl/top.v(215[9] 223[10])
    defparam wb_smpl_data_i13.GSR = "DISABLED";
    dynamic_pll lo_gen (.i_clk_2f_N_2249(i_clk_2f_N_2249), .lo_pll_out(lo_pll_out), 
            .i_ref_clk_c(i_ref_clk_c), .pll_clk(pll_clk), .pll_rst(pll_rst), 
            .pll_stb(pll_stb), .pll_we(pll_we), .pll_data_i({pll_data_i}), 
            .pll_addr({pll_addr}), .pll_data_o({pll_data_o}), .pll_ack(pll_ack), 
            .GND_net(GND_net)) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(167[13] 178[5])
    FD1S3IX wb_smpl_data_i12 (.D(n2150), .CK(dac_clk_p_c), .CD(n9474), 
            .Q(wb_smpl_data[12]));   // d:/documents/git_local/fm_modulator/rtl/top.v(215[9] 223[10])
    defparam wb_smpl_data_i12.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i11 (.D(n2151), .CK(dac_clk_p_c), .CD(n9474), 
            .Q(wb_smpl_data[11]));   // d:/documents/git_local/fm_modulator/rtl/top.v(215[9] 223[10])
    defparam wb_smpl_data_i11.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i10 (.D(n26696), .CK(dac_clk_p_c), .CD(n9474), 
            .Q(wb_smpl_data[10]));   // d:/documents/git_local/fm_modulator/rtl/top.v(215[9] 223[10])
    defparam wb_smpl_data_i10.GSR = "DISABLED";
    \txuartlite(TIMING_BITS=24,CLOCKS_PER_BAUD=10000)  txtransport (.dac_clk_p_c(dac_clk_p_c), 
            .dac_clk_p_c_enable_322(dac_clk_p_c_enable_322), .\lcl_data_7__N_511[0] (lcl_data_7__N_511[0]), 
            .zero_baud_counter(zero_baud_counter), .o_wbu_uart_tx_c(o_wbu_uart_tx_c), 
            .n26910(n26910), .GND_net(GND_net), .\state[0] (state_adj_3085[0]), 
            .\lcl_data[7] (lcl_data[7]), .n29502(n29502), .\lcl_data[6] (lcl_data[6]), 
            .\lcl_data_7__N_511[6] (lcl_data_7__N_511[6]), .\lcl_data[5] (lcl_data[5]), 
            .\lcl_data_7__N_511[5] (lcl_data_7__N_511[5]), .\lcl_data[4] (lcl_data[4]), 
            .\lcl_data_7__N_511[4] (lcl_data_7__N_511[4]), .\lcl_data[3] (lcl_data[3]), 
            .\lcl_data_7__N_511[3] (lcl_data_7__N_511[3]), .\lcl_data[2] (lcl_data[2]), 
            .\lcl_data_7__N_511[2] (lcl_data_7__N_511[2]), .\lcl_data[1] (lcl_data[1]), 
            .\lcl_data_7__N_511[1] (lcl_data_7__N_511[1]), .o_busy_N_536(o_busy_N_536), 
            .tx_busy(tx_busy), .n17844(n17844)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(62[58:115])
    FD1S3IX wb_smpl_data_i9 (.D(n26695), .CK(dac_clk_p_c), .CD(n9474), 
            .Q(wb_smpl_data[9]));   // d:/documents/git_local/fm_modulator/rtl/top.v(215[9] 223[10])
    defparam wb_smpl_data_i9.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i8 (.D(n2154), .CK(dac_clk_p_c), .CD(n9474), 
            .Q(wb_smpl_data[8]));   // d:/documents/git_local/fm_modulator/rtl/top.v(215[9] 223[10])
    defparam wb_smpl_data_i8.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i7 (.D(n2155), .CK(dac_clk_p_c), .CD(n9474), 
            .Q(wb_smpl_data[7]));   // d:/documents/git_local/fm_modulator/rtl/top.v(215[9] 223[10])
    defparam wb_smpl_data_i7.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i6 (.D(n2156), .CK(dac_clk_p_c), .CD(n9474), 
            .Q(wb_smpl_data[6]));   // d:/documents/git_local/fm_modulator/rtl/top.v(215[9] 223[10])
    defparam wb_smpl_data_i6.GSR = "DISABLED";
    FD1S3IX wb_smpl_data_i5 (.D(n26694), .CK(dac_clk_p_c), .CD(n9474), 
            .Q(wb_smpl_data[5]));   // d:/documents/git_local/fm_modulator/rtl/top.v(215[9] 223[10])
    defparam wb_smpl_data_i5.GSR = "DISABLED";
    LUT4 m0_lut (.Z(n29501)) /* synthesis lut_function=0, syn_instantiated=1 */ ;
    defparam m0_lut.init = 16'h0000;
    
endmodule
//
// Verilog Description of module \rxuartlite(CLOCKS_PER_BAUD=10000) 
//

module \rxuartlite(CLOCKS_PER_BAUD=10000)  (dac_clk_p_c, \rx_data[0] , rx_stb, 
            i_wbu_uart_rx_c, chg_counter, dac_clk_p_c_enable_175, chg_counter_23__N_406, 
            GND_net, \rx_data[6] , \rx_data[5] , \rx_data[4] , \rx_data[3] , 
            \rx_data[2] , \rx_data[1] ) /* synthesis syn_module_defined=1 */ ;
    input dac_clk_p_c;
    output \rx_data[0] ;
    output rx_stb;
    input i_wbu_uart_rx_c;
    output [23:0]chg_counter;
    input dac_clk_p_c_enable_175;
    output chg_counter_23__N_406;
    input GND_net;
    output \rx_data[6] ;
    output \rx_data[5] ;
    output \rx_data[4] ;
    output \rx_data[3] ;
    output \rx_data[2] ;
    output \rx_data[1] ;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(28[49:58])
    
    wire qq_uart, q_uart, ck_uart, o_data_7__N_418;
    wire [7:0]data_reg;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(142[12:20])
    wire [3:0]state;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(75[13:18])
    
    wire dac_clk_p_c_enable_348;
    wire [3:0]state_3__N_322;
    
    wire half_baud_time, half_baud_time_N_457;
    wire [23:0]baud_counter;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(78[17:29])
    
    wire dac_clk_p_c_enable_413, baud_counter_23__N_445;
    wire [23:0]baud_counter_23__N_421;
    wire [23:0]n534;
    
    wire n17659;
    wire [23:0]n290;
    
    wire n17660;
    wire [3:0]n560;
    
    wire zero_baud_counter, dac_clk_p_c_enable_141, n14916, n17658, 
        n17657, n17656, n17590, n17589, n17588, n17587, n17586, 
        n17585, n26803, zero_baud_counter_N_454, n11685, n17584, state_3__N_415, 
        n17635, half_baud_time_N_458, n26782, n20490, n21083, n21275, 
        n21273, n21257, n21255, n21196, n21249, n21200, n26921, 
        n179, n17583, n17634, n17633, data_reg_7__N_416, n17582, 
        n17632, n17631, n17581, n17630, n17629, n17580, n17628, 
        n17627, n17626, n17625, n17579, n17624, n25928, n25929, 
        n172, n27166, n27165, dac_clk_p_c_enable_344, n17667, n17666, 
        n17665, n17664, n17663, n17662, n17661;
    
    FD1S3AY qq_uart_70 (.D(q_uart), .CK(dac_clk_p_c), .Q(qq_uart)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(90[9] 91[66])
    defparam qq_uart_70.GSR = "DISABLED";
    FD1S3AY ck_uart_71 (.D(qq_uart), .CK(dac_clk_p_c), .Q(ck_uart)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(90[9] 91[66])
    defparam ck_uart_71.GSR = "DISABLED";
    FD1P3AX o_data__i1 (.D(data_reg[0]), .SP(o_data_7__N_418), .CK(dac_clk_p_c), 
            .Q(\rx_data[0] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(155[9] 161[18])
    defparam o_data__i1.GSR = "DISABLED";
    FD1P3AY state_i0 (.D(state_3__N_322[0]), .SP(dac_clk_p_c_enable_348), 
            .CK(dac_clk_p_c), .Q(state[0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(116[9] 134[5])
    defparam state_i0.GSR = "DISABLED";
    FD1S3AX half_baud_time_73 (.D(half_baud_time_N_457), .CK(dac_clk_p_c), 
            .Q(half_baud_time)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(111[9] 112[70])
    defparam half_baud_time_73.GSR = "DISABLED";
    FD1S3AX o_wr_76 (.D(o_data_7__N_418), .CK(dac_clk_p_c), .Q(rx_stb)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(155[9] 161[18])
    defparam o_wr_76.GSR = "DISABLED";
    FD1S3AY q_uart_69 (.D(i_wbu_uart_rx_c), .CK(dac_clk_p_c), .Q(q_uart)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(90[9] 91[66])
    defparam q_uart_69.GSR = "DISABLED";
    FD1P3JX baud_counter_i1 (.D(baud_counter_23__N_421[1]), .SP(dac_clk_p_c_enable_413), 
            .PD(baud_counter_23__N_445), .CK(dac_clk_p_c), .Q(baud_counter[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i1.GSR = "DISABLED";
    FD1P3IX chg_counter__i0 (.D(n534[0]), .SP(dac_clk_p_c_enable_175), .CD(chg_counter_23__N_406), 
            .CK(dac_clk_p_c), .Q(chg_counter[0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[34])
    defparam chg_counter__i0.GSR = "DISABLED";
    FD1P3JX baud_counter_i2 (.D(baud_counter_23__N_421[2]), .SP(dac_clk_p_c_enable_413), 
            .PD(baud_counter_23__N_445), .CK(dac_clk_p_c), .Q(baud_counter[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i2.GSR = "DISABLED";
    FD1P3JX baud_counter_i3 (.D(baud_counter_23__N_421[3]), .SP(dac_clk_p_c_enable_413), 
            .PD(baud_counter_23__N_445), .CK(dac_clk_p_c), .Q(baud_counter[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i3.GSR = "DISABLED";
    CCU2D sub_49_add_2_9 (.A0(baud_counter[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17659), .COUT(n17660), .S0(n290[7]), .S1(n290[8]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_9.INIT0 = 16'h5555;
    defparam sub_49_add_2_9.INIT1 = 16'h5555;
    defparam sub_49_add_2_9.INJECT1_0 = "NO";
    defparam sub_49_add_2_9.INJECT1_1 = "NO";
    LUT4 i779_2_lut_3_lut_4_lut (.A(state[0]), .B(state[3]), .C(state[2]), 
         .D(state[1]), .Z(n560[2])) /* synthesis lut_function=(A (B (C)+!B !(C (D)+!C !(D)))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(133[13:22])
    defparam i779_2_lut_3_lut_4_lut.init = 16'hd2f0;
    FD1P3AY zero_baud_counter_79 (.D(n14916), .SP(dac_clk_p_c_enable_141), 
            .CK(dac_clk_p_c), .Q(zero_baud_counter)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(187[9] 195[29])
    defparam zero_baud_counter_79.GSR = "DISABLED";
    CCU2D sub_49_add_2_7 (.A0(baud_counter[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17658), .COUT(n17659), .S0(n290[5]), .S1(n290[6]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_7.INIT0 = 16'h5555;
    defparam sub_49_add_2_7.INIT1 = 16'h5555;
    defparam sub_49_add_2_7.INJECT1_0 = "NO";
    defparam sub_49_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_49_add_2_5 (.A0(baud_counter[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17657), .COUT(n17658), .S0(n290[3]), .S1(n290[4]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_5.INIT0 = 16'h5555;
    defparam sub_49_add_2_5.INIT1 = 16'h5555;
    defparam sub_49_add_2_5.INJECT1_0 = "NO";
    defparam sub_49_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_49_add_2_3 (.A0(baud_counter[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17656), .COUT(n17657), .S0(n290[1]), .S1(n290[2]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_3.INIT0 = 16'h5555;
    defparam sub_49_add_2_3.INIT1 = 16'h5555;
    defparam sub_49_add_2_3.INJECT1_0 = "NO";
    defparam sub_49_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_49_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(baud_counter[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n17656), .S1(n290[0]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_1.INIT0 = 16'hF000;
    defparam sub_49_add_2_1.INIT1 = 16'h5555;
    defparam sub_49_add_2_1.INJECT1_0 = "NO";
    defparam sub_49_add_2_1.INJECT1_1 = "NO";
    FD1P3IX chg_counter__i23 (.D(n534[23]), .SP(dac_clk_p_c_enable_175), 
            .CD(chg_counter_23__N_406), .CK(dac_clk_p_c), .Q(chg_counter[23])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[34])
    defparam chg_counter__i23.GSR = "DISABLED";
    FD1P3JX baud_counter_i8 (.D(baud_counter_23__N_421[8]), .SP(dac_clk_p_c_enable_413), 
            .PD(baud_counter_23__N_445), .CK(dac_clk_p_c), .Q(baud_counter[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i8.GSR = "DISABLED";
    FD1P3IX chg_counter__i22 (.D(n534[22]), .SP(dac_clk_p_c_enable_175), 
            .CD(chg_counter_23__N_406), .CK(dac_clk_p_c), .Q(chg_counter[22])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[34])
    defparam chg_counter__i22.GSR = "DISABLED";
    FD1P3IX chg_counter__i21 (.D(n534[21]), .SP(dac_clk_p_c_enable_175), 
            .CD(chg_counter_23__N_406), .CK(dac_clk_p_c), .Q(chg_counter[21])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[34])
    defparam chg_counter__i21.GSR = "DISABLED";
    FD1P3IX chg_counter__i20 (.D(n534[20]), .SP(dac_clk_p_c_enable_175), 
            .CD(chg_counter_23__N_406), .CK(dac_clk_p_c), .Q(chg_counter[20])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[34])
    defparam chg_counter__i20.GSR = "DISABLED";
    FD1P3IX chg_counter__i19 (.D(n534[19]), .SP(dac_clk_p_c_enable_175), 
            .CD(chg_counter_23__N_406), .CK(dac_clk_p_c), .Q(chg_counter[19])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[34])
    defparam chg_counter__i19.GSR = "DISABLED";
    FD1P3IX chg_counter__i18 (.D(n534[18]), .SP(dac_clk_p_c_enable_175), 
            .CD(chg_counter_23__N_406), .CK(dac_clk_p_c), .Q(chg_counter[18])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[34])
    defparam chg_counter__i18.GSR = "DISABLED";
    FD1P3IX chg_counter__i17 (.D(n534[17]), .SP(dac_clk_p_c_enable_175), 
            .CD(chg_counter_23__N_406), .CK(dac_clk_p_c), .Q(chg_counter[17])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[34])
    defparam chg_counter__i17.GSR = "DISABLED";
    FD1P3IX chg_counter__i16 (.D(n534[16]), .SP(dac_clk_p_c_enable_175), 
            .CD(chg_counter_23__N_406), .CK(dac_clk_p_c), .Q(chg_counter[16])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[34])
    defparam chg_counter__i16.GSR = "DISABLED";
    FD1P3IX chg_counter__i15 (.D(n534[15]), .SP(dac_clk_p_c_enable_175), 
            .CD(chg_counter_23__N_406), .CK(dac_clk_p_c), .Q(chg_counter[15])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[34])
    defparam chg_counter__i15.GSR = "DISABLED";
    FD1P3IX chg_counter__i14 (.D(n534[14]), .SP(dac_clk_p_c_enable_175), 
            .CD(chg_counter_23__N_406), .CK(dac_clk_p_c), .Q(chg_counter[14])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[34])
    defparam chg_counter__i14.GSR = "DISABLED";
    FD1P3IX chg_counter__i13 (.D(n534[13]), .SP(dac_clk_p_c_enable_175), 
            .CD(chg_counter_23__N_406), .CK(dac_clk_p_c), .Q(chg_counter[13])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[34])
    defparam chg_counter__i13.GSR = "DISABLED";
    FD1P3IX chg_counter__i12 (.D(n534[12]), .SP(dac_clk_p_c_enable_175), 
            .CD(chg_counter_23__N_406), .CK(dac_clk_p_c), .Q(chg_counter[12])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[34])
    defparam chg_counter__i12.GSR = "DISABLED";
    FD1P3IX chg_counter__i11 (.D(n534[11]), .SP(dac_clk_p_c_enable_175), 
            .CD(chg_counter_23__N_406), .CK(dac_clk_p_c), .Q(chg_counter[11])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[34])
    defparam chg_counter__i11.GSR = "DISABLED";
    FD1P3IX chg_counter__i10 (.D(n534[10]), .SP(dac_clk_p_c_enable_175), 
            .CD(chg_counter_23__N_406), .CK(dac_clk_p_c), .Q(chg_counter[10])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[34])
    defparam chg_counter__i10.GSR = "DISABLED";
    FD1P3IX chg_counter__i9 (.D(n534[9]), .SP(dac_clk_p_c_enable_175), .CD(chg_counter_23__N_406), 
            .CK(dac_clk_p_c), .Q(chg_counter[9])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[34])
    defparam chg_counter__i9.GSR = "DISABLED";
    FD1P3IX chg_counter__i8 (.D(n534[8]), .SP(dac_clk_p_c_enable_175), .CD(chg_counter_23__N_406), 
            .CK(dac_clk_p_c), .Q(chg_counter[8])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[34])
    defparam chg_counter__i8.GSR = "DISABLED";
    FD1P3IX chg_counter__i7 (.D(n534[7]), .SP(dac_clk_p_c_enable_175), .CD(chg_counter_23__N_406), 
            .CK(dac_clk_p_c), .Q(chg_counter[7])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[34])
    defparam chg_counter__i7.GSR = "DISABLED";
    FD1P3IX chg_counter__i6 (.D(n534[6]), .SP(dac_clk_p_c_enable_175), .CD(chg_counter_23__N_406), 
            .CK(dac_clk_p_c), .Q(chg_counter[6])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[34])
    defparam chg_counter__i6.GSR = "DISABLED";
    FD1P3IX chg_counter__i5 (.D(n534[5]), .SP(dac_clk_p_c_enable_175), .CD(chg_counter_23__N_406), 
            .CK(dac_clk_p_c), .Q(chg_counter[5])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[34])
    defparam chg_counter__i5.GSR = "DISABLED";
    FD1P3IX chg_counter__i4 (.D(n534[4]), .SP(dac_clk_p_c_enable_175), .CD(chg_counter_23__N_406), 
            .CK(dac_clk_p_c), .Q(chg_counter[4])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[34])
    defparam chg_counter__i4.GSR = "DISABLED";
    FD1P3IX chg_counter__i3 (.D(n534[3]), .SP(dac_clk_p_c_enable_175), .CD(chg_counter_23__N_406), 
            .CK(dac_clk_p_c), .Q(chg_counter[3])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[34])
    defparam chg_counter__i3.GSR = "DISABLED";
    FD1P3IX chg_counter__i2 (.D(n534[2]), .SP(dac_clk_p_c_enable_175), .CD(chg_counter_23__N_406), 
            .CK(dac_clk_p_c), .Q(chg_counter[2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[34])
    defparam chg_counter__i2.GSR = "DISABLED";
    FD1P3IX chg_counter__i1 (.D(n534[1]), .SP(dac_clk_p_c_enable_175), .CD(chg_counter_23__N_406), 
            .CK(dac_clk_p_c), .Q(chg_counter[1])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(99[9] 103[34])
    defparam chg_counter__i1.GSR = "DISABLED";
    FD1P3JX baud_counter_i9 (.D(baud_counter_23__N_421[9]), .SP(dac_clk_p_c_enable_413), 
            .PD(baud_counter_23__N_445), .CK(dac_clk_p_c), .Q(baud_counter[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i9.GSR = "DISABLED";
    FD1P3JX baud_counter_i10 (.D(baud_counter_23__N_421[10]), .SP(dac_clk_p_c_enable_413), 
            .PD(baud_counter_23__N_445), .CK(dac_clk_p_c), .Q(baud_counter[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i10.GSR = "DISABLED";
    FD1P3JX baud_counter_i13 (.D(baud_counter_23__N_421[13]), .SP(dac_clk_p_c_enable_413), 
            .PD(baud_counter_23__N_445), .CK(dac_clk_p_c), .Q(baud_counter[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i13.GSR = "DISABLED";
    CCU2D add_90_25 (.A0(chg_counter[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n17590), .S0(n534[23]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:33])
    defparam add_90_25.INIT0 = 16'h5aaa;
    defparam add_90_25.INIT1 = 16'h0000;
    defparam add_90_25.INJECT1_0 = "NO";
    defparam add_90_25.INJECT1_1 = "NO";
    CCU2D add_90_23 (.A0(chg_counter[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17589), .COUT(n17590), .S0(n534[21]), 
          .S1(n534[22]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:33])
    defparam add_90_23.INIT0 = 16'h5aaa;
    defparam add_90_23.INIT1 = 16'h5aaa;
    defparam add_90_23.INJECT1_0 = "NO";
    defparam add_90_23.INJECT1_1 = "NO";
    CCU2D add_90_21 (.A0(chg_counter[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17588), .COUT(n17589), .S0(n534[19]), 
          .S1(n534[20]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:33])
    defparam add_90_21.INIT0 = 16'h5aaa;
    defparam add_90_21.INIT1 = 16'h5aaa;
    defparam add_90_21.INJECT1_0 = "NO";
    defparam add_90_21.INJECT1_1 = "NO";
    CCU2D add_90_19 (.A0(chg_counter[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17587), .COUT(n17588), .S0(n534[17]), 
          .S1(n534[18]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:33])
    defparam add_90_19.INIT0 = 16'h5aaa;
    defparam add_90_19.INIT1 = 16'h5aaa;
    defparam add_90_19.INJECT1_0 = "NO";
    defparam add_90_19.INJECT1_1 = "NO";
    CCU2D add_90_17 (.A0(chg_counter[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17586), .COUT(n17587), .S0(n534[15]), 
          .S1(n534[16]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:33])
    defparam add_90_17.INIT0 = 16'h5aaa;
    defparam add_90_17.INIT1 = 16'h5aaa;
    defparam add_90_17.INJECT1_0 = "NO";
    defparam add_90_17.INJECT1_1 = "NO";
    CCU2D add_90_15 (.A0(chg_counter[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17585), .COUT(n17586), .S0(n534[13]), 
          .S1(n534[14]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:33])
    defparam add_90_15.INIT0 = 16'h5aaa;
    defparam add_90_15.INIT1 = 16'h5aaa;
    defparam add_90_15.INJECT1_0 = "NO";
    defparam add_90_15.INJECT1_1 = "NO";
    LUT4 i11537_3_lut_4_lut (.A(state[0]), .B(n26803), .C(zero_baud_counter_N_454), 
         .D(n290[1]), .Z(baud_counter_23__N_421[1])) /* synthesis lut_function=(A (B (C+(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(144[27:48])
    defparam i11537_3_lut_4_lut.init = 16'hddd0;
    LUT4 i1_2_lut_3_lut_4_lut (.A(state[0]), .B(n26803), .C(zero_baud_counter_N_454), 
         .D(baud_counter_23__N_445), .Z(n11685)) /* synthesis lut_function=(A ((C+(D))+!B)+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(144[27:48])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfff2;
    LUT4 i11536_3_lut_4_lut (.A(state[0]), .B(n26803), .C(zero_baud_counter_N_454), 
         .D(n290[2]), .Z(baud_counter_23__N_421[2])) /* synthesis lut_function=(A (B (C+(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(144[27:48])
    defparam i11536_3_lut_4_lut.init = 16'hddd0;
    LUT4 i11535_3_lut_4_lut (.A(state[0]), .B(n26803), .C(zero_baud_counter_N_454), 
         .D(n290[3]), .Z(baud_counter_23__N_421[3])) /* synthesis lut_function=(A (B (C+(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(144[27:48])
    defparam i11535_3_lut_4_lut.init = 16'hddd0;
    LUT4 i22713_3_lut_4_lut (.A(state[0]), .B(n26803), .C(baud_counter_23__N_445), 
         .D(zero_baud_counter_N_454), .Z(n14916)) /* synthesis lut_function=(!(A (B (C+(D))+!B (C))+!A (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(144[27:48])
    defparam i22713_3_lut_4_lut.init = 16'h020f;
    LUT4 i11534_3_lut_4_lut (.A(state[0]), .B(n26803), .C(zero_baud_counter_N_454), 
         .D(n290[8]), .Z(baud_counter_23__N_421[8])) /* synthesis lut_function=(A (B (C+(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(144[27:48])
    defparam i11534_3_lut_4_lut.init = 16'hddd0;
    LUT4 i11533_3_lut_4_lut (.A(state[0]), .B(n26803), .C(zero_baud_counter_N_454), 
         .D(n290[9]), .Z(baud_counter_23__N_421[9])) /* synthesis lut_function=(A (B (C+(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(144[27:48])
    defparam i11533_3_lut_4_lut.init = 16'hddd0;
    LUT4 i11532_3_lut_4_lut (.A(state[0]), .B(n26803), .C(zero_baud_counter_N_454), 
         .D(n290[10]), .Z(baud_counter_23__N_421[10])) /* synthesis lut_function=(A (B (C+(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(144[27:48])
    defparam i11532_3_lut_4_lut.init = 16'hddd0;
    LUT4 i11531_3_lut_4_lut (.A(state[0]), .B(n26803), .C(zero_baud_counter_N_454), 
         .D(n290[13]), .Z(baud_counter_23__N_421[13])) /* synthesis lut_function=(A (B (C+(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(144[27:48])
    defparam i11531_3_lut_4_lut.init = 16'hddd0;
    LUT4 i11000_3_lut_4_lut (.A(state[0]), .B(n26803), .C(zero_baud_counter_N_454), 
         .D(n290[0]), .Z(baud_counter_23__N_421[0])) /* synthesis lut_function=(A (B (C+(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(144[27:48])
    defparam i11000_3_lut_4_lut.init = 16'hddd0;
    CCU2D add_90_13 (.A0(chg_counter[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17584), .COUT(n17585), .S0(n534[11]), 
          .S1(n534[12]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:33])
    defparam add_90_13.INIT0 = 16'h5aaa;
    defparam add_90_13.INIT1 = 16'h5aaa;
    defparam add_90_13.INJECT1_0 = "NO";
    defparam add_90_13.INJECT1_1 = "NO";
    LUT4 i1_3_lut (.A(ck_uart), .B(state_3__N_415), .C(half_baud_time), 
         .Z(baud_counter_23__N_445)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(171[6:57])
    defparam i1_3_lut.init = 16'h4040;
    LUT4 zero_baud_counter_I_0_2_lut (.A(zero_baud_counter), .B(state[3]), 
         .Z(zero_baud_counter_N_454)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(175[11:52])
    defparam zero_baud_counter_I_0_2_lut.init = 16'h2222;
    LUT4 qq_uart_I_0_2_lut (.A(qq_uart), .B(ck_uart), .Z(chg_counter_23__N_406)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(100[6:24])
    defparam qq_uart_I_0_2_lut.init = 16'h6666;
    CCU2D sub_394_add_2_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n17635), .S0(half_baud_time_N_458));
    defparam sub_394_add_2_cout.INIT0 = 16'h0000;
    defparam sub_394_add_2_cout.INIT1 = 16'h0000;
    defparam sub_394_add_2_cout.INJECT1_0 = "NO";
    defparam sub_394_add_2_cout.INJECT1_1 = "NO";
    LUT4 i1_4_lut (.A(zero_baud_counter_N_454), .B(n26782), .C(baud_counter_23__N_445), 
         .D(n20490), .Z(dac_clk_p_c_enable_141)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;
    defparam i1_4_lut.init = 16'hfffb;
    LUT4 i1_4_lut_adj_133 (.A(n21083), .B(n21275), .C(n21273), .D(n21257), 
         .Z(n20490)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_4_lut_adj_133.init = 16'h0002;
    LUT4 i1_4_lut_adj_134 (.A(baud_counter[16]), .B(baud_counter[14]), .C(baud_counter[2]), 
         .D(baud_counter[0]), .Z(n21083)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut_adj_134.init = 16'h0100;
    LUT4 i18913_4_lut (.A(baud_counter[23]), .B(n21255), .C(n21196), .D(baud_counter[11]), 
         .Z(n21275)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18913_4_lut.init = 16'hfffe;
    LUT4 i18911_4_lut (.A(baud_counter[10]), .B(n21249), .C(n21200), .D(baud_counter[17]), 
         .Z(n21273)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18911_4_lut.init = 16'hfffe;
    LUT4 i1_3_lut_4_lut (.A(state[0]), .B(n26921), .C(ck_uart), .D(state[3]), 
         .Z(n179)) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;
    defparam i1_3_lut_4_lut.init = 16'he000;
    LUT4 i18895_4_lut (.A(baud_counter[22]), .B(baud_counter[8]), .C(baud_counter[15]), 
         .D(baud_counter[5]), .Z(n21257)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18895_4_lut.init = 16'hfffe;
    LUT4 i18893_4_lut (.A(baud_counter[20]), .B(baud_counter[9]), .C(baud_counter[13]), 
         .D(baud_counter[19]), .Z(n21255)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18893_4_lut.init = 16'hfffe;
    LUT4 i18835_2_lut (.A(baud_counter[7]), .B(baud_counter[4]), .Z(n21196)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i18835_2_lut.init = 16'heeee;
    LUT4 i18887_4_lut (.A(baud_counter[21]), .B(baud_counter[3]), .C(baud_counter[1]), 
         .D(baud_counter[18]), .Z(n21249)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i18887_4_lut.init = 16'hfffe;
    LUT4 i18839_2_lut (.A(baud_counter[6]), .B(baud_counter[12]), .Z(n21200)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i18839_2_lut.init = 16'heeee;
    CCU2D add_90_11 (.A0(chg_counter[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17583), .COUT(n17584), .S0(n534[9]), .S1(n534[10]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:33])
    defparam add_90_11.INIT0 = 16'h5aaa;
    defparam add_90_11.INIT1 = 16'h5aaa;
    defparam add_90_11.INJECT1_0 = "NO";
    defparam add_90_11.INJECT1_1 = "NO";
    CCU2D sub_394_add_2_24 (.A0(chg_counter[22]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[23]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17634), .COUT(n17635));
    defparam sub_394_add_2_24.INIT0 = 16'h5555;
    defparam sub_394_add_2_24.INIT1 = 16'h5555;
    defparam sub_394_add_2_24.INJECT1_0 = "NO";
    defparam sub_394_add_2_24.INJECT1_1 = "NO";
    CCU2D sub_394_add_2_22 (.A0(chg_counter[20]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[21]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17633), .COUT(n17634));
    defparam sub_394_add_2_22.INIT0 = 16'h5555;
    defparam sub_394_add_2_22.INIT1 = 16'h5555;
    defparam sub_394_add_2_22.INJECT1_0 = "NO";
    defparam sub_394_add_2_22.INJECT1_1 = "NO";
    LUT4 zero_baud_counter_I_0_82_2_lut_3_lut_4_lut (.A(state[3]), .B(n26921), 
         .C(zero_baud_counter), .D(state[0]), .Z(data_reg_7__N_416)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(144[27:48])
    defparam zero_baud_counter_I_0_82_2_lut_3_lut_4_lut.init = 16'hf0d0;
    CCU2D add_90_9 (.A0(chg_counter[7]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(chg_counter[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n17582), .COUT(n17583), .S0(n534[7]), .S1(n534[8]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:33])
    defparam add_90_9.INIT0 = 16'h5aaa;
    defparam add_90_9.INIT1 = 16'h5aaa;
    defparam add_90_9.INJECT1_0 = "NO";
    defparam add_90_9.INJECT1_1 = "NO";
    CCU2D sub_394_add_2_20 (.A0(chg_counter[18]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[19]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17632), .COUT(n17633));
    defparam sub_394_add_2_20.INIT0 = 16'h5555;
    defparam sub_394_add_2_20.INIT1 = 16'h5555;
    defparam sub_394_add_2_20.INJECT1_0 = "NO";
    defparam sub_394_add_2_20.INJECT1_1 = "NO";
    CCU2D sub_394_add_2_18 (.A0(chg_counter[16]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[17]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17631), .COUT(n17632));
    defparam sub_394_add_2_18.INIT0 = 16'h5555;
    defparam sub_394_add_2_18.INIT1 = 16'h5555;
    defparam sub_394_add_2_18.INJECT1_0 = "NO";
    defparam sub_394_add_2_18.INJECT1_1 = "NO";
    CCU2D add_90_7 (.A0(chg_counter[5]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(chg_counter[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n17581), .COUT(n17582), .S0(n534[5]), .S1(n534[6]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:33])
    defparam add_90_7.INIT0 = 16'h5aaa;
    defparam add_90_7.INIT1 = 16'h5aaa;
    defparam add_90_7.INJECT1_0 = "NO";
    defparam add_90_7.INJECT1_1 = "NO";
    CCU2D sub_394_add_2_16 (.A0(chg_counter[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17630), .COUT(n17631));
    defparam sub_394_add_2_16.INIT0 = 16'h5555;
    defparam sub_394_add_2_16.INIT1 = 16'h5555;
    defparam sub_394_add_2_16.INJECT1_0 = "NO";
    defparam sub_394_add_2_16.INJECT1_1 = "NO";
    CCU2D sub_394_add_2_14 (.A0(chg_counter[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17629), .COUT(n17630));
    defparam sub_394_add_2_14.INIT0 = 16'h5aaa;
    defparam sub_394_add_2_14.INIT1 = 16'h5555;
    defparam sub_394_add_2_14.INJECT1_0 = "NO";
    defparam sub_394_add_2_14.INJECT1_1 = "NO";
    CCU2D add_90_5 (.A0(chg_counter[3]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(chg_counter[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n17580), .COUT(n17581), .S0(n534[3]), .S1(n534[4]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:33])
    defparam add_90_5.INIT0 = 16'h5aaa;
    defparam add_90_5.INIT1 = 16'h5aaa;
    defparam add_90_5.INJECT1_0 = "NO";
    defparam add_90_5.INJECT1_1 = "NO";
    CCU2D sub_394_add_2_12 (.A0(chg_counter[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17628), .COUT(n17629));
    defparam sub_394_add_2_12.INIT0 = 16'h5555;
    defparam sub_394_add_2_12.INIT1 = 16'h5555;
    defparam sub_394_add_2_12.INJECT1_0 = "NO";
    defparam sub_394_add_2_12.INJECT1_1 = "NO";
    CCU2D sub_394_add_2_10 (.A0(chg_counter[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17627), .COUT(n17628));
    defparam sub_394_add_2_10.INIT0 = 16'h5aaa;
    defparam sub_394_add_2_10.INIT1 = 16'h5aaa;
    defparam sub_394_add_2_10.INJECT1_0 = "NO";
    defparam sub_394_add_2_10.INJECT1_1 = "NO";
    CCU2D sub_394_add_2_8 (.A0(chg_counter[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17626), .COUT(n17627));
    defparam sub_394_add_2_8.INIT0 = 16'h5555;
    defparam sub_394_add_2_8.INIT1 = 16'h5aaa;
    defparam sub_394_add_2_8.INJECT1_0 = "NO";
    defparam sub_394_add_2_8.INJECT1_1 = "NO";
    CCU2D sub_394_add_2_6 (.A0(chg_counter[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17625), .COUT(n17626));
    defparam sub_394_add_2_6.INIT0 = 16'h5555;
    defparam sub_394_add_2_6.INIT1 = 16'h5555;
    defparam sub_394_add_2_6.INJECT1_0 = "NO";
    defparam sub_394_add_2_6.INJECT1_1 = "NO";
    CCU2D add_90_3 (.A0(chg_counter[1]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(chg_counter[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n17579), .COUT(n17580), .S0(n534[1]), .S1(n534[2]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:33])
    defparam add_90_3.INIT0 = 16'h5aaa;
    defparam add_90_3.INIT1 = 16'h5aaa;
    defparam add_90_3.INJECT1_0 = "NO";
    defparam add_90_3.INJECT1_1 = "NO";
    CCU2D add_90_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(chg_counter[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n17579), .S1(n534[0]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(103[18:33])
    defparam add_90_1.INIT0 = 16'hF000;
    defparam add_90_1.INIT1 = 16'h5555;
    defparam add_90_1.INJECT1_0 = "NO";
    defparam add_90_1.INJECT1_1 = "NO";
    CCU2D sub_394_add_2_4 (.A0(chg_counter[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(chg_counter[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17624), .COUT(n17625));
    defparam sub_394_add_2_4.INIT0 = 16'h5aaa;
    defparam sub_394_add_2_4.INIT1 = 16'h5555;
    defparam sub_394_add_2_4.INJECT1_0 = "NO";
    defparam sub_394_add_2_4.INJECT1_1 = "NO";
    LUT4 state_3__N_415_bdd_2_lut (.A(half_baud_time), .B(ck_uart), .Z(n25928)) /* synthesis lut_function=((B)+!A) */ ;
    defparam state_3__N_415_bdd_2_lut.init = 16'hdddd;
    CCU2D sub_394_add_2_2 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(chg_counter[1]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n17624));
    defparam sub_394_add_2_2.INIT0 = 16'h0000;
    defparam sub_394_add_2_2.INIT1 = 16'h5aaa;
    defparam sub_394_add_2_2.INJECT1_0 = "NO";
    defparam sub_394_add_2_2.INJECT1_1 = "NO";
    LUT4 state_3__N_415_bdd_4_lut (.A(state[0]), .B(state[3]), .C(n26921), 
         .D(ck_uart), .Z(n25929)) /* synthesis lut_function=(A (B)+!A (((D)+!C)+!B)) */ ;
    defparam state_3__N_415_bdd_4_lut.init = 16'hdd9d;
    LUT4 state_3__I_0_80_i4_4_lut_then_4_lut (.A(n172), .B(state[0]), .C(state[2]), 
         .D(state[1]), .Z(n27166)) /* synthesis lut_function=(!(A (B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(125[11] 134[5])
    defparam state_3__I_0_80_i4_4_lut_then_4_lut.init = 16'h7fff;
    LUT4 state_3__I_0_80_i4_4_lut_else_4_lut (.A(state[0]), .B(n179), .C(state[2]), 
         .D(state[1]), .Z(n27165)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(125[11] 134[5])
    defparam state_3__I_0_80_i4_4_lut_else_4_lut.init = 16'heccc;
    LUT4 i1_3_lut_4_lut_adj_135 (.A(state[0]), .B(n26803), .C(ck_uart), 
         .D(zero_baud_counter), .Z(o_data_7__N_418)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(144[27:48])
    defparam i1_3_lut_4_lut_adj_135.init = 16'h1000;
    LUT4 i1_3_lut_adj_136 (.A(state_3__N_415), .B(n179), .C(zero_baud_counter), 
         .Z(dac_clk_p_c_enable_348)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_3_lut_adj_136.init = 16'hfefe;
    LUT4 i21_2_lut (.A(ck_uart), .B(half_baud_time), .Z(n172)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(121[7:35])
    defparam i21_2_lut.init = 16'h4444;
    LUT4 i1_4_lut_adj_137 (.A(state[0]), .B(state[2]), .C(state[3]), .D(state[1]), 
         .Z(state_3__N_415)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_137.init = 16'h8000;
    LUT4 ck_uart_N_448_I_0_2_lut (.A(ck_uart), .B(half_baud_time_N_458), 
         .Z(half_baud_time_N_457)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(112[21:69])
    defparam ck_uart_N_448_I_0_2_lut.init = 16'h4444;
    LUT4 i1_3_lut_4_lut_adj_138 (.A(baud_counter_23__N_445), .B(n26782), 
         .C(state[3]), .D(zero_baud_counter), .Z(dac_clk_p_c_enable_413)) /* synthesis lut_function=(A+!(B (C (D)))) */ ;
    defparam i1_3_lut_4_lut_adj_138.init = 16'hbfff;
    FD1P3IX baud_counter_i23 (.D(n290[23]), .SP(dac_clk_p_c_enable_344), 
            .CD(n11685), .CK(dac_clk_p_c), .Q(baud_counter[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i23.GSR = "DISABLED";
    LUT4 i9648_1_lut (.A(zero_baud_counter), .Z(dac_clk_p_c_enable_344)) /* synthesis lut_function=(!(A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(187[9] 195[29])
    defparam i9648_1_lut.init = 16'h5555;
    FD1P3IX baud_counter_i22 (.D(n290[22]), .SP(dac_clk_p_c_enable_344), 
            .CD(n11685), .CK(dac_clk_p_c), .Q(baud_counter[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i22.GSR = "DISABLED";
    FD1P3IX baud_counter_i21 (.D(n290[21]), .SP(dac_clk_p_c_enable_344), 
            .CD(n11685), .CK(dac_clk_p_c), .Q(baud_counter[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i21.GSR = "DISABLED";
    FD1P3IX baud_counter_i20 (.D(n290[20]), .SP(dac_clk_p_c_enable_344), 
            .CD(n11685), .CK(dac_clk_p_c), .Q(baud_counter[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i20.GSR = "DISABLED";
    FD1P3IX baud_counter_i19 (.D(n290[19]), .SP(dac_clk_p_c_enable_344), 
            .CD(n11685), .CK(dac_clk_p_c), .Q(baud_counter[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i19.GSR = "DISABLED";
    FD1P3IX baud_counter_i18 (.D(n290[18]), .SP(dac_clk_p_c_enable_344), 
            .CD(n11685), .CK(dac_clk_p_c), .Q(baud_counter[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i18.GSR = "DISABLED";
    FD1P3IX baud_counter_i17 (.D(n290[17]), .SP(dac_clk_p_c_enable_344), 
            .CD(n11685), .CK(dac_clk_p_c), .Q(baud_counter[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i17.GSR = "DISABLED";
    LUT4 state_3__I_0_80_i3_4_lut (.A(n172), .B(n560[2]), .C(state_3__N_415), 
         .D(n179), .Z(state_3__N_322[2])) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A !(B+(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(125[11] 134[5])
    defparam state_3__I_0_80_i3_4_lut.init = 16'h5f5c;
    FD1P3IX baud_counter_i16 (.D(n290[16]), .SP(dac_clk_p_c_enable_344), 
            .CD(n11685), .CK(dac_clk_p_c), .Q(baud_counter[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i16.GSR = "DISABLED";
    FD1P3IX baud_counter_i15 (.D(n290[15]), .SP(dac_clk_p_c_enable_344), 
            .CD(n11685), .CK(dac_clk_p_c), .Q(baud_counter[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i15.GSR = "DISABLED";
    LUT4 state_3__I_0_80_i2_4_lut (.A(n172), .B(n560[1]), .C(state_3__N_415), 
         .D(n179), .Z(state_3__N_322[1])) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A !(B+(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(125[11] 134[5])
    defparam state_3__I_0_80_i2_4_lut.init = 16'h5f5c;
    FD1P3IX baud_counter_i14 (.D(n290[14]), .SP(dac_clk_p_c_enable_344), 
            .CD(n11685), .CK(dac_clk_p_c), .Q(baud_counter[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i14.GSR = "DISABLED";
    FD1P3IX baud_counter_i12 (.D(n290[12]), .SP(dac_clk_p_c_enable_344), 
            .CD(n11685), .CK(dac_clk_p_c), .Q(baud_counter[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i12.GSR = "DISABLED";
    FD1P3IX baud_counter_i11 (.D(n290[11]), .SP(dac_clk_p_c_enable_344), 
            .CD(n11685), .CK(dac_clk_p_c), .Q(baud_counter[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i11.GSR = "DISABLED";
    FD1P3IX baud_counter_i7 (.D(n290[7]), .SP(dac_clk_p_c_enable_344), .CD(n11685), 
            .CK(dac_clk_p_c), .Q(baud_counter[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i7.GSR = "DISABLED";
    FD1P3IX baud_counter_i6 (.D(n290[6]), .SP(dac_clk_p_c_enable_344), .CD(n11685), 
            .CK(dac_clk_p_c), .Q(baud_counter[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i6.GSR = "DISABLED";
    FD1P3IX baud_counter_i5 (.D(n290[5]), .SP(dac_clk_p_c_enable_344), .CD(n11685), 
            .CK(dac_clk_p_c), .Q(baud_counter[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i5.GSR = "DISABLED";
    FD1P3IX baud_counter_i4 (.D(n290[4]), .SP(dac_clk_p_c_enable_344), .CD(n11685), 
            .CK(dac_clk_p_c), .Q(baud_counter[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i4.GSR = "DISABLED";
    FD1P3AY state_i3 (.D(state_3__N_322[3]), .SP(dac_clk_p_c_enable_348), 
            .CK(dac_clk_p_c), .Q(state[3])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(116[9] 134[5])
    defparam state_i3.GSR = "DISABLED";
    FD1P3AY state_i2 (.D(state_3__N_322[2]), .SP(dac_clk_p_c_enable_348), 
            .CK(dac_clk_p_c), .Q(state[2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(116[9] 134[5])
    defparam state_i2.GSR = "DISABLED";
    FD1P3AY state_i1 (.D(state_3__N_322[1]), .SP(dac_clk_p_c_enable_348), 
            .CK(dac_clk_p_c), .Q(state[1])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(116[9] 134[5])
    defparam state_i1.GSR = "DISABLED";
    FD1P3AX o_data__i7 (.D(data_reg[6]), .SP(o_data_7__N_418), .CK(dac_clk_p_c), 
            .Q(\rx_data[6] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(155[9] 161[18])
    defparam o_data__i7.GSR = "DISABLED";
    FD1P3AX o_data__i6 (.D(data_reg[5]), .SP(o_data_7__N_418), .CK(dac_clk_p_c), 
            .Q(\rx_data[5] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(155[9] 161[18])
    defparam o_data__i6.GSR = "DISABLED";
    FD1P3AX o_data__i5 (.D(data_reg[4]), .SP(o_data_7__N_418), .CK(dac_clk_p_c), 
            .Q(\rx_data[4] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(155[9] 161[18])
    defparam o_data__i5.GSR = "DISABLED";
    FD1P3AX o_data__i4 (.D(data_reg[3]), .SP(o_data_7__N_418), .CK(dac_clk_p_c), 
            .Q(\rx_data[3] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(155[9] 161[18])
    defparam o_data__i4.GSR = "DISABLED";
    FD1P3AX o_data__i3 (.D(data_reg[2]), .SP(o_data_7__N_418), .CK(dac_clk_p_c), 
            .Q(\rx_data[2] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(155[9] 161[18])
    defparam o_data__i3.GSR = "DISABLED";
    FD1P3AX o_data__i2 (.D(data_reg[1]), .SP(o_data_7__N_418), .CK(dac_clk_p_c), 
            .Q(\rx_data[1] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(155[9] 161[18])
    defparam o_data__i2.GSR = "DISABLED";
    LUT4 i772_2_lut_3_lut (.A(state[0]), .B(state[3]), .C(state[1]), .Z(n560[1])) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(133[13:22])
    defparam i772_2_lut_3_lut.init = 16'hd2d2;
    LUT4 i6518_2_lut_rep_598 (.A(state[1]), .B(state[2]), .Z(n26921)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(129[7:26])
    defparam i6518_2_lut_rep_598.init = 16'heeee;
    LUT4 i1_2_lut_rep_480_3_lut (.A(state[1]), .B(state[2]), .C(state[3]), 
         .Z(n26803)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(129[7:26])
    defparam i1_2_lut_rep_480_3_lut.init = 16'hefef;
    LUT4 i1_2_lut_rep_459_3_lut_4_lut (.A(state[1]), .B(state[2]), .C(state[0]), 
         .D(state[3]), .Z(n26782)) /* synthesis lut_function=(A+(B+!(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(129[7:26])
    defparam i1_2_lut_rep_459_3_lut_4_lut.init = 16'hefff;
    PFUMX i24757 (.BLUT(n27165), .ALUT(n27166), .C0(state[3]), .Z(state_3__N_322[3]));
    PFUMX i24111 (.BLUT(n25929), .ALUT(n25928), .C0(state_3__N_415), .Z(state_3__N_322[0]));
    FD1P3JX baud_counter_i0 (.D(baud_counter_23__N_421[0]), .SP(dac_clk_p_c_enable_413), 
            .PD(baud_counter_23__N_445), .CK(dac_clk_p_c), .Q(baud_counter[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(170[9] 178[37])
    defparam baud_counter_i0.GSR = "DISABLED";
    FD1P3AX data_reg_i0_i0 (.D(data_reg[1]), .SP(data_reg_7__N_416), .CK(dac_clk_p_c), 
            .Q(data_reg[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(143[9] 145[42])
    defparam data_reg_i0_i0.GSR = "DISABLED";
    CCU2D sub_49_add_2_25 (.A0(baud_counter[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n17667), .S0(n290[23]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_25.INIT0 = 16'h5555;
    defparam sub_49_add_2_25.INIT1 = 16'h0000;
    defparam sub_49_add_2_25.INJECT1_0 = "NO";
    defparam sub_49_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_49_add_2_23 (.A0(baud_counter[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17666), .COUT(n17667), .S0(n290[21]), 
          .S1(n290[22]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_23.INIT0 = 16'h5555;
    defparam sub_49_add_2_23.INIT1 = 16'h5555;
    defparam sub_49_add_2_23.INJECT1_0 = "NO";
    defparam sub_49_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_49_add_2_21 (.A0(baud_counter[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17665), .COUT(n17666), .S0(n290[19]), 
          .S1(n290[20]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_21.INIT0 = 16'h5555;
    defparam sub_49_add_2_21.INIT1 = 16'h5555;
    defparam sub_49_add_2_21.INJECT1_0 = "NO";
    defparam sub_49_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_49_add_2_19 (.A0(baud_counter[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17664), .COUT(n17665), .S0(n290[17]), 
          .S1(n290[18]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_19.INIT0 = 16'h5555;
    defparam sub_49_add_2_19.INIT1 = 16'h5555;
    defparam sub_49_add_2_19.INJECT1_0 = "NO";
    defparam sub_49_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_49_add_2_17 (.A0(baud_counter[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17663), .COUT(n17664), .S0(n290[15]), 
          .S1(n290[16]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_17.INIT0 = 16'h5555;
    defparam sub_49_add_2_17.INIT1 = 16'h5555;
    defparam sub_49_add_2_17.INJECT1_0 = "NO";
    defparam sub_49_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_49_add_2_15 (.A0(baud_counter[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17662), .COUT(n17663), .S0(n290[13]), 
          .S1(n290[14]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_15.INIT0 = 16'h5555;
    defparam sub_49_add_2_15.INIT1 = 16'h5555;
    defparam sub_49_add_2_15.INJECT1_0 = "NO";
    defparam sub_49_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_49_add_2_13 (.A0(baud_counter[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17661), .COUT(n17662), .S0(n290[11]), 
          .S1(n290[12]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_13.INIT0 = 16'h5555;
    defparam sub_49_add_2_13.INIT1 = 16'h5555;
    defparam sub_49_add_2_13.INJECT1_0 = "NO";
    defparam sub_49_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_49_add_2_11 (.A0(baud_counter[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17660), .COUT(n17661), .S0(n290[9]), .S1(n290[10]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(178[19:36])
    defparam sub_49_add_2_11.INIT0 = 16'h5555;
    defparam sub_49_add_2_11.INIT1 = 16'h5555;
    defparam sub_49_add_2_11.INJECT1_0 = "NO";
    defparam sub_49_add_2_11.INJECT1_1 = "NO";
    FD1P3AX data_reg_i0_i7 (.D(qq_uart), .SP(data_reg_7__N_416), .CK(dac_clk_p_c), 
            .Q(data_reg[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(143[9] 145[42])
    defparam data_reg_i0_i7.GSR = "DISABLED";
    FD1P3AX data_reg_i0_i6 (.D(data_reg[7]), .SP(data_reg_7__N_416), .CK(dac_clk_p_c), 
            .Q(data_reg[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(143[9] 145[42])
    defparam data_reg_i0_i6.GSR = "DISABLED";
    FD1P3AX data_reg_i0_i5 (.D(data_reg[6]), .SP(data_reg_7__N_416), .CK(dac_clk_p_c), 
            .Q(data_reg[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(143[9] 145[42])
    defparam data_reg_i0_i5.GSR = "DISABLED";
    FD1P3AX data_reg_i0_i4 (.D(data_reg[5]), .SP(data_reg_7__N_416), .CK(dac_clk_p_c), 
            .Q(data_reg[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(143[9] 145[42])
    defparam data_reg_i0_i4.GSR = "DISABLED";
    FD1P3AX data_reg_i0_i3 (.D(data_reg[4]), .SP(data_reg_7__N_416), .CK(dac_clk_p_c), 
            .Q(data_reg[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(143[9] 145[42])
    defparam data_reg_i0_i3.GSR = "DISABLED";
    FD1P3AX data_reg_i0_i2 (.D(data_reg[3]), .SP(data_reg_7__N_416), .CK(dac_clk_p_c), 
            .Q(data_reg[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(143[9] 145[42])
    defparam data_reg_i0_i2.GSR = "DISABLED";
    FD1P3AX data_reg_i0_i1 (.D(data_reg[2]), .SP(data_reg_7__N_416), .CK(dac_clk_p_c), 
            .Q(data_reg[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=57, LSE_RCOL=105, LSE_LLINE=53, LSE_RLINE=53 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/rxuartlite.v(143[9] 145[42])
    defparam data_reg_i0_i1.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module hbbus
//

module hbbus (dac_clk_p_c, wb_we, wb_odata, wb_stb, wb_cyc, wb_err, 
            wb_ack, \wb_idata[0] , wb_addr, \wb_idata[2] , \wb_idata[3] , 
            \wb_idata[4] , \wb_idata[5] , \wb_idata[6] , \wb_idata[7] , 
            \wb_idata[8] , \wb_idata[9] , \wb_idata[10] , \wb_idata[11] , 
            \wb_idata[12] , \wb_idata[13] , \wb_idata[14] , \wb_idata[15] , 
            \wb_idata[16] , \wb_idata[17] , \wb_idata[18] , \wb_idata[19] , 
            \wb_idata[20] , \wb_idata[21] , \wb_idata[22] , \wb_idata[23] , 
            \wb_idata[24] , \wb_idata[25] , \wb_idata[26] , \wb_idata[27] , 
            \wb_idata[28] , \wb_idata[29] , \wb_idata[30] , \wb_idata[31] , 
            n2, GND_net, n12737, n29502, VCC_net, rx_stb, \rx_data[4] , 
            \rx_data[3] , \rx_data[1] , \rx_data[0] , \rx_data[5] , 
            \rx_data[2] , \rx_data[6] , tx_busy, n26910, \lcl_data[1] , 
            \lcl_data_7__N_511[0] , \lcl_data[4] , \lcl_data_7__N_511[3] , 
            \lcl_data[5] , \lcl_data_7__N_511[4] , \lcl_data[6] , \lcl_data_7__N_511[5] , 
            zero_baud_counter, dac_clk_p_c_enable_322, \lcl_data[7] , 
            \lcl_data_7__N_511[6] , \lcl_data[3] , \lcl_data_7__N_511[2] , 
            \lcl_data[2] , \lcl_data_7__N_511[1] , o_busy_N_536, \state[0] , 
            n17844) /* synthesis syn_module_defined=1 */ ;
    input dac_clk_p_c;
    output wb_we;
    output [31:0]wb_odata;
    output wb_stb;
    output wb_cyc;
    input wb_err;
    input wb_ack;
    input \wb_idata[0] ;
    output [29:0]wb_addr;
    input \wb_idata[2] ;
    input \wb_idata[3] ;
    input \wb_idata[4] ;
    input \wb_idata[5] ;
    input \wb_idata[6] ;
    input \wb_idata[7] ;
    input \wb_idata[8] ;
    input \wb_idata[9] ;
    input \wb_idata[10] ;
    input \wb_idata[11] ;
    input \wb_idata[12] ;
    input \wb_idata[13] ;
    input \wb_idata[14] ;
    input \wb_idata[15] ;
    input \wb_idata[16] ;
    input \wb_idata[17] ;
    input \wb_idata[18] ;
    input \wb_idata[19] ;
    input \wb_idata[20] ;
    input \wb_idata[21] ;
    input \wb_idata[22] ;
    input \wb_idata[23] ;
    input \wb_idata[24] ;
    input \wb_idata[25] ;
    input \wb_idata[26] ;
    input \wb_idata[27] ;
    input \wb_idata[28] ;
    input \wb_idata[29] ;
    input \wb_idata[30] ;
    input \wb_idata[31] ;
    output n2;
    input GND_net;
    input n12737;
    input n29502;
    input VCC_net;
    input rx_stb;
    input \rx_data[4] ;
    input \rx_data[3] ;
    input \rx_data[1] ;
    input \rx_data[0] ;
    input \rx_data[5] ;
    input \rx_data[2] ;
    input \rx_data[6] ;
    input tx_busy;
    output n26910;
    input \lcl_data[1] ;
    output \lcl_data_7__N_511[0] ;
    input \lcl_data[4] ;
    output \lcl_data_7__N_511[3] ;
    input \lcl_data[5] ;
    output \lcl_data_7__N_511[4] ;
    input \lcl_data[6] ;
    output \lcl_data_7__N_511[5] ;
    input zero_baud_counter;
    output dac_clk_p_c_enable_322;
    input \lcl_data[7] ;
    output \lcl_data_7__N_511[6] ;
    input \lcl_data[3] ;
    output \lcl_data_7__N_511[2] ;
    input \lcl_data[2] ;
    output \lcl_data_7__N_511[1] ;
    input o_busy_N_536;
    input \state[0] ;
    output n17844;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(28[49:58])
    
    wire inc, dac_clk_p_c_enable_132, i_cmd_wr;
    wire [33:0]iw_word;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(71[14:21])
    
    wire ow_stb;
    wire [33:0]ow_word;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(73[14:21])
    
    wire n29561, n22219, newaddr_N_990, n29560, n17451, n27112, 
        n27111, dac_clk_p_c_enable_446, dac_clk_p_c_enable_308, idl_stb, 
        hb_busy;
    wire [4:0]hb_bits;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(79[13:20])
    
    wire nl_busy, hx_stb;
    wire [33:0]idl_word;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(77[14:22])
    
    wire dac_clk_p_c_enable_194, w_reset, n26906, dac_clk_p_c_enable_381;
    wire [4:0]dec_bits;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(69[13:21])
    
    wire o_pck_stb_N_765, cmd_loaded, dac_clk_p_c_enable_196, cmd_loaded_N_768, 
        dac_clk_p_c_enable_350;
    wire [33:0]n14;
    wire [7:0]w_gx_char;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbgenhex.v(80[12:21])
    
    wire n11749;
    wire [33:0]int_word;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(75[14:22])
    
    wire dac_clk_p_c_enable_416, n12748, n26940, n26903, int_stb;
    
    hbexec wbexec (.inc(inc), .dac_clk_p_c(dac_clk_p_c), .dac_clk_p_c_enable_132(dac_clk_p_c_enable_132), 
           .wb_we(wb_we), .i_cmd_wr(i_cmd_wr), .wb_odata({wb_odata}), 
           .\iw_word[0] (iw_word[0]), .ow_stb(ow_stb), .ow_word({ow_word}), 
           .n29561(n29561), .wb_stb(wb_stb), .n22219(n22219), .wb_cyc(wb_cyc), 
           .newaddr_N_990(newaddr_N_990), .\iw_word[31] (iw_word[31]), .wb_err(wb_err), 
           .n29560(n29560), .wb_ack(wb_ack), .\wb_idata[0] (\wb_idata[0] ), 
           .wb_addr({wb_addr}), .\wb_idata[2] (\wb_idata[2] ), .\wb_idata[3] (\wb_idata[3] ), 
           .\wb_idata[4] (\wb_idata[4] ), .\wb_idata[5] (\wb_idata[5] ), 
           .\wb_idata[6] (\wb_idata[6] ), .\wb_idata[7] (\wb_idata[7] ), 
           .\wb_idata[8] (\wb_idata[8] ), .\wb_idata[9] (\wb_idata[9] ), 
           .\wb_idata[10] (\wb_idata[10] ), .\wb_idata[11] (\wb_idata[11] ), 
           .\wb_idata[12] (\wb_idata[12] ), .\wb_idata[13] (\wb_idata[13] ), 
           .\wb_idata[14] (\wb_idata[14] ), .\wb_idata[15] (\wb_idata[15] ), 
           .\wb_idata[16] (\wb_idata[16] ), .\iw_word[30] (iw_word[30]), 
           .\iw_word[29] (iw_word[29]), .\iw_word[28] (iw_word[28]), .\wb_idata[17] (\wb_idata[17] ), 
           .\iw_word[27] (iw_word[27]), .\iw_word[26] (iw_word[26]), .\iw_word[25] (iw_word[25]), 
           .\iw_word[24] (iw_word[24]), .\iw_word[23] (iw_word[23]), .\iw_word[22] (iw_word[22]), 
           .\iw_word[21] (iw_word[21]), .\iw_word[20] (iw_word[20]), .\iw_word[19] (iw_word[19]), 
           .\iw_word[18] (iw_word[18]), .\iw_word[17] (iw_word[17]), .\iw_word[16] (iw_word[16]), 
           .\iw_word[15] (iw_word[15]), .\iw_word[14] (iw_word[14]), .\iw_word[13] (iw_word[13]), 
           .\iw_word[12] (iw_word[12]), .\iw_word[11] (iw_word[11]), .\iw_word[10] (iw_word[10]), 
           .\iw_word[9] (iw_word[9]), .\iw_word[8] (iw_word[8]), .\iw_word[7] (iw_word[7]), 
           .\wb_idata[18] (\wb_idata[18] ), .\iw_word[6] (iw_word[6]), .\iw_word[5] (iw_word[5]), 
           .\iw_word[4] (iw_word[4]), .\iw_word[3] (iw_word[3]), .\iw_word[2] (iw_word[2]), 
           .\iw_word[1] (iw_word[1]), .\wb_idata[19] (\wb_idata[19] ), .\wb_idata[20] (\wb_idata[20] ), 
           .\wb_idata[21] (\wb_idata[21] ), .\wb_idata[22] (\wb_idata[22] ), 
           .\wb_idata[23] (\wb_idata[23] ), .\wb_idata[24] (\wb_idata[24] ), 
           .\wb_idata[25] (\wb_idata[25] ), .\wb_idata[26] (\wb_idata[26] ), 
           .\wb_idata[27] (\wb_idata[27] ), .\wb_idata[28] (\wb_idata[28] ), 
           .\wb_idata[29] (\wb_idata[29] ), .\wb_idata[30] (\wb_idata[30] ), 
           .\wb_idata[31] (\wb_idata[31] ), .n2(n2), .n17451(n17451), 
           .GND_net(GND_net), .n27112(n27112), .\iw_word[32] (iw_word[32]), 
           .n27111(n27111), .n12737(n12737), .dac_clk_p_c_enable_446(dac_clk_p_c_enable_446)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(105[15] 109[15])
    hbdeword unpackx (.dac_clk_p_c(dac_clk_p_c), .dac_clk_p_c_enable_308(dac_clk_p_c_enable_308), 
            .idl_stb(idl_stb), .hb_busy(hb_busy), .hb_bits({hb_bits}), 
            .n29560(n29560), .nl_busy(nl_busy), .hx_stb(hx_stb), .idl_word({idl_word}), 
            .dac_clk_p_c_enable_194(dac_clk_p_c_enable_194), .n29561(n29561), 
            .n29502(n29502), .w_reset(w_reset), .n26906(n26906)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(127[11] 129[29])
    hbpack packxi (.dac_clk_p_c(dac_clk_p_c), .dac_clk_p_c_enable_381(dac_clk_p_c_enable_381), 
           .n29561(n29561), .iw_word({Open_0, Open_1, Open_2, Open_3, 
           Open_4, Open_5, Open_6, Open_7, Open_8, Open_9, Open_10, 
           Open_11, Open_12, Open_13, Open_14, Open_15, Open_16, 
           Open_17, Open_18, Open_19, Open_20, Open_21, Open_22, 
           Open_23, Open_24, Open_25, Open_26, Open_27, Open_28, 
           Open_29, Open_30, iw_word[2], Open_31, iw_word[0]}), .\dec_bits[4] (dec_bits[4]), 
           .w_reset(w_reset), .o_pck_stb_N_765(o_pck_stb_N_765), .cmd_loaded(cmd_loaded), 
           .dac_clk_p_c_enable_196(dac_clk_p_c_enable_196), .cmd_loaded_N_768(cmd_loaded_N_768), 
           .\dec_bits[1] (dec_bits[1]), .wb_cyc(wb_cyc), .inc(inc), .n17451(n17451), 
           .\iw_word[32] (iw_word[32]), .\iw_word[31] (iw_word[31]), .\iw_word[30] (iw_word[30]), 
           .\iw_word[29] (iw_word[29]), .\iw_word[28] (iw_word[28]), .\iw_word[27] (iw_word[27]), 
           .\iw_word[26] (iw_word[26]), .\iw_word[25] (iw_word[25]), .\iw_word[24] (iw_word[24]), 
           .\iw_word[23] (iw_word[23]), .\iw_word[22] (iw_word[22]), .\iw_word[21] (iw_word[21]), 
           .\iw_word[20] (iw_word[20]), .\iw_word[19] (iw_word[19]), .\iw_word[18] (iw_word[18]), 
           .\iw_word[17] (iw_word[17]), .\iw_word[16] (iw_word[16]), .\iw_word[15] (iw_word[15]), 
           .\iw_word[14] (iw_word[14]), .\iw_word[13] (iw_word[13]), .\iw_word[12] (iw_word[12]), 
           .\iw_word[11] (iw_word[11]), .\iw_word[10] (iw_word[10]), .\iw_word[9] (iw_word[9]), 
           .\iw_word[8] (iw_word[8]), .\iw_word[7] (iw_word[7]), .\iw_word[6] (iw_word[6]), 
           .\iw_word[5] (iw_word[5]), .\iw_word[4] (iw_word[4]), .\iw_word[3] (iw_word[3]), 
           .\iw_word[1] (iw_word[1]), .n27111(n27111), .i_cmd_wr(i_cmd_wr), 
           .wb_stb(wb_stb), .n22219(n22219), .n27112(n27112), .dac_clk_p_c_enable_132(dac_clk_p_c_enable_132), 
           .n29560(n29560), .newaddr_N_990(newaddr_N_990), .\dec_bits[0] (dec_bits[0]), 
           .dac_clk_p_c_enable_350(dac_clk_p_c_enable_350), .n45(n14[3]), 
           .n46(n14[2]), .dac_clk_p_c_enable_446(dac_clk_p_c_enable_446)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(99[9] 100[38])
    hbgenhex genhex (.hb_bits({hb_bits}), .\w_gx_char[0] (w_gx_char[0]), 
            .\w_gx_char[1] (w_gx_char[1]), .\w_gx_char[2] (w_gx_char[2]), 
            .\w_gx_char[3] (w_gx_char[3]), .\w_gx_char[4] (w_gx_char[4]), 
            .\w_gx_char[5] (w_gx_char[5]), .\w_gx_char[6] (w_gx_char[6]), 
            .dac_clk_p_c(dac_clk_p_c), .dac_clk_p_c_enable_308(dac_clk_p_c_enable_308), 
            .GND_net(GND_net), .VCC_net(VCC_net), .hx_stb(hx_stb), .w_reset(w_reset), 
            .hb_busy(hb_busy), .nl_busy(nl_busy), .n29560(n29560), .n26906(n26906), 
            .dac_clk_p_c_enable_194(dac_clk_p_c_enable_194), .n11749(n11749)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(132[11] 133[29])
    hbdechex dechxi (.dac_clk_p_c(dac_clk_p_c), .dec_bits({dec_bits[4], 
            Open_32, Open_33, Open_34, dec_bits[0]}), .w_reset(w_reset), 
            .rx_stb(rx_stb), .\rx_data[4] (\rx_data[4] ), .\rx_data[3] (\rx_data[3] ), 
            .\rx_data[1] (\rx_data[1] ), .\rx_data[0] (\rx_data[0] ), .\rx_data[5] (\rx_data[5] ), 
            .n45(n14[3]), .n46(n14[2]), .\dec_bits[1] (dec_bits[1]), .\rx_data[2] (\rx_data[2] ), 
            .\rx_data[6] (\rx_data[6] ), .n29561(n29561), .n29560(n29560), 
            .dac_clk_p_c_enable_381(dac_clk_p_c_enable_381), .dac_clk_p_c_enable_350(dac_clk_p_c_enable_350), 
            .cmd_loaded(cmd_loaded), .o_pck_stb_N_765(o_pck_stb_N_765), 
            .dac_clk_p_c_enable_196(dac_clk_p_c_enable_196), .cmd_loaded_N_768(cmd_loaded_N_768)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(93[11] 95[30])
    hbnewline addnl (.hx_stb(hx_stb), .nl_busy(nl_busy), .\w_gx_char[5] (w_gx_char[5]), 
            .dac_clk_p_c(dac_clk_p_c), .n29561(n29561), .\w_gx_char[1] (w_gx_char[1]), 
            .\w_gx_char[6] (w_gx_char[6]), .n11749(n11749), .tx_busy(tx_busy), 
            .n26910(n26910), .\lcl_data[1] (\lcl_data[1] ), .\lcl_data_7__N_511[0] (\lcl_data_7__N_511[0] ), 
            .\lcl_data[4] (\lcl_data[4] ), .\lcl_data_7__N_511[3] (\lcl_data_7__N_511[3] ), 
            .w_reset(w_reset), .\lcl_data[5] (\lcl_data[5] ), .\lcl_data_7__N_511[4] (\lcl_data_7__N_511[4] ), 
            .\lcl_data[6] (\lcl_data[6] ), .\lcl_data_7__N_511[5] (\lcl_data_7__N_511[5] ), 
            .zero_baud_counter(zero_baud_counter), .dac_clk_p_c_enable_322(dac_clk_p_c_enable_322), 
            .\lcl_data[7] (\lcl_data[7] ), .\lcl_data_7__N_511[6] (\lcl_data_7__N_511[6] ), 
            .\lcl_data[3] (\lcl_data[3] ), .\lcl_data_7__N_511[2] (\lcl_data_7__N_511[2] ), 
            .\lcl_data[2] (\lcl_data[2] ), .\lcl_data_7__N_511[1] (\lcl_data_7__N_511[1] ), 
            .o_busy_N_536(o_busy_N_536), .\state[0] (\state[0] ), .n17844(n17844), 
            .\w_gx_char[2] (w_gx_char[2]), .\w_gx_char[0] (w_gx_char[0]), 
            .\w_gx_char[4] (w_gx_char[4]), .n29560(n29560), .\w_gx_char[3] (w_gx_char[3])) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(138[12] 139[40])
    hbints addints (.int_word({int_word}), .dac_clk_p_c(dac_clk_p_c), .dac_clk_p_c_enable_416(dac_clk_p_c_enable_416), 
           .n12748(n12748), .ow_word({ow_word}), .n29560(n29560), .n26940(n26940), 
           .n26903(n26903), .int_stb(int_stb), .ow_stb(ow_stb), .n29561(n29561)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(114[9] 116[32])
    hbidle addidles (.idl_word({idl_word}), .dac_clk_p_c(dac_clk_p_c), .int_word({int_word}), 
           .idl_stb(idl_stb), .w_reset(w_reset), .hb_busy(hb_busy), .n26903(n26903), 
           .int_stb(int_stb), .n29560(n29560), .n26940(n26940), .n12748(n12748), 
           .dac_clk_p_c_enable_416(dac_clk_p_c_enable_416)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(121[9] 123[31])
    
endmodule
//
// Verilog Description of module hbexec
//

module hbexec (inc, dac_clk_p_c, dac_clk_p_c_enable_132, wb_we, i_cmd_wr, 
            wb_odata, \iw_word[0] , ow_stb, ow_word, n29561, wb_stb, 
            n22219, wb_cyc, newaddr_N_990, \iw_word[31] , wb_err, 
            n29560, wb_ack, \wb_idata[0] , wb_addr, \wb_idata[2] , 
            \wb_idata[3] , \wb_idata[4] , \wb_idata[5] , \wb_idata[6] , 
            \wb_idata[7] , \wb_idata[8] , \wb_idata[9] , \wb_idata[10] , 
            \wb_idata[11] , \wb_idata[12] , \wb_idata[13] , \wb_idata[14] , 
            \wb_idata[15] , \wb_idata[16] , \iw_word[30] , \iw_word[29] , 
            \iw_word[28] , \wb_idata[17] , \iw_word[27] , \iw_word[26] , 
            \iw_word[25] , \iw_word[24] , \iw_word[23] , \iw_word[22] , 
            \iw_word[21] , \iw_word[20] , \iw_word[19] , \iw_word[18] , 
            \iw_word[17] , \iw_word[16] , \iw_word[15] , \iw_word[14] , 
            \iw_word[13] , \iw_word[12] , \iw_word[11] , \iw_word[10] , 
            \iw_word[9] , \iw_word[8] , \iw_word[7] , \wb_idata[18] , 
            \iw_word[6] , \iw_word[5] , \iw_word[4] , \iw_word[3] , 
            \iw_word[2] , \iw_word[1] , \wb_idata[19] , \wb_idata[20] , 
            \wb_idata[21] , \wb_idata[22] , \wb_idata[23] , \wb_idata[24] , 
            \wb_idata[25] , \wb_idata[26] , \wb_idata[27] , \wb_idata[28] , 
            \wb_idata[29] , \wb_idata[30] , \wb_idata[31] , n2, n17451, 
            GND_net, n27112, \iw_word[32] , n27111, n12737, dac_clk_p_c_enable_446) /* synthesis syn_module_defined=1 */ ;
    output inc;
    input dac_clk_p_c;
    input dac_clk_p_c_enable_132;
    output wb_we;
    input i_cmd_wr;
    output [31:0]wb_odata;
    input \iw_word[0] ;
    output ow_stb;
    output [33:0]ow_word;
    input n29561;
    output wb_stb;
    input n22219;
    output wb_cyc;
    input newaddr_N_990;
    input \iw_word[31] ;
    input wb_err;
    input n29560;
    input wb_ack;
    input \wb_idata[0] ;
    output [29:0]wb_addr;
    input \wb_idata[2] ;
    input \wb_idata[3] ;
    input \wb_idata[4] ;
    input \wb_idata[5] ;
    input \wb_idata[6] ;
    input \wb_idata[7] ;
    input \wb_idata[8] ;
    input \wb_idata[9] ;
    input \wb_idata[10] ;
    input \wb_idata[11] ;
    input \wb_idata[12] ;
    input \wb_idata[13] ;
    input \wb_idata[14] ;
    input \wb_idata[15] ;
    input \wb_idata[16] ;
    input \iw_word[30] ;
    input \iw_word[29] ;
    input \iw_word[28] ;
    input \wb_idata[17] ;
    input \iw_word[27] ;
    input \iw_word[26] ;
    input \iw_word[25] ;
    input \iw_word[24] ;
    input \iw_word[23] ;
    input \iw_word[22] ;
    input \iw_word[21] ;
    input \iw_word[20] ;
    input \iw_word[19] ;
    input \iw_word[18] ;
    input \iw_word[17] ;
    input \iw_word[16] ;
    input \iw_word[15] ;
    input \iw_word[14] ;
    input \iw_word[13] ;
    input \iw_word[12] ;
    input \iw_word[11] ;
    input \iw_word[10] ;
    input \iw_word[9] ;
    input \iw_word[8] ;
    input \iw_word[7] ;
    input \wb_idata[18] ;
    input \iw_word[6] ;
    input \iw_word[5] ;
    input \iw_word[4] ;
    input \iw_word[3] ;
    input \iw_word[2] ;
    input \iw_word[1] ;
    input \wb_idata[19] ;
    input \wb_idata[20] ;
    input \wb_idata[21] ;
    input \wb_idata[22] ;
    input \wb_idata[23] ;
    input \wb_idata[24] ;
    input \wb_idata[25] ;
    input \wb_idata[26] ;
    input \wb_idata[27] ;
    input \wb_idata[28] ;
    input \wb_idata[29] ;
    input \wb_idata[30] ;
    input \wb_idata[31] ;
    output n2;
    input n17451;
    input GND_net;
    input n27112;
    input \iw_word[32] ;
    input n27111;
    input n12737;
    input dac_clk_p_c_enable_446;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(28[49:58])
    
    wire i_cmd_word_0__N_995, o_cmd_busy_N_931, n9018, o_rsp_stb_N_987;
    wire [33:0]n338;
    wire [33:0]o_rsp_word_33__N_951;
    
    wire n19812, newaddr;
    wire [32:0]n2249;
    
    wire n17709, n17396, n17394;
    wire [29:0]n125;
    
    wire n17708, n17400, n17398, n17707, n17404, n17402, n17706, 
        n17408, n17406, n17705, n17412, n17410, n17704, n17416, 
        n17414, n17703, n17420, n17418, n17702, n17424, n17422, 
        n17701, n17428, n17426, n17700, n17432, n17430, n17699, 
        n17436, n17434, n17698, n17440, n17438, n17697, n17444, 
        n17442, n17696, n17448, n17446, n17695, n17450, n3, n20476, 
        o_cmd_busy_N_941, o_cmd_busy_N_933, dac_clk_p_c_enable_415;
    
    FD1P3AX inc_71 (.D(i_cmd_word_0__N_995), .SP(dac_clk_p_c_enable_132), 
            .CK(dac_clk_p_c), .Q(inc)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(192[9] 236[5])
    defparam inc_71.GSR = "DISABLED";
    FD1P3AX o_wb_we_69 (.D(i_cmd_wr), .SP(o_cmd_busy_N_931), .CK(dac_clk_p_c), 
            .Q(wb_we)) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(184[9] 186[26])
    defparam o_wb_we_69.GSR = "DISABLED";
    FD1S3AX o_wb_data_i0 (.D(\iw_word[0] ), .CK(dac_clk_p_c), .Q(wb_odata[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i0.GSR = "DISABLED";
    FD1S3JX o_rsp_stb_74 (.D(o_rsp_stb_N_987), .CK(dac_clk_p_c), .PD(n9018), 
            .Q(ow_stb)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_stb_74.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i0 (.D(n338[0]), .CK(dac_clk_p_c), .CD(n9018), 
            .Q(ow_word[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i0.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i2 (.D(n338[2]), .CK(dac_clk_p_c), .CD(n9018), 
            .Q(ow_word[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i2.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i3 (.D(n338[3]), .CK(dac_clk_p_c), .CD(n9018), 
            .Q(ow_word[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i3.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i4 (.D(n338[4]), .CK(dac_clk_p_c), .CD(n9018), 
            .Q(ow_word[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i4.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i5 (.D(n338[5]), .CK(dac_clk_p_c), .CD(n9018), 
            .Q(ow_word[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i5.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i6 (.D(n338[6]), .CK(dac_clk_p_c), .CD(n9018), 
            .Q(ow_word[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i6.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i7 (.D(n338[7]), .CK(dac_clk_p_c), .CD(n9018), 
            .Q(ow_word[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i7.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i8 (.D(n338[8]), .CK(dac_clk_p_c), .CD(n9018), 
            .Q(ow_word[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i8.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i9 (.D(n338[9]), .CK(dac_clk_p_c), .CD(n9018), 
            .Q(ow_word[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i9.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i10 (.D(n338[10]), .CK(dac_clk_p_c), .CD(n9018), 
            .Q(ow_word[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i10.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i11 (.D(n338[11]), .CK(dac_clk_p_c), .CD(n9018), 
            .Q(ow_word[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i11.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i12 (.D(n338[12]), .CK(dac_clk_p_c), .CD(n9018), 
            .Q(ow_word[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i12.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i13 (.D(n338[13]), .CK(dac_clk_p_c), .CD(n9018), 
            .Q(ow_word[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i13.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i14 (.D(n338[14]), .CK(dac_clk_p_c), .CD(n9018), 
            .Q(ow_word[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i14.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i15 (.D(n338[15]), .CK(dac_clk_p_c), .CD(n9018), 
            .Q(ow_word[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i15.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i16 (.D(n338[16]), .CK(dac_clk_p_c), .CD(n9018), 
            .Q(ow_word[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i16.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i17 (.D(n338[17]), .CK(dac_clk_p_c), .CD(n9018), 
            .Q(ow_word[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i17.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i18 (.D(n338[18]), .CK(dac_clk_p_c), .CD(n9018), 
            .Q(ow_word[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i18.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i19 (.D(n338[19]), .CK(dac_clk_p_c), .CD(n9018), 
            .Q(ow_word[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i19.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i20 (.D(n338[20]), .CK(dac_clk_p_c), .CD(n9018), 
            .Q(ow_word[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i20.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i21 (.D(n338[21]), .CK(dac_clk_p_c), .CD(n9018), 
            .Q(ow_word[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i21.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i22 (.D(n338[22]), .CK(dac_clk_p_c), .CD(n9018), 
            .Q(ow_word[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i22.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i23 (.D(n338[23]), .CK(dac_clk_p_c), .CD(n9018), 
            .Q(ow_word[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i23.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i24 (.D(n338[24]), .CK(dac_clk_p_c), .CD(n9018), 
            .Q(ow_word[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i24.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i25 (.D(n338[25]), .CK(dac_clk_p_c), .CD(n9018), 
            .Q(ow_word[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i25.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i26 (.D(n338[26]), .CK(dac_clk_p_c), .CD(n9018), 
            .Q(ow_word[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i26.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i27 (.D(n338[27]), .CK(dac_clk_p_c), .CD(n9018), 
            .Q(ow_word[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i27.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i28 (.D(n338[28]), .CK(dac_clk_p_c), .CD(n9018), 
            .Q(ow_word[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i28.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i29 (.D(o_rsp_word_33__N_951[29]), .CK(dac_clk_p_c), 
            .CD(n29561), .Q(ow_word[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i29.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i30 (.D(n338[30]), .CK(dac_clk_p_c), .CD(n9018), 
            .Q(ow_word[30])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i30.GSR = "DISABLED";
    FD1S3IX o_rsp_word_i31 (.D(n338[31]), .CK(dac_clk_p_c), .CD(n9018), 
            .Q(ow_word[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i31.GSR = "DISABLED";
    FD1S3JX o_rsp_word_i32 (.D(n338[32]), .CK(dac_clk_p_c), .PD(n9018), 
            .Q(ow_word[32])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i32.GSR = "DISABLED";
    FD1S3JX o_rsp_word_i33 (.D(o_cmd_busy_N_931), .CK(dac_clk_p_c), .PD(n9018), 
            .Q(ow_word[33])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i33.GSR = "DISABLED";
    FD1P3IX o_wb_stb_68 (.D(n22219), .SP(o_cmd_busy_N_931), .CD(n19812), 
            .CK(dac_clk_p_c), .Q(wb_stb)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(121[9] 168[5])
    defparam o_wb_stb_68.GSR = "DISABLED";
    FD1S3IX newaddr_72 (.D(newaddr_N_990), .CK(dac_clk_p_c), .CD(wb_cyc), 
            .Q(newaddr)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(192[9] 236[5])
    defparam newaddr_72.GSR = "DISABLED";
    FD1S3AX o_wb_data_i31 (.D(\iw_word[31] ), .CK(dac_clk_p_c), .Q(wb_odata[31])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i31.GSR = "DISABLED";
    LUT4 i_cmd_word_0__I_0_1_lut (.A(\iw_word[0] ), .Z(i_cmd_word_0__N_995)) /* synthesis lut_function=(!(A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(214[11:25])
    defparam i_cmd_word_0__I_0_1_lut.init = 16'h5555;
    LUT4 o_cmd_busy_I_0_1_lut (.A(wb_cyc), .Z(o_cmd_busy_N_931)) /* synthesis lut_function=(!(A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(194[21:34])
    defparam o_cmd_busy_I_0_1_lut.init = 16'h5555;
    LUT4 i6522_2_lut (.A(wb_err), .B(n29560), .Z(n9018)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(283[11] 309[5])
    defparam i6522_2_lut.init = 16'heeee;
    LUT4 newaddr_I_0_3_lut (.A(newaddr), .B(wb_ack), .C(wb_cyc), .Z(o_rsp_stb_N_987)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam newaddr_I_0_3_lut.init = 16'hcaca;
    LUT4 mux_59_i1_4_lut (.A(inc), .B(\wb_idata[0] ), .C(wb_cyc), .D(wb_we), 
         .Z(n338[0])) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A (B (C (D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i1_4_lut.init = 16'h05c5;
    LUT4 mux_59_i3_4_lut (.A(wb_addr[0]), .B(\wb_idata[2] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[2])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i3_4_lut.init = 16'h0aca;
    LUT4 mux_59_i4_4_lut (.A(wb_addr[1]), .B(\wb_idata[3] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[3])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i4_4_lut.init = 16'h0aca;
    LUT4 mux_59_i5_4_lut (.A(wb_addr[2]), .B(\wb_idata[4] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[4])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i5_4_lut.init = 16'h0aca;
    LUT4 mux_59_i6_4_lut (.A(wb_addr[3]), .B(\wb_idata[5] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[5])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i6_4_lut.init = 16'h0aca;
    LUT4 mux_59_i7_4_lut (.A(wb_addr[4]), .B(\wb_idata[6] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[6])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i7_4_lut.init = 16'h0aca;
    LUT4 mux_59_i8_4_lut (.A(wb_addr[5]), .B(\wb_idata[7] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[7])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i8_4_lut.init = 16'h0aca;
    LUT4 mux_59_i9_4_lut (.A(wb_addr[6]), .B(\wb_idata[8] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[8])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i9_4_lut.init = 16'h0aca;
    LUT4 mux_59_i10_4_lut (.A(wb_addr[7]), .B(\wb_idata[9] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[9])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i10_4_lut.init = 16'h0aca;
    LUT4 mux_59_i11_4_lut (.A(wb_addr[8]), .B(\wb_idata[10] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[10])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i11_4_lut.init = 16'h0aca;
    LUT4 mux_59_i12_4_lut (.A(wb_addr[9]), .B(\wb_idata[11] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[11])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i12_4_lut.init = 16'h0aca;
    LUT4 mux_59_i13_4_lut (.A(wb_addr[10]), .B(\wb_idata[12] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[12])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i13_4_lut.init = 16'h0aca;
    LUT4 mux_59_i14_4_lut (.A(wb_addr[11]), .B(\wb_idata[13] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[13])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i14_4_lut.init = 16'h0aca;
    LUT4 mux_59_i15_4_lut (.A(wb_addr[12]), .B(\wb_idata[14] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[14])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i15_4_lut.init = 16'h0aca;
    LUT4 mux_59_i16_4_lut (.A(wb_addr[13]), .B(\wb_idata[15] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[15])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i16_4_lut.init = 16'h0aca;
    LUT4 mux_59_i17_4_lut (.A(wb_addr[14]), .B(\wb_idata[16] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[16])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i17_4_lut.init = 16'h0aca;
    FD1S3AX o_wb_data_i30 (.D(\iw_word[30] ), .CK(dac_clk_p_c), .Q(wb_odata[30])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i30.GSR = "DISABLED";
    FD1S3AX o_wb_data_i29 (.D(\iw_word[29] ), .CK(dac_clk_p_c), .Q(wb_odata[29])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i29.GSR = "DISABLED";
    FD1S3AX o_wb_data_i28 (.D(\iw_word[28] ), .CK(dac_clk_p_c), .Q(wb_odata[28])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i28.GSR = "DISABLED";
    LUT4 mux_59_i18_4_lut (.A(wb_addr[15]), .B(\wb_idata[17] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[17])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i18_4_lut.init = 16'h0aca;
    FD1S3AX o_wb_data_i27 (.D(\iw_word[27] ), .CK(dac_clk_p_c), .Q(wb_odata[27])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i27.GSR = "DISABLED";
    FD1S3AX o_wb_data_i26 (.D(\iw_word[26] ), .CK(dac_clk_p_c), .Q(wb_odata[26])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i26.GSR = "DISABLED";
    FD1S3AX o_wb_data_i25 (.D(\iw_word[25] ), .CK(dac_clk_p_c), .Q(wb_odata[25])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i25.GSR = "DISABLED";
    FD1S3AX o_wb_data_i24 (.D(\iw_word[24] ), .CK(dac_clk_p_c), .Q(wb_odata[24])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i24.GSR = "DISABLED";
    FD1S3AX o_wb_data_i23 (.D(\iw_word[23] ), .CK(dac_clk_p_c), .Q(wb_odata[23])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i23.GSR = "DISABLED";
    FD1S3AX o_wb_data_i22 (.D(\iw_word[22] ), .CK(dac_clk_p_c), .Q(wb_odata[22])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i22.GSR = "DISABLED";
    FD1S3AX o_wb_data_i21 (.D(\iw_word[21] ), .CK(dac_clk_p_c), .Q(wb_odata[21])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i21.GSR = "DISABLED";
    FD1S3AX o_wb_data_i20 (.D(\iw_word[20] ), .CK(dac_clk_p_c), .Q(wb_odata[20])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i20.GSR = "DISABLED";
    FD1S3AX o_wb_data_i19 (.D(\iw_word[19] ), .CK(dac_clk_p_c), .Q(wb_odata[19])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i19.GSR = "DISABLED";
    FD1S3AX o_wb_data_i18 (.D(\iw_word[18] ), .CK(dac_clk_p_c), .Q(wb_odata[18])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i18.GSR = "DISABLED";
    FD1S3AX o_wb_data_i17 (.D(\iw_word[17] ), .CK(dac_clk_p_c), .Q(wb_odata[17])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i17.GSR = "DISABLED";
    FD1S3AX o_wb_data_i16 (.D(\iw_word[16] ), .CK(dac_clk_p_c), .Q(wb_odata[16])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i16.GSR = "DISABLED";
    FD1S3AX o_wb_data_i15 (.D(\iw_word[15] ), .CK(dac_clk_p_c), .Q(wb_odata[15])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i15.GSR = "DISABLED";
    FD1S3AX o_wb_data_i14 (.D(\iw_word[14] ), .CK(dac_clk_p_c), .Q(wb_odata[14])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i14.GSR = "DISABLED";
    FD1S3AX o_wb_data_i13 (.D(\iw_word[13] ), .CK(dac_clk_p_c), .Q(wb_odata[13])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i13.GSR = "DISABLED";
    FD1S3AX o_wb_data_i12 (.D(\iw_word[12] ), .CK(dac_clk_p_c), .Q(wb_odata[12])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i12.GSR = "DISABLED";
    FD1S3AX o_wb_data_i11 (.D(\iw_word[11] ), .CK(dac_clk_p_c), .Q(wb_odata[11])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i11.GSR = "DISABLED";
    FD1S3AX o_wb_data_i10 (.D(\iw_word[10] ), .CK(dac_clk_p_c), .Q(wb_odata[10])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i10.GSR = "DISABLED";
    FD1S3AX o_wb_data_i9 (.D(\iw_word[9] ), .CK(dac_clk_p_c), .Q(wb_odata[9])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i9.GSR = "DISABLED";
    FD1S3AX o_wb_data_i8 (.D(\iw_word[8] ), .CK(dac_clk_p_c), .Q(wb_odata[8])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i8.GSR = "DISABLED";
    FD1S3AX o_wb_data_i7 (.D(\iw_word[7] ), .CK(dac_clk_p_c), .Q(wb_odata[7])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i7.GSR = "DISABLED";
    LUT4 mux_59_i19_4_lut (.A(wb_addr[16]), .B(\wb_idata[18] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[18])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i19_4_lut.init = 16'h0aca;
    FD1S3AX o_wb_data_i6 (.D(\iw_word[6] ), .CK(dac_clk_p_c), .Q(wb_odata[6])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i6.GSR = "DISABLED";
    FD1S3AX o_wb_data_i5 (.D(\iw_word[5] ), .CK(dac_clk_p_c), .Q(wb_odata[5])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i5.GSR = "DISABLED";
    FD1S3AX o_wb_data_i4 (.D(\iw_word[4] ), .CK(dac_clk_p_c), .Q(wb_odata[4])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i4.GSR = "DISABLED";
    FD1S3AX o_wb_data_i3 (.D(\iw_word[3] ), .CK(dac_clk_p_c), .Q(wb_odata[3])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i3.GSR = "DISABLED";
    FD1S3AX o_wb_data_i2 (.D(\iw_word[2] ), .CK(dac_clk_p_c), .Q(wb_odata[2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i2.GSR = "DISABLED";
    FD1S3AX o_wb_data_i1 (.D(\iw_word[1] ), .CK(dac_clk_p_c), .Q(wb_odata[1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(241[9] 261[5])
    defparam o_wb_data_i1.GSR = "DISABLED";
    LUT4 mux_59_i20_4_lut (.A(wb_addr[17]), .B(\wb_idata[19] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[19])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i20_4_lut.init = 16'h0aca;
    LUT4 mux_59_i21_4_lut (.A(wb_addr[18]), .B(\wb_idata[20] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[20])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i21_4_lut.init = 16'h0aca;
    LUT4 mux_59_i22_4_lut (.A(wb_addr[19]), .B(\wb_idata[21] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[21])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i22_4_lut.init = 16'h0aca;
    LUT4 mux_59_i23_4_lut (.A(wb_addr[20]), .B(\wb_idata[22] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[22])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i23_4_lut.init = 16'h0aca;
    LUT4 mux_59_i24_4_lut (.A(wb_addr[21]), .B(\wb_idata[23] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[23])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i24_4_lut.init = 16'h0aca;
    LUT4 mux_59_i25_4_lut (.A(wb_addr[22]), .B(\wb_idata[24] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[24])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i25_4_lut.init = 16'h0aca;
    LUT4 mux_59_i26_4_lut (.A(wb_addr[23]), .B(\wb_idata[25] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[25])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i26_4_lut.init = 16'h0aca;
    LUT4 mux_59_i27_4_lut (.A(wb_addr[24]), .B(\wb_idata[26] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[26])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i27_4_lut.init = 16'h0aca;
    LUT4 mux_59_i28_4_lut (.A(wb_addr[25]), .B(\wb_idata[27] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[27])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i28_4_lut.init = 16'h0aca;
    LUT4 mux_59_i29_4_lut (.A(wb_addr[26]), .B(\wb_idata[28] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[28])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i29_4_lut.init = 16'h0aca;
    LUT4 i11277_4_lut (.A(wb_addr[27]), .B(wb_err), .C(n2249[29]), .D(wb_cyc), 
         .Z(o_rsp_word_33__N_951[29])) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(287[11] 309[5])
    defparam i11277_4_lut.init = 16'hfcee;
    LUT4 i11325_2_lut (.A(\wb_idata[29] ), .B(wb_we), .Z(n2249[29])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(299[4:47])
    defparam i11325_2_lut.init = 16'h2222;
    LUT4 mux_59_i31_4_lut (.A(wb_addr[28]), .B(\wb_idata[30] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[30])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i31_4_lut.init = 16'h0aca;
    LUT4 mux_59_i32_4_lut (.A(wb_addr[29]), .B(\wb_idata[31] ), .C(wb_cyc), 
         .D(wb_we), .Z(n338[31])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam mux_59_i32_4_lut.init = 16'h0aca;
    LUT4 i11285_2_lut (.A(wb_we), .B(wb_cyc), .Z(n338[32])) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(300[11] 309[5])
    defparam i11285_2_lut.init = 16'h8888;
    LUT4 i2_1_lut (.A(wb_stb), .Z(n2)) /* synthesis lut_function=(!(A)) */ ;
    defparam i2_1_lut.init = 16'h5555;
    CCU2D o_wb_addr_548_add_4_31 (.A0(n17396), .B0(\iw_word[1] ), .C0(dac_clk_p_c_enable_132), 
          .D0(\iw_word[30] ), .A1(n17394), .B1(\iw_word[1] ), .C1(dac_clk_p_c_enable_132), 
          .D1(\iw_word[31] ), .CIN(n17709), .S0(n125[28]), .S1(n125[29]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_548_add_4_31.INIT0 = 16'h5aaa;
    defparam o_wb_addr_548_add_4_31.INIT1 = 16'h5aaa;
    defparam o_wb_addr_548_add_4_31.INJECT1_0 = "NO";
    defparam o_wb_addr_548_add_4_31.INJECT1_1 = "NO";
    CCU2D o_wb_addr_548_add_4_29 (.A0(n17400), .B0(\iw_word[1] ), .C0(dac_clk_p_c_enable_132), 
          .D0(\iw_word[28] ), .A1(n17398), .B1(\iw_word[1] ), .C1(dac_clk_p_c_enable_132), 
          .D1(\iw_word[29] ), .CIN(n17708), .COUT(n17709), .S0(n125[26]), 
          .S1(n125[27]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_548_add_4_29.INIT0 = 16'h5aaa;
    defparam o_wb_addr_548_add_4_29.INIT1 = 16'h5aaa;
    defparam o_wb_addr_548_add_4_29.INJECT1_0 = "NO";
    defparam o_wb_addr_548_add_4_29.INJECT1_1 = "NO";
    CCU2D o_wb_addr_548_add_4_27 (.A0(n17404), .B0(\iw_word[1] ), .C0(dac_clk_p_c_enable_132), 
          .D0(\iw_word[26] ), .A1(n17402), .B1(\iw_word[1] ), .C1(dac_clk_p_c_enable_132), 
          .D1(\iw_word[27] ), .CIN(n17707), .COUT(n17708), .S0(n125[24]), 
          .S1(n125[25]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_548_add_4_27.INIT0 = 16'h5aaa;
    defparam o_wb_addr_548_add_4_27.INIT1 = 16'h5aaa;
    defparam o_wb_addr_548_add_4_27.INJECT1_0 = "NO";
    defparam o_wb_addr_548_add_4_27.INJECT1_1 = "NO";
    CCU2D o_wb_addr_548_add_4_25 (.A0(n17408), .B0(\iw_word[1] ), .C0(dac_clk_p_c_enable_132), 
          .D0(\iw_word[24] ), .A1(n17406), .B1(\iw_word[1] ), .C1(dac_clk_p_c_enable_132), 
          .D1(\iw_word[25] ), .CIN(n17706), .COUT(n17707), .S0(n125[22]), 
          .S1(n125[23]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_548_add_4_25.INIT0 = 16'h5aaa;
    defparam o_wb_addr_548_add_4_25.INIT1 = 16'h5aaa;
    defparam o_wb_addr_548_add_4_25.INJECT1_0 = "NO";
    defparam o_wb_addr_548_add_4_25.INJECT1_1 = "NO";
    CCU2D o_wb_addr_548_add_4_23 (.A0(n17412), .B0(\iw_word[1] ), .C0(dac_clk_p_c_enable_132), 
          .D0(\iw_word[22] ), .A1(n17410), .B1(\iw_word[1] ), .C1(dac_clk_p_c_enable_132), 
          .D1(\iw_word[23] ), .CIN(n17705), .COUT(n17706), .S0(n125[20]), 
          .S1(n125[21]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_548_add_4_23.INIT0 = 16'h5aaa;
    defparam o_wb_addr_548_add_4_23.INIT1 = 16'h5aaa;
    defparam o_wb_addr_548_add_4_23.INJECT1_0 = "NO";
    defparam o_wb_addr_548_add_4_23.INJECT1_1 = "NO";
    CCU2D o_wb_addr_548_add_4_21 (.A0(n17416), .B0(\iw_word[1] ), .C0(dac_clk_p_c_enable_132), 
          .D0(\iw_word[20] ), .A1(n17414), .B1(\iw_word[1] ), .C1(dac_clk_p_c_enable_132), 
          .D1(\iw_word[21] ), .CIN(n17704), .COUT(n17705), .S0(n125[18]), 
          .S1(n125[19]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_548_add_4_21.INIT0 = 16'h5aaa;
    defparam o_wb_addr_548_add_4_21.INIT1 = 16'h5aaa;
    defparam o_wb_addr_548_add_4_21.INJECT1_0 = "NO";
    defparam o_wb_addr_548_add_4_21.INJECT1_1 = "NO";
    CCU2D o_wb_addr_548_add_4_19 (.A0(n17420), .B0(\iw_word[1] ), .C0(dac_clk_p_c_enable_132), 
          .D0(\iw_word[18] ), .A1(n17418), .B1(\iw_word[1] ), .C1(dac_clk_p_c_enable_132), 
          .D1(\iw_word[19] ), .CIN(n17703), .COUT(n17704), .S0(n125[16]), 
          .S1(n125[17]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_548_add_4_19.INIT0 = 16'h5aaa;
    defparam o_wb_addr_548_add_4_19.INIT1 = 16'h5aaa;
    defparam o_wb_addr_548_add_4_19.INJECT1_0 = "NO";
    defparam o_wb_addr_548_add_4_19.INJECT1_1 = "NO";
    CCU2D o_wb_addr_548_add_4_17 (.A0(n17424), .B0(\iw_word[1] ), .C0(dac_clk_p_c_enable_132), 
          .D0(\iw_word[16] ), .A1(n17422), .B1(\iw_word[1] ), .C1(dac_clk_p_c_enable_132), 
          .D1(\iw_word[17] ), .CIN(n17702), .COUT(n17703), .S0(n125[14]), 
          .S1(n125[15]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_548_add_4_17.INIT0 = 16'h5aaa;
    defparam o_wb_addr_548_add_4_17.INIT1 = 16'h5aaa;
    defparam o_wb_addr_548_add_4_17.INJECT1_0 = "NO";
    defparam o_wb_addr_548_add_4_17.INJECT1_1 = "NO";
    CCU2D o_wb_addr_548_add_4_15 (.A0(n17428), .B0(\iw_word[1] ), .C0(dac_clk_p_c_enable_132), 
          .D0(\iw_word[14] ), .A1(n17426), .B1(\iw_word[1] ), .C1(dac_clk_p_c_enable_132), 
          .D1(\iw_word[15] ), .CIN(n17701), .COUT(n17702), .S0(n125[12]), 
          .S1(n125[13]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_548_add_4_15.INIT0 = 16'h5aaa;
    defparam o_wb_addr_548_add_4_15.INIT1 = 16'h5aaa;
    defparam o_wb_addr_548_add_4_15.INJECT1_0 = "NO";
    defparam o_wb_addr_548_add_4_15.INJECT1_1 = "NO";
    CCU2D o_wb_addr_548_add_4_13 (.A0(n17432), .B0(\iw_word[1] ), .C0(dac_clk_p_c_enable_132), 
          .D0(\iw_word[12] ), .A1(n17430), .B1(\iw_word[1] ), .C1(dac_clk_p_c_enable_132), 
          .D1(\iw_word[13] ), .CIN(n17700), .COUT(n17701), .S0(n125[10]), 
          .S1(n125[11]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_548_add_4_13.INIT0 = 16'h5aaa;
    defparam o_wb_addr_548_add_4_13.INIT1 = 16'h5aaa;
    defparam o_wb_addr_548_add_4_13.INJECT1_0 = "NO";
    defparam o_wb_addr_548_add_4_13.INJECT1_1 = "NO";
    CCU2D o_wb_addr_548_add_4_11 (.A0(n17436), .B0(\iw_word[1] ), .C0(dac_clk_p_c_enable_132), 
          .D0(\iw_word[10] ), .A1(n17434), .B1(\iw_word[1] ), .C1(dac_clk_p_c_enable_132), 
          .D1(\iw_word[11] ), .CIN(n17699), .COUT(n17700), .S0(n125[8]), 
          .S1(n125[9]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_548_add_4_11.INIT0 = 16'h5aaa;
    defparam o_wb_addr_548_add_4_11.INIT1 = 16'h5aaa;
    defparam o_wb_addr_548_add_4_11.INJECT1_0 = "NO";
    defparam o_wb_addr_548_add_4_11.INJECT1_1 = "NO";
    CCU2D o_wb_addr_548_add_4_9 (.A0(n17440), .B0(\iw_word[1] ), .C0(dac_clk_p_c_enable_132), 
          .D0(\iw_word[8] ), .A1(n17438), .B1(\iw_word[1] ), .C1(dac_clk_p_c_enable_132), 
          .D1(\iw_word[9] ), .CIN(n17698), .COUT(n17699), .S0(n125[6]), 
          .S1(n125[7]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_548_add_4_9.INIT0 = 16'h5aaa;
    defparam o_wb_addr_548_add_4_9.INIT1 = 16'h5aaa;
    defparam o_wb_addr_548_add_4_9.INJECT1_0 = "NO";
    defparam o_wb_addr_548_add_4_9.INJECT1_1 = "NO";
    CCU2D o_wb_addr_548_add_4_7 (.A0(n17444), .B0(\iw_word[1] ), .C0(dac_clk_p_c_enable_132), 
          .D0(\iw_word[6] ), .A1(n17442), .B1(\iw_word[1] ), .C1(dac_clk_p_c_enable_132), 
          .D1(\iw_word[7] ), .CIN(n17697), .COUT(n17698), .S0(n125[4]), 
          .S1(n125[5]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_548_add_4_7.INIT0 = 16'h5aaa;
    defparam o_wb_addr_548_add_4_7.INIT1 = 16'h5aaa;
    defparam o_wb_addr_548_add_4_7.INJECT1_0 = "NO";
    defparam o_wb_addr_548_add_4_7.INJECT1_1 = "NO";
    CCU2D o_wb_addr_548_add_4_5 (.A0(n17448), .B0(\iw_word[1] ), .C0(dac_clk_p_c_enable_132), 
          .D0(\iw_word[4] ), .A1(n17446), .B1(\iw_word[1] ), .C1(dac_clk_p_c_enable_132), 
          .D1(\iw_word[5] ), .CIN(n17696), .COUT(n17697), .S0(n125[2]), 
          .S1(n125[3]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_548_add_4_5.INIT0 = 16'h5aaa;
    defparam o_wb_addr_548_add_4_5.INIT1 = 16'h5aaa;
    defparam o_wb_addr_548_add_4_5.INJECT1_0 = "NO";
    defparam o_wb_addr_548_add_4_5.INJECT1_1 = "NO";
    CCU2D o_wb_addr_548_add_4_3 (.A0(n17451), .B0(dac_clk_p_c_enable_132), 
          .C0(\iw_word[1] ), .D0(wb_addr[0]), .A1(n17450), .B1(\iw_word[1] ), 
          .C1(dac_clk_p_c_enable_132), .D1(\iw_word[3] ), .CIN(n17695), 
          .COUT(n17696), .S0(n125[0]), .S1(n125[1]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_548_add_4_3.INIT0 = 16'h59aa;
    defparam o_wb_addr_548_add_4_3.INIT1 = 16'h5aaa;
    defparam o_wb_addr_548_add_4_3.INJECT1_0 = "NO";
    defparam o_wb_addr_548_add_4_3.INJECT1_1 = "NO";
    CCU2D o_wb_addr_548_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\iw_word[1] ), .B1(dac_clk_p_c_enable_132), 
          .C1(GND_net), .D1(GND_net), .COUT(n17695));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_548_add_4_1.INIT0 = 16'hF000;
    defparam o_wb_addr_548_add_4_1.INIT1 = 16'hffff;
    defparam o_wb_addr_548_add_4_1.INJECT1_0 = "NO";
    defparam o_wb_addr_548_add_4_1.INJECT1_1 = "NO";
    LUT4 i15584_2_lut (.A(wb_addr[28]), .B(n3), .Z(n17396)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15584_2_lut.init = 16'h8888;
    LUT4 i15585_2_lut (.A(wb_addr[29]), .B(n3), .Z(n17394)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15585_2_lut.init = 16'h8888;
    LUT4 i1_4_lut (.A(\iw_word[1] ), .B(n27112), .C(wb_cyc), .D(\iw_word[32] ), 
         .Z(n3)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;
    defparam i1_4_lut.init = 16'hfffb;
    LUT4 i15579_2_lut (.A(wb_addr[26]), .B(n3), .Z(n17400)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15579_2_lut.init = 16'h8888;
    LUT4 i15583_2_lut (.A(wb_addr[27]), .B(n3), .Z(n17398)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15583_2_lut.init = 16'h8888;
    LUT4 i15577_2_lut (.A(wb_addr[24]), .B(n3), .Z(n17404)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15577_2_lut.init = 16'h8888;
    LUT4 i15578_2_lut (.A(wb_addr[25]), .B(n3), .Z(n17402)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15578_2_lut.init = 16'h8888;
    LUT4 i15568_2_lut (.A(wb_addr[22]), .B(n3), .Z(n17408)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15568_2_lut.init = 16'h8888;
    LUT4 i15572_2_lut (.A(wb_addr[23]), .B(n3), .Z(n17406)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15572_2_lut.init = 16'h8888;
    LUT4 i15582_2_lut (.A(wb_addr[20]), .B(n3), .Z(n17412)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15582_2_lut.init = 16'h8888;
    LUT4 i15539_2_lut (.A(wb_addr[21]), .B(n3), .Z(n17410)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15539_2_lut.init = 16'h8888;
    LUT4 i15554_2_lut (.A(wb_addr[18]), .B(n3), .Z(n17416)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15554_2_lut.init = 16'h8888;
    LUT4 i15567_2_lut (.A(wb_addr[19]), .B(n3), .Z(n17414)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15567_2_lut.init = 16'h8888;
    LUT4 i15540_2_lut (.A(wb_addr[16]), .B(n3), .Z(n17420)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15540_2_lut.init = 16'h8888;
    LUT4 i15553_2_lut (.A(wb_addr[17]), .B(n3), .Z(n17418)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15553_2_lut.init = 16'h8888;
    LUT4 i15521_2_lut (.A(wb_addr[14]), .B(n3), .Z(n17424)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15521_2_lut.init = 16'h8888;
    LUT4 i15538_2_lut (.A(wb_addr[15]), .B(n3), .Z(n17422)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15538_2_lut.init = 16'h8888;
    LUT4 i15569_2_lut (.A(wb_addr[12]), .B(n3), .Z(n17428)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15569_2_lut.init = 16'h8888;
    LUT4 i15581_2_lut (.A(wb_addr[13]), .B(n3), .Z(n17426)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15581_2_lut.init = 16'h8888;
    LUT4 i15556_2_lut (.A(wb_addr[10]), .B(n3), .Z(n17432)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15556_2_lut.init = 16'h8888;
    LUT4 i15557_2_lut (.A(wb_addr[11]), .B(n3), .Z(n17430)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15557_2_lut.init = 16'h8888;
    LUT4 i15543_2_lut (.A(wb_addr[8]), .B(n3), .Z(n17436)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15543_2_lut.init = 16'h8888;
    LUT4 i15555_2_lut (.A(wb_addr[9]), .B(n3), .Z(n17434)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15555_2_lut.init = 16'h8888;
    LUT4 i15541_2_lut (.A(wb_addr[6]), .B(n3), .Z(n17440)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15541_2_lut.init = 16'h8888;
    LUT4 i15542_2_lut (.A(wb_addr[7]), .B(n3), .Z(n17438)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15542_2_lut.init = 16'h8888;
    LUT4 i15536_2_lut (.A(wb_addr[4]), .B(n3), .Z(n17444)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15536_2_lut.init = 16'h8888;
    LUT4 i15537_2_lut (.A(wb_addr[5]), .B(n3), .Z(n17442)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15537_2_lut.init = 16'h8888;
    LUT4 i15534_2_lut (.A(wb_addr[2]), .B(n3), .Z(n17448)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15534_2_lut.init = 16'h8888;
    LUT4 i15535_2_lut (.A(wb_addr[3]), .B(n3), .Z(n17446)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15535_2_lut.init = 16'h8888;
    LUT4 i15533_2_lut (.A(wb_addr[1]), .B(n3), .Z(n17450)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam i15533_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_131 (.A(wb_err), .B(n29560), .C(wb_we), .D(wb_cyc), 
         .Z(n20476)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut_adj_131.init = 16'h0100;
    LUT4 i1_4_lut_adj_132 (.A(n27111), .B(o_cmd_busy_N_941), .C(wb_ack), 
         .D(o_cmd_busy_N_933), .Z(dac_clk_p_c_enable_415)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+!((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(122[6:41])
    defparam i1_4_lut_adj_132.init = 16'heefc;
    LUT4 i22636_2_lut (.A(wb_cyc), .B(wb_stb), .Z(o_cmd_busy_N_933)) /* synthesis lut_function=(!(A+(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(149[11] 168[5])
    defparam i22636_2_lut.init = 16'h1111;
    LUT4 i1_2_lut_3_lut_4_lut (.A(wb_err), .B(wb_cyc), .C(wb_stb), .D(n29560), 
         .Z(n19812)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(122[17:41])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfff8;
    LUT4 i1_2_lut_rep_546_3_lut (.A(wb_err), .B(wb_cyc), .C(n29560), .Z(o_cmd_busy_N_941)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(122[17:41])
    defparam i1_2_lut_rep_546_3_lut.init = 16'hf8f8;
    FD1S3IX o_rsp_word_i1 (.D(n20476), .CK(dac_clk_p_c), .CD(n12737), 
            .Q(ow_word[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(278[9] 309[5])
    defparam o_rsp_word_i1.GSR = "DISABLED";
    FD1P3IX o_wb_cyc_67 (.D(o_cmd_busy_N_933), .SP(dac_clk_p_c_enable_415), 
            .CD(o_cmd_busy_N_941), .CK(dac_clk_p_c), .Q(wb_cyc)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=15, LSE_RCOL=15, LSE_LLINE=105, LSE_RLINE=109 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(121[9] 168[5])
    defparam o_wb_cyc_67.GSR = "DISABLED";
    FD1P3AX o_wb_addr_548__i29 (.D(n125[29]), .SP(dac_clk_p_c_enable_446), 
            .CK(dac_clk_p_c), .Q(wb_addr[29])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_548__i29.GSR = "DISABLED";
    FD1P3AX o_wb_addr_548__i28 (.D(n125[28]), .SP(dac_clk_p_c_enable_446), 
            .CK(dac_clk_p_c), .Q(wb_addr[28])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_548__i28.GSR = "DISABLED";
    FD1P3AX o_wb_addr_548__i27 (.D(n125[27]), .SP(dac_clk_p_c_enable_446), 
            .CK(dac_clk_p_c), .Q(wb_addr[27])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_548__i27.GSR = "DISABLED";
    FD1P3AX o_wb_addr_548__i26 (.D(n125[26]), .SP(dac_clk_p_c_enable_446), 
            .CK(dac_clk_p_c), .Q(wb_addr[26])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_548__i26.GSR = "DISABLED";
    FD1P3AX o_wb_addr_548__i25 (.D(n125[25]), .SP(dac_clk_p_c_enable_446), 
            .CK(dac_clk_p_c), .Q(wb_addr[25])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_548__i25.GSR = "DISABLED";
    FD1P3AX o_wb_addr_548__i24 (.D(n125[24]), .SP(dac_clk_p_c_enable_446), 
            .CK(dac_clk_p_c), .Q(wb_addr[24])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_548__i24.GSR = "DISABLED";
    FD1P3AX o_wb_addr_548__i23 (.D(n125[23]), .SP(dac_clk_p_c_enable_446), 
            .CK(dac_clk_p_c), .Q(wb_addr[23])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_548__i23.GSR = "DISABLED";
    FD1P3AX o_wb_addr_548__i22 (.D(n125[22]), .SP(dac_clk_p_c_enable_446), 
            .CK(dac_clk_p_c), .Q(wb_addr[22])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_548__i22.GSR = "DISABLED";
    FD1P3AX o_wb_addr_548__i21 (.D(n125[21]), .SP(dac_clk_p_c_enable_446), 
            .CK(dac_clk_p_c), .Q(wb_addr[21])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_548__i21.GSR = "DISABLED";
    FD1P3AX o_wb_addr_548__i20 (.D(n125[20]), .SP(dac_clk_p_c_enable_446), 
            .CK(dac_clk_p_c), .Q(wb_addr[20])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_548__i20.GSR = "DISABLED";
    FD1P3AX o_wb_addr_548__i19 (.D(n125[19]), .SP(dac_clk_p_c_enable_446), 
            .CK(dac_clk_p_c), .Q(wb_addr[19])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_548__i19.GSR = "DISABLED";
    FD1P3AX o_wb_addr_548__i18 (.D(n125[18]), .SP(dac_clk_p_c_enable_446), 
            .CK(dac_clk_p_c), .Q(wb_addr[18])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_548__i18.GSR = "DISABLED";
    FD1P3AX o_wb_addr_548__i17 (.D(n125[17]), .SP(dac_clk_p_c_enable_446), 
            .CK(dac_clk_p_c), .Q(wb_addr[17])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_548__i17.GSR = "DISABLED";
    FD1P3AX o_wb_addr_548__i16 (.D(n125[16]), .SP(dac_clk_p_c_enable_446), 
            .CK(dac_clk_p_c), .Q(wb_addr[16])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_548__i16.GSR = "DISABLED";
    FD1P3AX o_wb_addr_548__i15 (.D(n125[15]), .SP(dac_clk_p_c_enable_446), 
            .CK(dac_clk_p_c), .Q(wb_addr[15])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_548__i15.GSR = "DISABLED";
    FD1P3AX o_wb_addr_548__i14 (.D(n125[14]), .SP(dac_clk_p_c_enable_446), 
            .CK(dac_clk_p_c), .Q(wb_addr[14])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_548__i14.GSR = "DISABLED";
    FD1P3AX o_wb_addr_548__i13 (.D(n125[13]), .SP(dac_clk_p_c_enable_446), 
            .CK(dac_clk_p_c), .Q(wb_addr[13])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_548__i13.GSR = "DISABLED";
    FD1P3AX o_wb_addr_548__i12 (.D(n125[12]), .SP(dac_clk_p_c_enable_446), 
            .CK(dac_clk_p_c), .Q(wb_addr[12])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_548__i12.GSR = "DISABLED";
    FD1P3AX o_wb_addr_548__i11 (.D(n125[11]), .SP(dac_clk_p_c_enable_446), 
            .CK(dac_clk_p_c), .Q(wb_addr[11])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_548__i11.GSR = "DISABLED";
    FD1P3AX o_wb_addr_548__i10 (.D(n125[10]), .SP(dac_clk_p_c_enable_446), 
            .CK(dac_clk_p_c), .Q(wb_addr[10])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_548__i10.GSR = "DISABLED";
    FD1P3AX o_wb_addr_548__i9 (.D(n125[9]), .SP(dac_clk_p_c_enable_446), 
            .CK(dac_clk_p_c), .Q(wb_addr[9])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_548__i9.GSR = "DISABLED";
    FD1P3AX o_wb_addr_548__i8 (.D(n125[8]), .SP(dac_clk_p_c_enable_446), 
            .CK(dac_clk_p_c), .Q(wb_addr[8])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_548__i8.GSR = "DISABLED";
    FD1P3AX o_wb_addr_548__i7 (.D(n125[7]), .SP(dac_clk_p_c_enable_446), 
            .CK(dac_clk_p_c), .Q(wb_addr[7])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_548__i7.GSR = "DISABLED";
    FD1P3AX o_wb_addr_548__i6 (.D(n125[6]), .SP(dac_clk_p_c_enable_446), 
            .CK(dac_clk_p_c), .Q(wb_addr[6])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_548__i6.GSR = "DISABLED";
    FD1P3AX o_wb_addr_548__i5 (.D(n125[5]), .SP(dac_clk_p_c_enable_446), 
            .CK(dac_clk_p_c), .Q(wb_addr[5])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_548__i5.GSR = "DISABLED";
    FD1P3AX o_wb_addr_548__i4 (.D(n125[4]), .SP(dac_clk_p_c_enable_446), 
            .CK(dac_clk_p_c), .Q(wb_addr[4])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_548__i4.GSR = "DISABLED";
    FD1P3AX o_wb_addr_548__i3 (.D(n125[3]), .SP(dac_clk_p_c_enable_446), 
            .CK(dac_clk_p_c), .Q(wb_addr[3])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_548__i3.GSR = "DISABLED";
    FD1P3AX o_wb_addr_548__i2 (.D(n125[2]), .SP(dac_clk_p_c_enable_446), 
            .CK(dac_clk_p_c), .Q(wb_addr[2])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_548__i2.GSR = "DISABLED";
    FD1P3AX o_wb_addr_548__i1 (.D(n125[1]), .SP(dac_clk_p_c_enable_446), 
            .CK(dac_clk_p_c), .Q(wb_addr[1])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_548__i1.GSR = "DISABLED";
    FD1P3AX o_wb_addr_548__i0 (.D(n125[0]), .SP(dac_clk_p_c_enable_446), 
            .CK(dac_clk_p_c), .Q(wb_addr[0])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbexec.v(215[12] 222[51])
    defparam o_wb_addr_548__i0.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module hbdeword
//

module hbdeword (dac_clk_p_c, dac_clk_p_c_enable_308, idl_stb, hb_busy, 
            hb_bits, n29560, nl_busy, hx_stb, idl_word, dac_clk_p_c_enable_194, 
            n29561, n29502, w_reset, n26906) /* synthesis syn_module_defined=1 */ ;
    input dac_clk_p_c;
    input dac_clk_p_c_enable_308;
    input idl_stb;
    output hb_busy;
    output [4:0]hb_bits;
    input n29560;
    input nl_busy;
    input hx_stb;
    input [33:0]idl_word;
    input dac_clk_p_c_enable_194;
    input n29561;
    input n29502;
    input w_reset;
    output n26906;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(28[49:58])
    wire [3:0]r_len;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(58[12:17])
    
    wire n26787;
    wire [3:0]n13;
    
    wire n26547;
    wire [31:0]r_word;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(59[13:19])
    wire [4:0]o_dw_bits_4__N_1188;
    
    wire dac_clk_p_c_enable_237, n12823;
    wire [31:0]r_word_31__N_1197;
    wire [3:0]r_len_3__N_1229;
    
    wire o_dw_busy_N_1269, n11571;
    wire [4:0]o_dw_bits_4__N_1279;
    
    wire n11569, n20214, n26108, n26905;
    
    FD1P3IX r_len__i0 (.D(n13[0]), .SP(dac_clk_p_c_enable_308), .CD(n26787), 
            .CK(dac_clk_p_c), .Q(r_len[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(64[9] 81[6])
    defparam r_len__i0.GSR = "DISABLED";
    LUT4 r_word_28__bdd_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(n26547), 
         .D(r_word[28]), .Z(o_dw_bits_4__N_1188[0])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_28__bdd_3_lut_4_lut.init = 16'hfd20;
    FD1P3AX o_dw_bits_i0 (.D(o_dw_bits_4__N_1188[0]), .SP(dac_clk_p_c_enable_237), 
            .CK(dac_clk_p_c), .Q(hb_bits[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(95[9] 103[41])
    defparam o_dw_bits_i0.GSR = "DISABLED";
    LUT4 i7071_2_lut_rep_464_3_lut (.A(idl_stb), .B(hb_busy), .C(n29560), 
         .Z(n26787)) /* synthesis lut_function=(A ((C)+!B)+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam i7071_2_lut_rep_464_3_lut.init = 16'hf2f2;
    LUT4 i22646_2_lut_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(nl_busy), 
         .D(hx_stb), .Z(n12823)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam i22646_2_lut_3_lut_4_lut.init = 16'h0ddd;
    LUT4 i1_2_lut_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(nl_busy), 
         .D(hx_stb), .Z(dac_clk_p_c_enable_237)) /* synthesis lut_function=(!(A (B (C (D)))+!A (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h2fff;
    LUT4 r_word_31__I_0_i32_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[31]), 
         .D(r_word[27]), .Z(r_word_31__N_1197[31])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i32_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i31_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[30]), 
         .D(r_word[26]), .Z(r_word_31__N_1197[30])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i31_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i30_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[29]), 
         .D(r_word[25]), .Z(r_word_31__N_1197[29])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i30_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i29_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[28]), 
         .D(r_word[24]), .Z(r_word_31__N_1197[28])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i29_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i28_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[27]), 
         .D(r_word[23]), .Z(r_word_31__N_1197[27])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i28_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i27_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[26]), 
         .D(r_word[22]), .Z(r_word_31__N_1197[26])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i27_3_lut_4_lut.init = 16'hfd20;
    FD1P3AX o_dw_bits_i3 (.D(o_dw_bits_4__N_1188[3]), .SP(dac_clk_p_c_enable_237), 
            .CK(dac_clk_p_c), .Q(hb_bits[3])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(95[9] 103[41])
    defparam o_dw_bits_i3.GSR = "DISABLED";
    FD1P3AX o_dw_bits_i2 (.D(o_dw_bits_4__N_1188[2]), .SP(dac_clk_p_c_enable_237), 
            .CK(dac_clk_p_c), .Q(hb_bits[2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(95[9] 103[41])
    defparam o_dw_bits_i2.GSR = "DISABLED";
    FD1P3AX o_dw_bits_i1 (.D(o_dw_bits_4__N_1188[1]), .SP(dac_clk_p_c_enable_237), 
            .CK(dac_clk_p_c), .Q(hb_bits[1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(95[9] 103[41])
    defparam o_dw_bits_i1.GSR = "DISABLED";
    FD1P3AX r_word_i31 (.D(r_word_31__N_1197[31]), .SP(dac_clk_p_c_enable_237), 
            .CK(dac_clk_p_c), .Q(r_word[31])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i31.GSR = "DISABLED";
    LUT4 r_word_31__I_0_i26_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[25]), 
         .D(r_word[21]), .Z(r_word_31__N_1197[25])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i26_3_lut_4_lut.init = 16'hfd20;
    FD1P3IX r_len__i3 (.D(r_len_3__N_1229[3]), .SP(dac_clk_p_c_enable_194), 
            .CD(n29561), .CK(dac_clk_p_c), .Q(r_len[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(64[9] 81[6])
    defparam r_len__i3.GSR = "DISABLED";
    FD1P3IX r_word_i1 (.D(idl_word[1]), .SP(dac_clk_p_c_enable_237), .CD(n12823), 
            .CK(dac_clk_p_c), .Q(r_word[1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i1.GSR = "DISABLED";
    FD1P3IX r_word_i2 (.D(idl_word[2]), .SP(dac_clk_p_c_enable_237), .CD(n12823), 
            .CK(dac_clk_p_c), .Q(r_word[2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i2.GSR = "DISABLED";
    FD1P3IX r_word_i3 (.D(idl_word[3]), .SP(dac_clk_p_c_enable_237), .CD(n12823), 
            .CK(dac_clk_p_c), .Q(r_word[3])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i3.GSR = "DISABLED";
    FD1P3IX o_dw_bits_i4 (.D(n29502), .SP(dac_clk_p_c_enable_237), .CD(n12823), 
            .CK(dac_clk_p_c), .Q(hb_bits[4])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(95[9] 103[41])
    defparam o_dw_bits_i4.GSR = "DISABLED";
    FD1P3IX o_dw_stb_36 (.D(o_dw_busy_N_1269), .SP(dac_clk_p_c_enable_194), 
            .CD(w_reset), .CK(dac_clk_p_c), .Q(hb_busy)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(64[9] 81[6])
    defparam o_dw_stb_36.GSR = "DISABLED";
    FD1P3IX r_word_i0 (.D(idl_word[0]), .SP(dac_clk_p_c_enable_237), .CD(n12823), 
            .CK(dac_clk_p_c), .Q(r_word[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i0.GSR = "DISABLED";
    FD1P3AX r_word_i30 (.D(r_word_31__N_1197[30]), .SP(dac_clk_p_c_enable_237), 
            .CK(dac_clk_p_c), .Q(r_word[30])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i30.GSR = "DISABLED";
    FD1P3AX r_word_i29 (.D(r_word_31__N_1197[29]), .SP(dac_clk_p_c_enable_237), 
            .CK(dac_clk_p_c), .Q(r_word[29])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i29.GSR = "DISABLED";
    FD1P3AX r_word_i28 (.D(r_word_31__N_1197[28]), .SP(dac_clk_p_c_enable_237), 
            .CK(dac_clk_p_c), .Q(r_word[28])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i28.GSR = "DISABLED";
    FD1P3AX r_word_i27 (.D(r_word_31__N_1197[27]), .SP(dac_clk_p_c_enable_237), 
            .CK(dac_clk_p_c), .Q(r_word[27])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i27.GSR = "DISABLED";
    FD1P3AX r_word_i26 (.D(r_word_31__N_1197[26]), .SP(dac_clk_p_c_enable_237), 
            .CK(dac_clk_p_c), .Q(r_word[26])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i26.GSR = "DISABLED";
    FD1P3AX r_word_i25 (.D(r_word_31__N_1197[25]), .SP(dac_clk_p_c_enable_237), 
            .CK(dac_clk_p_c), .Q(r_word[25])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i25.GSR = "DISABLED";
    FD1P3AX r_word_i24 (.D(r_word_31__N_1197[24]), .SP(dac_clk_p_c_enable_237), 
            .CK(dac_clk_p_c), .Q(r_word[24])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i24.GSR = "DISABLED";
    FD1P3AX r_word_i23 (.D(r_word_31__N_1197[23]), .SP(dac_clk_p_c_enable_237), 
            .CK(dac_clk_p_c), .Q(r_word[23])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i23.GSR = "DISABLED";
    FD1P3AX r_word_i22 (.D(r_word_31__N_1197[22]), .SP(dac_clk_p_c_enable_237), 
            .CK(dac_clk_p_c), .Q(r_word[22])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i22.GSR = "DISABLED";
    FD1P3AX r_word_i21 (.D(r_word_31__N_1197[21]), .SP(dac_clk_p_c_enable_237), 
            .CK(dac_clk_p_c), .Q(r_word[21])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i21.GSR = "DISABLED";
    FD1P3AX r_word_i20 (.D(r_word_31__N_1197[20]), .SP(dac_clk_p_c_enable_237), 
            .CK(dac_clk_p_c), .Q(r_word[20])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i20.GSR = "DISABLED";
    FD1P3AX r_word_i19 (.D(r_word_31__N_1197[19]), .SP(dac_clk_p_c_enable_237), 
            .CK(dac_clk_p_c), .Q(r_word[19])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i19.GSR = "DISABLED";
    FD1P3AX r_word_i18 (.D(r_word_31__N_1197[18]), .SP(dac_clk_p_c_enable_237), 
            .CK(dac_clk_p_c), .Q(r_word[18])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i18.GSR = "DISABLED";
    FD1P3AX r_word_i17 (.D(r_word_31__N_1197[17]), .SP(dac_clk_p_c_enable_237), 
            .CK(dac_clk_p_c), .Q(r_word[17])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i17.GSR = "DISABLED";
    FD1P3AX r_word_i16 (.D(r_word_31__N_1197[16]), .SP(dac_clk_p_c_enable_237), 
            .CK(dac_clk_p_c), .Q(r_word[16])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i16.GSR = "DISABLED";
    FD1P3AX r_word_i15 (.D(r_word_31__N_1197[15]), .SP(dac_clk_p_c_enable_237), 
            .CK(dac_clk_p_c), .Q(r_word[15])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i15.GSR = "DISABLED";
    FD1P3AX r_word_i14 (.D(r_word_31__N_1197[14]), .SP(dac_clk_p_c_enable_237), 
            .CK(dac_clk_p_c), .Q(r_word[14])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i14.GSR = "DISABLED";
    FD1P3AX r_word_i13 (.D(r_word_31__N_1197[13]), .SP(dac_clk_p_c_enable_237), 
            .CK(dac_clk_p_c), .Q(r_word[13])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i13.GSR = "DISABLED";
    FD1P3AX r_word_i12 (.D(r_word_31__N_1197[12]), .SP(dac_clk_p_c_enable_237), 
            .CK(dac_clk_p_c), .Q(r_word[12])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i12.GSR = "DISABLED";
    FD1P3AX r_word_i11 (.D(r_word_31__N_1197[11]), .SP(dac_clk_p_c_enable_237), 
            .CK(dac_clk_p_c), .Q(r_word[11])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i11.GSR = "DISABLED";
    FD1P3AX r_word_i10 (.D(r_word_31__N_1197[10]), .SP(dac_clk_p_c_enable_237), 
            .CK(dac_clk_p_c), .Q(r_word[10])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i10.GSR = "DISABLED";
    FD1P3AX r_word_i9 (.D(r_word_31__N_1197[9]), .SP(dac_clk_p_c_enable_237), 
            .CK(dac_clk_p_c), .Q(r_word[9])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i9.GSR = "DISABLED";
    FD1P3AX r_word_i8 (.D(r_word_31__N_1197[8]), .SP(dac_clk_p_c_enable_237), 
            .CK(dac_clk_p_c), .Q(r_word[8])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i8.GSR = "DISABLED";
    FD1P3AX r_word_i7 (.D(r_word_31__N_1197[7]), .SP(dac_clk_p_c_enable_237), 
            .CK(dac_clk_p_c), .Q(r_word[7])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i7.GSR = "DISABLED";
    FD1P3AX r_word_i6 (.D(r_word_31__N_1197[6]), .SP(dac_clk_p_c_enable_237), 
            .CK(dac_clk_p_c), .Q(r_word[6])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i6.GSR = "DISABLED";
    FD1P3AX r_word_i5 (.D(r_word_31__N_1197[5]), .SP(dac_clk_p_c_enable_237), 
            .CK(dac_clk_p_c), .Q(r_word[5])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i5.GSR = "DISABLED";
    FD1P3AX r_word_i4 (.D(r_word_31__N_1197[4]), .SP(dac_clk_p_c_enable_237), 
            .CK(dac_clk_p_c), .Q(r_word[4])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(83[9] 93[37])
    defparam r_word_i4.GSR = "DISABLED";
    LUT4 r_word_31__I_0_i25_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[24]), 
         .D(r_word[20]), .Z(r_word_31__N_1197[24])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i25_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i24_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[23]), 
         .D(r_word[19]), .Z(r_word_31__N_1197[23])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i24_3_lut_4_lut.init = 16'hfd20;
    LUT4 i1_3_lut_4_lut_3_lut_4_lut (.A(r_len[0]), .B(r_len[1]), .C(r_len[2]), 
         .D(r_len[3]), .Z(n11571)) /* synthesis lut_function=(A (B)+!A !(B+!(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(80[14:26])
    defparam i1_3_lut_4_lut_3_lut_4_lut.init = 16'h9998;
    LUT4 r_word_31__I_0_i20_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[19]), 
         .D(r_word[15]), .Z(r_word_31__N_1197[19])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i20_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i23_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[22]), 
         .D(r_word[18]), .Z(r_word_31__N_1197[22])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i23_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i19_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[18]), 
         .D(r_word[14]), .Z(r_word_31__N_1197[18])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i19_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i22_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[21]), 
         .D(r_word[17]), .Z(r_word_31__N_1197[21])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i22_3_lut_4_lut.init = 16'hfd20;
    LUT4 i11017_2_lut (.A(idl_word[32]), .B(idl_word[33]), .Z(o_dw_bits_4__N_1279[3])) /* synthesis lut_function=(A (B)) */ ;
    defparam i11017_2_lut.init = 16'h8888;
    LUT4 r_word_31__I_0_i21_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[20]), 
         .D(r_word[16]), .Z(r_word_31__N_1197[20])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i21_3_lut_4_lut.init = 16'hfd20;
    FD1P3IX r_len__i2 (.D(n11569), .SP(dac_clk_p_c_enable_308), .CD(n26787), 
            .CK(dac_clk_p_c), .Q(r_len[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(64[9] 81[6])
    defparam r_len__i2.GSR = "DISABLED";
    FD1P3IX r_len__i1 (.D(n11571), .SP(dac_clk_p_c_enable_308), .CD(n26787), 
            .CK(dac_clk_p_c), .Q(r_len[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=127, LSE_RLINE=129 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(64[9] 81[6])
    defparam r_len__i1.GSR = "DISABLED";
    LUT4 r_word_31__I_0_i18_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[17]), 
         .D(r_word[13]), .Z(r_word_31__N_1197[17])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i18_3_lut_4_lut.init = 16'hfd20;
    LUT4 o_dw_bits_4__I_0_i3_4_lut (.A(r_word[30]), .B(idl_word[31]), .C(n26906), 
         .D(o_dw_bits_4__N_1279[3]), .Z(o_dw_bits_4__N_1188[2])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(102[12] 103[41])
    defparam o_dw_bits_4__I_0_i3_4_lut.init = 16'hca0a;
    LUT4 mux_15_i4_4_lut (.A(r_len[3]), .B(o_dw_bits_4__N_1279[3]), .C(n26906), 
         .D(n20214), .Z(r_len_3__N_1229[3])) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(76[12] 81[6])
    defparam mux_15_i4_4_lut.init = 16'h3a35;
    LUT4 r_word_29__bdd_3_lut_24269 (.A(idl_word[30]), .B(idl_word[33]), 
         .C(idl_word[32]), .Z(n26108)) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam r_word_29__bdd_3_lut_24269.init = 16'h8c8c;
    LUT4 r_word_28__bdd_3_lut_24594 (.A(idl_word[29]), .B(idl_word[32]), 
         .C(idl_word[33]), .Z(n26547)) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;
    defparam r_word_28__bdd_3_lut_24594.init = 16'h8c8c;
    LUT4 r_word_31__I_0_i17_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[16]), 
         .D(r_word[12]), .Z(r_word_31__N_1197[16])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i17_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i14_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[13]), 
         .D(r_word[9]), .Z(r_word_31__N_1197[13])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i14_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i13_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[12]), 
         .D(r_word[8]), .Z(r_word_31__N_1197[12])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i13_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i12_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[11]), 
         .D(r_word[7]), .Z(r_word_31__N_1197[11])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i12_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i11_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[10]), 
         .D(r_word[6]), .Z(r_word_31__N_1197[10])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i11_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i10_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[9]), 
         .D(r_word[5]), .Z(r_word_31__N_1197[9])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i10_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i9_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[8]), 
         .D(r_word[4]), .Z(r_word_31__N_1197[8])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i9_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i8_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[7]), 
         .D(r_word[3]), .Z(r_word_31__N_1197[7])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i8_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i7_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[6]), 
         .D(r_word[2]), .Z(r_word_31__N_1197[6])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i7_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i6_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[5]), 
         .D(r_word[1]), .Z(r_word_31__N_1197[5])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i6_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i5_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[4]), 
         .D(r_word[0]), .Z(r_word_31__N_1197[4])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i5_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_29__bdd_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(n26108), 
         .D(r_word[29]), .Z(o_dw_bits_4__N_1188[1])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_29__bdd_3_lut_4_lut.init = 16'hfd20;
    LUT4 r_word_31__I_0_i16_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[15]), 
         .D(r_word[11]), .Z(r_word_31__N_1197[15])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i16_3_lut_4_lut.init = 16'hfd20;
    LUT4 i1_3_lut_3_lut_4_lut (.A(r_len[0]), .B(r_len[1]), .C(r_len[3]), 
         .D(r_len[2]), .Z(n11569)) /* synthesis lut_function=(A (D)+!A (B (D)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(80[14:26])
    defparam i1_3_lut_3_lut_4_lut.init = 16'hee10;
    LUT4 r_word_31__I_0_i15_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(idl_word[14]), 
         .D(r_word[10]), .Z(r_word_31__N_1197[14])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam r_word_31__I_0_i15_3_lut_4_lut.init = 16'hfd20;
    LUT4 i1_4_lut_4_lut (.A(r_len[0]), .B(r_len[1]), .C(r_len[3]), .D(r_len[2]), 
         .Z(n20214)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(80[14:26])
    defparam i1_4_lut_4_lut.init = 16'hffef;
    LUT4 i3_4_lut_rep_582 (.A(r_len[0]), .B(r_len[1]), .C(r_len[2]), .D(r_len[3]), 
         .Z(n26905)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(78[16:31])
    defparam i3_4_lut_rep_582.init = 16'hfffe;
    LUT4 i1_2_lut_4_lut (.A(r_len[0]), .B(r_len[1]), .C(r_len[2]), .D(r_len[3]), 
         .Z(n13[0])) /* synthesis lut_function=(!(A+!(B+(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(78[16:31])
    defparam i1_2_lut_4_lut.init = 16'h5554;
    LUT4 i_stb_I_0_2_lut_rep_583 (.A(idl_stb), .B(hb_busy), .Z(n26906)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam i_stb_I_0_2_lut_rep_583.init = 16'h2222;
    LUT4 o_dw_bits_4__I_0_i4_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(o_dw_bits_4__N_1279[3]), 
         .D(r_word[31]), .Z(o_dw_bits_4__N_1188[3])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam o_dw_bits_4__I_0_i4_3_lut_4_lut.init = 16'hfd20;
    LUT4 i11026_2_lut_3_lut (.A(idl_stb), .B(hb_busy), .C(n26905), .Z(o_dw_busy_N_1269)) /* synthesis lut_function=(A ((C)+!B)+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(69[16:37])
    defparam i11026_2_lut_3_lut.init = 16'hf2f2;
    
endmodule
//
// Verilog Description of module hbpack
//

module hbpack (dac_clk_p_c, dac_clk_p_c_enable_381, n29561, iw_word, 
            \dec_bits[4] , w_reset, o_pck_stb_N_765, cmd_loaded, dac_clk_p_c_enable_196, 
            cmd_loaded_N_768, \dec_bits[1] , wb_cyc, inc, n17451, 
            \iw_word[32] , \iw_word[31] , \iw_word[30] , \iw_word[29] , 
            \iw_word[28] , \iw_word[27] , \iw_word[26] , \iw_word[25] , 
            \iw_word[24] , \iw_word[23] , \iw_word[22] , \iw_word[21] , 
            \iw_word[20] , \iw_word[19] , \iw_word[18] , \iw_word[17] , 
            \iw_word[16] , \iw_word[15] , \iw_word[14] , \iw_word[13] , 
            \iw_word[12] , \iw_word[11] , \iw_word[10] , \iw_word[9] , 
            \iw_word[8] , \iw_word[7] , \iw_word[6] , \iw_word[5] , 
            \iw_word[4] , \iw_word[3] , \iw_word[1] , n27111, i_cmd_wr, 
            wb_stb, n22219, n27112, dac_clk_p_c_enable_132, n29560, 
            newaddr_N_990, \dec_bits[0] , dac_clk_p_c_enable_350, n45, 
            n46, dac_clk_p_c_enable_446) /* synthesis syn_module_defined=1 */ ;
    input dac_clk_p_c;
    input dac_clk_p_c_enable_381;
    input n29561;
    output [33:0]iw_word;
    input \dec_bits[4] ;
    input w_reset;
    input o_pck_stb_N_765;
    output cmd_loaded;
    input dac_clk_p_c_enable_196;
    input cmd_loaded_N_768;
    input \dec_bits[1] ;
    input wb_cyc;
    input inc;
    output n17451;
    output \iw_word[32] ;
    output \iw_word[31] ;
    output \iw_word[30] ;
    output \iw_word[29] ;
    output \iw_word[28] ;
    output \iw_word[27] ;
    output \iw_word[26] ;
    output \iw_word[25] ;
    output \iw_word[24] ;
    output \iw_word[23] ;
    output \iw_word[22] ;
    output \iw_word[21] ;
    output \iw_word[20] ;
    output \iw_word[19] ;
    output \iw_word[18] ;
    output \iw_word[17] ;
    output \iw_word[16] ;
    output \iw_word[15] ;
    output \iw_word[14] ;
    output \iw_word[13] ;
    output \iw_word[12] ;
    output \iw_word[11] ;
    output \iw_word[10] ;
    output \iw_word[9] ;
    output \iw_word[8] ;
    output \iw_word[7] ;
    output \iw_word[6] ;
    output \iw_word[5] ;
    output \iw_word[4] ;
    output \iw_word[3] ;
    output \iw_word[1] ;
    output n27111;
    output i_cmd_wr;
    input wb_stb;
    output n22219;
    output n27112;
    output dac_clk_p_c_enable_132;
    input n29560;
    output newaddr_N_990;
    input \dec_bits[0] ;
    input dac_clk_p_c_enable_350;
    input n45;
    input n46;
    output dac_clk_p_c_enable_446;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(28[49:58])
    wire [33:0]r_word;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(71[13:19])
    wire [33:0]n14;
    
    wire iw_stb, n26895;
    wire [33:0]iw_word_c;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(71[14:21])
    
    FD1P3IX r_word__i0 (.D(n14[0]), .SP(dac_clk_p_c_enable_381), .CD(n29561), 
            .CK(dac_clk_p_c), .Q(r_word[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i0.GSR = "DISABLED";
    FD1P3IX o_pck_word__i0 (.D(r_word[0]), .SP(dac_clk_p_c_enable_381), 
            .CD(n29561), .CK(dac_clk_p_c), .Q(iw_word[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i0.GSR = "DISABLED";
    LUT4 i11309_2_lut (.A(r_word[9]), .B(\dec_bits[4] ), .Z(n14[13])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11309_2_lut.init = 16'h2222;
    LUT4 i11310_2_lut (.A(r_word[8]), .B(\dec_bits[4] ), .Z(n14[12])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11310_2_lut.init = 16'h2222;
    FD1S3IX o_pck_stb_24 (.D(o_pck_stb_N_765), .CK(dac_clk_p_c), .CD(w_reset), 
            .Q(iw_stb)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(83[9] 84[65])
    defparam o_pck_stb_24.GSR = "DISABLED";
    LUT4 i11311_2_lut (.A(r_word[7]), .B(\dec_bits[4] ), .Z(n14[11])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11311_2_lut.init = 16'h2222;
    LUT4 i11312_2_lut (.A(r_word[6]), .B(\dec_bits[4] ), .Z(n14[10])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11312_2_lut.init = 16'h2222;
    LUT4 i11313_2_lut (.A(r_word[5]), .B(\dec_bits[4] ), .Z(n14[9])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11313_2_lut.init = 16'h2222;
    LUT4 i11315_2_lut (.A(r_word[4]), .B(\dec_bits[4] ), .Z(n14[8])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11315_2_lut.init = 16'h2222;
    LUT4 i11317_2_lut (.A(r_word[3]), .B(\dec_bits[4] ), .Z(n14[7])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11317_2_lut.init = 16'h2222;
    LUT4 i11318_2_lut (.A(r_word[2]), .B(\dec_bits[4] ), .Z(n14[6])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11318_2_lut.init = 16'h2222;
    LUT4 i11319_2_lut (.A(r_word[1]), .B(\dec_bits[4] ), .Z(n14[5])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11319_2_lut.init = 16'h2222;
    LUT4 i11320_2_lut (.A(r_word[0]), .B(\dec_bits[4] ), .Z(n14[4])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11320_2_lut.init = 16'h2222;
    FD1P3IX cmd_loaded_23 (.D(cmd_loaded_N_768), .SP(dac_clk_p_c_enable_196), 
            .CD(w_reset), .CK(dac_clk_p_c), .Q(cmd_loaded)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(74[9] 80[23])
    defparam cmd_loaded_23.GSR = "DISABLED";
    LUT4 i11321_2_lut (.A(\dec_bits[1] ), .B(\dec_bits[4] ), .Z(n14[1])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11321_2_lut.init = 16'h2222;
    LUT4 i15532_3_lut_4_lut (.A(n26895), .B(wb_cyc), .C(iw_word[2]), .D(inc), 
         .Z(n17451)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(83[9] 84[65])
    defparam i15532_3_lut_4_lut.init = 16'hfd20;
    FD1P3IX o_pck_word__i33 (.D(r_word[33]), .SP(dac_clk_p_c_enable_381), 
            .CD(w_reset), .CK(dac_clk_p_c), .Q(iw_word_c[33])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i33.GSR = "DISABLED";
    FD1P3IX o_pck_word__i32 (.D(r_word[32]), .SP(dac_clk_p_c_enable_381), 
            .CD(w_reset), .CK(dac_clk_p_c), .Q(\iw_word[32] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i32.GSR = "DISABLED";
    FD1P3IX o_pck_word__i31 (.D(r_word[31]), .SP(dac_clk_p_c_enable_381), 
            .CD(w_reset), .CK(dac_clk_p_c), .Q(\iw_word[31] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i31.GSR = "DISABLED";
    FD1P3IX o_pck_word__i30 (.D(r_word[30]), .SP(dac_clk_p_c_enable_381), 
            .CD(w_reset), .CK(dac_clk_p_c), .Q(\iw_word[30] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i30.GSR = "DISABLED";
    FD1P3IX o_pck_word__i29 (.D(r_word[29]), .SP(dac_clk_p_c_enable_381), 
            .CD(w_reset), .CK(dac_clk_p_c), .Q(\iw_word[29] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i29.GSR = "DISABLED";
    FD1P3IX o_pck_word__i28 (.D(r_word[28]), .SP(dac_clk_p_c_enable_381), 
            .CD(w_reset), .CK(dac_clk_p_c), .Q(\iw_word[28] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i28.GSR = "DISABLED";
    FD1P3IX o_pck_word__i27 (.D(r_word[27]), .SP(dac_clk_p_c_enable_381), 
            .CD(w_reset), .CK(dac_clk_p_c), .Q(\iw_word[27] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i27.GSR = "DISABLED";
    FD1P3IX o_pck_word__i26 (.D(r_word[26]), .SP(dac_clk_p_c_enable_381), 
            .CD(w_reset), .CK(dac_clk_p_c), .Q(\iw_word[26] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i26.GSR = "DISABLED";
    FD1P3IX o_pck_word__i25 (.D(r_word[25]), .SP(dac_clk_p_c_enable_381), 
            .CD(w_reset), .CK(dac_clk_p_c), .Q(\iw_word[25] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i25.GSR = "DISABLED";
    FD1P3IX o_pck_word__i24 (.D(r_word[24]), .SP(dac_clk_p_c_enable_381), 
            .CD(w_reset), .CK(dac_clk_p_c), .Q(\iw_word[24] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i24.GSR = "DISABLED";
    FD1P3IX o_pck_word__i23 (.D(r_word[23]), .SP(dac_clk_p_c_enable_381), 
            .CD(n29561), .CK(dac_clk_p_c), .Q(\iw_word[23] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i23.GSR = "DISABLED";
    FD1P3IX o_pck_word__i22 (.D(r_word[22]), .SP(dac_clk_p_c_enable_381), 
            .CD(n29561), .CK(dac_clk_p_c), .Q(\iw_word[22] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i22.GSR = "DISABLED";
    FD1P3IX o_pck_word__i21 (.D(r_word[21]), .SP(dac_clk_p_c_enable_381), 
            .CD(w_reset), .CK(dac_clk_p_c), .Q(\iw_word[21] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i21.GSR = "DISABLED";
    FD1P3IX o_pck_word__i20 (.D(r_word[20]), .SP(dac_clk_p_c_enable_381), 
            .CD(n29561), .CK(dac_clk_p_c), .Q(\iw_word[20] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i20.GSR = "DISABLED";
    FD1P3IX o_pck_word__i19 (.D(r_word[19]), .SP(dac_clk_p_c_enable_381), 
            .CD(n29561), .CK(dac_clk_p_c), .Q(\iw_word[19] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i19.GSR = "DISABLED";
    FD1P3IX o_pck_word__i18 (.D(r_word[18]), .SP(dac_clk_p_c_enable_381), 
            .CD(n29561), .CK(dac_clk_p_c), .Q(\iw_word[18] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i18.GSR = "DISABLED";
    FD1P3IX o_pck_word__i17 (.D(r_word[17]), .SP(dac_clk_p_c_enable_381), 
            .CD(n29561), .CK(dac_clk_p_c), .Q(\iw_word[17] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i17.GSR = "DISABLED";
    FD1P3IX o_pck_word__i16 (.D(r_word[16]), .SP(dac_clk_p_c_enable_381), 
            .CD(n29561), .CK(dac_clk_p_c), .Q(\iw_word[16] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i16.GSR = "DISABLED";
    FD1P3IX o_pck_word__i15 (.D(r_word[15]), .SP(dac_clk_p_c_enable_381), 
            .CD(n29561), .CK(dac_clk_p_c), .Q(\iw_word[15] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i15.GSR = "DISABLED";
    FD1P3IX o_pck_word__i14 (.D(r_word[14]), .SP(dac_clk_p_c_enable_381), 
            .CD(n29561), .CK(dac_clk_p_c), .Q(\iw_word[14] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i14.GSR = "DISABLED";
    FD1P3IX o_pck_word__i13 (.D(r_word[13]), .SP(dac_clk_p_c_enable_381), 
            .CD(n29561), .CK(dac_clk_p_c), .Q(\iw_word[13] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i13.GSR = "DISABLED";
    FD1P3IX o_pck_word__i12 (.D(r_word[12]), .SP(dac_clk_p_c_enable_381), 
            .CD(n29561), .CK(dac_clk_p_c), .Q(\iw_word[12] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i12.GSR = "DISABLED";
    FD1P3IX o_pck_word__i11 (.D(r_word[11]), .SP(dac_clk_p_c_enable_381), 
            .CD(n29561), .CK(dac_clk_p_c), .Q(\iw_word[11] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i11.GSR = "DISABLED";
    FD1P3IX o_pck_word__i10 (.D(r_word[10]), .SP(dac_clk_p_c_enable_381), 
            .CD(n29561), .CK(dac_clk_p_c), .Q(\iw_word[10] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i10.GSR = "DISABLED";
    FD1P3IX o_pck_word__i9 (.D(r_word[9]), .SP(dac_clk_p_c_enable_381), 
            .CD(n29561), .CK(dac_clk_p_c), .Q(\iw_word[9] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i9.GSR = "DISABLED";
    FD1P3IX o_pck_word__i8 (.D(r_word[8]), .SP(dac_clk_p_c_enable_381), 
            .CD(n29561), .CK(dac_clk_p_c), .Q(\iw_word[8] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i8.GSR = "DISABLED";
    FD1P3IX o_pck_word__i7 (.D(r_word[7]), .SP(dac_clk_p_c_enable_381), 
            .CD(n29561), .CK(dac_clk_p_c), .Q(\iw_word[7] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i7.GSR = "DISABLED";
    FD1P3IX o_pck_word__i6 (.D(r_word[6]), .SP(dac_clk_p_c_enable_381), 
            .CD(n29561), .CK(dac_clk_p_c), .Q(\iw_word[6] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i6.GSR = "DISABLED";
    FD1P3IX o_pck_word__i5 (.D(r_word[5]), .SP(dac_clk_p_c_enable_381), 
            .CD(n29561), .CK(dac_clk_p_c), .Q(\iw_word[5] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i5.GSR = "DISABLED";
    FD1P3IX o_pck_word__i4 (.D(r_word[4]), .SP(dac_clk_p_c_enable_381), 
            .CD(n29561), .CK(dac_clk_p_c), .Q(\iw_word[4] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i4.GSR = "DISABLED";
    FD1P3IX o_pck_word__i3 (.D(r_word[3]), .SP(dac_clk_p_c_enable_381), 
            .CD(n29561), .CK(dac_clk_p_c), .Q(\iw_word[3] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i3.GSR = "DISABLED";
    FD1P3IX o_pck_word__i2 (.D(r_word[2]), .SP(dac_clk_p_c_enable_381), 
            .CD(n29561), .CK(dac_clk_p_c), .Q(iw_word[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i2.GSR = "DISABLED";
    FD1P3IX o_pck_word__i1 (.D(r_word[1]), .SP(dac_clk_p_c_enable_381), 
            .CD(n29561), .CK(dac_clk_p_c), .Q(\iw_word[1] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(106[9] 110[25])
    defparam o_pck_word__i1.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_788 (.A(iw_stb), .B(iw_word_c[33]), .Z(n27111)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(83[9] 84[65])
    defparam i1_2_lut_rep_788.init = 16'h2222;
    LUT4 i1_2_lut_3_lut (.A(iw_stb), .B(iw_word_c[33]), .C(\iw_word[32] ), 
         .Z(i_cmd_wr)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(83[9] 84[65])
    defparam i1_2_lut_3_lut.init = 16'h2020;
    LUT4 i19782_3_lut_3_lut (.A(iw_stb), .B(iw_word_c[33]), .C(wb_stb), 
         .Z(n22219)) /* synthesis lut_function=(A ((C)+!B)+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(83[9] 84[65])
    defparam i19782_3_lut_3_lut.init = 16'hf2f2;
    LUT4 i1_2_lut_rep_789 (.A(iw_word_c[33]), .B(iw_stb), .Z(n27112)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(83[9] 84[65])
    defparam i1_2_lut_rep_789.init = 16'h8888;
    LUT4 i1_2_lut_rep_572_3_lut (.A(iw_word_c[33]), .B(iw_stb), .C(\iw_word[32] ), 
         .Z(n26895)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(83[9] 84[65])
    defparam i1_2_lut_rep_572_3_lut.init = 16'h0808;
    LUT4 i1_2_lut_rep_460_3_lut_4_lut (.A(iw_word_c[33]), .B(iw_stb), .C(wb_cyc), 
         .D(\iw_word[32] ), .Z(dac_clk_p_c_enable_132)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(83[9] 84[65])
    defparam i1_2_lut_rep_460_3_lut_4_lut.init = 16'h0008;
    LUT4 i1_2_lut_3_lut_4_lut (.A(iw_word_c[33]), .B(iw_stb), .C(n29560), 
         .D(\iw_word[32] ), .Z(newaddr_N_990)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(83[9] 84[65])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0008;
    LUT4 i11012_2_lut (.A(\dec_bits[0] ), .B(\dec_bits[4] ), .Z(n14[0])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11012_2_lut.init = 16'h2222;
    LUT4 i11288_2_lut (.A(r_word[27]), .B(\dec_bits[4] ), .Z(n14[31])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11288_2_lut.init = 16'h2222;
    LUT4 i11289_2_lut (.A(r_word[26]), .B(\dec_bits[4] ), .Z(n14[30])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11289_2_lut.init = 16'h2222;
    LUT4 i11290_2_lut (.A(r_word[25]), .B(\dec_bits[4] ), .Z(n14[29])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11290_2_lut.init = 16'h2222;
    LUT4 i11291_2_lut (.A(r_word[24]), .B(\dec_bits[4] ), .Z(n14[28])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11291_2_lut.init = 16'h2222;
    LUT4 i11293_2_lut (.A(r_word[23]), .B(\dec_bits[4] ), .Z(n14[27])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11293_2_lut.init = 16'h2222;
    LUT4 i11294_2_lut (.A(r_word[22]), .B(\dec_bits[4] ), .Z(n14[26])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11294_2_lut.init = 16'h2222;
    LUT4 i11295_2_lut (.A(r_word[21]), .B(\dec_bits[4] ), .Z(n14[25])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11295_2_lut.init = 16'h2222;
    LUT4 i11296_2_lut (.A(r_word[20]), .B(\dec_bits[4] ), .Z(n14[24])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11296_2_lut.init = 16'h2222;
    LUT4 i11297_2_lut (.A(r_word[19]), .B(\dec_bits[4] ), .Z(n14[23])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11297_2_lut.init = 16'h2222;
    LUT4 i11299_2_lut (.A(r_word[18]), .B(\dec_bits[4] ), .Z(n14[22])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11299_2_lut.init = 16'h2222;
    LUT4 i11300_2_lut (.A(r_word[17]), .B(\dec_bits[4] ), .Z(n14[21])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11300_2_lut.init = 16'h2222;
    LUT4 i11301_2_lut (.A(r_word[16]), .B(\dec_bits[4] ), .Z(n14[20])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11301_2_lut.init = 16'h2222;
    LUT4 i11303_2_lut (.A(r_word[15]), .B(\dec_bits[4] ), .Z(n14[19])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11303_2_lut.init = 16'h2222;
    LUT4 i11304_2_lut (.A(r_word[14]), .B(\dec_bits[4] ), .Z(n14[18])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11304_2_lut.init = 16'h2222;
    LUT4 i11305_2_lut (.A(r_word[13]), .B(\dec_bits[4] ), .Z(n14[17])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11305_2_lut.init = 16'h2222;
    LUT4 i11306_2_lut (.A(r_word[12]), .B(\dec_bits[4] ), .Z(n14[16])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11306_2_lut.init = 16'h2222;
    FD1P3IX r_word__i33 (.D(\dec_bits[1] ), .SP(dac_clk_p_c_enable_350), 
            .CD(n29561), .CK(dac_clk_p_c), .Q(r_word[33])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i33.GSR = "DISABLED";
    FD1P3IX r_word__i32 (.D(\dec_bits[0] ), .SP(dac_clk_p_c_enable_350), 
            .CD(n29561), .CK(dac_clk_p_c), .Q(r_word[32])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i32.GSR = "DISABLED";
    LUT4 i11307_2_lut (.A(r_word[11]), .B(\dec_bits[4] ), .Z(n14[15])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11307_2_lut.init = 16'h2222;
    FD1P3IX r_word__i31 (.D(n14[31]), .SP(dac_clk_p_c_enable_381), .CD(n29561), 
            .CK(dac_clk_p_c), .Q(r_word[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i31.GSR = "DISABLED";
    LUT4 i11308_2_lut (.A(r_word[10]), .B(\dec_bits[4] ), .Z(n14[14])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(102[5:51])
    defparam i11308_2_lut.init = 16'h2222;
    FD1P3IX r_word__i30 (.D(n14[30]), .SP(dac_clk_p_c_enable_381), .CD(n29561), 
            .CK(dac_clk_p_c), .Q(r_word[30])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i30.GSR = "DISABLED";
    FD1P3IX r_word__i29 (.D(n14[29]), .SP(dac_clk_p_c_enable_381), .CD(n29561), 
            .CK(dac_clk_p_c), .Q(r_word[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i29.GSR = "DISABLED";
    FD1P3IX r_word__i28 (.D(n14[28]), .SP(dac_clk_p_c_enable_381), .CD(n29561), 
            .CK(dac_clk_p_c), .Q(r_word[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i28.GSR = "DISABLED";
    FD1P3IX r_word__i27 (.D(n14[27]), .SP(dac_clk_p_c_enable_381), .CD(n29561), 
            .CK(dac_clk_p_c), .Q(r_word[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i27.GSR = "DISABLED";
    FD1P3IX r_word__i26 (.D(n14[26]), .SP(dac_clk_p_c_enable_381), .CD(n29561), 
            .CK(dac_clk_p_c), .Q(r_word[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i26.GSR = "DISABLED";
    FD1P3IX r_word__i25 (.D(n14[25]), .SP(dac_clk_p_c_enable_381), .CD(n29561), 
            .CK(dac_clk_p_c), .Q(r_word[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i25.GSR = "DISABLED";
    FD1P3IX r_word__i24 (.D(n14[24]), .SP(dac_clk_p_c_enable_381), .CD(n29561), 
            .CK(dac_clk_p_c), .Q(r_word[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i24.GSR = "DISABLED";
    FD1P3IX r_word__i23 (.D(n14[23]), .SP(dac_clk_p_c_enable_381), .CD(n29561), 
            .CK(dac_clk_p_c), .Q(r_word[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i23.GSR = "DISABLED";
    FD1P3IX r_word__i22 (.D(n14[22]), .SP(dac_clk_p_c_enable_381), .CD(n29561), 
            .CK(dac_clk_p_c), .Q(r_word[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i22.GSR = "DISABLED";
    FD1P3IX r_word__i21 (.D(n14[21]), .SP(dac_clk_p_c_enable_381), .CD(n29561), 
            .CK(dac_clk_p_c), .Q(r_word[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i21.GSR = "DISABLED";
    FD1P3IX r_word__i20 (.D(n14[20]), .SP(dac_clk_p_c_enable_381), .CD(n29561), 
            .CK(dac_clk_p_c), .Q(r_word[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i20.GSR = "DISABLED";
    FD1P3IX r_word__i19 (.D(n14[19]), .SP(dac_clk_p_c_enable_381), .CD(n29561), 
            .CK(dac_clk_p_c), .Q(r_word[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i19.GSR = "DISABLED";
    FD1P3IX r_word__i18 (.D(n14[18]), .SP(dac_clk_p_c_enable_381), .CD(n29561), 
            .CK(dac_clk_p_c), .Q(r_word[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i18.GSR = "DISABLED";
    FD1P3IX r_word__i17 (.D(n14[17]), .SP(dac_clk_p_c_enable_381), .CD(n29561), 
            .CK(dac_clk_p_c), .Q(r_word[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i17.GSR = "DISABLED";
    FD1P3IX r_word__i16 (.D(n14[16]), .SP(dac_clk_p_c_enable_381), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i16.GSR = "DISABLED";
    FD1P3IX r_word__i15 (.D(n14[15]), .SP(dac_clk_p_c_enable_381), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i15.GSR = "DISABLED";
    FD1P3IX r_word__i14 (.D(n14[14]), .SP(dac_clk_p_c_enable_381), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i14.GSR = "DISABLED";
    FD1P3IX r_word__i13 (.D(n14[13]), .SP(dac_clk_p_c_enable_381), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i13.GSR = "DISABLED";
    FD1P3IX r_word__i12 (.D(n14[12]), .SP(dac_clk_p_c_enable_381), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i12.GSR = "DISABLED";
    FD1P3IX r_word__i11 (.D(n14[11]), .SP(dac_clk_p_c_enable_381), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i11.GSR = "DISABLED";
    FD1P3IX r_word__i10 (.D(n14[10]), .SP(dac_clk_p_c_enable_381), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i10.GSR = "DISABLED";
    FD1P3IX r_word__i9 (.D(n14[9]), .SP(dac_clk_p_c_enable_381), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i9.GSR = "DISABLED";
    FD1P3IX r_word__i8 (.D(n14[8]), .SP(dac_clk_p_c_enable_381), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i8.GSR = "DISABLED";
    FD1P3IX r_word__i7 (.D(n14[7]), .SP(dac_clk_p_c_enable_381), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i7.GSR = "DISABLED";
    FD1P3IX r_word__i6 (.D(n14[6]), .SP(dac_clk_p_c_enable_381), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i6.GSR = "DISABLED";
    FD1P3IX r_word__i5 (.D(n14[5]), .SP(dac_clk_p_c_enable_381), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i5.GSR = "DISABLED";
    FD1P3IX r_word__i4 (.D(n14[4]), .SP(dac_clk_p_c_enable_381), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i4.GSR = "DISABLED";
    FD1P3IX r_word__i3 (.D(n45), .SP(dac_clk_p_c_enable_381), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i3.GSR = "DISABLED";
    FD1P3IX r_word__i2 (.D(n46), .SP(dac_clk_p_c_enable_381), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i2.GSR = "DISABLED";
    FD1P3IX r_word__i1 (.D(n14[1]), .SP(dac_clk_p_c_enable_381), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(r_word[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=38, LSE_LLINE=99, LSE_RLINE=100 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(87[9] 103[6])
    defparam r_word__i1.GSR = "DISABLED";
    LUT4 i11006_2_lut_3_lut_4_lut (.A(\iw_word[32] ), .B(n27112), .C(wb_stb), 
         .D(wb_cyc), .Z(dac_clk_p_c_enable_446)) /* synthesis lut_function=(A (C)+!A (B (C+!(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbpack.v(83[9] 84[65])
    defparam i11006_2_lut_3_lut_4_lut.init = 16'hf0f4;
    
endmodule
//
// Verilog Description of module hbgenhex
//

module hbgenhex (hb_bits, \w_gx_char[0] , \w_gx_char[1] , \w_gx_char[2] , 
            \w_gx_char[3] , \w_gx_char[4] , \w_gx_char[5] , \w_gx_char[6] , 
            dac_clk_p_c, dac_clk_p_c_enable_308, GND_net, VCC_net, hx_stb, 
            w_reset, hb_busy, nl_busy, n29560, n26906, dac_clk_p_c_enable_194, 
            n11749) /* synthesis syn_module_defined=1 */ ;
    input [4:0]hb_bits;
    output \w_gx_char[0] ;
    output \w_gx_char[1] ;
    output \w_gx_char[2] ;
    output \w_gx_char[3] ;
    output \w_gx_char[4] ;
    output \w_gx_char[5] ;
    output \w_gx_char[6] ;
    input dac_clk_p_c;
    output dac_clk_p_c_enable_308;
    input GND_net;
    input VCC_net;
    output hx_stb;
    input w_reset;
    input hb_busy;
    input nl_busy;
    input n29560;
    input n26906;
    output dac_clk_p_c_enable_194;
    output n11749;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(28[49:58])
    
    wire dac_clk_p_c_enable_143, n20569;
    
    SP8KC mux_105 (.DI0(GND_net), .DI1(GND_net), .DI2(GND_net), .DI3(GND_net), 
          .DI4(GND_net), .DI5(GND_net), .DI6(GND_net), .DI7(GND_net), 
          .DI8(GND_net), .AD0(GND_net), .AD1(GND_net), .AD2(GND_net), 
          .AD3(hb_bits[0]), .AD4(hb_bits[1]), .AD5(hb_bits[2]), .AD6(hb_bits[3]), 
          .AD7(hb_bits[4]), .AD8(GND_net), .AD9(GND_net), .AD10(GND_net), 
          .AD11(GND_net), .AD12(GND_net), .CE(dac_clk_p_c_enable_308), 
          .OCE(VCC_net), .CLK(dac_clk_p_c), .WE(GND_net), .CS0(GND_net), 
          .CS1(GND_net), .CS2(GND_net), .RST(GND_net), .DO0(\w_gx_char[0] ), 
          .DO1(\w_gx_char[1] ), .DO2(\w_gx_char[2] ), .DO3(\w_gx_char[3] ), 
          .DO4(\w_gx_char[4] ), .DO5(\w_gx_char[5] ), .DO6(\w_gx_char[6] ));
    defparam mux_105.DATA_WIDTH = 9;
    defparam mux_105.REGMODE = "NOREG";
    defparam mux_105.CSDECODE = "0b000";
    defparam mux_105.WRITEMODE = "NORMAL";
    defparam mux_105.GSR = "DISABLED";
    defparam mux_105.RESETMODE = "ASYNC";
    defparam mux_105.ASYNC_RESET_RELEASE = "SYNC";
    defparam mux_105.INIT_DATA = "STATIC";
    defparam mux_105.INITVAL_00 = "0x01A0D01A0D0B44908A5401A0D01A0D0A641096520CC650C8630C4610723806E3606A340663206230";
    defparam mux_105.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_105.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_105.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_105.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_105.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_105.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_105.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_105.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_105.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_105.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_105.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_105.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_105.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_105.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_105.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_105.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_105.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_105.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_105.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_105.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_105.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_105.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_105.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_105.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_105.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_105.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_105.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_105.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_105.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_105.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam mux_105.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    FD1P3IX o_gx_stb_13 (.D(hb_busy), .SP(dac_clk_p_c_enable_143), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(hx_stb)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=29, LSE_LLINE=132, LSE_RLINE=133 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbgenhex.v(74[9] 78[21])
    defparam o_gx_stb_13.GSR = "DISABLED";
    LUT4 i22632_2_lut_rep_465 (.A(hx_stb), .B(nl_busy), .Z(dac_clk_p_c_enable_308)) /* synthesis lut_function=(!(A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(76[16:26])
    defparam i22632_2_lut_rep_465.init = 16'h7777;
    LUT4 i634_2_lut_3_lut (.A(hx_stb), .B(nl_busy), .C(n29560), .Z(dac_clk_p_c_enable_143)) /* synthesis lut_function=(((C)+!B)+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(76[16:26])
    defparam i634_2_lut_3_lut.init = 16'hf7f7;
    LUT4 i1_2_lut_3_lut_4_lut (.A(hx_stb), .B(nl_busy), .C(n29560), .D(n26906), 
         .Z(dac_clk_p_c_enable_194)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdeword.v(76[16:26])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hfff7;
    LUT4 i1_4_lut (.A(\w_gx_char[3] ), .B(\w_gx_char[0] ), .C(\w_gx_char[2] ), 
         .D(n20569), .Z(n11749)) /* synthesis lut_function=((((D)+!C)+!B)+!A) */ ;
    defparam i1_4_lut.init = 16'hff7f;
    LUT4 i1_4_lut_adj_130 (.A(\w_gx_char[1] ), .B(\w_gx_char[6] ), .C(\w_gx_char[4] ), 
         .D(\w_gx_char[5] ), .Z(n20569)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_130.init = 16'hfffe;
    
endmodule
//
// Verilog Description of module hbdechex
//

module hbdechex (dac_clk_p_c, dec_bits, w_reset, rx_stb, \rx_data[4] , 
            \rx_data[3] , \rx_data[1] , \rx_data[0] , \rx_data[5] , 
            n45, n46, \dec_bits[1] , \rx_data[2] , \rx_data[6] , n29561, 
            n29560, dac_clk_p_c_enable_381, dac_clk_p_c_enable_350, cmd_loaded, 
            o_pck_stb_N_765, dac_clk_p_c_enable_196, cmd_loaded_N_768) /* synthesis syn_module_defined=1 */ ;
    input dac_clk_p_c;
    output [4:0]dec_bits;
    output w_reset;
    input rx_stb;
    input \rx_data[4] ;
    input \rx_data[3] ;
    input \rx_data[1] ;
    input \rx_data[0] ;
    input \rx_data[5] ;
    output n45;
    output n46;
    output \dec_bits[1] ;
    input \rx_data[2] ;
    input \rx_data[6] ;
    output n29561;
    output n29560;
    output dac_clk_p_c_enable_381;
    output dac_clk_p_c_enable_350;
    input cmd_loaded;
    output o_pck_stb_N_765;
    output dac_clk_p_c_enable_196;
    output cmd_loaded_N_768;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(28[49:58])
    
    wire dec_stb, o_dh_stb_N_623;
    wire [4:0]o_dh_bits_4__N_596;
    
    wire o_reset_N_625, n21107, n21099, n20545, n52, n26710, n29498, 
        n27203, n27204, n27205, n26680, n26679, n49;
    wire [4:0]dec_bits_c;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbbus.v(69[13:21])
    
    wire n25973, n25972, n26711, n28761, n28760, n29465, n64, 
        n9, n27110, n27113, n20492, n27114, n43, n27115, n25971, 
        n26677, n26676, n26678, n25976, n25994, n25995, n20599, 
        n25993, n20521, n26896, n62, n20517, n24, n20246, n47, 
        n20509;
    
    FD1S3AX o_dh_stb_35 (.D(o_dh_stb_N_623), .CK(dac_clk_p_c), .Q(dec_stb)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=30, LSE_LLINE=93, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(57[9] 58[47])
    defparam o_dh_stb_35.GSR = "DISABLED";
    FD1S3AX o_dh_bits_i0 (.D(o_dh_bits_4__N_596[0]), .CK(dac_clk_p_c), .Q(dec_bits[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=30, LSE_LLINE=93, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(60[9] 100[5])
    defparam o_dh_bits_i0.GSR = "DISABLED";
    FD1S3AY o_reset_34 (.D(o_reset_N_625), .CK(dac_clk_p_c), .Q(w_reset)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=30, LSE_LLINE=93, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(53[9] 54[46])
    defparam o_reset_34.GSR = "DISABLED";
    LUT4 i_stb_I_0_58_4_lut (.A(rx_stb), .B(n21107), .C(n21099), .D(\rx_data[4] ), 
         .Z(o_dh_stb_N_623)) /* synthesis lut_function=(!((B (C (D)))+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(58[15:46])
    defparam i_stb_I_0_58_4_lut.init = 16'h2aaa;
    LUT4 i1_2_lut (.A(\rx_data[3] ), .B(\rx_data[1] ), .Z(n21099)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i1_4_lut (.A(n20545), .B(n52), .C(n26710), .D(n29498), .Z(o_dh_bits_4__N_596[0])) /* synthesis lut_function=(A (B+(C))+!A (B+(C+!(D)))) */ ;
    defparam i1_4_lut.init = 16'hfcfd;
    PFUMX i24781 (.BLUT(n27203), .ALUT(n27204), .C0(\rx_data[0] ), .Z(n27205));
    LUT4 n26680_bdd_4_lut (.A(n26680), .B(n26679), .C(\rx_data[5] ), .D(n49), 
         .Z(n26710)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;
    defparam n26680_bdd_4_lut.init = 16'hffca;
    LUT4 i1_2_lut_adj_113 (.A(dec_bits[4]), .B(dec_bits_c[3]), .Z(n45)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(60[9] 100[5])
    defparam i1_2_lut_adj_113.init = 16'h4444;
    LUT4 i1_2_lut_adj_114 (.A(dec_bits[4]), .B(dec_bits_c[2]), .Z(n46)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(60[9] 100[5])
    defparam i1_2_lut_adj_114.init = 16'h4444;
    LUT4 n25973_bdd_4_lut (.A(n25973), .B(n25972), .C(\rx_data[5] ), .D(\rx_data[1] ), 
         .Z(n26711)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam n25973_bdd_4_lut.init = 16'h00ca;
    LUT4 n28761_bdd_4_lut (.A(n28761), .B(\rx_data[3] ), .C(n28760), .D(\rx_data[4] ), 
         .Z(n29465)) /* synthesis lut_function=(A (C+!(D))+!A (B (C+!(D))+!B (C (D)))) */ ;
    defparam n28761_bdd_4_lut.init = 16'hf0ee;
    FD1S3AX o_dh_bits_i4 (.D(o_dh_bits_4__N_596[4]), .CK(dac_clk_p_c), .Q(dec_bits[4])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=30, LSE_LLINE=93, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(60[9] 100[5])
    defparam o_dh_bits_i4.GSR = "DISABLED";
    FD1S3AX o_dh_bits_i3 (.D(o_dh_bits_4__N_596[3]), .CK(dac_clk_p_c), .Q(dec_bits_c[3])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=30, LSE_LLINE=93, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(60[9] 100[5])
    defparam o_dh_bits_i3.GSR = "DISABLED";
    FD1S3AX o_dh_bits_i2 (.D(o_dh_bits_4__N_596[2]), .CK(dac_clk_p_c), .Q(dec_bits_c[2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=30, LSE_LLINE=93, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(60[9] 100[5])
    defparam o_dh_bits_i2.GSR = "DISABLED";
    FD1S3AX o_dh_bits_i1 (.D(o_dh_bits_4__N_596[1]), .CK(dac_clk_p_c), .Q(\dec_bits[1] )) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=30, LSE_LLINE=93, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(60[9] 100[5])
    defparam o_dh_bits_i1.GSR = "DISABLED";
    LUT4 i1_4_lut_4_lut_rep_825 (.A(\rx_data[5] ), .B(\rx_data[2] ), .C(\rx_data[1] ), 
         .D(\rx_data[0] ), .Z(n29498)) /* synthesis lut_function=(!((B (C (D))+!B !(C+(D)))+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(65[3] 99[10])
    defparam i1_4_lut_4_lut_rep_825.init = 16'h2aa8;
    LUT4 i1_2_lut_4_lut_4_lut (.A(\rx_data[5] ), .B(\rx_data[2] ), .C(\rx_data[1] ), 
         .D(\rx_data[0] ), .Z(n64)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C+(D)))+!A (B+(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(65[3] 99[10])
    defparam i1_2_lut_4_lut_4_lut.init = 16'h2ba8;
    LUT4 i1_2_lut_3_lut (.A(\rx_data[1] ), .B(\rx_data[0] ), .C(\rx_data[2] ), 
         .Z(n9)) /* synthesis lut_function=(A+(B+!(C))) */ ;
    defparam i1_2_lut_3_lut.init = 16'hefef;
    LUT4 i1_3_lut_rep_787 (.A(\rx_data[5] ), .B(\rx_data[6] ), .C(\rx_data[3] ), 
         .Z(n27110)) /* synthesis lut_function=(A+((C)+!B)) */ ;
    defparam i1_3_lut_rep_787.init = 16'hfbfb;
    LUT4 i18821_2_lut_rep_790 (.A(\rx_data[5] ), .B(\rx_data[4] ), .Z(n27113)) /* synthesis lut_function=(A (B)) */ ;
    defparam i18821_2_lut_rep_790.init = 16'h8888;
    LUT4 i1_3_lut_4_lut (.A(\rx_data[2] ), .B(\rx_data[0] ), .C(\rx_data[1] ), 
         .D(\rx_data[5] ), .Z(n20492)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(65[3] 99[10])
    defparam i1_3_lut_4_lut.init = 16'h0002;
    LUT4 i1_2_lut_rep_791 (.A(\rx_data[2] ), .B(\rx_data[1] ), .Z(n27114)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(65[3] 99[10])
    defparam i1_2_lut_rep_791.init = 16'heeee;
    LUT4 i1_3_lut_4_lut_adj_115 (.A(\rx_data[2] ), .B(\rx_data[1] ), .C(\rx_data[6] ), 
         .D(\rx_data[3] ), .Z(n43)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(65[3] 99[10])
    defparam i1_3_lut_4_lut_adj_115.init = 16'hfe00;
    LUT4 i1_2_lut_4_lut (.A(\rx_data[1] ), .B(\rx_data[2] ), .C(\rx_data[0] ), 
         .D(\rx_data[4] ), .Z(n20545)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C+(D)))) */ ;
    defparam i1_2_lut_4_lut.init = 16'hff10;
    LUT4 i1_2_lut_rep_792 (.A(\rx_data[5] ), .B(\rx_data[2] ), .Z(n27115)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_792.init = 16'h8888;
    LUT4 i1_3_lut_4_lut_adj_116 (.A(\rx_data[5] ), .B(\rx_data[2] ), .C(\rx_data[6] ), 
         .D(\rx_data[0] ), .Z(n21107)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_3_lut_4_lut_adj_116.init = 16'h8000;
    LUT4 rx_data_3__bdd_4_lut_25508 (.A(\rx_data[3] ), .B(\rx_data[6] ), 
         .C(\rx_data[0] ), .D(\rx_data[4] ), .Z(n25971)) /* synthesis lut_function=(A+(B (C+(D))+!B !(D))) */ ;
    defparam rx_data_3__bdd_4_lut_25508.init = 16'heefb;
    LUT4 rx_data_0__bdd_4_lut_24272 (.A(\rx_data[0] ), .B(\rx_data[6] ), 
         .C(\rx_data[4] ), .D(\rx_data[3] ), .Z(n25972)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam rx_data_0__bdd_4_lut_24272.init = 16'h0008;
    LUT4 rx_data_0__bdd_3_lut_24273 (.A(\rx_data[0] ), .B(\rx_data[2] ), 
         .C(\rx_data[4] ), .Z(n25973)) /* synthesis lut_function=(!(A (B+(C))+!A !(B (C)))) */ ;
    defparam rx_data_0__bdd_3_lut_24273.init = 16'h4242;
    PFUMX i24713 (.BLUT(n26677), .ALUT(n26676), .C0(\rx_data[2] ), .Z(n26678));
    LUT4 rx_data_2__bdd_3_lut (.A(\rx_data[2] ), .B(\rx_data[0] ), .C(\rx_data[1] ), 
         .Z(n25976)) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;
    defparam rx_data_2__bdd_3_lut.init = 16'h6a6a;
    LUT4 n967_bdd_2_lut_24271 (.A(n25994), .B(\rx_data[5] ), .Z(n25995)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam n967_bdd_2_lut_24271.init = 16'hbbbb;
    LUT4 rx_data_4__bdd_4_lut_24826 (.A(\rx_data[4] ), .B(\rx_data[2] ), 
         .C(\rx_data[1] ), .D(\rx_data[3] ), .Z(n25994)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;
    defparam rx_data_4__bdd_4_lut_24826.init = 16'hfe00;
    LUT4 n20599_bdd_4_lut_24270 (.A(n20599), .B(\rx_data[0] ), .C(\rx_data[2] ), 
         .D(\rx_data[1] ), .Z(n25993)) /* synthesis lut_function=(!((B (C (D))+!B !(C+(D)))+!A)) */ ;
    defparam n20599_bdd_4_lut_24270.init = 16'h2aa8;
    LUT4 n967_bdd_2_lut_26259 (.A(n29465), .B(\rx_data[5] ), .Z(o_dh_bits_4__N_596[4])) /* synthesis lut_function=(A+!(B)) */ ;
    defparam n967_bdd_2_lut_26259.init = 16'hbbbb;
    LUT4 rx_data_1__bdd_4_lut_25932 (.A(\rx_data[1] ), .B(\rx_data[3] ), 
         .C(\rx_data[6] ), .D(\rx_data[2] ), .Z(n28760)) /* synthesis lut_function=(A (B+(C))+!A (B (C+(D))+!B (C))) */ ;
    defparam rx_data_1__bdd_4_lut_25932.init = 16'hfcf8;
    LUT4 rx_data_1__bdd_4_lut (.A(\rx_data[1] ), .B(\rx_data[0] ), .C(\rx_data[6] ), 
         .D(\rx_data[2] ), .Z(n28761)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A !(B (C)+!B (C (D)))) */ ;
    defparam rx_data_1__bdd_4_lut.init = 16'h8f1f;
    FD1S3AY o_reset_34_rep_827 (.D(o_reset_N_625), .CK(dac_clk_p_c), .Q(n29561)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=30, LSE_LLINE=93, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(53[9] 54[46])
    defparam o_reset_34_rep_827.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_117 (.A(n20521), .B(n25995), .C(n26896), .D(\rx_data[6] ), 
         .Z(o_dh_bits_4__N_596[3])) /* synthesis lut_function=(A+(B (C+!(D))+!B (C (D)))) */ ;
    defparam i1_4_lut_adj_117.init = 16'hfaee;
    LUT4 i1_4_lut_adj_118 (.A(\rx_data[4] ), .B(n25993), .C(n64), .D(\rx_data[6] ), 
         .Z(n20521)) /* synthesis lut_function=(A (B)+!A (B+!(C (D)))) */ ;
    defparam i1_4_lut_adj_118.init = 16'hcddd;
    LUT4 i1_4_lut_adj_119 (.A(n20599), .B(n62), .C(n20517), .D(n25976), 
         .Z(o_dh_bits_4__N_596[2])) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C))) */ ;
    defparam i1_4_lut_adj_119.init = 16'hfefc;
    LUT4 i65_4_lut (.A(n64), .B(n24), .C(\rx_data[4] ), .D(n20492), 
         .Z(n62)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (B+((D)+!C))) */ ;
    defparam i65_4_lut.init = 16'hf5c5;
    LUT4 i1_4_lut_adj_120 (.A(n43), .B(n20246), .C(\rx_data[6] ), .D(n27113), 
         .Z(n20517)) /* synthesis lut_function=(A+(B+!(C+(D)))) */ ;
    defparam i1_4_lut_adj_120.init = 16'heeef;
    LUT4 i1_2_lut_adj_121 (.A(\rx_data[6] ), .B(n47), .Z(n24)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i1_2_lut_adj_121.init = 16'h2222;
    LUT4 i1_4_lut_adj_122 (.A(n27205), .B(n52), .C(n26711), .D(n20509), 
         .Z(o_dh_bits_4__N_596[1])) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_122.init = 16'hfffe;
    LUT4 i1_4_lut_adj_123 (.A(\rx_data[1] ), .B(n49), .C(\rx_data[5] ), 
         .D(n25971), .Z(n20509)) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B)) */ ;
    defparam i1_4_lut_adj_123.init = 16'hccec;
    FD1S3AY o_reset_34_rep_826 (.D(o_reset_N_625), .CK(dac_clk_p_c), .Q(n29560)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=11, LSE_RCOL=30, LSE_LLINE=93, LSE_RLINE=95 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(53[9] 54[46])
    defparam o_reset_34_rep_826.GSR = "DISABLED";
    LUT4 rx_data_5__bdd_4_lut_25890 (.A(\rx_data[5] ), .B(\rx_data[0] ), 
         .C(\rx_data[1] ), .D(\rx_data[2] ), .Z(n47)) /* synthesis lut_function=(!(A+!(B (C)+!B !(C (D)+!C !(D))))) */ ;
    defparam rx_data_5__bdd_4_lut_25890.init = 16'h4150;
    LUT4 rx_data_0__bdd_4_lut_25891 (.A(\rx_data[0] ), .B(\rx_data[3] ), 
         .C(\rx_data[4] ), .D(\rx_data[6] ), .Z(n26676)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B+(C+!(D))))) */ ;
    defparam rx_data_0__bdd_4_lut_25891.init = 16'h0120;
    LUT4 rx_data_0__bdd_3_lut_24715 (.A(\rx_data[0] ), .B(\rx_data[4] ), 
         .C(\rx_data[6] ), .Z(n26677)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam rx_data_0__bdd_3_lut_24715.init = 16'h0808;
    LUT4 n26678_bdd_3_lut (.A(n26678), .B(n26676), .C(\rx_data[1] ), .Z(n26679)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n26678_bdd_3_lut.init = 16'hcaca;
    LUT4 rx_data_0__bdd_3_lut_25894 (.A(\rx_data[0] ), .B(\rx_data[1] ), 
         .C(\rx_data[4] ), .Z(n26680)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam rx_data_0__bdd_3_lut_25894.init = 16'h8080;
    LUT4 i1_3_lut_4_lut_adj_124 (.A(\rx_data[4] ), .B(n27110), .C(rx_stb), 
         .D(n9), .Z(o_reset_N_625)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(92[3:8])
    defparam i1_3_lut_4_lut_adj_124.init = 16'h0020;
    LUT4 i1_2_lut_rep_603 (.A(n29560), .B(dec_stb), .Z(dac_clk_p_c_enable_381)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(53[9] 54[46])
    defparam i1_2_lut_rep_603.init = 16'heeee;
    LUT4 i8107_2_lut_3_lut (.A(n29560), .B(dec_stb), .C(dec_bits[4]), 
         .Z(dac_clk_p_c_enable_350)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(53[9] 54[46])
    defparam i8107_2_lut_3_lut.init = 16'he0e0;
    LUT4 i1_3_lut_4_lut_adj_125 (.A(\rx_data[3] ), .B(n27114), .C(n27113), 
         .D(\rx_data[6] ), .Z(n49)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (C+(D)))) */ ;
    defparam i1_3_lut_4_lut_adj_125.init = 16'h008f;
    LUT4 i1_3_lut_rep_573 (.A(n47), .B(\rx_data[3] ), .C(\rx_data[4] ), 
         .Z(n26896)) /* synthesis lut_function=(A (B)+!A (B+(C))) */ ;
    defparam i1_3_lut_rep_573.init = 16'hdcdc;
    LUT4 i1_2_lut_4_lut_adj_126 (.A(n47), .B(\rx_data[3] ), .C(\rx_data[4] ), 
         .D(\rx_data[6] ), .Z(n52)) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C (D)))) */ ;
    defparam i1_2_lut_4_lut_adj_126.init = 16'hdc00;
    LUT4 i83_4_lut_then_4_lut (.A(\rx_data[2] ), .B(\rx_data[4] ), .C(\rx_data[5] ), 
         .D(\rx_data[1] ), .Z(n27204)) /* synthesis lut_function=(!(A (B+!((D)+!C))+!A (C+!(D)))) */ ;
    defparam i83_4_lut_then_4_lut.init = 16'h2702;
    LUT4 i83_4_lut_else_4_lut (.A(\rx_data[2] ), .B(\rx_data[4] ), .C(\rx_data[5] ), 
         .D(\rx_data[1] ), .Z(n27203)) /* synthesis lut_function=(!(A (B+(C))+!A (B+(C (D))))) */ ;
    defparam i83_4_lut_else_4_lut.init = 16'h0313;
    LUT4 i1_2_lut_3_lut_adj_127 (.A(dec_stb), .B(dec_bits[4]), .C(cmd_loaded), 
         .Z(o_pck_stb_N_765)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(60[9] 100[5])
    defparam i1_2_lut_3_lut_adj_127.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_128 (.A(dec_stb), .B(dec_bits[4]), .C(n29560), 
         .Z(dac_clk_p_c_enable_196)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(60[9] 100[5])
    defparam i1_2_lut_3_lut_adj_128.init = 16'hf8f8;
    LUT4 i2_3_lut_4_lut (.A(dec_stb), .B(dec_bits[4]), .C(dec_bits_c[2]), 
         .D(dec_bits_c[3]), .Z(cmd_loaded_N_768)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(60[9] 100[5])
    defparam i2_3_lut_4_lut.init = 16'h0008;
    LUT4 i1_3_lut_4_lut_adj_129 (.A(\rx_data[6] ), .B(\rx_data[3] ), .C(\rx_data[4] ), 
         .D(n27115), .Z(n20246)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbdechex.v(87[3:8])
    defparam i1_3_lut_4_lut_adj_129.init = 16'h1000;
    LUT4 rx_data_4__bdd_3_lut_4_lut (.A(\rx_data[5] ), .B(\rx_data[6] ), 
         .C(\rx_data[3] ), .D(\rx_data[4] ), .Z(n20599)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam rx_data_4__bdd_3_lut_4_lut.init = 16'h0008;
    
endmodule
//
// Verilog Description of module hbnewline
//

module hbnewline (hx_stb, nl_busy, \w_gx_char[5] , dac_clk_p_c, n29561, 
            \w_gx_char[1] , \w_gx_char[6] , n11749, tx_busy, n26910, 
            \lcl_data[1] , \lcl_data_7__N_511[0] , \lcl_data[4] , \lcl_data_7__N_511[3] , 
            w_reset, \lcl_data[5] , \lcl_data_7__N_511[4] , \lcl_data[6] , 
            \lcl_data_7__N_511[5] , zero_baud_counter, dac_clk_p_c_enable_322, 
            \lcl_data[7] , \lcl_data_7__N_511[6] , \lcl_data[3] , \lcl_data_7__N_511[2] , 
            \lcl_data[2] , \lcl_data_7__N_511[1] , o_busy_N_536, \state[0] , 
            n17844, \w_gx_char[2] , \w_gx_char[0] , \w_gx_char[4] , 
            n29560, \w_gx_char[3] ) /* synthesis syn_module_defined=1 */ ;
    input hx_stb;
    output nl_busy;
    input \w_gx_char[5] ;
    input dac_clk_p_c;
    input n29561;
    input \w_gx_char[1] ;
    input \w_gx_char[6] ;
    input n11749;
    input tx_busy;
    output n26910;
    input \lcl_data[1] ;
    output \lcl_data_7__N_511[0] ;
    input \lcl_data[4] ;
    output \lcl_data_7__N_511[3] ;
    input w_reset;
    input \lcl_data[5] ;
    output \lcl_data_7__N_511[4] ;
    input \lcl_data[6] ;
    output \lcl_data_7__N_511[5] ;
    input zero_baud_counter;
    output dac_clk_p_c_enable_322;
    input \lcl_data[7] ;
    output \lcl_data_7__N_511[6] ;
    input \lcl_data[3] ;
    output \lcl_data_7__N_511[2] ;
    input \lcl_data[2] ;
    output \lcl_data_7__N_511[1] ;
    input o_busy_N_536;
    input \state[0] ;
    output n17844;
    input \w_gx_char[2] ;
    input \w_gx_char[0] ;
    input \w_gx_char[4] ;
    input n29560;
    input \w_gx_char[3] ;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(28[49:58])
    wire [6:0]n32;
    wire [6:0]o_nl_byte_6__N_1302;
    
    wire last_cr, last_cr_N_1323, tx_stb, o_nl_stb_N_1315, cr_state_N_1331, 
        n27227, n27228;
    wire [7:0]tx_data;   // d:/documents/git_local/fm_modulator/rtl/top.v(59[12:19])
    
    wire dac_clk_p_c_enable_199;
    wire [6:0]o_nl_byte_6__N_1295;
    
    wire cr_state, loaded, n26763, n24528, n24527, n26883;
    
    LUT4 i10789_3_lut_4_lut (.A(hx_stb), .B(nl_busy), .C(\w_gx_char[5] ), 
         .D(n32[4]), .Z(o_nl_byte_6__N_1302[5])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(90[16:37])
    defparam i10789_3_lut_4_lut.init = 16'hfd20;
    FD1S3JX last_cr_45 (.D(last_cr_N_1323), .CK(dac_clk_p_c), .PD(n29561), 
            .Q(last_cr)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=12, LSE_RCOL=40, LSE_LLINE=138, LSE_RLINE=139 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam last_cr_45.GSR = "DISABLED";
    FD1S3IX o_nl_stb_46 (.D(o_nl_stb_N_1315), .CK(dac_clk_p_c), .CD(n29561), 
            .Q(tx_stb)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=12, LSE_RCOL=40, LSE_LLINE=138, LSE_RLINE=139 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam o_nl_stb_46.GSR = "DISABLED";
    LUT4 i10792_3_lut_4_lut (.A(hx_stb), .B(nl_busy), .C(\w_gx_char[1] ), 
         .D(last_cr), .Z(o_nl_byte_6__N_1302[1])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(90[16:37])
    defparam i10792_3_lut_4_lut.init = 16'hfd20;
    LUT4 mux_24_i7_3_lut_4_lut (.A(hx_stb), .B(nl_busy), .C(\w_gx_char[6] ), 
         .D(n32[4]), .Z(o_nl_byte_6__N_1302[6])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(90[16:37])
    defparam mux_24_i7_3_lut_4_lut.init = 16'hfd20;
    LUT4 cr_state_I_41_3_lut_4_lut (.A(hx_stb), .B(nl_busy), .C(n11749), 
         .D(last_cr), .Z(cr_state_N_1331)) /* synthesis lut_function=(!(A (B (D)+!B (C))+!A (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(90[16:37])
    defparam cr_state_I_41_3_lut_4_lut.init = 16'h02df;
    PFUMX i24797 (.BLUT(n27227), .ALUT(n27228), .C0(last_cr), .Z(last_cr_N_1323));
    LUT4 i1_2_lut_rep_587 (.A(tx_stb), .B(tx_busy), .Z(n26910)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam i1_2_lut_rep_587.init = 16'h2222;
    LUT4 lcl_data_7__I_0_i1_3_lut_4_lut (.A(tx_stb), .B(tx_busy), .C(tx_data[0]), 
         .D(\lcl_data[1] ), .Z(\lcl_data_7__N_511[0] )) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam lcl_data_7__I_0_i1_3_lut_4_lut.init = 16'hfd20;
    LUT4 lcl_data_7__I_0_i4_3_lut_4_lut (.A(tx_stb), .B(tx_busy), .C(tx_data[3]), 
         .D(\lcl_data[4] ), .Z(\lcl_data_7__N_511[3] )) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam lcl_data_7__I_0_i4_3_lut_4_lut.init = 16'hfd20;
    FD1P3JX o_nl_byte_i2 (.D(o_nl_byte_6__N_1302[1]), .SP(dac_clk_p_c_enable_199), 
            .PD(w_reset), .CK(dac_clk_p_c), .Q(tx_data[1])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=12, LSE_RCOL=40, LSE_LLINE=138, LSE_RLINE=139 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam o_nl_byte_i2.GSR = "DISABLED";
    FD1P3JX o_nl_byte_i3 (.D(o_nl_byte_6__N_1302[2]), .SP(dac_clk_p_c_enable_199), 
            .PD(w_reset), .CK(dac_clk_p_c), .Q(tx_data[2])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=12, LSE_RCOL=40, LSE_LLINE=138, LSE_RLINE=139 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam o_nl_byte_i3.GSR = "DISABLED";
    FD1P3AY o_nl_byte_i4 (.D(o_nl_byte_6__N_1295[3]), .SP(dac_clk_p_c_enable_199), 
            .CK(dac_clk_p_c), .Q(tx_data[3])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=12, LSE_RCOL=40, LSE_LLINE=138, LSE_RLINE=139 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam o_nl_byte_i4.GSR = "DISABLED";
    FD1P3JX o_nl_byte_i5 (.D(o_nl_byte_6__N_1302[4]), .SP(dac_clk_p_c_enable_199), 
            .PD(w_reset), .CK(dac_clk_p_c), .Q(tx_data[4])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=12, LSE_RCOL=40, LSE_LLINE=138, LSE_RLINE=139 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam o_nl_byte_i5.GSR = "DISABLED";
    FD1P3JX o_nl_byte_i6 (.D(o_nl_byte_6__N_1302[5]), .SP(dac_clk_p_c_enable_199), 
            .PD(w_reset), .CK(dac_clk_p_c), .Q(tx_data[5])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=12, LSE_RCOL=40, LSE_LLINE=138, LSE_RLINE=139 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam o_nl_byte_i6.GSR = "DISABLED";
    FD1P3JX o_nl_byte_i7 (.D(o_nl_byte_6__N_1302[6]), .SP(dac_clk_p_c_enable_199), 
            .PD(w_reset), .CK(dac_clk_p_c), .Q(tx_data[6])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=12, LSE_RCOL=40, LSE_LLINE=138, LSE_RLINE=139 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam o_nl_byte_i7.GSR = "DISABLED";
    FD1P3IX cr_state_44 (.D(cr_state_N_1331), .SP(dac_clk_p_c_enable_199), 
            .CD(n29561), .CK(dac_clk_p_c), .Q(cr_state)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=12, LSE_RCOL=40, LSE_LLINE=138, LSE_RLINE=139 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam cr_state_44.GSR = "DISABLED";
    FD1P3IX loaded_47 (.D(n26763), .SP(dac_clk_p_c_enable_199), .CD(n29561), 
            .CK(dac_clk_p_c), .Q(loaded)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=12, LSE_RCOL=40, LSE_LLINE=138, LSE_RLINE=139 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam loaded_47.GSR = "DISABLED";
    FD1P3JX o_nl_byte_i1 (.D(o_nl_byte_6__N_1302[0]), .SP(dac_clk_p_c_enable_199), 
            .PD(n29561), .CK(dac_clk_p_c), .Q(tx_data[0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=12, LSE_RCOL=40, LSE_LLINE=138, LSE_RLINE=139 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam o_nl_byte_i1.GSR = "DISABLED";
    LUT4 lcl_data_7__I_0_i5_3_lut_4_lut (.A(tx_stb), .B(tx_busy), .C(tx_data[4]), 
         .D(\lcl_data[5] ), .Z(\lcl_data_7__N_511[4] )) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam lcl_data_7__I_0_i5_3_lut_4_lut.init = 16'hfd20;
    LUT4 lcl_data_7__I_0_i6_3_lut_4_lut (.A(tx_stb), .B(tx_busy), .C(tx_data[5]), 
         .D(\lcl_data[6] ), .Z(\lcl_data_7__N_511[5] )) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam lcl_data_7__I_0_i6_3_lut_4_lut.init = 16'hfd20;
    LUT4 i561_2_lut_3_lut (.A(tx_stb), .B(tx_busy), .C(zero_baud_counter), 
         .Z(dac_clk_p_c_enable_322)) /* synthesis lut_function=(A ((C)+!B)+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam i561_2_lut_3_lut.init = 16'hf2f2;
    LUT4 lcl_data_7__I_0_i7_3_lut_4_lut (.A(tx_stb), .B(tx_busy), .C(tx_data[6]), 
         .D(\lcl_data[7] ), .Z(\lcl_data_7__N_511[6] )) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam lcl_data_7__I_0_i7_3_lut_4_lut.init = 16'hfd20;
    LUT4 lcl_data_7__I_0_i3_3_lut_4_lut (.A(tx_stb), .B(tx_busy), .C(tx_data[2]), 
         .D(\lcl_data[3] ), .Z(\lcl_data_7__N_511[2] )) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam lcl_data_7__I_0_i3_3_lut_4_lut.init = 16'hfd20;
    LUT4 lcl_data_7__I_0_i2_3_lut_4_lut (.A(tx_stb), .B(tx_busy), .C(tx_data[1]), 
         .D(\lcl_data[2] ), .Z(\lcl_data_7__N_511[1] )) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam lcl_data_7__I_0_i2_3_lut_4_lut.init = 16'hfd20;
    LUT4 tx_stb_bdd_3_lut (.A(hx_stb), .B(last_cr), .C(cr_state), .Z(n24528)) /* synthesis lut_function=(A (B+!(C))+!A ((C)+!B)) */ ;
    defparam tx_stb_bdd_3_lut.init = 16'hdbdb;
    LUT4 state_546_mux_6_i1_3_lut_4_lut (.A(tx_stb), .B(tx_busy), .C(o_busy_N_536), 
         .D(\state[0] ), .Z(n17844)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam state_546_mux_6_i1_3_lut_4_lut.init = 16'hd0df;
    LUT4 tx_stb_bdd_2_lut (.A(tx_stb), .B(hx_stb), .Z(n24527)) /* synthesis lut_function=(A+(B)) */ ;
    defparam tx_stb_bdd_2_lut.init = 16'heeee;
    LUT4 i1_2_lut (.A(last_cr), .B(cr_state), .Z(n32[4])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(82[9] 120[6])
    defparam i1_2_lut.init = 16'h2222;
    LUT4 i1_3_lut_4_lut (.A(last_cr), .B(n26883), .C(cr_state), .D(\w_gx_char[2] ), 
         .Z(o_nl_byte_6__N_1302[2])) /* synthesis lut_function=(A (B (D)+!B !(C))+!A ((D)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(97[12] 120[6])
    defparam i1_3_lut_4_lut.init = 16'hdf13;
    LUT4 i1_3_lut_4_lut_adj_110 (.A(last_cr), .B(n26883), .C(cr_state), 
         .D(\w_gx_char[0] ), .Z(o_nl_byte_6__N_1302[0])) /* synthesis lut_function=(A (B (D)+!B !(C))+!A ((D)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(97[12] 120[6])
    defparam i1_3_lut_4_lut_adj_110.init = 16'hdf13;
    LUT4 i_stb_I_0_2_lut_rep_560 (.A(hx_stb), .B(nl_busy), .Z(n26883)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(90[16:37])
    defparam i_stb_I_0_2_lut_rep_560.init = 16'h2222;
    LUT4 mux_24_i5_3_lut_4_lut (.A(hx_stb), .B(nl_busy), .C(\w_gx_char[4] ), 
         .D(n32[4]), .Z(o_nl_byte_6__N_1302[4])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(90[16:37])
    defparam mux_24_i5_3_lut_4_lut.init = 16'hfd20;
    LUT4 i1_3_lut_4_lut_adj_111 (.A(hx_stb), .B(nl_busy), .C(n29560), 
         .D(\w_gx_char[3] ), .Z(o_nl_byte_6__N_1295[3])) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(90[16:37])
    defparam i1_3_lut_4_lut_adj_111.init = 16'hfffd;
    LUT4 i1_3_lut_4_lut_adj_112 (.A(hx_stb), .B(nl_busy), .C(n29560), 
         .D(tx_busy), .Z(dac_clk_p_c_enable_199)) /* synthesis lut_function=(A ((C+!(D))+!B)+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(90[16:37])
    defparam i1_3_lut_4_lut_adj_112.init = 16'hf2ff;
    LUT4 i11027_3_lut_rep_440_4_lut (.A(hx_stb), .B(nl_busy), .C(cr_state), 
         .D(last_cr), .Z(n26763)) /* synthesis lut_function=(A ((C (D))+!B)+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(90[16:37])
    defparam i11027_3_lut_rep_440_4_lut.init = 16'hf222;
    LUT4 i21079_4_lut (.A(cr_state), .B(tx_stb), .C(tx_busy), .D(loaded), 
         .Z(nl_busy)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(123[21] 124[30])
    defparam i21079_4_lut.init = 16'hca0a;
    LUT4 last_cr_I_39_4_lut_then_3_lut (.A(n11749), .B(hx_stb), .C(nl_busy), 
         .Z(n27228)) /* synthesis lut_function=(((C)+!B)+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(97[12] 120[6])
    defparam last_cr_I_39_4_lut_then_3_lut.init = 16'hf7f7;
    LUT4 last_cr_I_39_4_lut_else_3_lut (.A(n11749), .B(tx_busy), .C(hx_stb), 
         .D(nl_busy), .Z(n27227)) /* synthesis lut_function=(!(A (B+(C))+!A (B ((D)+!C)+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbnewline.v(97[12] 120[6])
    defparam last_cr_I_39_4_lut_else_3_lut.init = 16'h0353;
    PFUMX i22878 (.BLUT(n24528), .ALUT(n24527), .C0(tx_busy), .Z(o_nl_stb_N_1315));
    
endmodule
//
// Verilog Description of module hbints
//

module hbints (int_word, dac_clk_p_c, dac_clk_p_c_enable_416, n12748, 
            ow_word, n29560, n26940, n26903, int_stb, ow_stb, n29561) /* synthesis syn_module_defined=1 */ ;
    output [33:0]int_word;
    input dac_clk_p_c;
    input dac_clk_p_c_enable_416;
    input n12748;
    input [33:0]ow_word;
    input n29560;
    output n26940;
    input n26903;
    output int_stb;
    input ow_stb;
    input n29561;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(28[49:58])
    
    wire dac_clk_p_c_enable_410, loaded, dac_clk_p_c_enable_409;
    
    FD1P3IX o_int_word_i9 (.D(ow_word[9]), .SP(dac_clk_p_c_enable_416), 
            .CD(n12748), .CK(dac_clk_p_c), .Q(int_word[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i9.GSR = "DISABLED";
    FD1P3JX o_int_word_i33 (.D(ow_word[33]), .SP(dac_clk_p_c_enable_416), 
            .PD(n12748), .CK(dac_clk_p_c), .Q(int_word[33])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i33.GSR = "DISABLED";
    FD1P3JX o_int_word_i32 (.D(ow_word[32]), .SP(dac_clk_p_c_enable_416), 
            .PD(n12748), .CK(dac_clk_p_c), .Q(int_word[32])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i32.GSR = "DISABLED";
    LUT4 i1_2_lut_3_lut_4_lut (.A(n29560), .B(n26940), .C(n26903), .D(int_stb), 
         .Z(dac_clk_p_c_enable_410)) /* synthesis lut_function=(A+(B+!(C+!(D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'hefee;
    LUT4 i1_3_lut_4_lut (.A(n29560), .B(n26940), .C(loaded), .D(n26903), 
         .Z(dac_clk_p_c_enable_409)) /* synthesis lut_function=(A+(B+!(C (D)))) */ ;
    defparam i1_3_lut_4_lut.init = 16'hefff;
    FD1P3IX o_int_word_i31 (.D(ow_word[31]), .SP(dac_clk_p_c_enable_416), 
            .CD(n12748), .CK(dac_clk_p_c), .Q(int_word[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i31.GSR = "DISABLED";
    FD1P3JX o_int_word_i30 (.D(ow_word[30]), .SP(dac_clk_p_c_enable_416), 
            .PD(n12748), .CK(dac_clk_p_c), .Q(int_word[30])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i30.GSR = "DISABLED";
    LUT4 i_stb_I_0_3_lut_rep_617 (.A(ow_stb), .B(int_stb), .C(loaded), 
         .Z(n26940)) /* synthesis lut_function=(!((B (C))+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(93[12:34])
    defparam i_stb_I_0_3_lut_rep_617.init = 16'h2a2a;
    FD1P3IX o_int_word_i8 (.D(ow_word[8]), .SP(dac_clk_p_c_enable_416), 
            .CD(n12748), .CK(dac_clk_p_c), .Q(int_word[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i8.GSR = "DISABLED";
    FD1P3IX o_int_word_i29 (.D(ow_word[29]), .SP(dac_clk_p_c_enable_416), 
            .CD(n12748), .CK(dac_clk_p_c), .Q(int_word[29])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i29.GSR = "DISABLED";
    FD1P3IX o_int_word_i28 (.D(ow_word[28]), .SP(dac_clk_p_c_enable_416), 
            .CD(n12748), .CK(dac_clk_p_c), .Q(int_word[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i28.GSR = "DISABLED";
    FD1P3IX o_int_word_i7 (.D(ow_word[7]), .SP(dac_clk_p_c_enable_416), 
            .CD(n12748), .CK(dac_clk_p_c), .Q(int_word[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i7.GSR = "DISABLED";
    FD1P3IX o_int_word_i27 (.D(ow_word[27]), .SP(dac_clk_p_c_enable_416), 
            .CD(n12748), .CK(dac_clk_p_c), .Q(int_word[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i27.GSR = "DISABLED";
    FD1P3IX o_int_word_i6 (.D(ow_word[6]), .SP(dac_clk_p_c_enable_416), 
            .CD(n12748), .CK(dac_clk_p_c), .Q(int_word[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i6.GSR = "DISABLED";
    FD1P3IX o_int_word_i26 (.D(ow_word[26]), .SP(dac_clk_p_c_enable_416), 
            .CD(n12748), .CK(dac_clk_p_c), .Q(int_word[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i26.GSR = "DISABLED";
    FD1P3IX o_int_word_i5 (.D(ow_word[5]), .SP(dac_clk_p_c_enable_416), 
            .CD(n12748), .CK(dac_clk_p_c), .Q(int_word[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i5.GSR = "DISABLED";
    FD1P3IX o_int_word_i4 (.D(ow_word[4]), .SP(dac_clk_p_c_enable_416), 
            .CD(n12748), .CK(dac_clk_p_c), .Q(int_word[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i4.GSR = "DISABLED";
    FD1P3IX o_int_word_i25 (.D(ow_word[25]), .SP(dac_clk_p_c_enable_416), 
            .CD(n12748), .CK(dac_clk_p_c), .Q(int_word[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i25.GSR = "DISABLED";
    FD1P3IX o_int_word_i24 (.D(ow_word[24]), .SP(dac_clk_p_c_enable_416), 
            .CD(n12748), .CK(dac_clk_p_c), .Q(int_word[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i24.GSR = "DISABLED";
    FD1P3IX o_int_word_i3 (.D(ow_word[3]), .SP(dac_clk_p_c_enable_416), 
            .CD(n12748), .CK(dac_clk_p_c), .Q(int_word[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i3.GSR = "DISABLED";
    FD1P3IX o_int_word_i23 (.D(ow_word[23]), .SP(dac_clk_p_c_enable_416), 
            .CD(n12748), .CK(dac_clk_p_c), .Q(int_word[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i23.GSR = "DISABLED";
    FD1P3IX o_int_word_i2 (.D(ow_word[2]), .SP(dac_clk_p_c_enable_416), 
            .CD(n12748), .CK(dac_clk_p_c), .Q(int_word[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i2.GSR = "DISABLED";
    FD1P3IX o_int_word_i22 (.D(ow_word[22]), .SP(dac_clk_p_c_enable_416), 
            .CD(n12748), .CK(dac_clk_p_c), .Q(int_word[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i22.GSR = "DISABLED";
    FD1P3IX o_int_word_i1 (.D(ow_word[1]), .SP(dac_clk_p_c_enable_416), 
            .CD(n12748), .CK(dac_clk_p_c), .Q(int_word[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i1.GSR = "DISABLED";
    FD1P3IX o_int_word_i0 (.D(ow_word[0]), .SP(dac_clk_p_c_enable_416), 
            .CD(n12748), .CK(dac_clk_p_c), .Q(int_word[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i0.GSR = "DISABLED";
    FD1P3IX o_int_word_i21 (.D(ow_word[21]), .SP(dac_clk_p_c_enable_416), 
            .CD(n12748), .CK(dac_clk_p_c), .Q(int_word[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i21.GSR = "DISABLED";
    FD1P3IX o_int_word_i20 (.D(ow_word[20]), .SP(dac_clk_p_c_enable_416), 
            .CD(n12748), .CK(dac_clk_p_c), .Q(int_word[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i20.GSR = "DISABLED";
    FD1P3IX o_int_word_i19 (.D(ow_word[19]), .SP(dac_clk_p_c_enable_416), 
            .CD(n12748), .CK(dac_clk_p_c), .Q(int_word[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i19.GSR = "DISABLED";
    FD1P3IX o_int_word_i18 (.D(ow_word[18]), .SP(dac_clk_p_c_enable_416), 
            .CD(n12748), .CK(dac_clk_p_c), .Q(int_word[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i18.GSR = "DISABLED";
    FD1P3IX o_int_word_i17 (.D(ow_word[17]), .SP(dac_clk_p_c_enable_416), 
            .CD(n12748), .CK(dac_clk_p_c), .Q(int_word[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i17.GSR = "DISABLED";
    FD1P3IX o_int_word_i16 (.D(ow_word[16]), .SP(dac_clk_p_c_enable_416), 
            .CD(n12748), .CK(dac_clk_p_c), .Q(int_word[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i16.GSR = "DISABLED";
    FD1P3IX o_int_word_i15 (.D(ow_word[15]), .SP(dac_clk_p_c_enable_416), 
            .CD(n12748), .CK(dac_clk_p_c), .Q(int_word[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i15.GSR = "DISABLED";
    FD1P3IX o_int_word_i14 (.D(ow_word[14]), .SP(dac_clk_p_c_enable_416), 
            .CD(n12748), .CK(dac_clk_p_c), .Q(int_word[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i14.GSR = "DISABLED";
    FD1P3IX o_int_stb_58 (.D(n26940), .SP(dac_clk_p_c_enable_409), .CD(n29561), 
            .CK(dac_clk_p_c), .Q(int_stb)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(90[9] 98[22])
    defparam o_int_stb_58.GSR = "DISABLED";
    FD1P3IX loaded_57 (.D(n26940), .SP(dac_clk_p_c_enable_410), .CD(n29561), 
            .CK(dac_clk_p_c), .Q(loaded)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(81[9] 87[19])
    defparam loaded_57.GSR = "DISABLED";
    FD1P3IX o_int_word_i13 (.D(ow_word[13]), .SP(dac_clk_p_c_enable_416), 
            .CD(n12748), .CK(dac_clk_p_c), .Q(int_word[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i13.GSR = "DISABLED";
    FD1P3IX o_int_word_i12 (.D(ow_word[12]), .SP(dac_clk_p_c_enable_416), 
            .CD(n12748), .CK(dac_clk_p_c), .Q(int_word[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i12.GSR = "DISABLED";
    FD1P3IX o_int_word_i11 (.D(ow_word[11]), .SP(dac_clk_p_c_enable_416), 
            .CD(n12748), .CK(dac_clk_p_c), .Q(int_word[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i11.GSR = "DISABLED";
    FD1P3IX o_int_word_i10 (.D(ow_word[10]), .SP(dac_clk_p_c_enable_416), 
            .CD(n12748), .CK(dac_clk_p_c), .Q(int_word[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=32, LSE_LLINE=114, LSE_RLINE=116 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbints.v(102[9] 112[6])
    defparam o_int_word_i10.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module hbidle
//

module hbidle (idl_word, dac_clk_p_c, int_word, idl_stb, w_reset, 
            hb_busy, n26903, int_stb, n29560, n26940, n12748, dac_clk_p_c_enable_416) /* synthesis syn_module_defined=1 */ ;
    output [33:0]idl_word;
    input dac_clk_p_c;
    input [33:0]int_word;
    output idl_stb;
    input w_reset;
    input hb_busy;
    output n26903;
    input int_stb;
    input n29560;
    input n26940;
    output n12748;
    output dac_clk_p_c_enable_416;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(28[49:58])
    
    wire dac_clk_p_c_enable_346, n12778, dac_clk_p_c_enable_195, n26785;
    
    FD1P3IX o_idl_word_i10 (.D(int_word[10]), .SP(dac_clk_p_c_enable_346), 
            .CD(n12778), .CK(dac_clk_p_c), .Q(idl_word[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i10.GSR = "DISABLED";
    FD1P3IX o_idl_word_i9 (.D(int_word[9]), .SP(dac_clk_p_c_enable_346), 
            .CD(n12778), .CK(dac_clk_p_c), .Q(idl_word[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i9.GSR = "DISABLED";
    FD1P3IX o_idl_word_i8 (.D(int_word[8]), .SP(dac_clk_p_c_enable_346), 
            .CD(n12778), .CK(dac_clk_p_c), .Q(idl_word[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i8.GSR = "DISABLED";
    FD1P3IX o_idl_word_i7 (.D(int_word[7]), .SP(dac_clk_p_c_enable_346), 
            .CD(n12778), .CK(dac_clk_p_c), .Q(idl_word[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i7.GSR = "DISABLED";
    FD1P3IX o_idl_word_i6 (.D(int_word[6]), .SP(dac_clk_p_c_enable_346), 
            .CD(n12778), .CK(dac_clk_p_c), .Q(idl_word[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i6.GSR = "DISABLED";
    FD1P3IX o_idl_word_i5 (.D(int_word[5]), .SP(dac_clk_p_c_enable_346), 
            .CD(n12778), .CK(dac_clk_p_c), .Q(idl_word[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i5.GSR = "DISABLED";
    FD1P3IX o_idl_word_i4 (.D(int_word[4]), .SP(dac_clk_p_c_enable_346), 
            .CD(n12778), .CK(dac_clk_p_c), .Q(idl_word[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i4.GSR = "DISABLED";
    FD1P3IX o_idl_stb_28 (.D(n26785), .SP(dac_clk_p_c_enable_195), .CD(w_reset), 
            .CK(dac_clk_p_c), .Q(idl_stb)) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(80[9] 88[22])
    defparam o_idl_stb_28.GSR = "DISABLED";
    FD1P3JX o_idl_word_i33 (.D(int_word[33]), .SP(dac_clk_p_c_enable_346), 
            .PD(n12778), .CK(dac_clk_p_c), .Q(idl_word[33])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i33.GSR = "DISABLED";
    FD1P3JX o_idl_word_i32 (.D(int_word[32]), .SP(dac_clk_p_c_enable_346), 
            .PD(n12778), .CK(dac_clk_p_c), .Q(idl_word[32])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i32.GSR = "DISABLED";
    FD1P3IX o_idl_word_i31 (.D(int_word[31]), .SP(dac_clk_p_c_enable_346), 
            .CD(n12778), .CK(dac_clk_p_c), .Q(idl_word[31])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i31.GSR = "DISABLED";
    FD1P3JX o_idl_word_i30 (.D(int_word[30]), .SP(dac_clk_p_c_enable_346), 
            .PD(n12778), .CK(dac_clk_p_c), .Q(idl_word[30])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i30.GSR = "DISABLED";
    FD1P3JX o_idl_word_i29 (.D(int_word[29]), .SP(dac_clk_p_c_enable_346), 
            .PD(n12778), .CK(dac_clk_p_c), .Q(idl_word[29])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i29.GSR = "DISABLED";
    FD1P3IX o_idl_word_i28 (.D(int_word[28]), .SP(dac_clk_p_c_enable_346), 
            .CD(n12778), .CK(dac_clk_p_c), .Q(idl_word[28])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i28.GSR = "DISABLED";
    FD1P3IX o_idl_word_i27 (.D(int_word[27]), .SP(dac_clk_p_c_enable_346), 
            .CD(n12778), .CK(dac_clk_p_c), .Q(idl_word[27])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i27.GSR = "DISABLED";
    FD1P3IX o_idl_word_i26 (.D(int_word[26]), .SP(dac_clk_p_c_enable_346), 
            .CD(n12778), .CK(dac_clk_p_c), .Q(idl_word[26])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i26.GSR = "DISABLED";
    FD1P3IX o_idl_word_i25 (.D(int_word[25]), .SP(dac_clk_p_c_enable_346), 
            .CD(n12778), .CK(dac_clk_p_c), .Q(idl_word[25])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i25.GSR = "DISABLED";
    FD1P3IX o_idl_word_i3 (.D(int_word[3]), .SP(dac_clk_p_c_enable_346), 
            .CD(n12778), .CK(dac_clk_p_c), .Q(idl_word[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i3.GSR = "DISABLED";
    FD1P3IX o_idl_word_i2 (.D(int_word[2]), .SP(dac_clk_p_c_enable_346), 
            .CD(n12778), .CK(dac_clk_p_c), .Q(idl_word[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i2.GSR = "DISABLED";
    FD1P3IX o_idl_word_i1 (.D(int_word[1]), .SP(dac_clk_p_c_enable_346), 
            .CD(n12778), .CK(dac_clk_p_c), .Q(idl_word[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i1.GSR = "DISABLED";
    FD1P3IX o_idl_word_i0 (.D(int_word[0]), .SP(dac_clk_p_c_enable_346), 
            .CD(n12778), .CK(dac_clk_p_c), .Q(idl_word[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i0.GSR = "DISABLED";
    FD1P3IX o_idl_word_i14 (.D(int_word[14]), .SP(dac_clk_p_c_enable_346), 
            .CD(n12778), .CK(dac_clk_p_c), .Q(idl_word[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i14.GSR = "DISABLED";
    FD1P3IX o_idl_word_i24 (.D(int_word[24]), .SP(dac_clk_p_c_enable_346), 
            .CD(n12778), .CK(dac_clk_p_c), .Q(idl_word[24])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i24.GSR = "DISABLED";
    FD1P3IX o_idl_word_i23 (.D(int_word[23]), .SP(dac_clk_p_c_enable_346), 
            .CD(n12778), .CK(dac_clk_p_c), .Q(idl_word[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i23.GSR = "DISABLED";
    FD1P3IX o_idl_word_i22 (.D(int_word[22]), .SP(dac_clk_p_c_enable_346), 
            .CD(n12778), .CK(dac_clk_p_c), .Q(idl_word[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i22.GSR = "DISABLED";
    FD1P3IX o_idl_word_i21 (.D(int_word[21]), .SP(dac_clk_p_c_enable_346), 
            .CD(n12778), .CK(dac_clk_p_c), .Q(idl_word[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i21.GSR = "DISABLED";
    FD1P3IX o_idl_word_i20 (.D(int_word[20]), .SP(dac_clk_p_c_enable_346), 
            .CD(n12778), .CK(dac_clk_p_c), .Q(idl_word[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i20.GSR = "DISABLED";
    FD1P3IX o_idl_word_i19 (.D(int_word[19]), .SP(dac_clk_p_c_enable_346), 
            .CD(n12778), .CK(dac_clk_p_c), .Q(idl_word[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i19.GSR = "DISABLED";
    FD1P3IX o_idl_word_i18 (.D(int_word[18]), .SP(dac_clk_p_c_enable_346), 
            .CD(n12778), .CK(dac_clk_p_c), .Q(idl_word[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i18.GSR = "DISABLED";
    FD1P3IX o_idl_word_i17 (.D(int_word[17]), .SP(dac_clk_p_c_enable_346), 
            .CD(n12778), .CK(dac_clk_p_c), .Q(idl_word[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i17.GSR = "DISABLED";
    FD1P3IX o_idl_word_i16 (.D(int_word[16]), .SP(dac_clk_p_c_enable_346), 
            .CD(n12778), .CK(dac_clk_p_c), .Q(idl_word[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i16.GSR = "DISABLED";
    FD1P3IX o_idl_word_i15 (.D(int_word[15]), .SP(dac_clk_p_c_enable_346), 
            .CD(n12778), .CK(dac_clk_p_c), .Q(idl_word[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i15.GSR = "DISABLED";
    FD1P3IX o_idl_word_i13 (.D(int_word[13]), .SP(dac_clk_p_c_enable_346), 
            .CD(n12778), .CK(dac_clk_p_c), .Q(idl_word[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i13.GSR = "DISABLED";
    FD1P3IX o_idl_word_i12 (.D(int_word[12]), .SP(dac_clk_p_c_enable_346), 
            .CD(n12778), .CK(dac_clk_p_c), .Q(idl_word[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i12.GSR = "DISABLED";
    FD1P3IX o_idl_word_i11 (.D(int_word[11]), .SP(dac_clk_p_c_enable_346), 
            .CD(n12778), .CK(dac_clk_p_c), .Q(idl_word[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=10, LSE_LCOL=9, LSE_RCOL=31, LSE_LLINE=121, LSE_RLINE=123 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(91[9] 95[29])
    defparam o_idl_word_i11.GSR = "DISABLED";
    LUT4 o_idl_stb_I_0_30_2_lut_rep_580 (.A(idl_stb), .B(hb_busy), .Z(n26903)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(97[22:43])
    defparam o_idl_stb_I_0_30_2_lut_rep_580.init = 16'h8888;
    LUT4 o_int_stb_I_0_66_2_lut_rep_462_3_lut (.A(idl_stb), .B(hb_busy), 
         .C(int_stb), .Z(n26785)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(97[22:43])
    defparam o_int_stb_I_0_66_2_lut_rep_462_3_lut.init = 16'h7070;
    LUT4 i1_3_lut_4_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(n29560), .D(int_stb), 
         .Z(dac_clk_p_c_enable_195)) /* synthesis lut_function=(A ((C)+!B)+!A ((C+(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(97[22:43])
    defparam i1_3_lut_4_lut_4_lut.init = 16'hf7f3;
    LUT4 i1_2_lut_3_lut_3_lut (.A(idl_stb), .B(hb_busy), .C(int_stb), 
         .Z(dac_clk_p_c_enable_346)) /* synthesis lut_function=(!(A (B)+!A !((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(97[22:43])
    defparam i1_2_lut_3_lut_3_lut.init = 16'h7373;
    LUT4 i22657_2_lut (.A(hb_busy), .B(int_stb), .Z(n12778)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i22657_2_lut.init = 16'h1111;
    LUT4 i22628_2_lut_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(n26940), 
         .D(int_stb), .Z(n12748)) /* synthesis lut_function=(!(A (B (C+(D))+!B (C))+!A (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(97[22:43])
    defparam i22628_2_lut_3_lut_4_lut.init = 16'h070f;
    LUT4 i1_2_lut_3_lut_4_lut (.A(idl_stb), .B(hb_busy), .C(n26940), .D(int_stb), 
         .Z(dac_clk_p_c_enable_416)) /* synthesis lut_function=(((C+!(D))+!B)+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/hbidle.v(97[22:43])
    defparam i1_2_lut_3_lut_4_lut.init = 16'hf7ff;
    
endmodule
//
// Verilog Description of module fm_generator_wb_slave
//

module fm_generator_wb_slave (dac_clk_p_c, wb_odata, i_resetb_N_301, wb_fm_data, 
            wb_fm_ack, wb_fm_data_31__N_63, GND_net, \wb_addr[0] , \wb_addr[1] , 
            \power_counter[1] , \smpl_register[1] , n2161, n26946, n38, 
            n34, \wb_addr[8] , \wb_addr[12] , n26947, \wb_addr[15] , 
            \wb_addr[9] , i_resetb_c, n20739, n2, \smpl_register[5] , 
            n26694, n2_adj_1, \smpl_register[20] , n26704, n2_adj_2, 
            \smpl_register[18] , n26703, n2_adj_3, \smpl_register[17] , 
            n26702, n2_adj_4, \smpl_register[16] , n26701, n2_adj_5, 
            \smpl_register[29] , n26699, n2_adj_6, \smpl_register[10] , 
            n26696, n2_adj_7, \smpl_register[9] , n26695, n20755, 
            n21184, n20749, n20719, o_baseband_q_c_7, o_baseband_i_c_7, 
            o_baseband_i_c_15, o_baseband_i_c_14, o_baseband_i_c_13, o_baseband_i_c_12, 
            o_baseband_i_c_11, o_baseband_i_c_10, n3655, o_baseband_i_c_8, 
            n29501, o_baseband_q_c_15, o_baseband_q_c_14, o_baseband_q_c_13, 
            o_baseband_q_c_12, o_baseband_q_c_11, o_baseband_q_c_10, n3656, 
            o_baseband_q_c_8) /* synthesis syn_module_defined=1 */ ;
    input dac_clk_p_c;
    input [31:0]wb_odata;
    input i_resetb_N_301;
    output [31:0]wb_fm_data;
    output wb_fm_ack;
    input wb_fm_data_31__N_63;
    input GND_net;
    input \wb_addr[0] ;
    input \wb_addr[1] ;
    input \power_counter[1] ;
    input \smpl_register[1] ;
    output n2161;
    input n26946;
    input n38;
    input n34;
    input \wb_addr[8] ;
    input \wb_addr[12] ;
    input n26947;
    input \wb_addr[15] ;
    input \wb_addr[9] ;
    input i_resetb_c;
    input n20739;
    input n2;
    input \smpl_register[5] ;
    output n26694;
    input n2_adj_1;
    input \smpl_register[20] ;
    output n26704;
    input n2_adj_2;
    input \smpl_register[18] ;
    output n26703;
    input n2_adj_3;
    input \smpl_register[17] ;
    output n26702;
    input n2_adj_4;
    input \smpl_register[16] ;
    output n26701;
    input n2_adj_5;
    input \smpl_register[29] ;
    output n26699;
    input n2_adj_6;
    input \smpl_register[10] ;
    output n26696;
    input n2_adj_7;
    input \smpl_register[9] ;
    output n26695;
    input n20755;
    input n21184;
    input n20749;
    input n20719;
    output o_baseband_q_c_7;
    output o_baseband_i_c_7;
    output o_baseband_i_c_15;
    output o_baseband_i_c_14;
    output o_baseband_i_c_13;
    output o_baseband_i_c_12;
    output o_baseband_i_c_11;
    output o_baseband_i_c_10;
    output n3655;
    output o_baseband_i_c_8;
    input n29501;
    output o_baseband_q_c_15;
    output o_baseband_q_c_14;
    output o_baseband_q_c_13;
    output o_baseband_q_c_12;
    output o_baseband_q_c_11;
    output o_baseband_q_c_10;
    output n3656;
    output o_baseband_q_c_8;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(28[49:58])
    wire [15:0]modulation_output /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(62[39:56])
    wire o_baseband_q_c_7 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[49:59])
    wire o_baseband_i_c_7 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[37:47])
    wire o_baseband_i_c_15 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[37:47])
    wire o_baseband_i_c_14 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[37:47])
    wire o_baseband_i_c_13 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[37:47])
    wire o_baseband_i_c_12 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[37:47])
    wire o_baseband_i_c_11 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[37:47])
    wire o_baseband_i_c_10 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[37:47])
    wire n3655 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[37:47])
    wire o_baseband_i_c_8 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[37:47])
    wire o_baseband_q_c_15 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[49:59])
    wire o_baseband_q_c_14 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[49:59])
    wire o_baseband_q_c_13 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[49:59])
    wire o_baseband_q_c_12 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[49:59])
    wire o_baseband_q_c_11 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[49:59])
    wire o_baseband_q_c_10 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[49:59])
    wire n3656 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[49:59])
    wire o_baseband_q_c_8 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[49:59])
    wire [31:0]\addr_space[3] ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(25[12:22])
    
    wire dac_clk_p_c_enable_147;
    wire [31:0]\addr_space[0] ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(25[12:22])
    
    wire dac_clk_p_c_enable_115;
    wire [31:0]\addr_space[1] ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(25[12:22])
    
    wire dac_clk_p_c_enable_76;
    wire [31:0]\addr_space[2] ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(25[12:22])
    
    wire dac_clk_p_c_enable_108;
    wire [30:0]carrier_center_increment_offset_ls;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(52[31:65])
    wire [30:0]n1;
    wire [31:0]o_wb_data_31__N_1337;
    wire [30:0]carrier_center_increment_offset_rs;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(52[67:101])
    wire [30:0]carrier_center_increment_offset_rs_30__N_1560;
    wire [30:0]carrier_increment;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(53[31:48])
    wire [30:0]carrier_increment_30__N_1591;
    wire [16:0]sine_lookup_width_minus_modulation_deviation_amount;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(74[27:78])
    wire [31:0]sine_lookup_width_minus_modulation_deviation_amount_16__N_1622;
    wire [16:0]modulation_deviation_amount_minus_sine_lookup_width;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(74[80:131])
    
    wire n63, n94, n22451, n64, n95, n17599, n26904, n26718, 
        n58, n89, n59, n55, n117, n88, n80, n103, n60, n56, 
        n118, n81, n104;
    wire [17:0]modulation_deviation_amount_minus_sine_lookup_width_16__N_1639;
    
    wire n26917, n72, n13522, n36_adj_2992, n13523, n40_adj_2993, 
        n44, n71, n9, n11, n13, n15, n13524, n7, n20382, n13521, 
        n26764, n13530, n37_adj_3000, n33_adj_3001, n41_adj_3002, 
        n45_adj_3003, n72_adj_3004, n14, n6, n8, n10, n12, n13529, 
        n38_adj_3005, n42_adj_3006, n46_adj_3007, n73, n22136, n24635, 
        n24636, n22135, n22127, n22126, n22121, n22120, n85, n26741, 
        n26742, n22118, n22117, n26726, n21389, n21388, n21386, 
        n21385, n17622, n14428, n26727, n21383, n79, n26757, n26728, 
        n21382, n26758, n26756, n21380, n78, n101, n102, n43_adj_3008, 
        n82, n26914, n105, n21379, n47_adj_3009, n74, n21377, 
        n21376, n83, n106, n48_adj_3010, n75, n20781, n21374, 
        n20775, n20773, n21373, n21371, n26690, n26689, n26691, 
        n21370, n21368, n73_adj_3013, n22285, n135, n134, n21367, 
        n21365, n21364, n178, n26672, n26671, n26673, n26786, 
        n26663, n26662, n26664, n21362, n20945, n20947, n20949, 
        n20935, n21361, n21359, n21358, n22217, n22216, n22214, 
        n22213, n26658, n39_adj_3014, n26659, n22211, n22210, n22208, 
        n22207, n22205, n22204, n22202, n22201, n22199, n22198, 
        n22196, n22195, n22193, n22192, n9080, n9078, n22190, 
        n70, n22189, n178_adj_3015, n52_adj_3016, n25, n27, n29, 
        n17, n19, n21, n23, n22187, n95_adj_3017, n26801, n49_adj_3018, 
        n53_adj_3019, n57_adj_3020, n30, n18, n20, n22, n24, n26, 
        n28, n22186, n96, n26916, n50_adj_3021, n54_adj_3022, n17621, 
        n97, n113, n16, n51_adj_3023, n98, n114, n17620, n99, 
        n115, n76, n45_adj_3024, n84, n26915, n22184, n100, n26725, 
        n77, n46_adj_3025, n22183, n22181, n22180, n17619, n132, 
        n133, n22172, n136, n137, n107, n123, n108, n22171, 
        n22163, n22162, n17618, n22154, n22153, n20665, n20679, 
        n20677, n20663, n20667, n22145, n22144, n17617, n17616, 
        n17615, n26660, n24637, n17614, n26657, n26939, n17613, 
        n17612, n17611, n17610, n17673, n17609, n17608, n17672, 
        n17671, n17670, n20879, n20881, n20883, n20869, n17606, 
        n17669, n17668, n17605, n17604, n17603, n17602, n17601, 
        n17600;
    wire [15:0]quarter_wave_sample_register_q;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(22[56:86])
    
    FD1P3AX \addr_space_3[[26__269  (.D(wb_odata[26]), .SP(dac_clk_p_c_enable_147), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[26__269 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[25__271  (.D(wb_odata[25]), .SP(dac_clk_p_c_enable_147), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[25__271 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[24__273  (.D(wb_odata[24]), .SP(dac_clk_p_c_enable_147), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[24__273 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[23__275  (.D(wb_odata[23]), .SP(dac_clk_p_c_enable_147), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[23__275 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[22__277  (.D(wb_odata[22]), .SP(dac_clk_p_c_enable_147), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[22__277 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[21__279  (.D(wb_odata[21]), .SP(dac_clk_p_c_enable_147), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[21__279 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[20__281  (.D(wb_odata[20]), .SP(dac_clk_p_c_enable_147), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[20__281 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[19__283  (.D(wb_odata[19]), .SP(dac_clk_p_c_enable_147), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[19__283 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[18__285  (.D(wb_odata[18]), .SP(dac_clk_p_c_enable_147), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[18__285 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[17__287  (.D(wb_odata[17]), .SP(dac_clk_p_c_enable_147), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[17__287 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[30__162  (.D(wb_odata[30]), .SP(dac_clk_p_c_enable_115), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[0] [30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[30__162 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[29__163  (.D(wb_odata[29]), .SP(dac_clk_p_c_enable_115), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[0] [29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[29__163 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[28__164  (.D(wb_odata[28]), .SP(dac_clk_p_c_enable_115), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[0] [28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[28__164 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[27__165  (.D(wb_odata[27]), .SP(dac_clk_p_c_enable_115), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[0] [27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[27__165 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[26__166  (.D(wb_odata[26]), .SP(dac_clk_p_c_enable_115), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[0] [26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[26__166 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[25__167  (.D(wb_odata[25]), .SP(dac_clk_p_c_enable_115), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[0] [25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[25__167 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[24__168  (.D(wb_odata[24]), .SP(dac_clk_p_c_enable_115), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[0] [24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[24__168 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[23__169  (.D(wb_odata[23]), .SP(dac_clk_p_c_enable_115), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[0] [23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[23__169 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[21__172  (.D(wb_odata[21]), .SP(dac_clk_p_c_enable_115), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[0] [21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[21__172 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[20__173  (.D(wb_odata[20]), .SP(dac_clk_p_c_enable_115), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[0] [20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[20__173 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[19__174  (.D(wb_odata[19]), .SP(dac_clk_p_c_enable_115), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[0] [19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[19__174 .GSR = "DISABLED";
    FD1P3BX \addr_space_0[[18__175  (.D(wb_odata[18]), .SP(dac_clk_p_c_enable_115), 
            .CK(dac_clk_p_c), .PD(i_resetb_N_301), .Q(\addr_space[0] [18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[18__175 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[17__176  (.D(wb_odata[17]), .SP(dac_clk_p_c_enable_115), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[0] [17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[17__176 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[16__177  (.D(wb_odata[16]), .SP(dac_clk_p_c_enable_115), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[0] [16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[16__177 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[15__178  (.D(wb_odata[15]), .SP(dac_clk_p_c_enable_115), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[0] [15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[15__178 .GSR = "DISABLED";
    FD1P3BX \addr_space_0[[14__179  (.D(wb_odata[14]), .SP(dac_clk_p_c_enable_115), 
            .CK(dac_clk_p_c), .PD(i_resetb_N_301), .Q(\addr_space[0] [14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[14__179 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[13__180  (.D(wb_odata[13]), .SP(dac_clk_p_c_enable_115), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[0] [13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[13__180 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[12__181  (.D(wb_odata[12]), .SP(dac_clk_p_c_enable_115), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[0] [12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[12__181 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[11__182  (.D(wb_odata[11]), .SP(dac_clk_p_c_enable_115), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[0] [11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[11__182 .GSR = "DISABLED";
    FD1P3BX \addr_space_0[[10__183  (.D(wb_odata[10]), .SP(dac_clk_p_c_enable_115), 
            .CK(dac_clk_p_c), .PD(i_resetb_N_301), .Q(\addr_space[0] [10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[10__183 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[9__184  (.D(wb_odata[9]), .SP(dac_clk_p_c_enable_115), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[0] [9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[9__184 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[8__185  (.D(wb_odata[8]), .SP(dac_clk_p_c_enable_115), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[0] [8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[8__185 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[7__186  (.D(wb_odata[7]), .SP(dac_clk_p_c_enable_115), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[0] [7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[7__186 .GSR = "DISABLED";
    FD1P3BX \addr_space_0[[6__187  (.D(wb_odata[6]), .SP(dac_clk_p_c_enable_115), 
            .CK(dac_clk_p_c), .PD(i_resetb_N_301), .Q(\addr_space[0] [6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[6__187 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[5__188  (.D(wb_odata[5]), .SP(dac_clk_p_c_enable_115), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[0] [5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[5__188 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[4__189  (.D(wb_odata[4]), .SP(dac_clk_p_c_enable_115), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[0] [4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[4__189 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[3__190  (.D(wb_odata[3]), .SP(dac_clk_p_c_enable_115), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[0] [3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[3__190 .GSR = "DISABLED";
    FD1P3BX \addr_space_0[[2__191  (.D(wb_odata[2]), .SP(dac_clk_p_c_enable_115), 
            .CK(dac_clk_p_c), .PD(i_resetb_N_301), .Q(\addr_space[0] [2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[2__191 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[1__192  (.D(wb_odata[1]), .SP(dac_clk_p_c_enable_115), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[0] [1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[1__192 .GSR = "DISABLED";
    FD1P3DX \addr_space_0[[0__193  (.D(wb_odata[0]), .SP(dac_clk_p_c_enable_115), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[0] [0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[0__193 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[31__194  (.D(wb_odata[31]), .SP(dac_clk_p_c_enable_76), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[1] [31])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[31__194 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[30__195  (.D(wb_odata[30]), .SP(dac_clk_p_c_enable_76), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[1] [30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[30__195 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[29__196  (.D(wb_odata[29]), .SP(dac_clk_p_c_enable_76), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[1] [29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[29__196 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[28__197  (.D(wb_odata[28]), .SP(dac_clk_p_c_enable_76), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[1] [28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[28__197 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[27__198  (.D(wb_odata[27]), .SP(dac_clk_p_c_enable_76), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[1] [27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[27__198 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[26__199  (.D(wb_odata[26]), .SP(dac_clk_p_c_enable_76), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[1] [26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[26__199 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[25__200  (.D(wb_odata[25]), .SP(dac_clk_p_c_enable_76), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[1] [25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[25__200 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[24__201  (.D(wb_odata[24]), .SP(dac_clk_p_c_enable_76), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[1] [24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[24__201 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[23__202  (.D(wb_odata[23]), .SP(dac_clk_p_c_enable_76), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[1] [23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[23__202 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[22__203  (.D(wb_odata[22]), .SP(dac_clk_p_c_enable_76), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[1] [22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[22__203 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[21__204  (.D(wb_odata[21]), .SP(dac_clk_p_c_enable_76), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[1] [21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[21__204 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[20__205  (.D(wb_odata[20]), .SP(dac_clk_p_c_enable_76), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[1] [20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[20__205 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[19__206  (.D(wb_odata[19]), .SP(dac_clk_p_c_enable_76), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[1] [19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[19__206 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[18__207  (.D(wb_odata[18]), .SP(dac_clk_p_c_enable_76), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[1] [18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[18__207 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[17__208  (.D(wb_odata[17]), .SP(dac_clk_p_c_enable_76), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[1] [17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[17__208 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[16__209  (.D(wb_odata[16]), .SP(dac_clk_p_c_enable_76), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[1] [16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[16__209 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[15__210  (.D(wb_odata[15]), .SP(dac_clk_p_c_enable_76), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[1] [15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[15__210 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[14__211  (.D(wb_odata[14]), .SP(dac_clk_p_c_enable_76), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[1] [14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[14__211 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[13__212  (.D(wb_odata[13]), .SP(dac_clk_p_c_enable_76), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[1] [13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[13__212 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[12__213  (.D(wb_odata[12]), .SP(dac_clk_p_c_enable_76), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[1] [12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[12__213 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[11__214  (.D(wb_odata[11]), .SP(dac_clk_p_c_enable_76), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[1] [11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[11__214 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[10__215  (.D(wb_odata[10]), .SP(dac_clk_p_c_enable_76), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[1] [10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[10__215 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[9__216  (.D(wb_odata[9]), .SP(dac_clk_p_c_enable_76), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[1] [9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[9__216 .GSR = "DISABLED";
    FD1P3BX \addr_space_1[[8__217  (.D(wb_odata[8]), .SP(dac_clk_p_c_enable_76), 
            .CK(dac_clk_p_c), .PD(i_resetb_N_301), .Q(\addr_space[1] [8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[8__217 .GSR = "DISABLED";
    FD1P3BX \addr_space_1[[7__218  (.D(wb_odata[7]), .SP(dac_clk_p_c_enable_76), 
            .CK(dac_clk_p_c), .PD(i_resetb_N_301), .Q(\addr_space[1] [7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[7__218 .GSR = "DISABLED";
    FD1P3DX \addr_space_1[[6__219  (.D(wb_odata[6]), .SP(dac_clk_p_c_enable_76), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[1] [6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[6__219 .GSR = "DISABLED";
    FD1P3BX \addr_space_1[[5__220  (.D(wb_odata[5]), .SP(dac_clk_p_c_enable_76), 
            .CK(dac_clk_p_c), .PD(i_resetb_N_301), .Q(\addr_space[1] [5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[5__220 .GSR = "DISABLED";
    FD1P3BX \addr_space_1[[4__221  (.D(wb_odata[4]), .SP(dac_clk_p_c_enable_76), 
            .CK(dac_clk_p_c), .PD(i_resetb_N_301), .Q(\addr_space[1] [4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[4__221 .GSR = "DISABLED";
    FD1P3BX \addr_space_1[[3__222  (.D(wb_odata[3]), .SP(dac_clk_p_c_enable_76), 
            .CK(dac_clk_p_c), .PD(i_resetb_N_301), .Q(\addr_space[1] [3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[3__222 .GSR = "DISABLED";
    FD1P3BX \addr_space_1[[2__223  (.D(wb_odata[2]), .SP(dac_clk_p_c_enable_76), 
            .CK(dac_clk_p_c), .PD(i_resetb_N_301), .Q(\addr_space[1] [2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[2__223 .GSR = "DISABLED";
    FD1P3BX \addr_space_1[[1__224  (.D(wb_odata[1]), .SP(dac_clk_p_c_enable_76), 
            .CK(dac_clk_p_c), .PD(i_resetb_N_301), .Q(\addr_space[1] [1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[1__224 .GSR = "DISABLED";
    FD1P3BX \addr_space_1[[0__225  (.D(wb_odata[0]), .SP(dac_clk_p_c_enable_76), 
            .CK(dac_clk_p_c), .PD(i_resetb_N_301), .Q(\addr_space[1] [0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_1[[0__225 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[31__226  (.D(wb_odata[31]), .SP(dac_clk_p_c_enable_108), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [31])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[31__226 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[30__227  (.D(wb_odata[30]), .SP(dac_clk_p_c_enable_108), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[30__227 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[29__228  (.D(wb_odata[29]), .SP(dac_clk_p_c_enable_108), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[29__228 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[28__229  (.D(wb_odata[28]), .SP(dac_clk_p_c_enable_108), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[28__229 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[27__230  (.D(wb_odata[27]), .SP(dac_clk_p_c_enable_108), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[27__230 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[26__231  (.D(wb_odata[26]), .SP(dac_clk_p_c_enable_108), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[26__231 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[25__232  (.D(wb_odata[25]), .SP(dac_clk_p_c_enable_108), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[25__232 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[24__233  (.D(wb_odata[24]), .SP(dac_clk_p_c_enable_108), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[24__233 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[23__234  (.D(wb_odata[23]), .SP(dac_clk_p_c_enable_108), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[23__234 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[22__235  (.D(wb_odata[22]), .SP(dac_clk_p_c_enable_108), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[22__235 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[21__236  (.D(wb_odata[21]), .SP(dac_clk_p_c_enable_108), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[21__236 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[20__237  (.D(wb_odata[20]), .SP(dac_clk_p_c_enable_108), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[20__237 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[19__238  (.D(wb_odata[19]), .SP(dac_clk_p_c_enable_108), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[19__238 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[18__239  (.D(wb_odata[18]), .SP(dac_clk_p_c_enable_108), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[18__239 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[17__240  (.D(wb_odata[17]), .SP(dac_clk_p_c_enable_108), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[17__240 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[16__241  (.D(wb_odata[16]), .SP(dac_clk_p_c_enable_108), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[16__241 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[15__242  (.D(wb_odata[15]), .SP(dac_clk_p_c_enable_108), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[15__242 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[14__243  (.D(wb_odata[14]), .SP(dac_clk_p_c_enable_108), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[14__243 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[13__244  (.D(wb_odata[13]), .SP(dac_clk_p_c_enable_108), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[13__244 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[12__245  (.D(wb_odata[12]), .SP(dac_clk_p_c_enable_108), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[12__245 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[11__246  (.D(wb_odata[11]), .SP(dac_clk_p_c_enable_108), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[11__246 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[10__247  (.D(wb_odata[10]), .SP(dac_clk_p_c_enable_108), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[10__247 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[9__248  (.D(wb_odata[9]), .SP(dac_clk_p_c_enable_108), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[9__248 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[8__249  (.D(wb_odata[8]), .SP(dac_clk_p_c_enable_108), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[8__249 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[7__250  (.D(wb_odata[7]), .SP(dac_clk_p_c_enable_108), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[7__250 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[6__251  (.D(wb_odata[6]), .SP(dac_clk_p_c_enable_108), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[6__251 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[5__252  (.D(wb_odata[5]), .SP(dac_clk_p_c_enable_108), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[5__252 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[4__253  (.D(wb_odata[4]), .SP(dac_clk_p_c_enable_108), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[4__253 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[3__254  (.D(wb_odata[3]), .SP(dac_clk_p_c_enable_108), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[3__254 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[2__255  (.D(wb_odata[2]), .SP(dac_clk_p_c_enable_108), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[2__255 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[1__256  (.D(wb_odata[1]), .SP(dac_clk_p_c_enable_108), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[1__256 .GSR = "DISABLED";
    FD1P3DX \addr_space_2[[0__257  (.D(wb_odata[0]), .SP(dac_clk_p_c_enable_108), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[2] [0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_2[[0__257 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[16__289  (.D(wb_odata[16]), .SP(dac_clk_p_c_enable_147), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[16__289 .GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i0 (.D(n1[0]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_ls[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_ls__i0.GSR = "DISABLED";
    FD1S3AX o_wb_data_i0 (.D(o_wb_data_31__N_1337[0]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i0.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_rs_i1 (.D(carrier_center_increment_offset_rs_30__N_1560[0]), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_rs[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_rs_i1.GSR = "DISABLED";
    FD1S3DX carrier_increment_i0 (.D(carrier_increment_30__N_1591[0]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(carrier_increment[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_increment_i0.GSR = "DISABLED";
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i0 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[0]), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(sine_lookup_width_minus_modulation_deviation_amount[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i0.GSR = "DISABLED";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i0 (.D(\addr_space[2] [0]), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(modulation_deviation_amount_minus_sine_lookup_width[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i0.GSR = "DISABLED";
    FD1P3DX \addr_space_0[[31__161  (.D(wb_odata[31]), .SP(dac_clk_p_c_enable_115), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(\addr_space[0] [31])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[31__161 .GSR = "DISABLED";
    FD1P3BX \addr_space_0[[22__171  (.D(wb_odata[22]), .SP(dac_clk_p_c_enable_115), 
            .CK(dac_clk_p_c), .PD(i_resetb_N_301), .Q(\addr_space[0] [22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_0[[22__171 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[15__291  (.D(wb_odata[15]), .SP(dac_clk_p_c_enable_147), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[15__291 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[14__293  (.D(wb_odata[14]), .SP(dac_clk_p_c_enable_147), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[14__293 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[13__295  (.D(wb_odata[13]), .SP(dac_clk_p_c_enable_147), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[13__295 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[12__297  (.D(wb_odata[12]), .SP(dac_clk_p_c_enable_147), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[12__297 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[11__299  (.D(wb_odata[11]), .SP(dac_clk_p_c_enable_147), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[11__299 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[10__301  (.D(wb_odata[10]), .SP(dac_clk_p_c_enable_147), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[10__301 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[9__303  (.D(wb_odata[9]), .SP(dac_clk_p_c_enable_147), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[9__303 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[8__305  (.D(wb_odata[8]), .SP(dac_clk_p_c_enable_147), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[8__305 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[7__307  (.D(wb_odata[7]), .SP(dac_clk_p_c_enable_147), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[7__307 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[6__309  (.D(wb_odata[6]), .SP(dac_clk_p_c_enable_147), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[6__309 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[5__311  (.D(wb_odata[5]), .SP(dac_clk_p_c_enable_147), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[5__311 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[4__313  (.D(wb_odata[4]), .SP(dac_clk_p_c_enable_147), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[4__313 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[3__315  (.D(wb_odata[3]), .SP(dac_clk_p_c_enable_147), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[3__315 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[2__317  (.D(wb_odata[2]), .SP(dac_clk_p_c_enable_147), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[2__317 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[1__319  (.D(wb_odata[1]), .SP(dac_clk_p_c_enable_147), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[1__319 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[0__321  (.D(wb_odata[0]), .SP(dac_clk_p_c_enable_147), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[0__321 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[31__259  (.D(wb_odata[31]), .SP(dac_clk_p_c_enable_147), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [31])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[31__259 .GSR = "DISABLED";
    FD1S3IX o_wb_ack_323 (.D(wb_fm_data_31__N_63), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(wb_fm_ack)) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(43[8] 48[4])
    defparam o_wb_ack_323.GSR = "DISABLED";
    FD1P3AX \addr_space_3[[30__261  (.D(wb_odata[30]), .SP(dac_clk_p_c_enable_147), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[30__261 .GSR = "DISABLED";
    PFUMX i6614 (.BLUT(n63), .ALUT(n94), .C0(n22451), .Z(carrier_center_increment_offset_rs_30__N_1560[0]));
    PFUMX i6616 (.BLUT(n64), .ALUT(n95), .C0(n22451), .Z(carrier_center_increment_offset_rs_30__N_1560[1]));
    FD1P3AX \addr_space_3[[29__263  (.D(wb_odata[29]), .SP(dac_clk_p_c_enable_147), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[29__263 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[28__265  (.D(wb_odata[28]), .SP(dac_clk_p_c_enable_147), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[28__265 .GSR = "DISABLED";
    FD1P3AX \addr_space_3[[27__267  (.D(wb_odata[27]), .SP(dac_clk_p_c_enable_147), 
            .CK(dac_clk_p_c), .Q(\addr_space[3] [27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(32[11] 36[5])
    defparam \addr_space_3[[27__267 .GSR = "DISABLED";
    CCU2D sub_396_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\addr_space[2] [0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n17599));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(85[58:109])
    defparam sub_396_add_2_1.INIT0 = 16'h0000;
    defparam sub_396_add_2_1.INIT1 = 16'h0aaa;
    defparam sub_396_add_2_1.INJECT1_0 = "NO";
    defparam sub_396_add_2_1.INJECT1_1 = "NO";
    LUT4 mux_393_Mux_1_i3_4_lut_4_lut_4_lut (.A(\wb_addr[0] ), .B(\wb_addr[1] ), 
         .C(\power_counter[1] ), .D(\smpl_register[1] ), .Z(n2161)) /* synthesis lut_function=(A (B (C)+!B (D))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(34[4:25])
    defparam mux_393_Mux_1_i3_4_lut_4_lut_4_lut.init = 16'hb391;
    LUT4 i1_2_lut_rep_395_3_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .B(n26904), .C(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .D(modulation_deviation_amount_minus_sine_lookup_width[2]), .Z(n26718)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i1_2_lut_rep_395_3_lut_4_lut.init = 16'h0004;
    LUT4 i10879_3_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .B(n26904), .C(modulation_deviation_amount_minus_sine_lookup_width[2]), 
         .D(n58), .Z(n89)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i10879_3_lut_4_lut.init = 16'h4f40;
    LUT4 i11032_2_lut_4_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[2]), .C(n59), 
         .D(n55), .Z(n117)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i11032_2_lut_4_lut_4_lut.init = 16'h5140;
    LUT4 modulation_output_15__I_0_332_i103_4_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[4]), .C(n88), 
         .D(n80), .Z(n103)) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C)+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam modulation_output_15__I_0_332_i103_4_lut_4_lut.init = 16'h7340;
    LUT4 i11033_2_lut_4_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[2]), .C(n60), 
         .D(n56), .Z(n118)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i11033_2_lut_4_lut_4_lut.init = 16'h5140;
    LUT4 modulation_output_15__I_0_332_i104_4_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[4]), .C(n89), 
         .D(n81), .Z(n104)) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C)+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam modulation_output_15__I_0_332_i104_4_lut_4_lut.init = 16'h7340;
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i16 (.D(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[16]), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(modulation_deviation_amount_minus_sine_lookup_width[16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i16.GSR = "DISABLED";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i15 (.D(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[15]), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(modulation_deviation_amount_minus_sine_lookup_width[15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i15.GSR = "DISABLED";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i14 (.D(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[14]), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(modulation_deviation_amount_minus_sine_lookup_width[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i14.GSR = "DISABLED";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i13 (.D(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[13]), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(modulation_deviation_amount_minus_sine_lookup_width[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i13.GSR = "DISABLED";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i12 (.D(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[12]), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(modulation_deviation_amount_minus_sine_lookup_width[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i12.GSR = "DISABLED";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i11 (.D(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[11]), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(modulation_deviation_amount_minus_sine_lookup_width[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i11.GSR = "DISABLED";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i10 (.D(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[10]), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(modulation_deviation_amount_minus_sine_lookup_width[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i10.GSR = "DISABLED";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i9 (.D(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[9]), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(modulation_deviation_amount_minus_sine_lookup_width[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i9.GSR = "DISABLED";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i8 (.D(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[8]), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(modulation_deviation_amount_minus_sine_lookup_width[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i8.GSR = "DISABLED";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i7 (.D(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[7]), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(modulation_deviation_amount_minus_sine_lookup_width[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i7.GSR = "DISABLED";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i6 (.D(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[6]), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(modulation_deviation_amount_minus_sine_lookup_width[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i6.GSR = "DISABLED";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i5 (.D(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[5]), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(modulation_deviation_amount_minus_sine_lookup_width[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i5.GSR = "DISABLED";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i4 (.D(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[4]), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(modulation_deviation_amount_minus_sine_lookup_width[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i4.GSR = "DISABLED";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i3 (.D(\addr_space[2] [3]), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(modulation_deviation_amount_minus_sine_lookup_width[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i3.GSR = "DISABLED";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i2 (.D(\addr_space[2] [2]), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(modulation_deviation_amount_minus_sine_lookup_width[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i2.GSR = "DISABLED";
    FD1S3DX modulation_deviation_amount_minus_sine_lookup_width_i1 (.D(\addr_space[2] [1]), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(modulation_deviation_amount_minus_sine_lookup_width[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam modulation_deviation_amount_minus_sine_lookup_width_i1.GSR = "DISABLED";
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i16 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[16]), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(sine_lookup_width_minus_modulation_deviation_amount[16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i16.GSR = "DISABLED";
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i15 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[15]), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(sine_lookup_width_minus_modulation_deviation_amount[15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i15.GSR = "DISABLED";
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i14 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[14]), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(sine_lookup_width_minus_modulation_deviation_amount[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i14.GSR = "DISABLED";
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i13 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[13]), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(sine_lookup_width_minus_modulation_deviation_amount[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i13.GSR = "DISABLED";
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i12 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[12]), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(sine_lookup_width_minus_modulation_deviation_amount[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i12.GSR = "DISABLED";
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i11 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[11]), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(sine_lookup_width_minus_modulation_deviation_amount[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i11.GSR = "DISABLED";
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i10 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[10]), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(sine_lookup_width_minus_modulation_deviation_amount[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i10.GSR = "DISABLED";
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i9 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[9]), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(sine_lookup_width_minus_modulation_deviation_amount[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i9.GSR = "DISABLED";
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i8 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[8]), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(sine_lookup_width_minus_modulation_deviation_amount[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i8.GSR = "DISABLED";
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i7 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[7]), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(sine_lookup_width_minus_modulation_deviation_amount[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i7.GSR = "DISABLED";
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i6 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[6]), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(sine_lookup_width_minus_modulation_deviation_amount[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i6.GSR = "DISABLED";
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i5 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[5]), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(sine_lookup_width_minus_modulation_deviation_amount[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i5.GSR = "DISABLED";
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i4 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[4]), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(sine_lookup_width_minus_modulation_deviation_amount[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i4.GSR = "DISABLED";
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i3 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[3]), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(sine_lookup_width_minus_modulation_deviation_amount[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i3.GSR = "DISABLED";
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i2 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[2]), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(sine_lookup_width_minus_modulation_deviation_amount[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i2.GSR = "DISABLED";
    FD1S3DX sine_lookup_width_minus_modulation_deviation_amount_i1 (.D(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[1]), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(sine_lookup_width_minus_modulation_deviation_amount[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam sine_lookup_width_minus_modulation_deviation_amount_i1.GSR = "DISABLED";
    FD1S3DX carrier_increment_i30 (.D(carrier_increment_30__N_1591[30]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(carrier_increment[30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_increment_i30.GSR = "DISABLED";
    FD1S3DX carrier_increment_i29 (.D(carrier_increment_30__N_1591[29]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(carrier_increment[29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_increment_i29.GSR = "DISABLED";
    FD1S3DX carrier_increment_i28 (.D(carrier_increment_30__N_1591[28]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(carrier_increment[28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_increment_i28.GSR = "DISABLED";
    FD1S3DX carrier_increment_i27 (.D(carrier_increment_30__N_1591[27]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(carrier_increment[27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_increment_i27.GSR = "DISABLED";
    FD1S3DX carrier_increment_i26 (.D(carrier_increment_30__N_1591[26]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(carrier_increment[26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_increment_i26.GSR = "DISABLED";
    FD1S3DX carrier_increment_i25 (.D(carrier_increment_30__N_1591[25]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(carrier_increment[25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_increment_i25.GSR = "DISABLED";
    LUT4 i6541_3_lut_4_lut (.A(n26917), .B(modulation_deviation_amount_minus_sine_lookup_width[2]), 
         .C(modulation_output[14]), .D(modulation_output[15]), .Z(n72)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam i6541_3_lut_4_lut.init = 16'hf780;
    FD1S3DX carrier_increment_i24 (.D(carrier_increment_30__N_1591[24]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(carrier_increment[24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_increment_i24.GSR = "DISABLED";
    FD1S3DX carrier_increment_i23 (.D(carrier_increment_30__N_1591[23]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(carrier_increment[23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_increment_i23.GSR = "DISABLED";
    FD1S3DX carrier_increment_i22 (.D(carrier_increment_30__N_1591[22]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(carrier_increment[22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_increment_i22.GSR = "DISABLED";
    FD1S3DX carrier_increment_i21 (.D(carrier_increment_30__N_1591[21]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(carrier_increment[21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_increment_i21.GSR = "DISABLED";
    FD1S3DX carrier_increment_i20 (.D(carrier_increment_30__N_1591[20]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(carrier_increment[20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_increment_i20.GSR = "DISABLED";
    FD1S3DX carrier_increment_i19 (.D(carrier_increment_30__N_1591[19]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(carrier_increment[19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_increment_i19.GSR = "DISABLED";
    FD1S3DX carrier_increment_i18 (.D(carrier_increment_30__N_1591[18]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(carrier_increment[18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_increment_i18.GSR = "DISABLED";
    FD1S3DX carrier_increment_i17 (.D(carrier_increment_30__N_1591[17]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(carrier_increment[17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_increment_i17.GSR = "DISABLED";
    FD1S3DX carrier_increment_i16 (.D(carrier_increment_30__N_1591[16]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(carrier_increment[16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_increment_i16.GSR = "DISABLED";
    FD1S3DX carrier_increment_i15 (.D(carrier_increment_30__N_1591[15]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(carrier_increment[15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_increment_i15.GSR = "DISABLED";
    FD1S3DX carrier_increment_i14 (.D(carrier_increment_30__N_1591[14]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(carrier_increment[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_increment_i14.GSR = "DISABLED";
    FD1S3DX carrier_increment_i13 (.D(carrier_increment_30__N_1591[13]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(carrier_increment[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_increment_i13.GSR = "DISABLED";
    FD1S3DX carrier_increment_i12 (.D(carrier_increment_30__N_1591[12]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(carrier_increment[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_increment_i12.GSR = "DISABLED";
    FD1S3DX carrier_increment_i11 (.D(carrier_increment_30__N_1591[11]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(carrier_increment[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_increment_i11.GSR = "DISABLED";
    FD1S3DX carrier_increment_i10 (.D(carrier_increment_30__N_1591[10]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(carrier_increment[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_increment_i10.GSR = "DISABLED";
    FD1S3DX carrier_increment_i9 (.D(carrier_increment_30__N_1591[9]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(carrier_increment[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_increment_i9.GSR = "DISABLED";
    FD1S3DX carrier_increment_i8 (.D(carrier_increment_30__N_1591[8]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(carrier_increment[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_increment_i8.GSR = "DISABLED";
    FD1S3DX carrier_increment_i7 (.D(carrier_increment_30__N_1591[7]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(carrier_increment[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_increment_i7.GSR = "DISABLED";
    FD1S3DX carrier_increment_i6 (.D(carrier_increment_30__N_1591[6]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(carrier_increment[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_increment_i6.GSR = "DISABLED";
    FD1S3DX carrier_increment_i5 (.D(carrier_increment_30__N_1591[5]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(carrier_increment[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_increment_i5.GSR = "DISABLED";
    FD1S3DX carrier_increment_i4 (.D(carrier_increment_30__N_1591[4]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(carrier_increment[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_increment_i4.GSR = "DISABLED";
    FD1S3DX carrier_increment_i3 (.D(carrier_increment_30__N_1591[3]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(carrier_increment[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_increment_i3.GSR = "DISABLED";
    FD1S3DX carrier_increment_i2 (.D(carrier_increment_30__N_1591[2]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(carrier_increment[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_increment_i2.GSR = "DISABLED";
    FD1S3DX carrier_increment_i1 (.D(carrier_increment_30__N_1591[1]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(carrier_increment[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_increment_i1.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_rs_i16 (.D(modulation_output[15]), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_rs[30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_rs_i16.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_rs_i15 (.D(carrier_center_increment_offset_rs_30__N_1560[14]), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_rs[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_rs_i15.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_rs_i14 (.D(carrier_center_increment_offset_rs_30__N_1560[13]), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_rs[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_rs_i14.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_rs_i13 (.D(carrier_center_increment_offset_rs_30__N_1560[12]), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_rs[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_rs_i13.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_rs_i12 (.D(carrier_center_increment_offset_rs_30__N_1560[11]), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_rs[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_rs_i12.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_rs_i11 (.D(carrier_center_increment_offset_rs_30__N_1560[10]), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_rs[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_rs_i11.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_rs_i10 (.D(carrier_center_increment_offset_rs_30__N_1560[9]), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_rs[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_rs_i10.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_rs_i9 (.D(carrier_center_increment_offset_rs_30__N_1560[8]), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_rs[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_rs_i9.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_rs_i8 (.D(carrier_center_increment_offset_rs_30__N_1560[7]), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_rs[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_rs_i8.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_rs_i7 (.D(carrier_center_increment_offset_rs_30__N_1560[6]), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_rs[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_rs_i7.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_rs_i6 (.D(carrier_center_increment_offset_rs_30__N_1560[5]), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_rs[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_rs_i6.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_rs_i5 (.D(carrier_center_increment_offset_rs_30__N_1560[4]), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_rs[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_rs_i5.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_rs_i4 (.D(carrier_center_increment_offset_rs_30__N_1560[3]), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_rs[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_rs_i4.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_rs_i3 (.D(carrier_center_increment_offset_rs_30__N_1560[2]), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_rs[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_rs_i3.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_rs_i2 (.D(carrier_center_increment_offset_rs_30__N_1560[1]), 
            .CK(dac_clk_p_c), .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_rs[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_rs_i2.GSR = "DISABLED";
    FD1S3AX o_wb_data_i31 (.D(o_wb_data_31__N_1337[31]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[31])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i31.GSR = "DISABLED";
    FD1S3AX o_wb_data_i30 (.D(o_wb_data_31__N_1337[30]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i30.GSR = "DISABLED";
    FD1S3AX o_wb_data_i29 (.D(o_wb_data_31__N_1337[29]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i29.GSR = "DISABLED";
    FD1S3AX o_wb_data_i28 (.D(o_wb_data_31__N_1337[28]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i28.GSR = "DISABLED";
    FD1S3AX o_wb_data_i27 (.D(o_wb_data_31__N_1337[27]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i27.GSR = "DISABLED";
    FD1S3AX o_wb_data_i26 (.D(o_wb_data_31__N_1337[26]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i26.GSR = "DISABLED";
    FD1S3AX o_wb_data_i25 (.D(o_wb_data_31__N_1337[25]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i25.GSR = "DISABLED";
    FD1S3AX o_wb_data_i24 (.D(o_wb_data_31__N_1337[24]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i24.GSR = "DISABLED";
    FD1S3AX o_wb_data_i23 (.D(o_wb_data_31__N_1337[23]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i23.GSR = "DISABLED";
    FD1S3AX o_wb_data_i22 (.D(o_wb_data_31__N_1337[22]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i22.GSR = "DISABLED";
    FD1S3AX o_wb_data_i21 (.D(o_wb_data_31__N_1337[21]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i21.GSR = "DISABLED";
    FD1S3AX o_wb_data_i20 (.D(o_wb_data_31__N_1337[20]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i20.GSR = "DISABLED";
    FD1S3AX o_wb_data_i19 (.D(o_wb_data_31__N_1337[19]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i19.GSR = "DISABLED";
    FD1S3AX o_wb_data_i18 (.D(o_wb_data_31__N_1337[18]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i18.GSR = "DISABLED";
    FD1S3AX o_wb_data_i17 (.D(o_wb_data_31__N_1337[17]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i17.GSR = "DISABLED";
    FD1S3AX o_wb_data_i16 (.D(o_wb_data_31__N_1337[16]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i16.GSR = "DISABLED";
    FD1S3AX o_wb_data_i15 (.D(o_wb_data_31__N_1337[15]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i15.GSR = "DISABLED";
    FD1S3AX o_wb_data_i14 (.D(o_wb_data_31__N_1337[14]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i14.GSR = "DISABLED";
    FD1S3AX o_wb_data_i13 (.D(o_wb_data_31__N_1337[13]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i13.GSR = "DISABLED";
    FD1S3AX o_wb_data_i12 (.D(o_wb_data_31__N_1337[12]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i12.GSR = "DISABLED";
    FD1S3AX o_wb_data_i11 (.D(o_wb_data_31__N_1337[11]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i11.GSR = "DISABLED";
    FD1S3AX o_wb_data_i10 (.D(o_wb_data_31__N_1337[10]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i10.GSR = "DISABLED";
    FD1S3AX o_wb_data_i9 (.D(o_wb_data_31__N_1337[9]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i9.GSR = "DISABLED";
    FD1S3AX o_wb_data_i8 (.D(o_wb_data_31__N_1337[8]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i8.GSR = "DISABLED";
    FD1S3AX o_wb_data_i7 (.D(o_wb_data_31__N_1337[7]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i7.GSR = "DISABLED";
    FD1S3AX o_wb_data_i6 (.D(o_wb_data_31__N_1337[6]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i6.GSR = "DISABLED";
    FD1S3AX o_wb_data_i5 (.D(o_wb_data_31__N_1337[5]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i5.GSR = "DISABLED";
    FD1S3AX o_wb_data_i4 (.D(o_wb_data_31__N_1337[4]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i4.GSR = "DISABLED";
    FD1S3AX o_wb_data_i3 (.D(o_wb_data_31__N_1337[3]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i3.GSR = "DISABLED";
    FD1S3AX o_wb_data_i2 (.D(o_wb_data_31__N_1337[2]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i2.GSR = "DISABLED";
    FD1S3AX o_wb_data_i1 (.D(o_wb_data_31__N_1337[1]), .CK(dac_clk_p_c), 
            .Q(wb_fm_data[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(39[8] 41[4])
    defparam o_wb_data_i1.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i30 (.D(n1[30]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_ls[30])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_ls__i30.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i29 (.D(n1[29]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_ls[29])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_ls__i29.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i28 (.D(n1[28]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_ls[28])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_ls__i28.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i27 (.D(n1[27]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_ls[27])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_ls__i27.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i26 (.D(n1[26]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_ls[26])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_ls__i26.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i25 (.D(n1[25]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_ls[25])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_ls__i25.GSR = "DISABLED";
    LUT4 i10866_3_lut (.A(n13522), .B(n36_adj_2992), .C(sine_lookup_width_minus_modulation_deviation_amount[2]), 
         .Z(n13523)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(74[27:78])
    defparam i10866_3_lut.init = 16'hcaca;
    FD1S3DX carrier_center_increment_offset_ls__i24 (.D(n1[24]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_ls[24])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_ls__i24.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i23 (.D(n1[23]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_ls[23])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_ls__i23.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i22 (.D(n1[22]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_ls[22])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_ls__i22.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i21 (.D(n1[21]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_ls[21])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_ls__i21.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i20 (.D(n1[20]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_ls[20])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_ls__i20.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i19 (.D(n1[19]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_ls[19])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_ls__i19.GSR = "DISABLED";
    LUT4 modulation_output_15__I_0_i71_3_lut (.A(n40_adj_2993), .B(n44), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[2]), .Z(n71)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam modulation_output_15__I_0_i71_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i40_3_lut (.A(n9), .B(n11), .C(sine_lookup_width_minus_modulation_deviation_amount[1]), 
         .Z(n40_adj_2993)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam modulation_output_15__I_0_i40_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i44_3_lut (.A(n13), .B(n15), .C(sine_lookup_width_minus_modulation_deviation_amount[1]), 
         .Z(n44)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam modulation_output_15__I_0_i44_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i15_3_lut (.A(modulation_output[14]), .B(modulation_output[15]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[0]), .Z(n15)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam modulation_output_15__I_0_i15_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i13_3_lut (.A(modulation_output[12]), .B(modulation_output[13]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[0]), .Z(n13)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam modulation_output_15__I_0_i13_3_lut.init = 16'hcaca;
    LUT4 i10865_3_lut (.A(modulation_output[2]), .B(modulation_output[3]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[0]), .Z(n13522)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(74[27:78])
    defparam i10865_3_lut.init = 16'hcaca;
    FD1S3DX carrier_center_increment_offset_ls__i18 (.D(n1[18]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_ls[18])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_ls__i18.GSR = "DISABLED";
    LUT4 i10869_3_lut (.A(n13524), .B(n7), .C(sine_lookup_width_minus_modulation_deviation_amount[1]), 
         .Z(n36_adj_2992)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(74[27:78])
    defparam i10869_3_lut.init = 16'hcaca;
    FD1S3DX carrier_center_increment_offset_ls__i17 (.D(n1[17]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_ls[17])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_ls__i17.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i16 (.D(n1[16]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_ls[16])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_ls__i16.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i15 (.D(n1[15]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_ls[15])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_ls__i15.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i14 (.D(n1[14]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_ls[14])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_ls__i14.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i13 (.D(n1[13]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_ls[13])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_ls__i13.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i12 (.D(n1[12]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_ls[12])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_ls__i12.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i11 (.D(n1[11]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_ls[11])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_ls__i11.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i10 (.D(n1[10]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_ls[10])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_ls__i10.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i9 (.D(n1[9]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_ls[9])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_ls__i9.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i8 (.D(n1[8]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_ls[8])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_ls__i8.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i7 (.D(n1[7]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_ls[7])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_ls__i7.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i6 (.D(n1[6]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_ls[6])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_ls__i6.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i5 (.D(n1[5]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_ls[5])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_ls__i5.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i4 (.D(n1[4]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_ls[4])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_ls__i4.GSR = "DISABLED";
    LUT4 i10867_3_lut (.A(modulation_output[4]), .B(modulation_output[5]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[0]), .Z(n13524)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(74[27:78])
    defparam i10867_3_lut.init = 16'hcaca;
    FD1S3DX carrier_center_increment_offset_ls__i3 (.D(n1[3]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_ls[3])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_ls__i3.GSR = "DISABLED";
    FD1S3DX carrier_center_increment_offset_ls__i2 (.D(n1[2]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_ls[2])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_ls__i2.GSR = "DISABLED";
    LUT4 i10868_3_lut (.A(modulation_output[6]), .B(modulation_output[7]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[0]), .Z(n7)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(74[27:78])
    defparam i10868_3_lut.init = 16'hcaca;
    FD1S3DX carrier_center_increment_offset_ls__i1 (.D(n20382), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(carrier_center_increment_offset_ls[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam carrier_center_increment_offset_ls__i1.GSR = "DISABLED";
    LUT4 modulation_output_15__I_0_i9_3_lut (.A(modulation_output[8]), .B(modulation_output[9]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[0]), .Z(n9)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam modulation_output_15__I_0_i9_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i11_3_lut (.A(modulation_output[10]), .B(modulation_output[11]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[0]), .Z(n11)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam modulation_output_15__I_0_i11_3_lut.init = 16'hcaca;
    LUT4 i10864_3_lut (.A(modulation_output[0]), .B(modulation_output[1]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[0]), .Z(n13521)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(74[27:78])
    defparam i10864_3_lut.init = 16'hcaca;
    LUT4 i22658_4_lut (.A(n26764), .B(sine_lookup_width_minus_modulation_deviation_amount[3]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[2]), .D(sine_lookup_width_minus_modulation_deviation_amount[1]), 
         .Z(n22451)) /* synthesis lut_function=(A+!(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam i22658_4_lut.init = 16'haaab;
    LUT4 i10874_3_lut (.A(n13530), .B(n37_adj_3000), .C(sine_lookup_width_minus_modulation_deviation_amount[2]), 
         .Z(n33_adj_3001)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(74[27:78])
    defparam i10874_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i72_3_lut (.A(n41_adj_3002), .B(n45_adj_3003), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[2]), .Z(n72_adj_3004)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam modulation_output_15__I_0_i72_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i45_3_lut (.A(n14), .B(modulation_output[15]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[1]), .Z(n45_adj_3003)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam modulation_output_15__I_0_i45_3_lut.init = 16'hcaca;
    LUT4 i10873_3_lut (.A(modulation_output[3]), .B(modulation_output[4]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[0]), .Z(n13530)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(74[27:78])
    defparam i10873_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i37_3_lut (.A(n6), .B(n8), .C(sine_lookup_width_minus_modulation_deviation_amount[1]), 
         .Z(n37_adj_3000)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam modulation_output_15__I_0_i37_3_lut.init = 16'hcaca;
    LUT4 i10875_3_lut (.A(modulation_output[5]), .B(modulation_output[6]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[0]), .Z(n6)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(74[27:78])
    defparam i10875_3_lut.init = 16'hcaca;
    LUT4 i10881_3_lut (.A(modulation_output[7]), .B(modulation_output[8]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[0]), .Z(n8)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(74[27:78])
    defparam i10881_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i14_3_lut (.A(modulation_output[13]), .B(modulation_output[14]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[0]), .Z(n14)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam modulation_output_15__I_0_i14_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i41_3_lut (.A(n10), .B(n12), .C(sine_lookup_width_minus_modulation_deviation_amount[1]), 
         .Z(n41_adj_3002)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam modulation_output_15__I_0_i41_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i10_3_lut (.A(modulation_output[9]), .B(modulation_output[10]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[0]), .Z(n10)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam modulation_output_15__I_0_i10_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i12_3_lut (.A(modulation_output[11]), .B(modulation_output[12]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[0]), .Z(n12)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam modulation_output_15__I_0_i12_3_lut.init = 16'hcaca;
    LUT4 i10872_3_lut (.A(modulation_output[1]), .B(modulation_output[2]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[0]), .Z(n13529)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(74[27:78])
    defparam i10872_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i38_3_lut (.A(n7), .B(n9), .C(sine_lookup_width_minus_modulation_deviation_amount[1]), 
         .Z(n38_adj_3005)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam modulation_output_15__I_0_i38_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i73_3_lut (.A(n42_adj_3006), .B(n46_adj_3007), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[2]), .Z(n73)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam modulation_output_15__I_0_i73_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i42_3_lut (.A(n11), .B(n13), .C(sine_lookup_width_minus_modulation_deviation_amount[1]), 
         .Z(n42_adj_3006)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam modulation_output_15__I_0_i42_3_lut.init = 16'hcaca;
    LUT4 i19699_3_lut (.A(\addr_space[2] [29]), .B(\addr_space[3] [29]), 
         .C(\wb_addr[0] ), .Z(n22136)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19699_3_lut.init = 16'hcaca;
    PFUMX i22950 (.BLUT(n24635), .ALUT(n38_adj_3005), .C0(sine_lookup_width_minus_modulation_deviation_amount[2]), 
          .Z(n24636));
    LUT4 i19698_3_lut (.A(\addr_space[0] [29]), .B(\addr_space[1] [29]), 
         .C(\wb_addr[0] ), .Z(n22135)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19698_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i64_3_lut (.A(n33_adj_3001), .B(n72_adj_3004), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[3]), .Z(n64)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam modulation_output_15__I_0_i64_3_lut.init = 16'hcaca;
    LUT4 i19690_3_lut (.A(\addr_space[2] [30]), .B(\addr_space[3] [30]), 
         .C(\wb_addr[0] ), .Z(n22127)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19690_3_lut.init = 16'hcaca;
    LUT4 i19689_3_lut (.A(\addr_space[0] [30]), .B(\addr_space[1] [30]), 
         .C(\wb_addr[0] ), .Z(n22126)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19689_3_lut.init = 16'hcaca;
    LUT4 i19684_3_lut (.A(\addr_space[2] [31]), .B(\addr_space[3] [31]), 
         .C(\wb_addr[0] ), .Z(n22121)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19684_3_lut.init = 16'hcaca;
    LUT4 i19683_3_lut (.A(\addr_space[0] [31]), .B(\addr_space[1] [31]), 
         .C(\wb_addr[0] ), .Z(n22120)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19683_3_lut.init = 16'hcaca;
    LUT4 i11847_2_lut_4_lut (.A(n85), .B(n26741), .C(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .D(n26742), .Z(n1[8])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(74[80:131])
    defparam i11847_2_lut_4_lut.init = 16'h00ca;
    LUT4 i19681_3_lut (.A(\addr_space[2] [0]), .B(\addr_space[3] [0]), .C(\wb_addr[0] ), 
         .Z(n22118)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19681_3_lut.init = 16'hcaca;
    LUT4 i19680_3_lut (.A(\addr_space[0] [0]), .B(\addr_space[1] [0]), .C(\wb_addr[0] ), 
         .Z(n22117)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19680_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_332_i112_3_lut_rep_403 (.A(n81), .B(n89), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[3]), .Z(n26726)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i112_3_lut_rep_403.init = 16'hcaca;
    LUT4 i18952_3_lut (.A(\addr_space[2] [1]), .B(\addr_space[3] [1]), .C(\wb_addr[0] ), 
         .Z(n21389)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18952_3_lut.init = 16'hcaca;
    LUT4 i18951_3_lut (.A(\addr_space[0] [1]), .B(\addr_space[1] [1]), .C(\wb_addr[0] ), 
         .Z(n21388)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18951_3_lut.init = 16'hcaca;
    LUT4 i18949_3_lut (.A(\addr_space[2] [2]), .B(\addr_space[3] [2]), .C(\wb_addr[0] ), 
         .Z(n21386)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18949_3_lut.init = 16'hcaca;
    LUT4 i11855_2_lut_4_lut (.A(n81), .B(n89), .C(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .D(n26742), .Z(n1[12])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam i11855_2_lut_4_lut.init = 16'h00ca;
    LUT4 i18948_3_lut (.A(\addr_space[0] [2]), .B(\addr_space[1] [2]), .C(\wb_addr[0] ), 
         .Z(n21385)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18948_3_lut.init = 16'hcaca;
    CCU2D add_384_31 (.A0(\addr_space[0] [29]), .B0(n14428), .C0(carrier_center_increment_offset_rs[30]), 
          .D0(carrier_center_increment_offset_ls[29]), .A1(\addr_space[0] [30]), 
          .B1(n14428), .C1(carrier_center_increment_offset_rs[30]), .D1(carrier_center_increment_offset_ls[30]), 
          .CIN(n17622), .S0(carrier_increment_30__N_1591[29]), .S1(carrier_increment_30__N_1591[30]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(92[4:87])
    defparam add_384_31.INIT0 = 16'h569a;
    defparam add_384_31.INIT1 = 16'h569a;
    defparam add_384_31.INJECT1_0 = "NO";
    defparam add_384_31.INJECT1_1 = "NO";
    LUT4 modulation_output_15__I_0_332_i111_3_lut_rep_404 (.A(n80), .B(n88), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[3]), .Z(n26727)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i111_3_lut_rep_404.init = 16'hcaca;
    LUT4 i18946_3_lut (.A(\addr_space[2] [3]), .B(\addr_space[3] [3]), .C(\wb_addr[0] ), 
         .Z(n21383)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18946_3_lut.init = 16'hcaca;
    LUT4 i11858_2_lut_4_lut (.A(n80), .B(n88), .C(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .D(n26742), .Z(n1[13])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam i11858_2_lut_4_lut.init = 16'h00ca;
    LUT4 modulation_output_15__I_0_332_i110_3_lut_rep_405 (.A(n79), .B(n26757), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[3]), .Z(n26728)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i110_3_lut_rep_405.init = 16'hcaca;
    LUT4 i18945_3_lut (.A(\addr_space[0] [3]), .B(\addr_space[1] [3]), .C(\wb_addr[0] ), 
         .Z(n21382)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18945_3_lut.init = 16'hcaca;
    LUT4 i11859_2_lut_4_lut (.A(n79), .B(n26757), .C(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .D(n26742), .Z(n1[14])) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam i11859_2_lut_4_lut.init = 16'h00ca;
    LUT4 i6638_3_lut_4_lut (.A(sine_lookup_width_minus_modulation_deviation_amount[2]), 
         .B(n26758), .C(modulation_output[15]), .D(n44), .Z(carrier_center_increment_offset_rs_30__N_1560[12])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam i6638_3_lut_4_lut.init = 16'hf1e0;
    LUT4 modulation_output_15__I_0_332_i86_3_lut_rep_433 (.A(n55), .B(n59), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[2]), .Z(n26756)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i86_3_lut_rep_433.init = 16'hcaca;
    LUT4 i18943_3_lut (.A(\addr_space[2] [4]), .B(\addr_space[3] [4]), .C(\wb_addr[0] ), 
         .Z(n21380)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18943_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_332_i101_3_lut (.A(modulation_output[15]), 
         .B(n78), .C(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .Z(n101)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i101_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_332_i102_3_lut (.A(modulation_output[15]), 
         .B(n79), .C(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .Z(n102)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i102_3_lut.init = 16'hcaca;
    LUT4 i6636_3_lut_4_lut (.A(sine_lookup_width_minus_modulation_deviation_amount[2]), 
         .B(n26758), .C(modulation_output[15]), .D(n43_adj_3008), .Z(carrier_center_increment_offset_rs_30__N_1560[11])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam i6636_3_lut_4_lut.init = 16'hf1e0;
    LUT4 modulation_output_15__I_0_332_i105_4_lut (.A(n82), .B(n59), .C(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .D(n26914), .Z(n105)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i105_4_lut.init = 16'hca0a;
    LUT4 i18942_3_lut (.A(\addr_space[0] [4]), .B(\addr_space[1] [4]), .C(\wb_addr[0] ), 
         .Z(n21379)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18942_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_332_i74_3_lut (.A(modulation_output[15]), 
         .B(n47_adj_3009), .C(modulation_deviation_amount_minus_sine_lookup_width[2]), 
         .Z(n74)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i74_3_lut.init = 16'hcaca;
    LUT4 i18940_3_lut (.A(\addr_space[2] [5]), .B(\addr_space[3] [5]), .C(\wb_addr[0] ), 
         .Z(n21377)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18940_3_lut.init = 16'hcaca;
    LUT4 i18939_3_lut (.A(\addr_space[0] [5]), .B(\addr_space[1] [5]), .C(\wb_addr[0] ), 
         .Z(n21376)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18939_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_332_i106_4_lut (.A(n83), .B(n60), .C(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .D(n26914), .Z(n106)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i106_4_lut.init = 16'hca0a;
    LUT4 modulation_output_15__I_0_332_i75_3_lut (.A(modulation_output[15]), 
         .B(n48_adj_3010), .C(modulation_deviation_amount_minus_sine_lookup_width[2]), 
         .Z(n75)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i75_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_332_i87_3_lut_rep_434 (.A(n56), .B(n60), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[2]), .Z(n26757)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i87_3_lut_rep_434.init = 16'hcaca;
    LUT4 i10870_3_lut (.A(n13523), .B(n71), .C(sine_lookup_width_minus_modulation_deviation_amount[3]), 
         .Z(n63)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(74[27:78])
    defparam i10870_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut (.A(n26946), .B(n38), .C(n34), .D(n20781), .Z(dac_clk_p_c_enable_147)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_4_lut.init = 16'h0100;
    LUT4 i18937_3_lut (.A(\addr_space[2] [6]), .B(\addr_space[3] [6]), .C(\wb_addr[0] ), 
         .Z(n21374)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18937_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_92 (.A(n20775), .B(\wb_addr[8] ), .C(\wb_addr[12] ), 
         .D(n20773), .Z(n20781)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_4_lut_adj_92.init = 16'h0200;
    LUT4 i18936_3_lut (.A(\addr_space[0] [6]), .B(\addr_space[1] [6]), .C(\wb_addr[0] ), 
         .Z(n21373)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18936_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_93 (.A(n26947), .B(\wb_addr[15] ), .C(\wb_addr[9] ), 
         .D(i_resetb_c), .Z(n20775)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_93.init = 16'h8000;
    LUT4 i18934_3_lut (.A(\addr_space[2] [7]), .B(\addr_space[3] [7]), .C(\wb_addr[0] ), 
         .Z(n21371)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18934_3_lut.init = 16'hcaca;
    PFUMX i24724 (.BLUT(n26690), .ALUT(n26689), .C0(sine_lookup_width_minus_modulation_deviation_amount[3]), 
          .Z(n26691));
    LUT4 i1_2_lut (.A(\wb_addr[0] ), .B(\wb_addr[1] ), .Z(n20773)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i18933_3_lut (.A(\addr_space[0] [7]), .B(\addr_space[1] [7]), .C(\wb_addr[0] ), 
         .Z(n21370)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18933_3_lut.init = 16'hcaca;
    LUT4 i18931_3_lut (.A(\addr_space[2] [8]), .B(\addr_space[3] [8]), .C(\wb_addr[0] ), 
         .Z(n21368)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18931_3_lut.init = 16'hcaca;
    PFUMX modulation_output_15__I_0_332_i135 (.BLUT(n73_adj_3013), .ALUT(n104), 
          .C0(n22285), .Z(n135)) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;
    PFUMX modulation_output_15__I_0_332_i134 (.BLUT(n72), .ALUT(n103), .C0(n22285), 
          .Z(n134)) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;
    LUT4 i18930_3_lut (.A(\addr_space[0] [8]), .B(\addr_space[1] [8]), .C(\wb_addr[0] ), 
         .Z(n21367)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18930_3_lut.init = 16'hcaca;
    LUT4 i18928_3_lut (.A(\addr_space[2] [9]), .B(\addr_space[3] [9]), .C(\wb_addr[0] ), 
         .Z(n21365)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18928_3_lut.init = 16'hcaca;
    LUT4 i18927_3_lut (.A(\addr_space[0] [9]), .B(\addr_space[1] [9]), .C(\wb_addr[0] ), 
         .Z(n21364)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18927_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_rep_435 (.A(sine_lookup_width_minus_modulation_deviation_amount[3]), 
         .B(n178), .C(sine_lookup_width_minus_modulation_deviation_amount[4]), 
         .Z(n26758)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam i1_3_lut_rep_435.init = 16'hfefe;
    PFUMX i24710 (.BLUT(n26672), .ALUT(n26671), .C0(sine_lookup_width_minus_modulation_deviation_amount[3]), 
          .Z(n26673));
    LUT4 i1_2_lut_rep_463_3_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .B(modulation_output[0]), .C(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .Z(n26786)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i1_2_lut_rep_463_3_lut.init = 16'h0404;
    PFUMX i24704 (.BLUT(n26663), .ALUT(n26662), .C0(sine_lookup_width_minus_modulation_deviation_amount[3]), 
          .Z(n26664));
    LUT4 i18925_3_lut (.A(\addr_space[2] [10]), .B(\addr_space[3] [10]), 
         .C(\wb_addr[0] ), .Z(n21362)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18925_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_94 (.A(n20945), .B(n20947), .C(n20949), .D(n20935), 
         .Z(n178)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam i1_4_lut_adj_94.init = 16'hfffe;
    LUT4 i1_2_lut_adj_95 (.A(sine_lookup_width_minus_modulation_deviation_amount[14]), 
         .B(sine_lookup_width_minus_modulation_deviation_amount[5]), .Z(n20945)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam i1_2_lut_adj_95.init = 16'heeee;
    LUT4 i1_4_lut_adj_96 (.A(sine_lookup_width_minus_modulation_deviation_amount[6]), 
         .B(sine_lookup_width_minus_modulation_deviation_amount[15]), .C(sine_lookup_width_minus_modulation_deviation_amount[16]), 
         .D(sine_lookup_width_minus_modulation_deviation_amount[9]), .Z(n20947)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam i1_4_lut_adj_96.init = 16'hfffe;
    LUT4 i1_4_lut_adj_97 (.A(sine_lookup_width_minus_modulation_deviation_amount[12]), 
         .B(sine_lookup_width_minus_modulation_deviation_amount[8]), .C(sine_lookup_width_minus_modulation_deviation_amount[11]), 
         .D(sine_lookup_width_minus_modulation_deviation_amount[13]), .Z(n20949)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam i1_4_lut_adj_97.init = 16'hfffe;
    LUT4 i18924_3_lut (.A(\addr_space[0] [10]), .B(\addr_space[1] [10]), 
         .C(\wb_addr[0] ), .Z(n21361)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18924_3_lut.init = 16'hcaca;
    LUT4 i18922_3_lut (.A(\addr_space[2] [11]), .B(\addr_space[3] [11]), 
         .C(\wb_addr[0] ), .Z(n21359)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18922_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_98 (.A(sine_lookup_width_minus_modulation_deviation_amount[7]), 
         .B(sine_lookup_width_minus_modulation_deviation_amount[10]), .Z(n20935)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam i1_2_lut_adj_98.init = 16'heeee;
    LUT4 i18921_3_lut (.A(\addr_space[0] [11]), .B(\addr_space[1] [11]), 
         .C(\wb_addr[0] ), .Z(n21358)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18921_3_lut.init = 16'hcaca;
    LUT4 i19780_3_lut (.A(\addr_space[2] [12]), .B(\addr_space[3] [12]), 
         .C(\wb_addr[0] ), .Z(n22217)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19780_3_lut.init = 16'hcaca;
    LUT4 i19779_3_lut (.A(\addr_space[0] [12]), .B(\addr_space[1] [12]), 
         .C(\wb_addr[0] ), .Z(n22216)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19779_3_lut.init = 16'hcaca;
    LUT4 i19777_3_lut (.A(\addr_space[2] [13]), .B(\addr_space[3] [13]), 
         .C(\wb_addr[0] ), .Z(n22214)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19777_3_lut.init = 16'hcaca;
    LUT4 i19776_3_lut (.A(\addr_space[0] [13]), .B(\addr_space[1] [13]), 
         .C(\wb_addr[0] ), .Z(n22213)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19776_3_lut.init = 16'hcaca;
    PFUMX i24701 (.BLUT(n26658), .ALUT(n39_adj_3014), .C0(sine_lookup_width_minus_modulation_deviation_amount[2]), 
          .Z(n26659));
    LUT4 i19774_3_lut (.A(\addr_space[2] [14]), .B(\addr_space[3] [14]), 
         .C(\wb_addr[0] ), .Z(n22211)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19774_3_lut.init = 16'hcaca;
    LUT4 i19773_3_lut (.A(\addr_space[0] [14]), .B(\addr_space[1] [14]), 
         .C(\wb_addr[0] ), .Z(n22210)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19773_3_lut.init = 16'hcaca;
    LUT4 i19771_3_lut (.A(\addr_space[2] [15]), .B(\addr_space[3] [15]), 
         .C(\wb_addr[0] ), .Z(n22208)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19771_3_lut.init = 16'hcaca;
    LUT4 i19770_3_lut (.A(\addr_space[0] [15]), .B(\addr_space[1] [15]), 
         .C(\wb_addr[0] ), .Z(n22207)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19770_3_lut.init = 16'hcaca;
    LUT4 i19768_3_lut (.A(\addr_space[2] [16]), .B(\addr_space[3] [16]), 
         .C(\wb_addr[0] ), .Z(n22205)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19768_3_lut.init = 16'hcaca;
    LUT4 i19767_3_lut (.A(\addr_space[0] [16]), .B(\addr_space[1] [16]), 
         .C(\wb_addr[0] ), .Z(n22204)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19767_3_lut.init = 16'hcaca;
    LUT4 i19765_3_lut (.A(\addr_space[2] [17]), .B(\addr_space[3] [17]), 
         .C(\wb_addr[0] ), .Z(n22202)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19765_3_lut.init = 16'hcaca;
    LUT4 i19764_3_lut (.A(\addr_space[0] [17]), .B(\addr_space[1] [17]), 
         .C(\wb_addr[0] ), .Z(n22201)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19764_3_lut.init = 16'hcaca;
    LUT4 i19762_3_lut (.A(\addr_space[2] [18]), .B(\addr_space[3] [18]), 
         .C(\wb_addr[0] ), .Z(n22199)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19762_3_lut.init = 16'hcaca;
    LUT4 i19761_3_lut (.A(\addr_space[0] [18]), .B(\addr_space[1] [18]), 
         .C(\wb_addr[0] ), .Z(n22198)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19761_3_lut.init = 16'hcaca;
    LUT4 i19759_3_lut (.A(\addr_space[2] [19]), .B(\addr_space[3] [19]), 
         .C(\wb_addr[0] ), .Z(n22196)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19759_3_lut.init = 16'hcaca;
    LUT4 i19758_3_lut (.A(\addr_space[0] [19]), .B(\addr_space[1] [19]), 
         .C(\wb_addr[0] ), .Z(n22195)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19758_3_lut.init = 16'hcaca;
    LUT4 i19756_3_lut (.A(\addr_space[2] [20]), .B(\addr_space[3] [20]), 
         .C(\wb_addr[0] ), .Z(n22193)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19756_3_lut.init = 16'hcaca;
    LUT4 i19755_3_lut (.A(\addr_space[0] [20]), .B(\addr_space[1] [20]), 
         .C(\wb_addr[0] ), .Z(n22192)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19755_3_lut.init = 16'hcaca;
    LUT4 i6642_4_lut (.A(modulation_output[14]), .B(modulation_output[15]), 
         .C(n9080), .D(n26758), .Z(carrier_center_increment_offset_rs_30__N_1560[14])) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam i6642_4_lut.init = 16'hccca;
    LUT4 i6640_4_lut (.A(n14), .B(modulation_output[15]), .C(n9078), .D(n26758), 
         .Z(carrier_center_increment_offset_rs_30__N_1560[13])) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam i6640_4_lut.init = 16'hccca;
    LUT4 i6582_2_lut (.A(sine_lookup_width_minus_modulation_deviation_amount[1]), 
         .B(sine_lookup_width_minus_modulation_deviation_amount[2]), .Z(n9078)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam i6582_2_lut.init = 16'heeee;
    LUT4 modulation_output_15__I_0_i43_3_lut (.A(n12), .B(n14), .C(sine_lookup_width_minus_modulation_deviation_amount[1]), 
         .Z(n43_adj_3008)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam modulation_output_15__I_0_i43_3_lut.init = 16'hcaca;
    LUT4 i6634_3_lut (.A(n73), .B(modulation_output[15]), .C(n26758), 
         .Z(carrier_center_increment_offset_rs_30__N_1560[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam i6634_3_lut.init = 16'hcaca;
    LUT4 i6632_3_lut (.A(n72_adj_3004), .B(modulation_output[15]), .C(n26758), 
         .Z(carrier_center_increment_offset_rs_30__N_1560[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam i6632_3_lut.init = 16'hcaca;
    LUT4 i6630_3_lut (.A(n71), .B(modulation_output[15]), .C(n26758), 
         .Z(carrier_center_increment_offset_rs_30__N_1560[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam i6630_3_lut.init = 16'hcaca;
    LUT4 i19753_3_lut (.A(\addr_space[2] [21]), .B(\addr_space[3] [21]), 
         .C(\wb_addr[0] ), .Z(n22190)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19753_3_lut.init = 16'hcaca;
    LUT4 i6628_3_lut (.A(n70), .B(modulation_output[15]), .C(n26758), 
         .Z(carrier_center_increment_offset_rs_30__N_1560[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam i6628_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i70_3_lut (.A(n39_adj_3014), .B(n43_adj_3008), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[2]), .Z(n70)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam modulation_output_15__I_0_i70_3_lut.init = 16'hcaca;
    LUT4 i19752_3_lut (.A(\addr_space[0] [21]), .B(\addr_space[1] [21]), 
         .C(\wb_addr[0] ), .Z(n22189)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19752_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_i39_3_lut (.A(n8), .B(n10), .C(sine_lookup_width_minus_modulation_deviation_amount[1]), 
         .Z(n39_adj_3014)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam modulation_output_15__I_0_i39_3_lut.init = 16'hcaca;
    LUT4 i11039_4_lut (.A(modulation_output[15]), .B(n178_adj_3015), .C(n26728), 
         .D(modulation_deviation_amount_minus_sine_lookup_width[4]), .Z(n1[30])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i11039_4_lut.init = 16'h3022;
    LUT4 modulation_output_15__I_0_332_i79_3_lut (.A(n48_adj_3010), .B(n52_adj_3016), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[2]), .Z(n79)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i79_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_332_i56_3_lut (.A(n25), .B(n27), .C(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .Z(n56)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i56_3_lut.init = 16'hcaca;
    LUT4 i10882_3_lut (.A(modulation_output[2]), .B(modulation_output[1]), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[0]), .Z(n29)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(74[80:131])
    defparam i10882_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_332_i48_3_lut (.A(n17), .B(n19), .C(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .Z(n48_adj_3010)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i48_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_332_i52_3_lut (.A(n21), .B(n23), .C(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .Z(n52_adj_3016)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i52_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_332_i21_3_lut (.A(modulation_output[10]), 
         .B(modulation_output[9]), .C(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .Z(n21)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i21_3_lut.init = 16'hcaca;
    LUT4 i10880_3_lut (.A(modulation_output[8]), .B(modulation_output[7]), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[0]), .Z(n23)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(74[80:131])
    defparam i10880_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_332_i17_3_lut (.A(modulation_output[14]), 
         .B(modulation_output[13]), .C(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .Z(n17)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i17_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_332_i19_3_lut (.A(modulation_output[12]), 
         .B(modulation_output[11]), .C(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .Z(n19)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i19_3_lut.init = 16'hcaca;
    LUT4 i19750_3_lut (.A(\addr_space[2] [22]), .B(\addr_space[3] [22]), 
         .C(\wb_addr[0] ), .Z(n22187)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19750_3_lut.init = 16'hcaca;
    LUT4 i10883_3_lut (.A(modulation_output[6]), .B(modulation_output[5]), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[0]), .Z(n25)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(74[80:131])
    defparam i10883_3_lut.init = 16'hcaca;
    LUT4 i10888_3_lut (.A(modulation_output[4]), .B(modulation_output[3]), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[0]), .Z(n27)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(74[80:131])
    defparam i10888_3_lut.init = 16'hcaca;
    LUT4 i11040_4_lut (.A(n95_adj_3017), .B(n178_adj_3015), .C(n26727), 
         .D(modulation_deviation_amount_minus_sine_lookup_width[4]), .Z(n1[29])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i11040_4_lut.init = 16'h3022;
    LUT4 i6549_4_lut (.A(modulation_output[15]), .B(modulation_output[14]), 
         .C(n26801), .D(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .Z(n95_adj_3017)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C (D)))) */ ;
    defparam i6549_4_lut.init = 16'hcaaa;
    LUT4 modulation_output_15__I_0_332_i80_3_lut (.A(n49_adj_3018), .B(n53_adj_3019), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[2]), .Z(n80)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i80_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_332_i88_4_lut (.A(n57_adj_3020), .B(n30), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[2]), .D(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .Z(n88)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i88_4_lut.init = 16'h0aca;
    LUT4 modulation_output_15__I_0_332_i49_3_lut (.A(n18), .B(n20), .C(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .Z(n49_adj_3018)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i49_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_332_i53_3_lut (.A(n22), .B(n24), .C(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .Z(n53_adj_3019)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i53_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_332_i22_3_lut (.A(modulation_output[9]), 
         .B(modulation_output[8]), .C(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .Z(n22)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i22_3_lut.init = 16'hcaca;
    LUT4 i10885_3_lut (.A(modulation_output[7]), .B(modulation_output[6]), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[0]), .Z(n24)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(74[80:131])
    defparam i10885_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_332_i18_3_lut (.A(modulation_output[13]), 
         .B(modulation_output[12]), .C(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .Z(n18)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i18_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_332_i20_3_lut (.A(modulation_output[11]), 
         .B(modulation_output[10]), .C(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .Z(n20)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i20_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_332_i57_3_lut (.A(n26), .B(n28), .C(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .Z(n57_adj_3020)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i57_3_lut.init = 16'hcaca;
    LUT4 i10884_3_lut (.A(modulation_output[1]), .B(modulation_output[0]), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[0]), .Z(n30)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(74[80:131])
    defparam i10884_3_lut.init = 16'hcaca;
    LUT4 i10886_3_lut (.A(modulation_output[5]), .B(modulation_output[4]), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[0]), .Z(n26)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(74[80:131])
    defparam i10886_3_lut.init = 16'hcaca;
    LUT4 i10887_3_lut (.A(modulation_output[3]), .B(modulation_output[2]), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[0]), .Z(n28)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(74[80:131])
    defparam i10887_3_lut.init = 16'hcaca;
    LUT4 i19749_3_lut (.A(\addr_space[0] [22]), .B(\addr_space[1] [22]), 
         .C(\wb_addr[0] ), .Z(n22186)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19749_3_lut.init = 16'hcaca;
    LUT4 i11044_4_lut (.A(n96), .B(n178_adj_3015), .C(n26726), .D(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .Z(n1[28])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i11044_4_lut.init = 16'h3022;
    LUT4 i6551_4_lut (.A(modulation_output[15]), .B(n17), .C(n26916), 
         .D(modulation_deviation_amount_minus_sine_lookup_width[3]), .Z(n96)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C (D)))) */ ;
    defparam i6551_4_lut.init = 16'hcaaa;
    LUT4 modulation_output_15__I_0_332_i81_3_lut (.A(n50_adj_3021), .B(n54_adj_3022), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[2]), .Z(n81)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i81_3_lut.init = 16'hcaca;
    CCU2D add_384_29 (.A0(\addr_space[0] [27]), .B0(n14428), .C0(carrier_center_increment_offset_rs[30]), 
          .D0(carrier_center_increment_offset_ls[27]), .A1(\addr_space[0] [28]), 
          .B1(n14428), .C1(carrier_center_increment_offset_rs[30]), .D1(carrier_center_increment_offset_ls[28]), 
          .CIN(n17621), .COUT(n17622), .S0(carrier_increment_30__N_1591[27]), 
          .S1(carrier_increment_30__N_1591[28]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(92[4:87])
    defparam add_384_29.INIT0 = 16'h569a;
    defparam add_384_29.INIT1 = 16'h569a;
    defparam add_384_29.INJECT1_0 = "NO";
    defparam add_384_29.INJECT1_1 = "NO";
    LUT4 modulation_output_15__I_0_332_i50_3_lut (.A(n19), .B(n21), .C(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .Z(n50_adj_3021)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i50_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_332_i54_3_lut (.A(n23), .B(n25), .C(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .Z(n54_adj_3022)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i54_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_332_i58_3_lut (.A(n27), .B(n29), .C(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .Z(n58)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i58_3_lut.init = 16'hcaca;
    LUT4 i11046_4_lut (.A(n97), .B(n178_adj_3015), .C(n113), .D(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .Z(n1[27])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i11046_4_lut.init = 16'h3022;
    LUT4 modulation_output_15__I_0_332_i47_3_lut (.A(n16), .B(n18), .C(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .Z(n47_adj_3009)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i47_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_332_i16_3_lut (.A(modulation_output[15]), 
         .B(modulation_output[14]), .C(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .Z(n16)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i16_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_332_i113_4_lut (.A(n82), .B(n59), .C(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .D(modulation_deviation_amount_minus_sine_lookup_width[2]), .Z(n113)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i113_4_lut.init = 16'h0aca;
    LUT4 modulation_output_15__I_0_332_i82_3_lut (.A(n51_adj_3023), .B(n55), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[2]), .Z(n82)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i82_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_332_i59_3_lut (.A(n28), .B(n30), .C(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .Z(n59)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i59_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_332_i51_3_lut (.A(n20), .B(n22), .C(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .Z(n51_adj_3023)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i51_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_332_i55_3_lut (.A(n24), .B(n26), .C(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .Z(n55)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i55_3_lut.init = 16'hcaca;
    LUT4 i11047_4_lut (.A(n98), .B(n178_adj_3015), .C(n114), .D(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .Z(n1[26])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i11047_4_lut.init = 16'h3022;
    LUT4 modulation_output_15__I_0_332_i114_4_lut (.A(n83), .B(n60), .C(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .D(modulation_deviation_amount_minus_sine_lookup_width[2]), .Z(n114)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i114_4_lut.init = 16'h0aca;
    CCU2D add_384_27 (.A0(\addr_space[0] [25]), .B0(n14428), .C0(carrier_center_increment_offset_rs[30]), 
          .D0(carrier_center_increment_offset_ls[25]), .A1(\addr_space[0] [26]), 
          .B1(n14428), .C1(carrier_center_increment_offset_rs[30]), .D1(carrier_center_increment_offset_ls[26]), 
          .CIN(n17620), .COUT(n17621), .S0(carrier_increment_30__N_1591[25]), 
          .S1(carrier_increment_30__N_1591[26]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(92[4:87])
    defparam add_384_27.INIT0 = 16'h569a;
    defparam add_384_27.INIT1 = 16'h569a;
    defparam add_384_27.INJECT1_0 = "NO";
    defparam add_384_27.INJECT1_1 = "NO";
    LUT4 modulation_output_15__I_0_332_i83_3_lut (.A(n52_adj_3016), .B(n56), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[2]), .Z(n83)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i83_3_lut.init = 16'hcaca;
    LUT4 i11049_4_lut (.A(n99), .B(n178_adj_3015), .C(n115), .D(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .Z(n1[25])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i11049_4_lut.init = 16'h3022;
    LUT4 modulation_output_15__I_0_332_i99_3_lut (.A(modulation_output[15]), 
         .B(n76), .C(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .Z(n99)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i99_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_332_i76_3_lut (.A(n45_adj_3024), .B(n49_adj_3018), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[2]), .Z(n76)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i76_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_332_i115_4_lut (.A(n84), .B(n30), .C(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .D(n26915), .Z(n115)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i115_4_lut.init = 16'h0aca;
    LUT4 modulation_output_15__I_0_332_i84_3_lut (.A(n53_adj_3019), .B(n57_adj_3020), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[2]), .Z(n84)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i84_3_lut.init = 16'hcaca;
    LUT4 i19747_3_lut (.A(\addr_space[2] [23]), .B(\addr_space[3] [23]), 
         .C(\wb_addr[0] ), .Z(n22184)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19747_3_lut.init = 16'hcaca;
    LUT4 i11050_4_lut (.A(n100), .B(n178_adj_3015), .C(n26725), .D(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .Z(n1[24])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i11050_4_lut.init = 16'h3022;
    LUT4 modulation_output_15__I_0_332_i100_3_lut (.A(modulation_output[15]), 
         .B(n77), .C(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .Z(n100)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i100_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_332_i77_3_lut (.A(n46_adj_3025), .B(n50_adj_3021), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[2]), .Z(n77)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i77_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_332_i46_3_lut (.A(modulation_output[15]), 
         .B(n17), .C(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .Z(n46_adj_3025)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i46_3_lut.init = 16'hcaca;
    LUT4 i19746_3_lut (.A(\addr_space[0] [23]), .B(\addr_space[1] [23]), 
         .C(\wb_addr[0] ), .Z(n22183)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19746_3_lut.init = 16'hcaca;
    LUT4 modulation_output_15__I_0_332_i85_3_lut (.A(n54_adj_3022), .B(n58), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[2]), .Z(n85)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i85_3_lut.init = 16'hcaca;
    LUT4 i19744_3_lut (.A(\addr_space[2] [24]), .B(\addr_space[3] [24]), 
         .C(\wb_addr[0] ), .Z(n22181)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19744_3_lut.init = 16'hcaca;
    LUT4 i19743_3_lut (.A(\addr_space[0] [24]), .B(\addr_space[1] [24]), 
         .C(\wb_addr[0] ), .Z(n22180)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19743_3_lut.init = 16'hcaca;
    CCU2D add_384_25 (.A0(\addr_space[0] [23]), .B0(n14428), .C0(carrier_center_increment_offset_rs[30]), 
          .D0(carrier_center_increment_offset_ls[23]), .A1(\addr_space[0] [24]), 
          .B1(n14428), .C1(carrier_center_increment_offset_rs[30]), .D1(carrier_center_increment_offset_ls[24]), 
          .CIN(n17619), .COUT(n17620), .S0(carrier_increment_30__N_1591[23]), 
          .S1(carrier_increment_30__N_1591[24]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(92[4:87])
    defparam add_384_25.INIT0 = 16'h569a;
    defparam add_384_25.INIT1 = 16'h569a;
    defparam add_384_25.INJECT1_0 = "NO";
    defparam add_384_25.INJECT1_1 = "NO";
    LUT4 i11051_2_lut (.A(n132), .B(n178_adj_3015), .Z(n1[23])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i11051_2_lut.init = 16'h2222;
    LUT4 i11052_2_lut (.A(n133), .B(n178_adj_3015), .Z(n1[22])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i11052_2_lut.init = 16'h2222;
    LUT4 i19735_3_lut (.A(\addr_space[2] [25]), .B(\addr_space[3] [25]), 
         .C(\wb_addr[0] ), .Z(n22172)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19735_3_lut.init = 16'hcaca;
    LUT4 i11053_2_lut (.A(n134), .B(n178_adj_3015), .Z(n1[21])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i11053_2_lut.init = 16'h2222;
    LUT4 i11054_2_lut (.A(n135), .B(n178_adj_3015), .Z(n1[20])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i11054_2_lut.init = 16'h2222;
    LUT4 i11057_2_lut (.A(n136), .B(n178_adj_3015), .Z(n1[19])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i11057_2_lut.init = 16'h2222;
    LUT4 i11059_2_lut (.A(n137), .B(n178_adj_3015), .Z(n1[18])) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i11059_2_lut.init = 16'h2222;
    LUT4 i11062_4_lut (.A(n107), .B(n178_adj_3015), .C(n123), .D(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .Z(n1[17])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i11062_4_lut.init = 16'h3022;
    LUT4 modulation_output_15__I_0_332_i107_3_lut (.A(n76), .B(n84), .C(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .Z(n107)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i107_3_lut.init = 16'hcaca;
    LUT4 i11063_4_lut (.A(n108), .B(n178_adj_3015), .C(n26718), .D(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .Z(n1[16])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i11063_4_lut.init = 16'h3022;
    LUT4 modulation_output_15__I_0_332_i108_3_lut (.A(n77), .B(n85), .C(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .Z(n108)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i108_3_lut.init = 16'hcaca;
    LUT4 i11860_4_lut (.A(n78), .B(n26742), .C(n26756), .D(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .Z(n1[15])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i11860_4_lut.init = 16'h3022;
    LUT4 modulation_output_15__I_0_332_i78_3_lut (.A(n47_adj_3009), .B(n51_adj_3023), 
         .C(modulation_deviation_amount_minus_sine_lookup_width[2]), .Z(n78)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam modulation_output_15__I_0_332_i78_3_lut.init = 16'hcaca;
    LUT4 i19734_3_lut (.A(\addr_space[0] [25]), .B(\addr_space[1] [25]), 
         .C(\wb_addr[0] ), .Z(n22171)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19734_3_lut.init = 16'hcaca;
    LUT4 i19726_3_lut (.A(\addr_space[2] [26]), .B(\addr_space[3] [26]), 
         .C(\wb_addr[0] ), .Z(n22163)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19726_3_lut.init = 16'hcaca;
    LUT4 i19725_3_lut (.A(\addr_space[0] [26]), .B(\addr_space[1] [26]), 
         .C(\wb_addr[0] ), .Z(n22162)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19725_3_lut.init = 16'hcaca;
    CCU2D add_384_23 (.A0(\addr_space[0] [21]), .B0(n14428), .C0(carrier_center_increment_offset_rs[30]), 
          .D0(carrier_center_increment_offset_ls[21]), .A1(\addr_space[0] [22]), 
          .B1(n14428), .C1(carrier_center_increment_offset_rs[30]), .D1(carrier_center_increment_offset_ls[22]), 
          .CIN(n17618), .COUT(n17619), .S0(carrier_increment_30__N_1591[21]), 
          .S1(carrier_increment_30__N_1591[22]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(92[4:87])
    defparam add_384_23.INIT0 = 16'h569a;
    defparam add_384_23.INIT1 = 16'h569a;
    defparam add_384_23.INJECT1_0 = "NO";
    defparam add_384_23.INJECT1_1 = "NO";
    LUT4 i19717_3_lut (.A(\addr_space[2] [27]), .B(\addr_space[3] [27]), 
         .C(\wb_addr[0] ), .Z(n22154)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19717_3_lut.init = 16'hcaca;
    LUT4 i19716_3_lut (.A(\addr_space[0] [27]), .B(\addr_space[1] [27]), 
         .C(\wb_addr[0] ), .Z(n22153)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19716_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_99 (.A(n20665), .B(n20679), .C(n20677), .D(\addr_space[2] [4]), 
         .Z(n14428)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_99.init = 16'hfffe;
    LUT4 i1_2_lut_adj_100 (.A(\addr_space[2] [7]), .B(\addr_space[2] [13]), 
         .Z(n20665)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_100.init = 16'heeee;
    LUT4 i1_4_lut_adj_101 (.A(\addr_space[2] [16]), .B(n20663), .C(n20667), 
         .D(\addr_space[2] [9]), .Z(n20679)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_101.init = 16'hfffe;
    LUT4 i1_4_lut_adj_102 (.A(\addr_space[2] [6]), .B(\addr_space[2] [10]), 
         .C(\addr_space[2] [15]), .D(\addr_space[2] [8]), .Z(n20677)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_4_lut_adj_102.init = 16'hfffe;
    LUT4 i1_2_lut_adj_103 (.A(\addr_space[2] [5]), .B(\addr_space[2] [14]), 
         .Z(n20663)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_103.init = 16'heeee;
    LUT4 i1_2_lut_adj_104 (.A(\addr_space[2] [12]), .B(\addr_space[2] [11]), 
         .Z(n20667)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_104.init = 16'heeee;
    LUT4 i19708_3_lut (.A(\addr_space[2] [28]), .B(\addr_space[3] [28]), 
         .C(\wb_addr[0] ), .Z(n22145)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19708_3_lut.init = 16'hcaca;
    LUT4 i19707_3_lut (.A(\addr_space[0] [28]), .B(\addr_space[1] [28]), 
         .C(\wb_addr[0] ), .Z(n22144)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19707_3_lut.init = 16'hcaca;
    CCU2D add_384_21 (.A0(\addr_space[0] [19]), .B0(n14428), .C0(carrier_center_increment_offset_rs[30]), 
          .D0(carrier_center_increment_offset_ls[19]), .A1(\addr_space[0] [20]), 
          .B1(n14428), .C1(carrier_center_increment_offset_rs[30]), .D1(carrier_center_increment_offset_ls[20]), 
          .CIN(n17617), .COUT(n17618), .S0(carrier_increment_30__N_1591[19]), 
          .S1(carrier_increment_30__N_1591[20]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(92[4:87])
    defparam add_384_21.INIT0 = 16'h569a;
    defparam add_384_21.INIT1 = 16'h569a;
    defparam add_384_21.INJECT1_0 = "NO";
    defparam add_384_21.INJECT1_1 = "NO";
    LUT4 i22725_2_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[3]), .Z(n22285)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam i22725_2_lut.init = 16'heeee;
    CCU2D add_384_19 (.A0(\addr_space[0] [17]), .B0(n14428), .C0(carrier_center_increment_offset_rs[30]), 
          .D0(carrier_center_increment_offset_ls[17]), .A1(\addr_space[0] [18]), 
          .B1(n14428), .C1(carrier_center_increment_offset_rs[30]), .D1(carrier_center_increment_offset_ls[18]), 
          .CIN(n17616), .COUT(n17617), .S0(carrier_increment_30__N_1591[17]), 
          .S1(carrier_increment_30__N_1591[18]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(92[4:87])
    defparam add_384_19.INIT0 = 16'h569a;
    defparam add_384_19.INIT1 = 16'h569a;
    defparam add_384_19.INJECT1_0 = "NO";
    defparam add_384_19.INJECT1_1 = "NO";
    CCU2D add_384_17 (.A0(\addr_space[0] [15]), .B0(n14428), .C0(carrier_center_increment_offset_rs[30]), 
          .D0(carrier_center_increment_offset_ls[15]), .A1(\addr_space[0] [16]), 
          .B1(n14428), .C1(carrier_center_increment_offset_rs[30]), .D1(carrier_center_increment_offset_ls[16]), 
          .CIN(n17615), .COUT(n17616), .S0(carrier_increment_30__N_1591[15]), 
          .S1(carrier_increment_30__N_1591[16]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(92[4:87])
    defparam add_384_17.INIT0 = 16'h569a;
    defparam add_384_17.INIT1 = 16'h569a;
    defparam add_384_17.INJECT1_0 = "NO";
    defparam add_384_17.INJECT1_1 = "NO";
    LUT4 i6623_2_lut_rep_441 (.A(sine_lookup_width_minus_modulation_deviation_amount[4]), 
         .B(n178), .Z(n26764)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam i6623_2_lut_rep_441.init = 16'heeee;
    LUT4 i1_2_lut_3_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[2]), 
         .B(n26786), .C(n26742), .D(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .Z(n1[0])) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0004;
    LUT4 n26660_bdd_3_lut_4_lut (.A(sine_lookup_width_minus_modulation_deviation_amount[4]), 
         .B(n178), .C(modulation_output[15]), .D(n26660), .Z(carrier_center_increment_offset_rs_30__N_1560[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam n26660_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n26673_bdd_3_lut_4_lut (.A(sine_lookup_width_minus_modulation_deviation_amount[4]), 
         .B(n178), .C(modulation_output[15]), .D(n26673), .Z(carrier_center_increment_offset_rs_30__N_1560[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam n26673_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n26664_bdd_3_lut_4_lut (.A(sine_lookup_width_minus_modulation_deviation_amount[4]), 
         .B(n178), .C(modulation_output[15]), .D(n26664), .Z(carrier_center_increment_offset_rs_30__N_1560[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam n26664_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n26691_bdd_3_lut_4_lut (.A(sine_lookup_width_minus_modulation_deviation_amount[4]), 
         .B(n178), .C(modulation_output[15]), .D(n26691), .Z(carrier_center_increment_offset_rs_30__N_1560[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam n26691_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n24637_bdd_3_lut_4_lut (.A(sine_lookup_width_minus_modulation_deviation_amount[4]), 
         .B(n178), .C(modulation_output[15]), .D(n24637), .Z(carrier_center_increment_offset_rs_30__N_1560[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam n24637_bdd_3_lut_4_lut.init = 16'hf1e0;
    LUT4 modulation_output_15__I_0_i94_3_lut_4_lut (.A(sine_lookup_width_minus_modulation_deviation_amount[4]), 
         .B(n178), .C(modulation_output[15]), .D(n13521), .Z(n94)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam modulation_output_15__I_0_i94_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i10871_3_lut_rep_402_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[2]), 
         .B(n26786), .C(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .D(n85), .Z(n26725)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i10871_3_lut_rep_402_4_lut.init = 16'h4f40;
    LUT4 modulation_output_15__I_0_i95_3_lut_4_lut (.A(sine_lookup_width_minus_modulation_deviation_amount[4]), 
         .B(n178), .C(modulation_output[15]), .D(n13529), .Z(n95)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam modulation_output_15__I_0_i95_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i6678_2_lut_rep_419 (.A(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .B(n178_adj_3015), .Z(n26742)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i6678_2_lut_rep_419.init = 16'heeee;
    LUT4 i11846_2_lut_3_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .B(n178_adj_3015), .C(n26756), .D(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .Z(n1[7])) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i11846_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 i11845_2_lut_3_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .B(n178_adj_3015), .C(n26757), .D(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .Z(n1[6])) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i11845_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 i11836_2_lut_3_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .B(n178_adj_3015), .C(n60), .D(n26914), .Z(n1[2])) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i11836_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 i11839_2_lut_3_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .B(n178_adj_3015), .C(n59), .D(n26914), .Z(n1[3])) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i11839_2_lut_3_lut_4_lut.init = 16'h1000;
    LUT4 i11844_2_lut_3_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .B(n178_adj_3015), .C(n88), .D(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .Z(n1[5])) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i11844_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 i11852_2_lut_3_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .B(n178_adj_3015), .C(n113), .Z(n1[11])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i11852_2_lut_3_lut.init = 16'h1010;
    LUT4 i11841_2_lut_3_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .B(n178_adj_3015), .C(n89), .D(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .Z(n1[4])) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i11841_2_lut_3_lut_4_lut.init = 16'h0010;
    CCU2D add_384_15 (.A0(\addr_space[0] [13]), .B0(n14428), .C0(carrier_center_increment_offset_rs[13]), 
          .D0(carrier_center_increment_offset_ls[13]), .A1(\addr_space[0] [14]), 
          .B1(n14428), .C1(carrier_center_increment_offset_rs[14]), .D1(carrier_center_increment_offset_ls[14]), 
          .CIN(n17614), .COUT(n17615), .S0(carrier_increment_30__N_1591[13]), 
          .S1(carrier_increment_30__N_1591[14]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(92[4:87])
    defparam add_384_15.INIT0 = 16'h569a;
    defparam add_384_15.INIT1 = 16'h569a;
    defparam add_384_15.INJECT1_0 = "NO";
    defparam add_384_15.INJECT1_1 = "NO";
    LUT4 i11851_2_lut_3_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .B(n178_adj_3015), .C(n114), .Z(n1[10])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i11851_2_lut_3_lut.init = 16'h1010;
    LUT4 i11848_2_lut_3_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .B(n178_adj_3015), .C(n115), .Z(n1[9])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i11848_2_lut_3_lut.init = 16'h1010;
    LUT4 i1_2_lut_3_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[4]), 
         .B(n178_adj_3015), .C(n123), .Z(n20382)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i1_2_lut_3_lut.init = 16'h1010;
    PFUMX i19709 (.BLUT(n22144), .ALUT(n22145), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[28]));
    PFUMX i19718 (.BLUT(n22153), .ALUT(n22154), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[27]));
    LUT4 n26659_bdd_3_lut (.A(n26659), .B(n26657), .C(sine_lookup_width_minus_modulation_deviation_amount[3]), 
         .Z(n26660)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n26659_bdd_3_lut.init = 16'hcaca;
    PFUMX i19727 (.BLUT(n22162), .ALUT(n22163), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[26]));
    LUT4 n39_bdd_3_lut_25561 (.A(n13530), .B(n6), .C(sine_lookup_width_minus_modulation_deviation_amount[1]), 
         .Z(n26658)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n39_bdd_3_lut_25561.init = 16'hcaca;
    LUT4 n39_bdd_3_lut_24700 (.A(n43_adj_3008), .B(modulation_output[15]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[2]), .Z(n26657)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n39_bdd_3_lut_24700.init = 16'hcaca;
    LUT4 n36_bdd_3_lut_24703 (.A(n44), .B(modulation_output[15]), .C(sine_lookup_width_minus_modulation_deviation_amount[2]), 
         .Z(n26662)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n36_bdd_3_lut_24703.init = 16'hcaca;
    LUT4 n36_bdd_3_lut_24894 (.A(n36_adj_2992), .B(n40_adj_2993), .C(sine_lookup_width_minus_modulation_deviation_amount[2]), 
         .Z(n26663)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n36_bdd_3_lut_24894.init = 16'hcaca;
    LUT4 n37_bdd_3_lut_24897 (.A(n37_adj_3000), .B(n41_adj_3002), .C(sine_lookup_width_minus_modulation_deviation_amount[2]), 
         .Z(n26672)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n37_bdd_3_lut_24897.init = 16'hcaca;
    LUT4 n37_bdd_4_lut (.A(n14), .B(modulation_output[15]), .C(sine_lookup_width_minus_modulation_deviation_amount[2]), 
         .D(sine_lookup_width_minus_modulation_deviation_amount[1]), .Z(n26671)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;
    defparam n37_bdd_4_lut.init = 16'hccca;
    PFUMX i19736 (.BLUT(n22171), .ALUT(n22172), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[25]));
    LUT4 i22727_4_lut (.A(n20739), .B(n26947), .C(n38), .D(\wb_addr[15] ), 
         .Z(dac_clk_p_c_enable_115)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(33[3] 35[6])
    defparam i22727_4_lut.init = 16'h0400;
    LUT4 n38_bdd_3_lut_25503 (.A(n38_adj_3005), .B(n42_adj_3006), .C(sine_lookup_width_minus_modulation_deviation_amount[2]), 
         .Z(n26690)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n38_bdd_3_lut_25503.init = 16'hcaca;
    LUT4 n38_bdd_4_lut (.A(modulation_output[14]), .B(modulation_output[15]), 
         .C(sine_lookup_width_minus_modulation_deviation_amount[2]), .D(n26939), 
         .Z(n26689)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;
    defparam n38_bdd_4_lut.init = 16'hccca;
    LUT4 n38_bdd_3_lut_23485 (.A(n13522), .B(n13524), .C(sine_lookup_width_minus_modulation_deviation_amount[1]), 
         .Z(n24635)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n38_bdd_3_lut_23485.init = 16'hcaca;
    LUT4 sub_396_inv_0_i1_1_lut (.A(\addr_space[2] [0]), .Z(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[0])) /* synthesis lut_function=(!(A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(85[58:109])
    defparam sub_396_inv_0_i1_1_lut.init = 16'h5555;
    CCU2D add_384_13 (.A0(\addr_space[0] [11]), .B0(n14428), .C0(carrier_center_increment_offset_rs[11]), 
          .D0(carrier_center_increment_offset_ls[11]), .A1(\addr_space[0] [12]), 
          .B1(n14428), .C1(carrier_center_increment_offset_rs[12]), .D1(carrier_center_increment_offset_ls[12]), 
          .CIN(n17613), .COUT(n17614), .S0(carrier_increment_30__N_1591[11]), 
          .S1(carrier_increment_30__N_1591[12]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(92[4:87])
    defparam add_384_13.INIT0 = 16'h569a;
    defparam add_384_13.INIT1 = 16'h569a;
    defparam add_384_13.INJECT1_0 = "NO";
    defparam add_384_13.INJECT1_1 = "NO";
    PFUMX i19745 (.BLUT(n22180), .ALUT(n22181), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[24]));
    PFUMX i19748 (.BLUT(n22183), .ALUT(n22184), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[23]));
    LUT4 i22752_2_lut_rep_591 (.A(modulation_deviation_amount_minus_sine_lookup_width[2]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[3]), .Z(n26914)) /* synthesis lut_function=(!(A+(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam i22752_2_lut_rep_591.init = 16'h1111;
    LUT4 i6544_2_lut_rep_592 (.A(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[2]), .Z(n26915)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam i6544_2_lut_rep_592.init = 16'heeee;
    LUT4 i11884_3_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[2]), .C(modulation_deviation_amount_minus_sine_lookup_width[3]), 
         .D(n30), .Z(n123)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam i11884_3_lut_4_lut.init = 16'h0100;
    LUT4 i6553_3_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[2]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[3]), .C(n47_adj_3009), 
         .D(modulation_output[15]), .Z(n97)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam i6553_3_lut_4_lut.init = 16'hf780;
    LUT4 i6555_3_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[2]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[3]), .C(n48_adj_3010), 
         .D(modulation_output[15]), .Z(n98)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam i6555_3_lut_4_lut.init = 16'hf780;
    LUT4 i6542_2_lut_rep_593 (.A(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[2]), .Z(n26916)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam i6542_2_lut_rep_593.init = 16'h8888;
    LUT4 i6543_3_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[2]), .C(n17), 
         .D(modulation_output[15]), .Z(n73_adj_3013)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam i6543_3_lut_4_lut.init = 16'hf780;
    LUT4 i6536_2_lut_rep_594 (.A(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[1]), .Z(n26917)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam i6536_2_lut_rep_594.init = 16'h8888;
    LUT4 i6540_2_lut_rep_478_3_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[1]), .C(modulation_deviation_amount_minus_sine_lookup_width[2]), 
         .Z(n26801)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam i6540_2_lut_rep_478_3_lut.init = 16'h8080;
    PFUMX i19751 (.BLUT(n22186), .ALUT(n22187), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[22]));
    LUT4 i6537_3_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[1]), .C(modulation_output[14]), 
         .D(modulation_output[15]), .Z(n45_adj_3024)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam i6537_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_rep_418_3_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .B(modulation_output[0]), .C(modulation_deviation_amount_minus_sine_lookup_width[2]), 
         .D(modulation_deviation_amount_minus_sine_lookup_width[1]), .Z(n26741)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i1_2_lut_rep_418_3_lut_4_lut.init = 16'h0004;
    PFUMX i19754 (.BLUT(n22189), .ALUT(n22190), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[21]));
    LUT4 n24636_bdd_3_lut (.A(n24636), .B(n73), .C(sine_lookup_width_minus_modulation_deviation_amount[3]), 
         .Z(n24637)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n24636_bdd_3_lut.init = 16'hcaca;
    PFUMX i19757 (.BLUT(n22192), .ALUT(n22193), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[20]));
    PFUMX i19760 (.BLUT(n22195), .ALUT(n22196), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[19]));
    LUT4 smpl_register_5__bdd_4_lut_4_lut (.A(\wb_addr[0] ), .B(\wb_addr[1] ), 
         .C(n2), .D(\smpl_register[5] ), .Z(n26694)) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(34[4:25])
    defparam smpl_register_5__bdd_4_lut_4_lut.init = 16'hf3d1;
    LUT4 smpl_register_20__bdd_4_lut_4_lut (.A(\wb_addr[0] ), .B(\wb_addr[1] ), 
         .C(n2_adj_1), .D(\smpl_register[20] ), .Z(n26704)) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(34[4:25])
    defparam smpl_register_20__bdd_4_lut_4_lut.init = 16'hf3d1;
    LUT4 smpl_register_18__bdd_4_lut_4_lut (.A(\wb_addr[0] ), .B(\wb_addr[1] ), 
         .C(n2_adj_2), .D(\smpl_register[18] ), .Z(n26703)) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(34[4:25])
    defparam smpl_register_18__bdd_4_lut_4_lut.init = 16'hf3d1;
    LUT4 smpl_register_17__bdd_4_lut_4_lut (.A(\wb_addr[0] ), .B(\wb_addr[1] ), 
         .C(n2_adj_3), .D(\smpl_register[17] ), .Z(n26702)) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(34[4:25])
    defparam smpl_register_17__bdd_4_lut_4_lut.init = 16'hf3d1;
    LUT4 smpl_register_16__bdd_4_lut_4_lut (.A(\wb_addr[0] ), .B(\wb_addr[1] ), 
         .C(n2_adj_4), .D(\smpl_register[16] ), .Z(n26701)) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(34[4:25])
    defparam smpl_register_16__bdd_4_lut_4_lut.init = 16'hf3d1;
    CCU2D add_384_11 (.A0(\addr_space[0] [9]), .B0(n14428), .C0(carrier_center_increment_offset_rs[9]), 
          .D0(carrier_center_increment_offset_ls[9]), .A1(\addr_space[0] [10]), 
          .B1(n14428), .C1(carrier_center_increment_offset_rs[10]), .D1(carrier_center_increment_offset_ls[10]), 
          .CIN(n17612), .COUT(n17613), .S0(carrier_increment_30__N_1591[9]), 
          .S1(carrier_increment_30__N_1591[10]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(92[4:87])
    defparam add_384_11.INIT0 = 16'h569a;
    defparam add_384_11.INIT1 = 16'h569a;
    defparam add_384_11.INJECT1_0 = "NO";
    defparam add_384_11.INJECT1_1 = "NO";
    PFUMX i19763 (.BLUT(n22198), .ALUT(n22199), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[18]));
    LUT4 smpl_register_29__bdd_4_lut_4_lut (.A(\wb_addr[0] ), .B(\wb_addr[1] ), 
         .C(n2_adj_5), .D(\smpl_register[29] ), .Z(n26699)) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(34[4:25])
    defparam smpl_register_29__bdd_4_lut_4_lut.init = 16'hf3d1;
    LUT4 smpl_register_10__bdd_4_lut_4_lut (.A(\wb_addr[0] ), .B(\wb_addr[1] ), 
         .C(n2_adj_6), .D(\smpl_register[10] ), .Z(n26696)) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(34[4:25])
    defparam smpl_register_10__bdd_4_lut_4_lut.init = 16'hf3d1;
    LUT4 smpl_register_9__bdd_4_lut_4_lut (.A(\wb_addr[0] ), .B(\wb_addr[1] ), 
         .C(n2_adj_7), .D(\smpl_register[9] ), .Z(n26695)) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(34[4:25])
    defparam smpl_register_9__bdd_4_lut_4_lut.init = 16'hf3d1;
    CCU2D add_384_9 (.A0(\addr_space[0] [7]), .B0(n14428), .C0(carrier_center_increment_offset_rs[7]), 
          .D0(carrier_center_increment_offset_ls[7]), .A1(\addr_space[0] [8]), 
          .B1(n14428), .C1(carrier_center_increment_offset_rs[8]), .D1(carrier_center_increment_offset_ls[8]), 
          .CIN(n17611), .COUT(n17612), .S0(carrier_increment_30__N_1591[7]), 
          .S1(carrier_increment_30__N_1591[8]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(92[4:87])
    defparam add_384_9.INIT0 = 16'h569a;
    defparam add_384_9.INIT1 = 16'h569a;
    defparam add_384_9.INJECT1_0 = "NO";
    defparam add_384_9.INJECT1_1 = "NO";
    CCU2D add_384_7 (.A0(\addr_space[0] [5]), .B0(n14428), .C0(carrier_center_increment_offset_rs[5]), 
          .D0(carrier_center_increment_offset_ls[5]), .A1(\addr_space[0] [6]), 
          .B1(n14428), .C1(carrier_center_increment_offset_rs[6]), .D1(carrier_center_increment_offset_ls[6]), 
          .CIN(n17610), .COUT(n17611), .S0(carrier_increment_30__N_1591[5]), 
          .S1(carrier_increment_30__N_1591[6]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(92[4:87])
    defparam add_384_7.INIT0 = 16'h569a;
    defparam add_384_7.INIT1 = 16'h569a;
    defparam add_384_7.INJECT1_0 = "NO";
    defparam add_384_7.INJECT1_1 = "NO";
    CCU2D sub_113_add_2_13 (.A0(\addr_space[2] [15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\addr_space[2] [16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17673), .S0(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[15]), 
          .S1(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[16]));
    defparam sub_113_add_2_13.INIT0 = 16'h5555;
    defparam sub_113_add_2_13.INIT1 = 16'h5555;
    defparam sub_113_add_2_13.INJECT1_0 = "NO";
    defparam sub_113_add_2_13.INJECT1_1 = "NO";
    CCU2D add_384_5 (.A0(\addr_space[0] [3]), .B0(n14428), .C0(carrier_center_increment_offset_rs[3]), 
          .D0(carrier_center_increment_offset_ls[3]), .A1(\addr_space[0] [4]), 
          .B1(n14428), .C1(carrier_center_increment_offset_rs[4]), .D1(carrier_center_increment_offset_ls[4]), 
          .CIN(n17609), .COUT(n17610), .S0(carrier_increment_30__N_1591[3]), 
          .S1(carrier_increment_30__N_1591[4]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(92[4:87])
    defparam add_384_5.INIT0 = 16'h569a;
    defparam add_384_5.INIT1 = 16'h569a;
    defparam add_384_5.INJECT1_0 = "NO";
    defparam add_384_5.INJECT1_1 = "NO";
    PFUMX i19766 (.BLUT(n22201), .ALUT(n22202), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[17]));
    PFUMX i19769 (.BLUT(n22204), .ALUT(n22205), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[16]));
    PFUMX i19772 (.BLUT(n22207), .ALUT(n22208), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[15]));
    PFUMX i19775 (.BLUT(n22210), .ALUT(n22211), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[14]));
    PFUMX i19778 (.BLUT(n22213), .ALUT(n22214), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[13]));
    PFUMX i19781 (.BLUT(n22216), .ALUT(n22217), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[12]));
    CCU2D add_384_3 (.A0(\addr_space[0] [1]), .B0(n14428), .C0(carrier_center_increment_offset_rs[1]), 
          .D0(carrier_center_increment_offset_ls[1]), .A1(\addr_space[0] [2]), 
          .B1(n14428), .C1(carrier_center_increment_offset_rs[2]), .D1(carrier_center_increment_offset_ls[2]), 
          .CIN(n17608), .COUT(n17609), .S0(carrier_increment_30__N_1591[1]), 
          .S1(carrier_increment_30__N_1591[2]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(92[4:87])
    defparam add_384_3.INIT0 = 16'h569a;
    defparam add_384_3.INIT1 = 16'h569a;
    defparam add_384_3.INJECT1_0 = "NO";
    defparam add_384_3.INJECT1_1 = "NO";
    LUT4 modulation_output_15__I_0_332_i60_3_lut_4_lut (.A(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .B(modulation_output[0]), .C(modulation_deviation_amount_minus_sine_lookup_width[1]), 
         .D(n29), .Z(n60)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam modulation_output_15__I_0_332_i60_3_lut_4_lut.init = 16'h4f40;
    CCU2D sub_113_add_2_11 (.A0(\addr_space[2] [13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\addr_space[2] [14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17672), .COUT(n17673), .S0(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[13]), 
          .S1(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[14]));
    defparam sub_113_add_2_11.INIT0 = 16'h5555;
    defparam sub_113_add_2_11.INIT1 = 16'h5555;
    defparam sub_113_add_2_11.INJECT1_0 = "NO";
    defparam sub_113_add_2_11.INJECT1_1 = "NO";
    PFUMX i18923 (.BLUT(n21358), .ALUT(n21359), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[11]));
    PFUMX i18926 (.BLUT(n21361), .ALUT(n21362), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[10]));
    PFUMX i18929 (.BLUT(n21364), .ALUT(n21365), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[9]));
    LUT4 i6580_2_lut_rep_616 (.A(sine_lookup_width_minus_modulation_deviation_amount[0]), 
         .B(sine_lookup_width_minus_modulation_deviation_amount[1]), .Z(n26939)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam i6580_2_lut_rep_616.init = 16'heeee;
    LUT4 i6584_2_lut_3_lut (.A(sine_lookup_width_minus_modulation_deviation_amount[0]), 
         .B(sine_lookup_width_minus_modulation_deviation_amount[1]), .C(sine_lookup_width_minus_modulation_deviation_amount[2]), 
         .Z(n9080)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam i6584_2_lut_3_lut.init = 16'hfefe;
    LUT4 i6581_3_lut_4_lut (.A(sine_lookup_width_minus_modulation_deviation_amount[0]), 
         .B(sine_lookup_width_minus_modulation_deviation_amount[1]), .C(modulation_output[15]), 
         .D(modulation_output[14]), .Z(n46_adj_3007)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(88[41:116])
    defparam i6581_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i18932 (.BLUT(n21367), .ALUT(n21368), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[8]));
    PFUMX i18935 (.BLUT(n21370), .ALUT(n21371), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[7]));
    PFUMX i18938 (.BLUT(n21373), .ALUT(n21374), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[6]));
    CCU2D sub_113_add_2_9 (.A0(\addr_space[2] [11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\addr_space[2] [12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17671), .COUT(n17672), .S0(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[11]), 
          .S1(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[12]));
    defparam sub_113_add_2_9.INIT0 = 16'h5555;
    defparam sub_113_add_2_9.INIT1 = 16'h5555;
    defparam sub_113_add_2_9.INJECT1_0 = "NO";
    defparam sub_113_add_2_9.INJECT1_1 = "NO";
    PFUMX i18941 (.BLUT(n21376), .ALUT(n21377), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[5]));
    PFUMX modulation_output_15__I_0_332_i137 (.BLUT(n75), .ALUT(n106), .C0(n22285), 
          .Z(n137)) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;
    PFUMX modulation_output_15__I_0_332_i136 (.BLUT(n74), .ALUT(n105), .C0(n22285), 
          .Z(n136)) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;
    PFUMX i18944 (.BLUT(n21379), .ALUT(n21380), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[4]));
    PFUMX modulation_output_15__I_0_332_i133 (.BLUT(n102), .ALUT(n118), 
          .C0(modulation_deviation_amount_minus_sine_lookup_width[4]), .Z(n133)) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;
    PFUMX modulation_output_15__I_0_332_i132 (.BLUT(n101), .ALUT(n117), 
          .C0(modulation_deviation_amount_minus_sine_lookup_width[4]), .Z(n132)) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=2, LSE_LLINE=124, LSE_RLINE=135 */ ;
    PFUMX i18947 (.BLUT(n21382), .ALUT(n21383), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[3]));
    PFUMX i18950 (.BLUT(n21385), .ALUT(n21386), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[2]));
    CCU2D sub_113_add_2_7 (.A0(\addr_space[2] [9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\addr_space[2] [10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17670), .COUT(n17671), .S0(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[9]), 
          .S1(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[10]));
    defparam sub_113_add_2_7.INIT0 = 16'h5555;
    defparam sub_113_add_2_7.INIT1 = 16'h5555;
    defparam sub_113_add_2_7.INJECT1_0 = "NO";
    defparam sub_113_add_2_7.INJECT1_1 = "NO";
    PFUMX i18953 (.BLUT(n21388), .ALUT(n21389), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[1]));
    PFUMX i19682 (.BLUT(n22117), .ALUT(n22118), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[0]));
    PFUMX i19685 (.BLUT(n22120), .ALUT(n22121), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[31]));
    LUT4 i22721_4_lut (.A(n26947), .B(n20755), .C(n38), .D(\wb_addr[1] ), 
         .Z(dac_clk_p_c_enable_108)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(33[3] 35[6])
    defparam i22721_4_lut.init = 16'h0200;
    PFUMX i19691 (.BLUT(n22126), .ALUT(n22127), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[30]));
    PFUMX i19700 (.BLUT(n22135), .ALUT(n22136), .C0(\wb_addr[1] ), .Z(o_wb_data_31__N_1337[29]));
    CCU2D add_384_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\addr_space[0] [0]), .B1(n14428), .C1(carrier_center_increment_offset_rs[0]), 
          .D1(carrier_center_increment_offset_ls[0]), .COUT(n17608), .S1(carrier_increment_30__N_1591[0]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(92[4:87])
    defparam add_384_1.INIT0 = 16'hF000;
    defparam add_384_1.INIT1 = 16'h569a;
    defparam add_384_1.INJECT1_0 = "NO";
    defparam add_384_1.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_105 (.A(n20879), .B(n20881), .C(n20883), .D(n20869), 
         .Z(n178_adj_3015)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam i1_4_lut_adj_105.init = 16'hfffe;
    LUT4 i1_2_lut_adj_106 (.A(modulation_deviation_amount_minus_sine_lookup_width[14]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[5]), .Z(n20879)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam i1_2_lut_adj_106.init = 16'heeee;
    LUT4 i1_4_lut_adj_107 (.A(modulation_deviation_amount_minus_sine_lookup_width[6]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[15]), .C(modulation_deviation_amount_minus_sine_lookup_width[16]), 
         .D(modulation_deviation_amount_minus_sine_lookup_width[9]), .Z(n20881)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam i1_4_lut_adj_107.init = 16'hfffe;
    LUT4 i1_4_lut_adj_108 (.A(modulation_deviation_amount_minus_sine_lookup_width[12]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[8]), .C(modulation_deviation_amount_minus_sine_lookup_width[11]), 
         .D(modulation_deviation_amount_minus_sine_lookup_width[13]), .Z(n20883)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam i1_4_lut_adj_108.init = 16'hfffe;
    LUT4 i1_2_lut_adj_109 (.A(modulation_deviation_amount_minus_sine_lookup_width[7]), 
         .B(modulation_deviation_amount_minus_sine_lookup_width[10]), .Z(n20869)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(87[41:116])
    defparam i1_2_lut_adj_109.init = 16'heeee;
    CCU2D sub_396_add_2_17 (.A0(\addr_space[2] [15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\addr_space[2] [16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17606), .S0(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[15]), 
          .S1(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[16]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(85[58:109])
    defparam sub_396_add_2_17.INIT0 = 16'hf555;
    defparam sub_396_add_2_17.INIT1 = 16'hf555;
    defparam sub_396_add_2_17.INJECT1_0 = "NO";
    defparam sub_396_add_2_17.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_581 (.A(modulation_deviation_amount_minus_sine_lookup_width[0]), 
         .B(modulation_output[0]), .Z(n26904)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(84[11] 94[5])
    defparam i1_2_lut_rep_581.init = 16'h4444;
    LUT4 i22723_4_lut (.A(n21184), .B(n20749), .C(n20719), .D(n38), 
         .Z(dac_clk_p_c_enable_76)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(33[3] 35[6])
    defparam i22723_4_lut.init = 16'h0002;
    CCU2D sub_113_add_2_5 (.A0(\addr_space[2] [7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\addr_space[2] [8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17669), .COUT(n17670), .S0(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[7]), 
          .S1(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[8]));
    defparam sub_113_add_2_5.INIT0 = 16'h5555;
    defparam sub_113_add_2_5.INIT1 = 16'h5555;
    defparam sub_113_add_2_5.INJECT1_0 = "NO";
    defparam sub_113_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_113_add_2_3 (.A0(\addr_space[2] [5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\addr_space[2] [6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17668), .COUT(n17669), .S0(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[5]), 
          .S1(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[6]));
    defparam sub_113_add_2_3.INIT0 = 16'h5555;
    defparam sub_113_add_2_3.INIT1 = 16'h5555;
    defparam sub_113_add_2_3.INJECT1_0 = "NO";
    defparam sub_113_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_113_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(\addr_space[2] [4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n17668), .S1(modulation_deviation_amount_minus_sine_lookup_width_16__N_1639[4]));
    defparam sub_113_add_2_1.INIT0 = 16'hF000;
    defparam sub_113_add_2_1.INIT1 = 16'h5555;
    defparam sub_113_add_2_1.INJECT1_0 = "NO";
    defparam sub_113_add_2_1.INJECT1_1 = "NO";
    CCU2D sub_396_add_2_15 (.A0(\addr_space[2] [13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\addr_space[2] [14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17605), .COUT(n17606), .S0(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[13]), 
          .S1(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[14]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(85[58:109])
    defparam sub_396_add_2_15.INIT0 = 16'hf555;
    defparam sub_396_add_2_15.INIT1 = 16'hf555;
    defparam sub_396_add_2_15.INJECT1_0 = "NO";
    defparam sub_396_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_396_add_2_13 (.A0(\addr_space[2] [11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\addr_space[2] [12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17604), .COUT(n17605), .S0(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[11]), 
          .S1(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[12]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(85[58:109])
    defparam sub_396_add_2_13.INIT0 = 16'hf555;
    defparam sub_396_add_2_13.INIT1 = 16'hf555;
    defparam sub_396_add_2_13.INJECT1_0 = "NO";
    defparam sub_396_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_396_add_2_11 (.A0(\addr_space[2] [9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\addr_space[2] [10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17603), .COUT(n17604), .S0(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[9]), 
          .S1(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[10]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(85[58:109])
    defparam sub_396_add_2_11.INIT0 = 16'hf555;
    defparam sub_396_add_2_11.INIT1 = 16'hf555;
    defparam sub_396_add_2_11.INJECT1_0 = "NO";
    defparam sub_396_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_396_add_2_9 (.A0(\addr_space[2] [7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\addr_space[2] [8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17602), .COUT(n17603), .S0(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[7]), 
          .S1(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[8]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(85[58:109])
    defparam sub_396_add_2_9.INIT0 = 16'hf555;
    defparam sub_396_add_2_9.INIT1 = 16'hf555;
    defparam sub_396_add_2_9.INJECT1_0 = "NO";
    defparam sub_396_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_396_add_2_7 (.A0(\addr_space[2] [5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\addr_space[2] [6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17601), .COUT(n17602), .S0(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[5]), 
          .S1(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[6]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(85[58:109])
    defparam sub_396_add_2_7.INIT0 = 16'hf555;
    defparam sub_396_add_2_7.INIT1 = 16'hf555;
    defparam sub_396_add_2_7.INJECT1_0 = "NO";
    defparam sub_396_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_396_add_2_5 (.A0(\addr_space[2] [3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\addr_space[2] [4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17600), .COUT(n17601), .S0(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[3]), 
          .S1(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[4]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(85[58:109])
    defparam sub_396_add_2_5.INIT0 = 16'hf555;
    defparam sub_396_add_2_5.INIT1 = 16'h0aaa;
    defparam sub_396_add_2_5.INJECT1_0 = "NO";
    defparam sub_396_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_396_add_2_3 (.A0(\addr_space[2] [1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\addr_space[2] [2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17599), .COUT(n17600), .S0(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[1]), 
          .S1(sine_lookup_width_minus_modulation_deviation_amount_16__N_1622[2]));   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(85[58:109])
    defparam sub_396_add_2_3.INIT0 = 16'hf555;
    defparam sub_396_add_2_3.INIT1 = 16'hf555;
    defparam sub_396_add_2_3.INJECT1_0 = "NO";
    defparam sub_396_add_2_3.INJECT1_1 = "NO";
    dds modulation (.dac_clk_p_c(dac_clk_p_c), .i_resetb_N_301(i_resetb_N_301), 
        .\addr_space[1][0] (\addr_space[1] [0]), .\addr_space[1][30] (\addr_space[1] [30]), 
        .\addr_space[1][29] (\addr_space[1] [29]), .\addr_space[1][28] (\addr_space[1] [28]), 
        .\addr_space[1][27] (\addr_space[1] [27]), .\addr_space[1][26] (\addr_space[1] [26]), 
        .\addr_space[1][25] (\addr_space[1] [25]), .\addr_space[1][24] (\addr_space[1] [24]), 
        .\addr_space[1][23] (\addr_space[1] [23]), .\addr_space[1][22] (\addr_space[1] [22]), 
        .\addr_space[1][21] (\addr_space[1] [21]), .\addr_space[1][20] (\addr_space[1] [20]), 
        .\addr_space[1][19] (\addr_space[1] [19]), .\addr_space[1][18] (\addr_space[1] [18]), 
        .\addr_space[1][17] (\addr_space[1] [17]), .\addr_space[1][16] (\addr_space[1] [16]), 
        .\addr_space[1][15] (\addr_space[1] [15]), .\addr_space[1][14] (\addr_space[1] [14]), 
        .\addr_space[1][13] (\addr_space[1] [13]), .\addr_space[1][12] (\addr_space[1] [12]), 
        .\addr_space[1][11] (\addr_space[1] [11]), .\addr_space[1][10] (\addr_space[1] [10]), 
        .\addr_space[1][9] (\addr_space[1] [9]), .\addr_space[1][8] (\addr_space[1] [8]), 
        .\addr_space[1][7] (\addr_space[1] [7]), .\addr_space[1][6] (\addr_space[1] [6]), 
        .\addr_space[1][5] (\addr_space[1] [5]), .\addr_space[1][4] (\addr_space[1] [4]), 
        .\addr_space[1][3] (\addr_space[1] [3]), .\addr_space[1][2] (\addr_space[1] [2]), 
        .\addr_space[1][1] (\addr_space[1] [1]), .modulation_output({modulation_output}), 
        .i_resetb_c(i_resetb_c), .\quarter_wave_sample_register_q[15] (quarter_wave_sample_register_q[15]), 
        .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(72[4:161])
    dds_U2 carrier (.dac_clk_p_c(dac_clk_p_c), .i_resetb_N_301(i_resetb_N_301), 
           .carrier_increment({carrier_increment}), .i_resetb_c(i_resetb_c), 
           .o_baseband_q_c_7(o_baseband_q_c_7), .o_baseband_i_c_7(o_baseband_i_c_7), 
           .o_baseband_i_c_15(o_baseband_i_c_15), .o_baseband_i_c_14(o_baseband_i_c_14), 
           .o_baseband_i_c_13(o_baseband_i_c_13), .o_baseband_i_c_12(o_baseband_i_c_12), 
           .o_baseband_i_c_11(o_baseband_i_c_11), .o_baseband_i_c_10(o_baseband_i_c_10), 
           .n3655(n3655), .o_baseband_i_c_8(o_baseband_i_c_8), .\quarter_wave_sample_register_q[15] (quarter_wave_sample_register_q[15]), 
           .n29501(n29501), .o_baseband_q_c_15(o_baseband_q_c_15), .o_baseband_q_c_14(o_baseband_q_c_14), 
           .o_baseband_q_c_13(o_baseband_q_c_13), .o_baseband_q_c_12(o_baseband_q_c_12), 
           .o_baseband_q_c_11(o_baseband_q_c_11), .o_baseband_q_c_10(o_baseband_q_c_10), 
           .n3656(n3656), .o_baseband_q_c_8(o_baseband_q_c_8), .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(67[4:158])
    
endmodule
//
// Verilog Description of module dds
//

module dds (dac_clk_p_c, i_resetb_N_301, \addr_space[1][0] , \addr_space[1][30] , 
            \addr_space[1][29] , \addr_space[1][28] , \addr_space[1][27] , 
            \addr_space[1][26] , \addr_space[1][25] , \addr_space[1][24] , 
            \addr_space[1][23] , \addr_space[1][22] , \addr_space[1][21] , 
            \addr_space[1][20] , \addr_space[1][19] , \addr_space[1][18] , 
            \addr_space[1][17] , \addr_space[1][16] , \addr_space[1][15] , 
            \addr_space[1][14] , \addr_space[1][13] , \addr_space[1][12] , 
            \addr_space[1][11] , \addr_space[1][10] , \addr_space[1][9] , 
            \addr_space[1][8] , \addr_space[1][7] , \addr_space[1][6] , 
            \addr_space[1][5] , \addr_space[1][4] , \addr_space[1][3] , 
            \addr_space[1][2] , \addr_space[1][1] , modulation_output, 
            i_resetb_c, \quarter_wave_sample_register_q[15] , GND_net) /* synthesis syn_module_defined=1 */ ;
    input dac_clk_p_c;
    input i_resetb_N_301;
    input \addr_space[1][0] ;
    input \addr_space[1][30] ;
    input \addr_space[1][29] ;
    input \addr_space[1][28] ;
    input \addr_space[1][27] ;
    input \addr_space[1][26] ;
    input \addr_space[1][25] ;
    input \addr_space[1][24] ;
    input \addr_space[1][23] ;
    input \addr_space[1][22] ;
    input \addr_space[1][21] ;
    input \addr_space[1][20] ;
    input \addr_space[1][19] ;
    input \addr_space[1][18] ;
    input \addr_space[1][17] ;
    input \addr_space[1][16] ;
    input \addr_space[1][15] ;
    input \addr_space[1][14] ;
    input \addr_space[1][13] ;
    input \addr_space[1][12] ;
    input \addr_space[1][11] ;
    input \addr_space[1][10] ;
    input \addr_space[1][9] ;
    input \addr_space[1][8] ;
    input \addr_space[1][7] ;
    input \addr_space[1][6] ;
    input \addr_space[1][5] ;
    input \addr_space[1][4] ;
    input \addr_space[1][3] ;
    input \addr_space[1][2] ;
    input \addr_space[1][1] ;
    output [15:0]modulation_output;
    input i_resetb_c;
    input \quarter_wave_sample_register_q[15] ;
    input GND_net;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(28[49:58])
    wire [15:0]modulation_output_c /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(62[39:56])
    wire [30:0]increment;   // d:/documents/git_local/fm_modulator/rtl/dds.v(14[31:40])
    wire [11:0]o_phase;   // d:/documents/git_local/fm_modulator/rtl/dds.v(18[26:33])
    
    FD1S3DX increment_i0 (.D(\addr_space[1][0] ), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(increment[0])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i0.GSR = "DISABLED";
    FD1S3DX increment_i30 (.D(\addr_space[1][30] ), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(increment[30])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i30.GSR = "DISABLED";
    FD1S3DX increment_i29 (.D(\addr_space[1][29] ), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(increment[29])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i29.GSR = "DISABLED";
    FD1S3DX increment_i28 (.D(\addr_space[1][28] ), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(increment[28])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i28.GSR = "DISABLED";
    FD1S3DX increment_i27 (.D(\addr_space[1][27] ), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(increment[27])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i27.GSR = "DISABLED";
    FD1S3DX increment_i26 (.D(\addr_space[1][26] ), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(increment[26])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i26.GSR = "DISABLED";
    FD1S3DX increment_i25 (.D(\addr_space[1][25] ), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(increment[25])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i25.GSR = "DISABLED";
    FD1S3DX increment_i24 (.D(\addr_space[1][24] ), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(increment[24])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i24.GSR = "DISABLED";
    FD1S3DX increment_i23 (.D(\addr_space[1][23] ), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(increment[23])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i23.GSR = "DISABLED";
    FD1S3DX increment_i22 (.D(\addr_space[1][22] ), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(increment[22])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i22.GSR = "DISABLED";
    FD1S3DX increment_i21 (.D(\addr_space[1][21] ), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(increment[21])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i21.GSR = "DISABLED";
    FD1S3DX increment_i20 (.D(\addr_space[1][20] ), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(increment[20])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i20.GSR = "DISABLED";
    FD1S3DX increment_i19 (.D(\addr_space[1][19] ), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(increment[19])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i19.GSR = "DISABLED";
    FD1S3DX increment_i18 (.D(\addr_space[1][18] ), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(increment[18])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i18.GSR = "DISABLED";
    FD1S3DX increment_i17 (.D(\addr_space[1][17] ), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(increment[17])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i17.GSR = "DISABLED";
    FD1S3DX increment_i16 (.D(\addr_space[1][16] ), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(increment[16])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i16.GSR = "DISABLED";
    FD1S3DX increment_i15 (.D(\addr_space[1][15] ), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(increment[15])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i15.GSR = "DISABLED";
    FD1S3DX increment_i14 (.D(\addr_space[1][14] ), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(increment[14])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i14.GSR = "DISABLED";
    FD1S3DX increment_i13 (.D(\addr_space[1][13] ), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(increment[13])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i13.GSR = "DISABLED";
    FD1S3DX increment_i12 (.D(\addr_space[1][12] ), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(increment[12])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i12.GSR = "DISABLED";
    FD1S3DX increment_i11 (.D(\addr_space[1][11] ), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(increment[11])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i11.GSR = "DISABLED";
    FD1S3DX increment_i10 (.D(\addr_space[1][10] ), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(increment[10])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i10.GSR = "DISABLED";
    FD1S3DX increment_i9 (.D(\addr_space[1][9] ), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(increment[9])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i9.GSR = "DISABLED";
    FD1S3DX increment_i8 (.D(\addr_space[1][8] ), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(increment[8])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i8.GSR = "DISABLED";
    FD1S3DX increment_i7 (.D(\addr_space[1][7] ), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(increment[7])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i7.GSR = "DISABLED";
    FD1S3DX increment_i6 (.D(\addr_space[1][6] ), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(increment[6])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i6.GSR = "DISABLED";
    FD1S3DX increment_i5 (.D(\addr_space[1][5] ), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(increment[5])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i5.GSR = "DISABLED";
    FD1S3DX increment_i4 (.D(\addr_space[1][4] ), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(increment[4])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i4.GSR = "DISABLED";
    FD1S3DX increment_i3 (.D(\addr_space[1][3] ), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(increment[3])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i3.GSR = "DISABLED";
    FD1S3DX increment_i2 (.D(\addr_space[1][2] ), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(increment[2])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i2.GSR = "DISABLED";
    FD1S3DX increment_i1 (.D(\addr_space[1][1] ), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(increment[1])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=161, LSE_LLINE=72, LSE_RLINE=72 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i1.GSR = "DISABLED";
    quarter_wave_sine_lookup qtr_inst (.modulation_output({modulation_output}), 
            .dac_clk_p_c(dac_clk_p_c), .i_resetb_N_301(i_resetb_N_301), 
            .i_resetb_c(i_resetb_c), .o_phase({o_phase}), .\quarter_wave_sample_register_q[15] (\quarter_wave_sample_register_q[15] ), 
            .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(21[70:134])
    \nco(OW=12)  nco_inst (.dac_clk_p_c(dac_clk_p_c), .i_resetb_N_301(i_resetb_N_301), 
            .increment({increment}), .o_phase({o_phase}), .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(20[49:100])
    
endmodule
//
// Verilog Description of module quarter_wave_sine_lookup
//

module quarter_wave_sine_lookup (modulation_output, dac_clk_p_c, i_resetb_N_301, 
            i_resetb_c, o_phase, \quarter_wave_sample_register_q[15] , 
            GND_net) /* synthesis syn_module_defined=1 */ ;
    output [15:0]modulation_output;
    input dac_clk_p_c;
    input i_resetb_N_301;
    input i_resetb_c;
    input [11:0]o_phase;
    input \quarter_wave_sample_register_q[15] ;
    input GND_net;
    
    wire [15:0]modulation_output_c /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/fm_generator_wb_slave.v(62[39:56])
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(28[49:58])
    wire [15:0]\o_val_pipeline_i[0]  /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(15[24:40])
    wire [9:0]index_i;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(31[17:24])
    
    wire n21808, n157, n23248, n23249, n23250, n23395, n23396, 
        n23400;
    wire [9:0]index_i_9__N_2106;
    
    wire n23463, n23464, n23465;
    wire [1:0]phase_negation_i;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(23[12:28])
    
    wire n22590, n22591, n22594;
    wire [11:0]phase_i;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(11[17:24])
    
    wire n22592, n22593, n22595;
    wire [15:0]quarter_wave_sample_register_i;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(22[24:54])
    wire [14:0]quarter_wave_sample_register_i_15__N_2126;
    
    wire n23166, n23167, n23171, n844, n11925, n23445, n26958, 
        n27013, n21899, n27007, n27008, n27233, n27234, n62, n25360, 
        n25357, n25361, n27004, n27138, n27139, n27140, n23362, 
        n23363, n23368, n23383, n23384, n23394, n23385, n23386, 
        n23391, n23392, n23398, n22457, n22458, n22463, n22459, 
        n22460, n22464, n23039, n23040, n23047, n23041, n23042, 
        n23048, n22503, n22504, n22505, n22531, n22532, n22538, 
        n22533, n22534, n22539, n21893, n22535, n22536, n22540, 
        n382, n509, n22545, n635, n22586, n22587, n22588, n22589, 
        n21556, n21557, n21558, n23156, n23157, n23160, n23161, 
        n23168, n23162, n23163, n23169, n27224, n27225, n27226, 
        n27221, n27222, n27223, n221, n252, n23026, n27132, n27133, 
        n27134, n21796, n21797, n476, n21814, n21815, n21816, 
        n17643;
    wire [15:0]o_val_pipeline_i_0__15__N_2157;
    
    wire n29466, n27018, n21884, n21493, n17642, n25656, n21653, 
        n21654, n173, n70, n24686, n29481, n17641, n17640, n21829, 
        n21830, n21831, n844_adj_2785, n11922, n21490, n21491, n21492, 
        n21887, n747, n475, n25655, n27146, n762, n21494, n21495, 
        n23236, n23237, n23244, n25512, n316, n443, n17639, n21869, 
        n25515, n251, n17638, n26880, n24717, n23242, n23243, 
        n23247, n15054, n252_adj_2786, n26845, n62_adj_2787, n860, 
        n17792, n12012, n26723, n955, n428, n604, n364, n22876, 
        n26800, n189, n26881, n26778, n637, n26879, n22874, n9308, 
        n765, n317, n93, n21629, n94, n26838, n700, n379, n890, 
        n891, n443_adj_2788, n17637, n21499, n21500, n21501, n251_adj_2789, 
        n109, n26868, n24714, n460, n26750, n22939, n22937, n27038, 
        n29496, n25553, n22938, n21502, n21503, n21504, n316_adj_2790, 
        n325, n22877, n22878, n747_adj_2791, n21904, n22884, n22885, 
        n412, n684, n716, n890_adj_2792, n26837, n445, n699, n731, 
        n141, n26950, n22960, n85, n26972, n22959, n27126, n27127, 
        n27128, n124, n29484, n27039, n22958, n27042, n22957, 
        n17636, n29482, n924, n26951, n22953, n108, n22952, n25049, 
        n23246, n29483, n541, n27015, n526, n22951, n645, n27012, 
        n22950, n27041, n22946, n27052, n526_adj_2793, n542, n23245, 
        n635_adj_2794, n21626, n1001, n22945, n26839, n26949, n25132, 
        n491, n22943, n27149, n27151, n21892, n29499, n21865, 
        n21866, n21867, n27036, n763, n24540, n762_adj_2795, n27150, 
        n25517, n22942, n22455, n27005, n26912, n700_adj_2796, n15034, 
        n1022, n26760, n24772, n26755, n24771, n25290, n25286, 
        n25291, n26961, n27019, n17790, n17789, n19786, n173_adj_2797, 
        n189_adj_2798, n508, n620, n13928, n21644, n27010, n25750, 
        n21868, n21870, n27037, n21902, n731_adj_2799, n23350, n23351, 
        n21877, n21878, n21879, n23352, n23353, n23354, n23355, 
        n23364, n23356, n23357, n23365, n557, n572, n23436, n732, 
        n763_adj_2800, n190, n26093, n22583, n22963, n21633, n22584, 
        n26919, n475_adj_2801, n27011, n491_adj_2802, n491_adj_2803, 
        n506, n21638, n26712, n21906, n891_adj_2804, n23373, n23374, 
        n23389, n23377, n23378, n27020, n25765, n21872, n24719, 
        n21526, n23379, n23380, n93_adj_2805, n23222, n25123, n22548, 
        n589, n23437, n23387, n23388, n22542, n21827, n29479, 
        n397, n620_adj_2806, n23438, n22537, n22541, n21609, n21612, 
        n22453, n21621, n21624, n22456, n574, n21627, n21630, 
        n764, n653, n668, n23439, n26969, n21641, n21509, n475_adj_2807, 
        n653_adj_2808, n684_adj_2809, n23023, n23024, n23025, n23027, 
        n23028, n684_adj_2810, n699_adj_2811, n23440, n27194, n27195, 
        n27196, n21643, n23029, n23030, n23031, n23032, n23043, 
        n716_adj_2812, n23441, n23035, n23036, n23045, n21524, n101, 
        n188, n460_adj_2813, n285, n24688, n23050, n21863, n23442, 
        n22499, n22500, n23044, n23049, n26963, n25030, n890_adj_2814, 
        n22501, n22502, n23052, n348, n22461, n22462, n22465, 
        n26340, n23223, n781, n796, n23443, n812, n23444, n985, 
        n986, n221_adj_2815, n27050, n573, n125, n22515, n22516, 
        n22530, n22517, n22518, n285_adj_2816, n22873, n22519, n22520, 
        n22521, n22522, n22523, n22524, n460_adj_2817, n573_adj_2818, 
        n23451, n23452, n23459, n23453, n23454, n23460, n23455, 
        n23456, n23461, n557_adj_2819, n573_adj_2820, n124_adj_2821, 
        n21611, n220, n23226, n46, n23221, n875, n23446, n23457, 
        n23458, n23462, n23170, n23173, n23172, n908, n923, n23447, 
        n574_adj_2822, n21559, n939, n954, n23448, n23051, n23399, 
        n23402, n23397, n23401, n21880, n21881, n21882, n21905, 
        n21636, n21639, n22585, n971, n23449, n26824, n892, n23113, 
        n23114, n23129, n23115, n23116, n23130, n21642, n21645, 
        n1002, n1017, n23450, n21648, n21651, n892_adj_2823, n21875, 
        n21883, n21885, n21886, n21888, n270, n21581, n21894, 
        n23117, n23118, n23131, n28288, n28289, n28290, n21898, 
        n21900, n26966, n286, n318, n381, n21901, n21903, n15052, 
        n26959, n27049, n444, n24548, n24541, n24549, n747_adj_2824, 
        n251_adj_2825, n26042, n26953, n25022, n23121, n23122, n23133, 
        n668_adj_2826, n23123, n23124, n23134, n23125, n23126, n23135, 
        n23127, n23128, n23136, n22949, n22956, n22582, n763_adj_2827, 
        n21826, n491_adj_2828, n25356, n26948, n21508, n797, n828, 
        n443_adj_2829, n859, n860_adj_2830, n23144, n23145, n23146, 
        n23147, n23148, n23149, n23150, n23151, n23152, n23153, 
        n23164, n23158, n23159, n21835, n27142, n21837, n908_adj_2831, 
        n924_adj_2832, n541_adj_2833, n891_adj_2834, n653_adj_2835, 
        n669, n12026, n21823, n21824, n21825, n620_adj_2836, n635_adj_2837, 
        n636, n476_adj_2838, n397_adj_2839, n26944, n413, n27009, 
        n27053, n404, n21515, n93_adj_2840, n14831, n286_adj_2841, 
        n27017, n173_adj_2842, n732_adj_2843, n22508, n875_adj_2844, 
        n890_adj_2845, n891_adj_2846, n859_adj_2847, n860_adj_2848, 
        n27163, n588, n12038, n26954, n26964, n21832, n21514, 
        n21516, n142, n26761, n158, n46_adj_2849, n526_adj_2850, 
        n125_adj_2851, n27016, n316_adj_2852, n21403, n21404, n21405, 
        n747_adj_2853, n762_adj_2854, n763_adj_2855, n28615, n252_adj_2856, 
        n28613, n397_adj_2857, n28616, n26034, n21607, n21608, n27162, 
        n21610, n26957, n26043, n1002_adj_2858, n506_adj_2859, n15, 
        n860_adj_2860, n21805, n21806, n21807, n26045, n21802, n21803, 
        n21804, n28754, n28755, n684_adj_2861, n700_adj_2862, n781_adj_2863, 
        n668_adj_2864, n669_adj_2865, n506_adj_2866, n542_adj_2867, 
        n892_adj_2868, n26814, n26970, n844_adj_2869, n24773, n270_adj_2870, 
        n15_adj_2871, n286_adj_2872, n15_adj_2873, n61, n26945, n94_adj_2874, 
        n301, n954_adj_2875, n21517, n21518, n21519, n21895, n24774, 
        n26089, n26968, n26735, n19863, n1018, n700_adj_2876, n21619, 
        n21620, n27051, n62_adj_2877, n26802, n31, n30, n31_adj_2878, 
        n890_adj_2879, n475_adj_2880, n27169, n27168, n21520, n21521, 
        n21522, n24542, n26705, n716_adj_2881, n732_adj_2882, n22882, 
        n653_adj_2883, n669_adj_2884, n21622, n21623, n604_adj_2885, 
        n605, n413_adj_2886, n21854, n21855, n14956, n26708, n21625, 
        n412_adj_2887, n22880, n21850, n21851, n21852, n413_adj_2888, 
        n317_adj_2889, n286_adj_2890, n142_adj_2891, n14052, n158_adj_2892, 
        n158_adj_2893, n189_adj_2894, n23220, n23224, n23225, n23238, 
        n22124, n23227, n23239, n21523, n21525, n25025, n23230, 
        n23231, n23241, n731_adj_2895, n732_adj_2896, n26715, n701, 
        n26236, n23232, n23233, n23234, n23235, n21628, n25029, 
        n28618, n26240, n25032, n21631, n21632, n875_adj_2897, n379_adj_2898, 
        n891_adj_2899, n15_adj_2900, n859_adj_2901, n860_adj_2902, n22123, 
        n22125, n157_adj_2903, n26829, n636_adj_2904, n25047, n17793, 
        n17794, n29467, n25050, n507, n460_adj_2905, n476_adj_2906, 
        n25133, n397_adj_2907, n413_adj_2908, n25054, n157_adj_2909, 
        n25055, n17825, n17826, n17827, n109_adj_2910, n124_adj_2911, 
        n125_adj_2912, n653_adj_2913, n635_adj_2914, n94_adj_2915, n26765, 
        n26771, n26271, n30_adj_2916, n31_adj_2917, n14825, n21634, 
        n21635, n26272, n26277, n12039, n21637, n21640, n26971, 
        n25122, n25120, n26519, n26516, n26518, n26517, n26515, 
        n23140, n25034, n23347, n26324, n924_adj_2918, n22129, n21896, 
        n21897, n21646, n21647, n25121, n700_adj_2919, n21649, n21650, 
        n25119, n23348, n25052, n26323, n25028, n23343, n26326, 
        n731_adj_2920, n348_adj_2921, n349, n21871, n21873, n93_adj_2922, 
        n94_adj_2923, n26780, n891_adj_2924, n812_adj_2925, n13955, 
        n828_adj_2926, n26722, n797_adj_2927, n668_adj_2928, n669_adj_2929, 
        n26956, n542_adj_2930, n11191, n252_adj_2931, n25714, n23345, 
        n22875, n22881, n22883, n26942, n24775, n26878, n766, 
        n21527, n27170, n716_adj_2932, n14798, n93_adj_2933, n11109, 
        n30_adj_2934, n526_adj_2935, n15_adj_2936, n397_adj_2937, n348_adj_2938, 
        n333, n17791, n364_adj_2939, n11988, n20356, n22940, n22941, 
        n573_adj_2940, n605_adj_2941, n636_adj_2942, n700_adj_2943, 
        n732_adj_2944, n21510, n860_adj_2945, n22947, n22948, n26965, 
        n22954, n22955, n21864, n23375, n28291, n25139, n142_adj_2946, 
        n22961, n22962, n22944, n317_adj_2947, n21876, n1021, n26237, 
        n26238, n491_adj_2948, n26339, n26327, n26325, n26328, n23359, 
        n23382, n27014, n684_adj_2949, n21847, n26844, n19848, n24684, 
        n22130, n22131, n986_adj_2950, n20685, n11940, n21909, n24545, 
        n26739, n987, n21921, n11941, n24546, n254, n62_adj_2951, 
        n332, n29480, n511, n26941, n25056, n21513, n254_adj_2952, 
        n14449, n26955, n25053, n25051, n25048, n573_adj_2953, n21919, 
        n21920, n605_adj_2954, n23033, n21506, n23034, n797_adj_2955, 
        n828_adj_2956, n20563, n21907, n21908, n22547, n25033, n25031, 
        n348_adj_2957, n221_adj_2958, n11942, n796_adj_2959, n27164, 
        n908_adj_2960, n22527, n25027, n25024, n25023, n26047, n22297, 
        n348_adj_2961, n23435, n684_adj_2962, n700_adj_2963, n26920, 
        n26962, n23390, n25755, n23393, n25767, n23165, n23154, 
        n23155, n21843, n349_adj_2964, n21846, n21849, n507_adj_2965, 
        n21858, n763_adj_2966, n22526, n882, n890_adj_2967, n26033, 
        n21874, n62_adj_2968, n301_adj_2969, n23371, n23369;
    wire [15:0]n1212;
    
    wire n26092, n26090, n25285, n26091, n21842, n27152, n25287, 
        n21512, n21407, n572_adj_2970, n924_adj_2971, n21511, n21786, 
        n221_adj_2972, n252_adj_2973, n21789, n349_adj_2974, n21792, 
        n25764, n900, n25762, n21844, n22466, n26046, n26044, 
        n142_adj_2975, n572_adj_2976, n828_adj_2977, n21810, n956, 
        n20328, n26035, n26032, n26036, n173_adj_2978, n21856, n21857, 
        n28617, n28614, n26779, n638, n26729, n26031, n12155, 
        n94_adj_2979, n364_adj_2980, n14450, n22412, n716_adj_2981, 
        n812_adj_2982, n22936, n27148, n21819, n349_adj_2983, n21822, 
        n444_adj_2984, n507_adj_2985, n21828, n21848, n25751, n21845, 
        n26754, n12030, n21834, n21841, n25554, n205, n21787, 
        n348_adj_2986, n21833, n491_adj_2987, n24547, n20196, n21821, 
        n21820, n21818, n21817, n444_adj_2988, n21785, n21809, n21784, 
        n12154, n25654, n333_adj_2989, n21791, n21790, n21788, n491_adj_2990, 
        n25551, n25713, n27147, n22549, n25753, n25556, n21586, 
        n25766, n25763, n25754, n25752, n924_adj_2991, n25514, n24718, 
        n25555, n25552, n25516, n25513, n24687, n24685;
    
    FD1S3DX o_val_pipeline_i_1__i13 (.D(\o_val_pipeline_i[0] [12]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(modulation_output[12])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i13.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i12 (.D(\o_val_pipeline_i[0] [11]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(modulation_output[11])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i12.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i11 (.D(\o_val_pipeline_i[0] [10]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(modulation_output[10])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i11.GSR = "DISABLED";
    LUT4 i19371_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21808)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19371_3_lut_4_lut_4_lut.init = 16'hda5a;
    FD1S3DX o_val_pipeline_i_1__i10 (.D(\o_val_pipeline_i[0] [9]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(modulation_output[9])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i10.GSR = "DISABLED";
    LUT4 mux_198_Mux_0_i157_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n157)) /* synthesis lut_function=(A (B (C+!(D))+!B !(D))+!A (B (D)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i157_3_lut_4_lut.init = 16'hd4aa;
    FD1S3DX o_val_pipeline_i_1__i9 (.D(\o_val_pipeline_i[0] [8]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(modulation_output[8])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i9.GSR = "DISABLED";
    PFUMX i20794 (.BLUT(n23248), .ALUT(n23249), .C0(index_i[8]), .Z(n23250));
    FD1S3DX o_val_pipeline_i_1__i8 (.D(\o_val_pipeline_i[0] [7]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(modulation_output[7])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i8.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i7 (.D(\o_val_pipeline_i[0] [6]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(modulation_output[6])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i7.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i6 (.D(\o_val_pipeline_i[0] [5]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(modulation_output[5])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i6.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i5 (.D(\o_val_pipeline_i[0] [4]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(modulation_output[4])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i5.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i4 (.D(\o_val_pipeline_i[0] [3]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(modulation_output[3])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i4.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i3 (.D(\o_val_pipeline_i[0] [2]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(modulation_output[2])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i3.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i2 (.D(\o_val_pipeline_i[0] [1]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(modulation_output[1])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i2.GSR = "DISABLED";
    L6MUX21 i20944 (.D0(n23395), .D1(n23396), .SD(index_i[7]), .Z(n23400));
    FD1S3DX index_i_i9 (.D(index_i_9__N_2106[9]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(index_i[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_i_i9.GSR = "DISABLED";
    FD1S3DX index_i_i8 (.D(index_i_9__N_2106[8]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(index_i[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_i_i8.GSR = "DISABLED";
    FD1S3DX index_i_i7 (.D(index_i_9__N_2106[7]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(index_i[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_i_i7.GSR = "DISABLED";
    FD1S3DX index_i_i6 (.D(index_i_9__N_2106[6]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(index_i[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_i_i6.GSR = "DISABLED";
    PFUMX i21009 (.BLUT(n23463), .ALUT(n23464), .C0(index_i[8]), .Z(n23465));
    FD1S3DX index_i_i5 (.D(index_i_9__N_2106[5]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(index_i[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_i_i5.GSR = "DISABLED";
    FD1S3DX index_i_i4 (.D(index_i_9__N_2106[4]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(index_i[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_i_i4.GSR = "DISABLED";
    FD1S3DX index_i_i3 (.D(index_i_9__N_2106[3]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(index_i[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_i_i3.GSR = "DISABLED";
    FD1S3DX index_i_i2 (.D(index_i_9__N_2106[2]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(index_i[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_i_i2.GSR = "DISABLED";
    FD1S3DX index_i_i1 (.D(index_i_9__N_2106[1]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(index_i[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_i_i1.GSR = "DISABLED";
    FD1S3DX phase_negation_i_i1 (.D(phase_negation_i[0]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(phase_negation_i[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_negation_i_i1.GSR = "DISABLED";
    PFUMX i20138 (.BLUT(n22590), .ALUT(n22591), .C0(index_i[8]), .Z(n22594));
    FD1P3AX phase_i_i0_i0 (.D(o_phase[0]), .SP(i_resetb_c), .CK(dac_clk_p_c), 
            .Q(phase_i[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i0.GSR = "DISABLED";
    L6MUX21 i20139 (.D0(n22592), .D1(n22593), .SD(index_i[8]), .Z(n22595));
    FD1S3DX phase_negation_i_i0 (.D(phase_i[11]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(phase_negation_i[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_negation_i_i0.GSR = "DISABLED";
    FD1S3DX index_i_i0 (.D(index_i_9__N_2106[0]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(index_i[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_i_i0.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i1 (.D(\o_val_pipeline_i[0] [0]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(modulation_output[0])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i1.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i0 (.D(quarter_wave_sample_register_i_15__N_2126[0]), 
            .CK(dac_clk_p_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_i[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i0.GSR = "DISABLED";
    L6MUX21 i20715 (.D0(n23166), .D1(n23167), .SD(index_i[7]), .Z(n23171));
    PFUMX i20989 (.BLUT(n844), .ALUT(n11925), .C0(index_i[4]), .Z(n23445));
    LUT4 i19462_3_lut (.A(n26958), .B(n27013), .C(index_i[3]), .Z(n21899)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19462_3_lut.init = 16'hcaca;
    FD1P3AX phase_i_i0_i11 (.D(o_phase[11]), .SP(i_resetb_c), .CK(dac_clk_p_c), 
            .Q(phase_i[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i11.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i10 (.D(o_phase[10]), .SP(i_resetb_c), .CK(dac_clk_p_c), 
            .Q(phase_i[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i10.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i9 (.D(o_phase[9]), .SP(i_resetb_c), .CK(dac_clk_p_c), 
            .Q(phase_i[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i9.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i8 (.D(o_phase[8]), .SP(i_resetb_c), .CK(dac_clk_p_c), 
            .Q(phase_i[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i8.GSR = "DISABLED";
    LUT4 mux_198_Mux_0_i363_3_lut_4_lut_3_lut_rep_684 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27007)) /* synthesis lut_function=(A (B+!(C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i363_3_lut_4_lut_3_lut_rep_684.init = 16'hdbdb;
    FD1P3AX phase_i_i0_i7 (.D(o_phase[7]), .SP(i_resetb_c), .CK(dac_clk_p_c), 
            .Q(phase_i[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i7.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i6 (.D(o_phase[6]), .SP(i_resetb_c), .CK(dac_clk_p_c), 
            .Q(phase_i[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i6.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i5 (.D(o_phase[5]), .SP(i_resetb_c), .CK(dac_clk_p_c), 
            .Q(phase_i[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i5.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i4 (.D(o_phase[4]), .SP(i_resetb_c), .CK(dac_clk_p_c), 
            .Q(phase_i[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i4.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i3 (.D(o_phase[3]), .SP(i_resetb_c), .CK(dac_clk_p_c), 
            .Q(phase_i[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i3.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i2 (.D(o_phase[2]), .SP(i_resetb_c), .CK(dac_clk_p_c), 
            .Q(phase_i[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i2.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i1 (.D(o_phase[1]), .SP(i_resetb_c), .CK(dac_clk_p_c), 
            .Q(phase_i[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i1.GSR = "DISABLED";
    LUT4 mux_198_Mux_6_i7_3_lut_4_lut_3_lut_rep_685 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27008)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_6_i7_3_lut_4_lut_3_lut_rep_685.init = 16'hd6d6;
    PFUMX i24801 (.BLUT(n27233), .ALUT(n27234), .C0(index_i[3]), .Z(n62));
    PFUMX i23597 (.BLUT(n25360), .ALUT(n25357), .C0(index_i[6]), .Z(n25361));
    LUT4 i11084_2_lut_rep_681 (.A(index_i[0]), .B(index_i[1]), .Z(n27004)) /* synthesis lut_function=((B)+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11084_2_lut_rep_681.init = 16'hdddd;
    PFUMX i24740 (.BLUT(n27138), .ALUT(n27139), .C0(index_i[1]), .Z(n27140));
    L6MUX21 i20912 (.D0(n23362), .D1(n23363), .SD(index_i[7]), .Z(n23368));
    L6MUX21 i20938 (.D0(n23383), .D1(n23384), .SD(index_i[6]), .Z(n23394));
    L6MUX21 i20939 (.D0(n23385), .D1(n23386), .SD(index_i[6]), .Z(n23395));
    L6MUX21 i20942 (.D0(n23391), .D1(n23392), .SD(index_i[7]), .Z(n23398));
    L6MUX21 i20007 (.D0(n22457), .D1(n22458), .SD(index_i[7]), .Z(n22463));
    PFUMX i20008 (.BLUT(n22459), .ALUT(n22460), .C0(index_i[7]), .Z(n22464));
    L6MUX21 i20591 (.D0(n23039), .D1(n23040), .SD(index_i[7]), .Z(n23047));
    L6MUX21 i20592 (.D0(n23041), .D1(n23042), .SD(index_i[7]), .Z(n23048));
    L6MUX21 i20049 (.D0(n22503), .D1(n22504), .SD(index_i[7]), .Z(n22505));
    L6MUX21 i20082 (.D0(n22531), .D1(n22532), .SD(index_i[7]), .Z(n22538));
    L6MUX21 i20083 (.D0(n22533), .D1(n22534), .SD(index_i[7]), .Z(n22539));
    LUT4 i19456_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21893)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C))+!A !(B (C)+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19456_3_lut_4_lut_4_lut.init = 16'h5ad3;
    PFUMX i20084 (.BLUT(n22535), .ALUT(n22536), .C0(index_i[7]), .Z(n22540));
    L6MUX21 i20089 (.D0(n382), .D1(n509), .SD(index_i[7]), .Z(n22545));
    LUT4 mux_198_Mux_0_i635_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n635)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i635_3_lut_4_lut_4_lut.init = 16'hfd0a;
    L6MUX21 i20136 (.D0(n22586), .D1(n22587), .SD(index_i[7]), .Z(n22592));
    L6MUX21 i20137 (.D0(n22588), .D1(n22589), .SD(index_i[7]), .Z(n22593));
    L6MUX21 i19121 (.D0(n21556), .D1(n21557), .SD(index_i[7]), .Z(n21558));
    L6MUX21 i20710 (.D0(n23156), .D1(n23157), .SD(index_i[6]), .Z(n23166));
    L6MUX21 i20712 (.D0(n23160), .D1(n23161), .SD(index_i[7]), .Z(n23168));
    L6MUX21 i20713 (.D0(n23162), .D1(n23163), .SD(index_i[7]), .Z(n23169));
    PFUMX i24795 (.BLUT(n27224), .ALUT(n27225), .C0(index_i[1]), .Z(n27226));
    PFUMX i24793 (.BLUT(n27221), .ALUT(n27222), .C0(index_i[3]), .Z(n27223));
    PFUMX i20570 (.BLUT(n221), .ALUT(n252), .C0(index_i[5]), .Z(n23026));
    PFUMX i24736 (.BLUT(n27132), .ALUT(n27133), .C0(index_i[1]), .Z(n27134));
    PFUMX i19361 (.BLUT(n21796), .ALUT(n21797), .C0(index_i[4]), .Z(n476));
    PFUMX i19379 (.BLUT(n21814), .ALUT(n21815), .C0(index_i[4]), .Z(n21816));
    CCU2D unary_minus_10_add_3_17 (.A0(\quarter_wave_sample_register_q[15] ), 
          .B0(GND_net), .C0(GND_net), .D0(GND_net), .A1(GND_net), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n17643), .S0(o_val_pipeline_i_0__15__N_2157[15]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam unary_minus_10_add_3_17.INIT0 = 16'hf555;
    defparam unary_minus_10_add_3_17.INIT1 = 16'h0000;
    defparam unary_minus_10_add_3_17.INJECT1_0 = "NO";
    defparam unary_minus_10_add_3_17.INJECT1_1 = "NO";
    LUT4 i19447_3_lut (.A(n29466), .B(n27018), .C(index_i[3]), .Z(n21884)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19447_3_lut.init = 16'hcaca;
    LUT4 i19056_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n21493)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (D))+!A !(D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19056_3_lut_4_lut_4_lut_4_lut.init = 16'ha25d;
    CCU2D unary_minus_10_add_3_15 (.A0(quarter_wave_sample_register_i[13]), 
          .B0(GND_net), .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[14]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17642), .COUT(n17643), 
          .S0(o_val_pipeline_i_0__15__N_2157[13]), .S1(o_val_pipeline_i_0__15__N_2157[14]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam unary_minus_10_add_3_15.INIT0 = 16'hf555;
    defparam unary_minus_10_add_3_15.INIT1 = 16'hf555;
    defparam unary_minus_10_add_3_15.INJECT1_0 = "NO";
    defparam unary_minus_10_add_3_15.INJECT1_1 = "NO";
    LUT4 i22128_3_lut (.A(n25656), .B(n21653), .C(index_i[5]), .Z(n21654)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22128_3_lut.init = 16'hcaca;
    LUT4 n173_bdd_4_lut (.A(n173), .B(n70), .C(index_i[4]), .D(index_i[3]), 
         .Z(n24686)) /* synthesis lut_function=(A (B+(C+!(D)))+!A !((C+!(D))+!B)) */ ;
    defparam n173_bdd_4_lut.init = 16'hacaa;
    LUT4 mux_198_Mux_0_i123_3_lut_3_lut_rep_808 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29481)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i123_3_lut_3_lut_rep_808.init = 16'h6c6c;
    CCU2D unary_minus_10_add_3_13 (.A0(quarter_wave_sample_register_i[11]), 
          .B0(GND_net), .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[12]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17641), .COUT(n17642), 
          .S0(o_val_pipeline_i_0__15__N_2157[11]), .S1(o_val_pipeline_i_0__15__N_2157[12]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam unary_minus_10_add_3_13.INIT0 = 16'hf555;
    defparam unary_minus_10_add_3_13.INIT1 = 16'hf555;
    defparam unary_minus_10_add_3_13.INJECT1_0 = "NO";
    defparam unary_minus_10_add_3_13.INJECT1_1 = "NO";
    CCU2D unary_minus_10_add_3_11 (.A0(quarter_wave_sample_register_i[9]), 
          .B0(GND_net), .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[10]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17640), .COUT(n17641), 
          .S0(o_val_pipeline_i_0__15__N_2157[9]), .S1(o_val_pipeline_i_0__15__N_2157[10]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam unary_minus_10_add_3_11.INIT0 = 16'hf555;
    defparam unary_minus_10_add_3_11.INIT1 = 16'hf555;
    defparam unary_minus_10_add_3_11.INJECT1_0 = "NO";
    defparam unary_minus_10_add_3_11.INJECT1_1 = "NO";
    PFUMX i19394 (.BLUT(n21829), .ALUT(n21830), .C0(index_i[4]), .Z(n21831));
    LUT4 i9472_3_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[3]), .C(index_i[0]), 
         .D(index_i[1]), .Z(n844_adj_2785)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9472_3_lut_4_lut_4_lut.init = 16'hf00e;
    LUT4 i9361_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n11922)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))+!A !(B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9361_3_lut_4_lut_4_lut.init = 16'hb5b3;
    LUT4 mux_198_Mux_5_i252_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[4]), .Z(n252)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+(D)))+!A (B (C (D))+!B !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_5_i252_3_lut_4_lut.init = 16'hc993;
    PFUMX i19055 (.BLUT(n21490), .ALUT(n21491), .C0(index_i[4]), .Z(n21492));
    LUT4 i19450_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n21887)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B (C+!(D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19450_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h1c18;
    LUT4 mux_198_Mux_7_i747_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), 
         .B(index_i[2]), .C(index_i[3]), .D(index_i[0]), .Z(n747)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))+!A (B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_7_i747_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'he1e3;
    LUT4 mux_198_Mux_5_i475_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n475)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_5_i475_3_lut_4_lut_4_lut.init = 16'hd4a5;
    LUT4 n172_bdd_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n25655)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n172_bdd_3_lut_4_lut_4_lut_4_lut.init = 16'h1e1c;
    LUT4 n17999_bdd_4_lut_else_4_lut (.A(index_i[3]), .B(index_i[4]), .C(index_i[1]), 
         .D(index_i[2]), .Z(n27146)) /* synthesis lut_function=(!(A (B (D)+!B ((D)+!C))+!A !(B+!((D)+!C)))) */ ;
    defparam n17999_bdd_4_lut_else_4_lut.init = 16'h44fc;
    LUT4 mux_198_Mux_7_i762_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), 
         .B(index_i[2]), .C(index_i[3]), .D(index_i[0]), .Z(n762)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B ((D)+!C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_7_i762_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h3878;
    PFUMX i19058 (.BLUT(n21493), .ALUT(n21494), .C0(index_i[4]), .Z(n21495));
    L6MUX21 i20788 (.D0(n23236), .D1(n23237), .SD(index_i[6]), .Z(n23244));
    LUT4 n301_bdd_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n25512)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A !((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n301_bdd_3_lut_4_lut_4_lut_4_lut.init = 16'h7173;
    LUT4 mux_198_Mux_9_i316_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), 
         .B(index_i[2]), .C(index_i[3]), .D(index_i[0]), .Z(n316)) /* synthesis lut_function=(!(A (B (C)+!B !(C+(D)))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_9_i316_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h7e7c;
    LUT4 mux_198_Mux_0_i443_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .D(index_i[3]), .Z(n443)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C (D))+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i443_3_lut_4_lut_4_lut_4_lut.init = 16'h0ed5;
    CCU2D unary_minus_10_add_3_9 (.A0(quarter_wave_sample_register_i[7]), 
          .B0(GND_net), .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[8]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17639), .COUT(n17640), 
          .S0(o_val_pipeline_i_0__15__N_2157[7]), .S1(o_val_pipeline_i_0__15__N_2157[8]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam unary_minus_10_add_3_9.INIT0 = 16'hf555;
    defparam unary_minus_10_add_3_9.INIT1 = 16'hf555;
    defparam unary_minus_10_add_3_9.INJECT1_0 = "NO";
    defparam unary_minus_10_add_3_9.INJECT1_1 = "NO";
    LUT4 i19432_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n21869)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B (C+(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19432_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h7c78;
    LUT4 n22_bdd_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n25515)) /* synthesis lut_function=(A (B (C)+!B ((D)+!C))+!A (B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n22_bdd_3_lut_4_lut_4_lut_4_lut.init = 16'he7c7;
    LUT4 mux_198_Mux_0_i251_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n251)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A !(B ((D)+!C)+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i251_3_lut_4_lut_4_lut_4_lut.init = 16'h543c;
    CCU2D unary_minus_10_add_3_7 (.A0(quarter_wave_sample_register_i[5]), 
          .B0(GND_net), .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[6]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17638), .COUT(n17639), 
          .S0(o_val_pipeline_i_0__15__N_2157[5]), .S1(o_val_pipeline_i_0__15__N_2157[6]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam unary_minus_10_add_3_7.INIT0 = 16'hf555;
    defparam unary_minus_10_add_3_7.INIT1 = 16'hf555;
    defparam unary_minus_10_add_3_7.INJECT1_0 = "NO";
    defparam unary_minus_10_add_3_7.INJECT1_1 = "NO";
    LUT4 index_i_4__bdd_3_lut_23019_4_lut (.A(n26880), .B(index_i[3]), .C(index_i[5]), 
         .D(index_i[4]), .Z(n24717)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam index_i_4__bdd_3_lut_23019_4_lut.init = 16'hf080;
    L6MUX21 i20791 (.D0(n23242), .D1(n23243), .SD(index_i[6]), .Z(n23247));
    LUT4 mux_198_Mux_3_i252_3_lut_4_lut (.A(n26880), .B(index_i[3]), .C(index_i[4]), 
         .D(n15054), .Z(n252_adj_2786)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_3_i252_3_lut_4_lut.init = 16'h08f8;
    LUT4 mux_198_Mux_10_i62_3_lut_3_lut_4_lut (.A(n26880), .B(index_i[3]), 
         .C(n26845), .D(index_i[4]), .Z(n62_adj_2787)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_10_i62_3_lut_3_lut_4_lut.init = 16'hf077;
    LUT4 mux_198_Mux_8_i860_3_lut_4_lut (.A(n26880), .B(index_i[3]), .C(index_i[4]), 
         .D(n26845), .Z(n860)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_8_i860_3_lut_4_lut.init = 16'h08f8;
    LUT4 i15528_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[1]), .Z(n17792)) /* synthesis lut_function=(A (B (C (D))+!B !(C))+!A (B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i15528_3_lut_4_lut_4_lut_4_lut.init = 16'hd656;
    LUT4 i9451_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n12012)) /* synthesis lut_function=(!(A (B (C)+!B ((D)+!C))+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9451_3_lut_4_lut_4_lut.init = 16'h4969;
    LUT4 mux_198_Mux_6_i955_3_lut_4_lut (.A(n26880), .B(index_i[3]), .C(index_i[4]), 
         .D(n26723), .Z(n955)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_6_i955_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_198_Mux_0_i428_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[2]), 
         .B(index_i[0]), .C(index_i[1]), .D(index_i[3]), .Z(n428)) /* synthesis lut_function=(A (B (C+!(D))+!B !((D)+!C))+!A (B (D)+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i428_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hd5a9;
    LUT4 mux_198_Mux_0_i604_3_lut_4_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[1]), .D(index_i[3]), .Z(n604)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A !(B (D)+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i604_3_lut_4_lut_4_lut_4_lut.init = 16'h5439;
    LUT4 i20420_3_lut_4_lut (.A(n26880), .B(index_i[3]), .C(index_i[4]), 
         .D(n364), .Z(n22876)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20420_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_198_Mux_3_i189_3_lut_3_lut_4_lut (.A(n26880), .B(index_i[3]), 
         .C(index_i[4]), .D(n26800), .Z(n189)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_3_i189_3_lut_3_lut_4_lut.init = 16'h08f8;
    LUT4 mux_198_Mux_10_i637_3_lut_4_lut_4_lut (.A(n26881), .B(index_i[4]), 
         .C(index_i[5]), .D(n26778), .Z(n637)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_10_i637_3_lut_4_lut_4_lut.init = 16'h1f1c;
    LUT4 i20418_3_lut_3_lut_4_lut (.A(n26879), .B(index_i[3]), .C(n316), 
         .D(index_i[4]), .Z(n22874)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20418_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 i11177_3_lut_4_lut (.A(n26879), .B(index_i[3]), .C(n9308), .D(index_i[6]), 
         .Z(n765)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11177_3_lut_4_lut.init = 16'hffe0;
    LUT4 mux_198_Mux_10_i317_3_lut_3_lut_4_lut (.A(n26879), .B(index_i[3]), 
         .C(n26800), .D(index_i[4]), .Z(n317)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_10_i317_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 i19192_3_lut_3_lut_4_lut (.A(n26879), .B(index_i[3]), .C(n93), 
         .D(index_i[4]), .Z(n21629)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19192_3_lut_3_lut_4_lut.init = 16'h11f0;
    LUT4 mux_198_Mux_9_i94_3_lut_4_lut (.A(n26879), .B(index_i[3]), .C(index_i[4]), 
         .D(n93), .Z(n94)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_9_i94_3_lut_4_lut.init = 16'hfe0e;
    LUT4 mux_198_Mux_9_i700_3_lut_4_lut (.A(n26879), .B(index_i[3]), .C(index_i[4]), 
         .D(n26838), .Z(n700)) /* synthesis lut_function=(!(A (C+!(D))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_9_i700_3_lut_4_lut.init = 16'h1f10;
    LUT4 mux_198_Mux_0_i379_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n379)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !((D)+!C))+!A !(B ((D)+!C)+!B (D))) */ ;
    defparam mux_198_Mux_0_i379_3_lut_4_lut_4_lut.init = 16'h8079;
    LUT4 mux_198_Mux_7_i891_3_lut_4_lut (.A(n26879), .B(index_i[3]), .C(index_i[4]), 
         .D(n890), .Z(n891)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_7_i891_3_lut_4_lut.init = 16'hfe0e;
    LUT4 mux_198_Mux_8_i443_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n443_adj_2788)) /* synthesis lut_function=(A (B (C+!(D))+!B !((D)+!C))+!A !(B (D)+!B ((D)+!C))) */ ;
    defparam mux_198_Mux_8_i443_3_lut_4_lut_4_lut.init = 16'h80fc;
    CCU2D unary_minus_10_add_3_5 (.A0(quarter_wave_sample_register_i[3]), 
          .B0(GND_net), .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[4]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17637), .COUT(n17638), 
          .S0(o_val_pipeline_i_0__15__N_2157[3]), .S1(o_val_pipeline_i_0__15__N_2157[4]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam unary_minus_10_add_3_5.INIT0 = 16'hf555;
    defparam unary_minus_10_add_3_5.INIT1 = 16'hf555;
    defparam unary_minus_10_add_3_5.INJECT1_0 = "NO";
    defparam unary_minus_10_add_3_5.INJECT1_1 = "NO";
    PFUMX i19064 (.BLUT(n21499), .ALUT(n21500), .C0(index_i[4]), .Z(n21501));
    LUT4 mux_198_Mux_8_i251_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[2]), .D(index_i[3]), .Z(n251_adj_2789)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_8_i251_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h07e0;
    LUT4 mux_198_Mux_8_i109_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n109)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C+!(D)))+!A (B (C (D)+!C !(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_8_i109_3_lut_4_lut_4_lut.init = 16'hf83e;
    LUT4 index_i_4__bdd_4_lut_23184 (.A(index_i[4]), .B(n26868), .C(index_i[7]), 
         .D(n26838), .Z(n24714)) /* synthesis lut_function=(A (C+!(D))+!A (B+!(C))) */ ;
    defparam index_i_4__bdd_4_lut_23184.init = 16'he5ef;
    LUT4 mux_198_Mux_0_i460_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n460)) /* synthesis lut_function=(A (B+(C (D)+!C !(D)))+!A (B (C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i460_3_lut_4_lut_4_lut.init = 16'hf8cb;
    LUT4 mux_198_Mux_8_i61_3_lut_rep_427_4_lut_4_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[2]), .D(index_i[3]), .Z(n26750)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A (B (C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_8_i61_3_lut_rep_427_4_lut_4_lut_4_lut.init = 16'he0f8;
    LUT4 i20483_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n22939)) /* synthesis lut_function=(A (B (C+!(D))+!B !((D)+!C))+!A !(B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20483_3_lut_4_lut_4_lut.init = 16'h81f8;
    LUT4 i20481_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n22937)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20481_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hf81f;
    LUT4 n262_bdd_3_lut_23759 (.A(n27038), .B(n29496), .C(index_i[3]), 
         .Z(n25553)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n262_bdd_3_lut_23759.init = 16'hcaca;
    LUT4 i20482_3_lut_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n22938)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C+!(D))+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20482_3_lut_3_lut_4_lut_4_lut.init = 16'h1f81;
    LUT4 i19378_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n21815)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C))+!A (B (C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19378_3_lut_4_lut_4_lut_4_lut.init = 16'he078;
    PFUMX i19067 (.BLUT(n21502), .ALUT(n21503), .C0(index_i[4]), .Z(n21504));
    LUT4 mux_198_Mux_0_i316_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n316_adj_2790)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+(D)))+!A (B (C+(D))+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i316_3_lut_4_lut_4_lut_4_lut.init = 16'h332d;
    LUT4 mux_198_Mux_6_i325_3_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n325)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_6_i325_3_lut_4_lut_3_lut.init = 16'h6d6d;
    L6MUX21 i20423 (.D0(n22877), .D1(n22878), .SD(index_i[6]), .Z(n382));
    LUT4 mux_198_Mux_0_i747_3_lut_3_lut_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n747_adj_2791)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (D))+!A (B (D)+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i747_3_lut_3_lut_3_lut_4_lut.init = 16'h09f6;
    LUT4 i19467_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n21904)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B+(C+(D))))) */ ;
    defparam i19467_3_lut_4_lut_4_lut_4_lut.init = 16'h2aab;
    L6MUX21 i20430 (.D0(n22884), .D1(n22885), .SD(index_i[6]), .Z(n509));
    LUT4 mux_198_Mux_0_i412_3_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[1]), .D(index_i[3]), .Z(n412)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C (D)))+!A (B (C+!(D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i412_3_lut_4_lut_4_lut.init = 16'hf14c;
    LUT4 i19057_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21494)) /* synthesis lut_function=(A (C)+!A !(B (C)+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19057_3_lut_4_lut_4_lut.init = 16'hb4b5;
    LUT4 mux_198_Mux_1_i684_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n684)) /* synthesis lut_function=(A (B ((D)+!C)+!B !((D)+!C))+!A !(B (C+(D))+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_1_i684_3_lut_4_lut_4_lut.init = 16'h992d;
    LUT4 mux_198_Mux_1_i716_3_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[1]), .D(index_i[3]), .Z(n716)) /* synthesis lut_function=(!(A (B (D)+!B !(C))+!A !(B (C (D))+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_1_i716_3_lut_4_lut_4_lut.init = 16'h70a9;
    LUT4 mux_198_Mux_0_i890_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n890_adj_2792)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)+!C !(D)))+!A !(B (C)+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i890_3_lut_4_lut_4_lut.init = 16'h70ca;
    LUT4 mux_198_Mux_11_i445_3_lut_4_lut_4_lut_4_lut (.A(index_i[3]), .B(index_i[4]), 
         .C(index_i[5]), .D(n26837), .Z(n445)) /* synthesis lut_function=(!(A (B (C))+!A !(B+(C+(D))))) */ ;
    defparam mux_198_Mux_11_i445_3_lut_4_lut_4_lut_4_lut.init = 16'h7f7e;
    LUT4 mux_198_Mux_7_i699_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n699)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C+!(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_7_i699_3_lut_4_lut_4_lut.init = 16'hf07e;
    LUT4 mux_198_Mux_2_i731_3_lut_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n731)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(B (C)+!B !(C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_2_i731_3_lut_3_lut_4_lut.init = 16'h69f0;
    LUT4 i20504_3_lut (.A(n141), .B(n26950), .C(index_i[3]), .Z(n22960)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20504_3_lut.init = 16'hcaca;
    LUT4 i20503_3_lut (.A(n85), .B(n26972), .C(index_i[3]), .Z(n22959)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20503_3_lut.init = 16'hcaca;
    PFUMX i24732 (.BLUT(n27126), .ALUT(n27127), .C0(index_i[0]), .Z(n27128));
    LUT4 mux_198_Mux_0_i124_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n124)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A !(B (D)+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i124_3_lut_4_lut_4_lut.init = 16'h6c99;
    LUT4 i20502_3_lut (.A(n29484), .B(n27039), .C(index_i[3]), .Z(n22958)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20502_3_lut.init = 16'hcaca;
    LUT4 i20501_3_lut (.A(n26950), .B(n27042), .C(index_i[3]), .Z(n22957)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20501_3_lut.init = 16'hcaca;
    CCU2D unary_minus_10_add_3_3 (.A0(quarter_wave_sample_register_i[1]), 
          .B0(GND_net), .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[2]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17636), .COUT(n17637), 
          .S0(o_val_pipeline_i_0__15__N_2157[1]), .S1(o_val_pipeline_i_0__15__N_2157[2]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam unary_minus_10_add_3_3.INIT0 = 16'hf555;
    defparam unary_minus_10_add_3_3.INIT1 = 16'hf555;
    defparam unary_minus_10_add_3_3.INJECT1_0 = "NO";
    defparam unary_minus_10_add_3_3.INJECT1_1 = "NO";
    LUT4 mux_198_Mux_0_i963_3_lut_3_lut_3_lut_rep_809 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29482)) /* synthesis lut_function=(!(A (B)+!A (B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i963_3_lut_3_lut_3_lut_rep_809.init = 16'h3636;
    LUT4 mux_198_Mux_6_i924_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[4]), .D(n762), .Z(n924)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_6_i924_3_lut_4_lut.init = 16'h6f60;
    LUT4 i20497_3_lut (.A(n26951), .B(n27042), .C(index_i[3]), .Z(n22953)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20497_3_lut.init = 16'hcaca;
    LUT4 i20496_3_lut (.A(n29484), .B(n108), .C(index_i[3]), .Z(n22952)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20496_3_lut.init = 16'hcaca;
    LUT4 n308_bdd_3_lut_23313_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n25049)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A !(B (C+(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n308_bdd_3_lut_23313_4_lut_4_lut.init = 16'h9936;
    LUT4 i20793_3_lut (.A(n23246), .B(n23247), .C(index_i[7]), .Z(n23249)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20793_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_6_i22_rep_810 (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .Z(n29483)) /* synthesis lut_function=(!(A (C)+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_6_i22_rep_810.init = 16'h4a4a;
    LUT4 i12084_2_lut (.A(index_i[1]), .B(index_i[3]), .Z(n541)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i12084_2_lut.init = 16'h1111;
    LUT4 mux_198_Mux_0_i526_3_lut (.A(n27015), .B(n26958), .C(index_i[3]), 
         .Z(n526)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i526_3_lut.init = 16'hcaca;
    LUT4 i20495_3_lut (.A(n85), .B(n27039), .C(index_i[3]), .Z(n22951)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20495_3_lut.init = 16'hcaca;
    LUT4 i20494_3_lut (.A(n645), .B(n27012), .C(index_i[3]), .Z(n22950)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20494_3_lut.init = 16'hcaca;
    LUT4 i20490_3_lut (.A(n27042), .B(n27041), .C(index_i[3]), .Z(n22946)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20490_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_8_i542_3_lut_4_lut (.A(n27052), .B(index_i[3]), .C(index_i[4]), 
         .D(n526_adj_2793), .Z(n542)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_8_i542_3_lut_4_lut.init = 16'h6f60;
    LUT4 i20792_3_lut (.A(n23244), .B(n23245), .C(index_i[7]), .Z(n23248)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20792_3_lut.init = 16'hcaca;
    LUT4 i19189_3_lut_4_lut (.A(n27052), .B(index_i[3]), .C(index_i[4]), 
         .D(n635_adj_2794), .Z(n21626)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19189_3_lut_4_lut.init = 16'hf606;
    LUT4 i20489_3_lut (.A(n1001), .B(n26951), .C(index_i[3]), .Z(n22945)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20489_3_lut.init = 16'hcaca;
    LUT4 index_i_6__bdd_4_lut_4_lut (.A(n26839), .B(index_i[5]), .C(n26949), 
         .D(index_i[6]), .Z(n25132)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C))+!A !(B (C+(D))+!B (C)))) */ ;
    defparam index_i_6__bdd_4_lut_4_lut.init = 16'h74f0;
    LUT4 mux_198_Mux_5_i491_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n491)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A !(B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_5_i491_3_lut_4_lut_4_lut.init = 16'ha54a;
    LUT4 i20487_3_lut (.A(n27041), .B(n645), .C(index_i[3]), .Z(n22943)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20487_3_lut.init = 16'hcaca;
    LUT4 index_i_1__bdd_4_lut_24960 (.A(index_i[1]), .B(index_i[0]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n27149)) /* synthesis lut_function=(!(A (B (D)+!B (C+!(D)))+!A !(B (C (D)+!C !(D))+!B !((D)+!C)))) */ ;
    defparam index_i_1__bdd_4_lut_24960.init = 16'h429c;
    LUT4 i23525_then_3_lut (.A(index_i[0]), .B(index_i[4]), .C(index_i[3]), 
         .Z(n27151)) /* synthesis lut_function=(A (B)+!A (B (C)+!B !(C))) */ ;
    defparam i23525_then_3_lut.init = 16'hc9c9;
    LUT4 i11284_3_lut_3_lut_3_lut_rep_811 (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .Z(n29484)) /* synthesis lut_function=(!(A+!(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11284_3_lut_3_lut_3_lut_rep_811.init = 16'h4545;
    LUT4 i19455_3_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[0]), 
         .D(index_i[3]), .Z(n21892)) /* synthesis lut_function=(!(A ((D)+!B)+!A !(B (D)+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19455_3_lut_4_lut_4_lut.init = 16'h4588;
    LUT4 index_i_0__bdd_4_lut (.A(index_i[0]), .B(index_i[3]), .C(index_i[1]), 
         .D(index_i[2]), .Z(n29499)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C (D)))+!A !(B (C+!(D))+!B !(C+(D))))) */ ;
    defparam index_i_0__bdd_4_lut.init = 16'h4ae7;
    PFUMX i19430 (.BLUT(n21865), .ALUT(n21866), .C0(index_i[4]), .Z(n21867));
    LUT4 n21586_bdd_4_lut_24303 (.A(n27036), .B(n763), .C(index_i[5]), 
         .D(index_i[4]), .Z(n24540)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam n21586_bdd_4_lut_24303.init = 16'hcfca;
    LUT4 mux_198_Mux_0_i762_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n762_adj_2795)) /* synthesis lut_function=(A (B+!((D)+!C))+!A !(B (D)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i762_3_lut_4_lut_4_lut.init = 16'h98fc;
    CCU2D unary_minus_10_add_3_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(quarter_wave_sample_register_i[0]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .COUT(n17636), .S1(o_val_pipeline_i_0__15__N_2157[0]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam unary_minus_10_add_3_1.INIT0 = 16'hF000;
    defparam unary_minus_10_add_3_1.INIT1 = 16'h0aaa;
    defparam unary_minus_10_add_3_1.INJECT1_0 = "NO";
    defparam unary_minus_10_add_3_1.INJECT1_1 = "NO";
    LUT4 i23525_else_3_lut (.A(index_i[0]), .B(index_i[2]), .C(index_i[4]), 
         .D(index_i[3]), .Z(n27150)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C (D)+!C !(D))+!B !(C)))) */ ;
    defparam i23525_else_3_lut.init = 16'h1e58;
    LUT4 i19999_3_lut (.A(n25517), .B(n22942), .C(index_i[6]), .Z(n22455)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19999_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_0_i627_3_lut_rep_682 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27005)) /* synthesis lut_function=(A (B+!(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i627_3_lut_rep_682.init = 16'hdada;
    LUT4 mux_198_Mux_1_i700_3_lut_4_lut (.A(n26912), .B(index_i[3]), .C(index_i[4]), 
         .D(n684), .Z(n700_adj_2796)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_1_i700_3_lut_4_lut.init = 16'hefe0;
    LUT4 i6421_2_lut (.A(phase_i[9]), .B(phase_i[10]), .Z(index_i_9__N_2106[9])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i6421_2_lut.init = 16'h6666;
    LUT4 i6422_2_lut (.A(phase_i[8]), .B(phase_i[10]), .Z(index_i_9__N_2106[8])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i6422_2_lut.init = 16'h6666;
    LUT4 i11178_4_lut (.A(n15034), .B(index_i[8]), .C(n765), .D(index_i[7]), 
         .Z(n1022)) /* synthesis lut_function=(A (B+(C (D)))+!A (B+(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11178_4_lut.init = 16'hfcdd;
    LUT4 index_i_6__bdd_4_lut_23331 (.A(index_i[6]), .B(n26760), .C(n26879), 
         .D(index_i[5]), .Z(n24772)) /* synthesis lut_function=(!(A (B (C+(D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C (D))))) */ ;
    defparam index_i_6__bdd_4_lut_23331.init = 16'h724e;
    LUT4 index_i_6__bdd_4_lut_23064 (.A(index_i[6]), .B(n26881), .C(index_i[5]), 
         .D(n26755), .Z(n24771)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A (B (C)+!B !(C)))) */ ;
    defparam index_i_6__bdd_4_lut_23064.init = 16'h1cbc;
    LUT4 i6423_2_lut (.A(phase_i[7]), .B(phase_i[10]), .Z(index_i_9__N_2106[7])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i6423_2_lut.init = 16'h6666;
    PFUMX i23527 (.BLUT(n25290), .ALUT(n25286), .C0(index_i[6]), .Z(n25291));
    LUT4 i6424_2_lut (.A(phase_i[6]), .B(phase_i[10]), .Z(index_i_9__N_2106[6])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i6424_2_lut.init = 16'h6666;
    LUT4 i6425_2_lut (.A(phase_i[5]), .B(phase_i[10]), .Z(index_i_9__N_2106[5])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i6425_2_lut.init = 16'h6666;
    LUT4 i15526_3_lut (.A(n26961), .B(n27019), .C(index_i[3]), .Z(n17790)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15526_3_lut.init = 16'hcaca;
    LUT4 i6812_2_lut (.A(index_i[4]), .B(index_i[5]), .Z(n9308)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i6812_2_lut.init = 16'h8888;
    LUT4 i15525_3_lut (.A(n27019), .B(n27015), .C(index_i[3]), .Z(n17789)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15525_3_lut.init = 16'hcaca;
    LUT4 i6426_2_lut (.A(phase_i[4]), .B(phase_i[10]), .Z(index_i_9__N_2106[4])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i6426_2_lut.init = 16'h6666;
    LUT4 i1_2_lut (.A(index_i[6]), .B(index_i[7]), .Z(n19786)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i6427_2_lut (.A(phase_i[3]), .B(phase_i[10]), .Z(index_i_9__N_2106[3])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i6427_2_lut.init = 16'h6666;
    LUT4 mux_198_Mux_2_i189_3_lut_3_lut_4_lut (.A(index_i[1]), .B(n27036), 
         .C(n173_adj_2797), .D(index_i[4]), .Z(n189_adj_2798)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(C+(D)))) */ ;
    defparam mux_198_Mux_2_i189_3_lut_3_lut_4_lut.init = 16'h77f0;
    LUT4 i6428_2_lut (.A(phase_i[2]), .B(phase_i[10]), .Z(index_i_9__N_2106[2])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i6428_2_lut.init = 16'h6666;
    LUT4 i11184_2_lut_3_lut_4_lut (.A(index_i[1]), .B(n27036), .C(index_i[5]), 
         .D(index_i[4]), .Z(n508)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;
    defparam i11184_2_lut_3_lut_4_lut.init = 16'hf080;
    LUT4 i21911_3_lut (.A(n620), .B(n13928), .C(index_i[4]), .Z(n21644)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21911_3_lut.init = 16'hcaca;
    LUT4 i6429_2_lut (.A(phase_i[1]), .B(phase_i[10]), .Z(index_i_9__N_2106[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i6429_2_lut.init = 16'h6666;
    LUT4 n77_bdd_3_lut_23951 (.A(n27010), .B(n29482), .C(index_i[3]), 
         .Z(n25750)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n77_bdd_3_lut_23951.init = 16'hacac;
    PFUMX i19433 (.BLUT(n21868), .ALUT(n21869), .C0(index_i[4]), .Z(n21870));
    LUT4 i19465_3_lut_4_lut (.A(n27037), .B(index_i[2]), .C(index_i[3]), 
         .D(n29481), .Z(n21902)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19465_3_lut_4_lut.init = 16'hf404;
    LUT4 mux_198_Mux_0_i731_3_lut_4_lut (.A(n27037), .B(index_i[2]), .C(index_i[3]), 
         .D(n26972), .Z(n731_adj_2799)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i731_3_lut_4_lut.init = 16'h4f40;
    L6MUX21 i20906 (.D0(n23350), .D1(n23351), .SD(index_i[6]), .Z(n23362));
    PFUMX i19442 (.BLUT(n21877), .ALUT(n21878), .C0(index_i[4]), .Z(n21879));
    L6MUX21 i20907 (.D0(n23352), .D1(n23353), .SD(index_i[6]), .Z(n23363));
    L6MUX21 i20908 (.D0(n23354), .D1(n23355), .SD(index_i[6]), .Z(n23364));
    PFUMX i20909 (.BLUT(n23356), .ALUT(n23357), .C0(index_i[6]), .Z(n23365));
    PFUMX i20980 (.BLUT(n557), .ALUT(n572), .C0(index_i[4]), .Z(n23436));
    PFUMX i20928 (.BLUT(n732), .ALUT(n763_adj_2800), .C0(index_i[5]), 
          .Z(n23384));
    LUT4 i20127_3_lut (.A(n190), .B(n26093), .C(index_i[6]), .Z(n22583)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20127_3_lut.init = 16'hcaca;
    LUT4 i20128_3_lut (.A(n22963), .B(n21633), .C(index_i[6]), .Z(n22584)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20128_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_0_i475_3_lut_4_lut (.A(n26919), .B(index_i[1]), .C(index_i[3]), 
         .D(n26839), .Z(n475_adj_2801)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i475_3_lut_4_lut.init = 16'h4f40;
    LUT4 mux_198_Mux_3_i491_3_lut_4_lut (.A(n26919), .B(index_i[1]), .C(index_i[3]), 
         .D(n27011), .Z(n491_adj_2802)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_3_i491_3_lut_4_lut.init = 16'h4f40;
    LUT4 i21923_3_lut (.A(n491_adj_2803), .B(n506), .C(index_i[4]), .Z(n21638)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21923_3_lut.init = 16'hcaca;
    LUT4 i11146_2_lut_rep_389_3_lut_4_lut (.A(n26760), .B(index_i[4]), .C(index_i[6]), 
         .D(index_i[5]), .Z(n26712)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11146_2_lut_rep_389_3_lut_4_lut.init = 16'hf080;
    LUT4 i22564_2_lut_rep_589 (.A(index_i[1]), .B(index_i[2]), .Z(n26912)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i22564_2_lut_rep_589.init = 16'h9999;
    L6MUX21 i20930 (.D0(n21906), .D1(n891_adj_2804), .SD(index_i[5]), 
            .Z(n23386));
    L6MUX21 i20933 (.D0(n23373), .D1(n23374), .SD(index_i[6]), .Z(n23389));
    L6MUX21 i20935 (.D0(n23377), .D1(n23378), .SD(index_i[6]), .Z(n23391));
    LUT4 i6432_2_lut (.A(phase_i[0]), .B(phase_i[10]), .Z(index_i_9__N_2106[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i6432_2_lut.init = 16'h6666;
    LUT4 n284_bdd_3_lut_24512 (.A(n27039), .B(n27020), .C(index_i[3]), 
         .Z(n25765)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n284_bdd_3_lut_24512.init = 16'hcaca;
    LUT4 i19435_3_lut_4_lut (.A(index_i[0]), .B(n27052), .C(index_i[3]), 
         .D(n27008), .Z(n21872)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19435_3_lut_4_lut.init = 16'hfb0b;
    LUT4 i19089_3_lut (.A(n24719), .B(n21558), .C(index_i[8]), .Z(n21526)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19089_3_lut.init = 16'hcaca;
    L6MUX21 i20936 (.D0(n23379), .D1(n23380), .SD(index_i[6]), .Z(n23392));
    LUT4 i20766_3_lut_3_lut_4_lut (.A(n26839), .B(index_i[3]), .C(n93_adj_2805), 
         .D(index_i[4]), .Z(n23222)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20766_3_lut_3_lut_4_lut.init = 16'hf077;
    LUT4 i12080_3_lut_rep_823 (.A(index_i[2]), .B(index_i[1]), .C(index_i[0]), 
         .Z(n29496)) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i12080_3_lut_rep_823.init = 16'hc4c4;
    LUT4 i20092_3_lut (.A(n25123), .B(n22545), .C(index_i[8]), .Z(n22548)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20092_3_lut.init = 16'hcaca;
    PFUMX i20981 (.BLUT(n589), .ALUT(n604), .C0(index_i[4]), .Z(n23437));
    L6MUX21 i20940 (.D0(n23387), .D1(n23388), .SD(index_i[6]), .Z(n23396));
    LUT4 i20086_3_lut (.A(n22539), .B(n22540), .C(index_i[8]), .Z(n22542)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20086_3_lut.init = 16'hcaca;
    LUT4 i19390_3_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[1]), .C(index_i[0]), 
         .D(index_i[3]), .Z(n21827)) /* synthesis lut_function=(A (B (C)+!B !(C+!(D)))+!A (B (C+!(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19390_3_lut_4_lut_4_lut.init = 16'hc3c4;
    LUT4 mux_198_Mux_0_i397_3_lut (.A(n27042), .B(n29479), .C(index_i[3]), 
         .Z(n397)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i397_3_lut.init = 16'hcaca;
    PFUMX i20982 (.BLUT(n620_adj_2806), .ALUT(n635), .C0(index_i[4]), 
          .Z(n23438));
    LUT4 i20085_3_lut (.A(n22537), .B(n22538), .C(index_i[8]), .Z(n22541)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20085_3_lut.init = 16'hcaca;
    L6MUX21 i19997 (.D0(n21609), .D1(n21612), .SD(index_i[6]), .Z(n22453));
    L6MUX21 i20000 (.D0(n21621), .D1(n21624), .SD(index_i[6]), .Z(n22456));
    L6MUX21 i20001 (.D0(n574), .D1(n21627), .SD(index_i[6]), .Z(n22457));
    L6MUX21 i20002 (.D0(n21630), .D1(n764), .SD(index_i[6]), .Z(n22458));
    PFUMX i20983 (.BLUT(n653), .ALUT(n668), .C0(index_i[4]), .Z(n23439));
    LUT4 i19204_3_lut_4_lut_4_lut_4_lut (.A(n26969), .B(index_i[2]), .C(index_i[3]), 
         .D(index_i[4]), .Z(n21641)) /* synthesis lut_function=(A (B)+!A (B (C (D))+!B !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19204_3_lut_4_lut_4_lut_4_lut.init = 16'hc999;
    LUT4 i19072_3_lut_4_lut (.A(n26969), .B(index_i[2]), .C(index_i[3]), 
         .D(n26950), .Z(n21509)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19072_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_198_Mux_7_i475_3_lut_4_lut (.A(n26969), .B(index_i[2]), .C(index_i[3]), 
         .D(n27042), .Z(n475_adj_2807)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_7_i475_3_lut_4_lut.init = 16'h9f90;
    LUT4 mux_198_Mux_7_i653_3_lut_4_lut (.A(n26969), .B(index_i[2]), .C(index_i[3]), 
         .D(n70), .Z(n653_adj_2808)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_7_i653_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_198_Mux_2_i684_3_lut_4_lut (.A(n26969), .B(index_i[2]), .C(index_i[3]), 
         .D(n29484), .Z(n684_adj_2809)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_2_i684_3_lut_4_lut.init = 16'h6f60;
    L6MUX21 i20583 (.D0(n23023), .D1(n23024), .SD(index_i[6]), .Z(n23039));
    L6MUX21 i20584 (.D0(n23025), .D1(n23026), .SD(index_i[6]), .Z(n23040));
    L6MUX21 i20585 (.D0(n23027), .D1(n23028), .SD(index_i[6]), .Z(n23041));
    PFUMX i20984 (.BLUT(n684_adj_2810), .ALUT(n699_adj_2811), .C0(index_i[4]), 
          .Z(n23440));
    PFUMX i24775 (.BLUT(n27194), .ALUT(n27195), .C0(index_i[8]), .Z(n27196));
    LUT4 i19206_4_lut_4_lut_4_lut (.A(n26969), .B(index_i[2]), .C(index_i[4]), 
         .D(index_i[3]), .Z(n21643)) /* synthesis lut_function=(A (B)+!A !(B (C+(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19206_4_lut_4_lut_4_lut.init = 16'h999c;
    L6MUX21 i20586 (.D0(n23029), .D1(n23030), .SD(index_i[6]), .Z(n23042));
    L6MUX21 i20587 (.D0(n23031), .D1(n23032), .SD(index_i[6]), .Z(n23043));
    PFUMX i20985 (.BLUT(n716_adj_2812), .ALUT(n731_adj_2799), .C0(index_i[4]), 
          .Z(n23441));
    L6MUX21 i20589 (.D0(n23035), .D1(n23036), .SD(index_i[6]), .Z(n23045));
    LUT4 i19087_3_lut_4_lut (.A(n27004), .B(index_i[2]), .C(index_i[3]), 
         .D(n29479), .Z(n21524)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19087_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_198_Mux_0_i188_3_lut (.A(n27041), .B(n101), .C(index_i[3]), 
         .Z(n188)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i188_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_3_i460_3_lut_4_lut (.A(n27004), .B(index_i[2]), .C(index_i[3]), 
         .D(n26958), .Z(n460_adj_2813)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_3_i460_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_198_Mux_6_i285_3_lut_4_lut (.A(n27004), .B(index_i[2]), .C(index_i[3]), 
         .D(n27010), .Z(n285)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_6_i285_3_lut_4_lut.init = 16'hf606;
    LUT4 i20594_3_lut (.A(n23045), .B(n24688), .C(index_i[7]), .Z(n23050)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20594_3_lut.init = 16'hcaca;
    LUT4 i19426_3_lut_4_lut (.A(n27004), .B(index_i[2]), .C(index_i[3]), 
         .D(n27019), .Z(n21863)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19426_3_lut_4_lut.init = 16'hf606;
    PFUMX i20986 (.BLUT(n747_adj_2791), .ALUT(n762_adj_2795), .C0(index_i[4]), 
          .Z(n23442));
    PFUMX i20047 (.BLUT(n22499), .ALUT(n22500), .C0(index_i[6]), .Z(n22503));
    LUT4 i20593_3_lut (.A(n23043), .B(n23044), .C(index_i[7]), .Z(n23049)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20593_3_lut.init = 16'hcaca;
    LUT4 n953_bdd_3_lut_23542_4_lut (.A(n26963), .B(index_i[2]), .C(index_i[3]), 
         .D(n27005), .Z(n25030)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n953_bdd_3_lut_23542_4_lut.init = 16'hf606;
    LUT4 mux_198_Mux_3_i890_3_lut_4_lut (.A(n26963), .B(index_i[2]), .C(index_i[3]), 
         .D(n325), .Z(n890_adj_2814)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_3_i890_3_lut_4_lut.init = 16'h6f60;
    PFUMX i20048 (.BLUT(n22501), .ALUT(n22502), .C0(index_i[6]), .Z(n22504));
    LUT4 i22531_3_lut (.A(n23049), .B(n23050), .C(index_i[8]), .Z(n23052)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22531_3_lut.init = 16'hcaca;
    LUT4 i19054_3_lut_4_lut (.A(n26963), .B(index_i[2]), .C(index_i[3]), 
         .D(n27010), .Z(n21491)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19054_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_198_Mux_0_i348_3_lut_4_lut (.A(n26963), .B(index_i[2]), .C(index_i[3]), 
         .D(n29484), .Z(n348)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i348_3_lut_4_lut.init = 16'h6f60;
    LUT4 i22502_3_lut (.A(n22461), .B(n22462), .C(index_i[8]), .Z(n22465)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22502_3_lut.init = 16'hcaca;
    LUT4 i21979_3_lut (.A(n26340), .B(n124), .C(index_i[4]), .Z(n23223)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21979_3_lut.init = 16'hcaca;
    PFUMX i20987 (.BLUT(n781), .ALUT(n796), .C0(index_i[4]), .Z(n23443));
    PFUMX i20988 (.BLUT(n812), .ALUT(n11922), .C0(index_i[4]), .Z(n23444));
    LUT4 mux_198_Mux_0_i986_3_lut (.A(n29481), .B(n985), .C(index_i[3]), 
         .Z(n986)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i986_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_3_i221_3_lut_4_lut (.A(n26839), .B(index_i[3]), .C(index_i[4]), 
         .D(n26868), .Z(n221_adj_2815)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_3_i221_3_lut_4_lut.init = 16'h08f8;
    LUT4 mux_198_Mux_4_i573_3_lut_4_lut_4_lut_4_lut (.A(n27050), .B(index_i[3]), 
         .C(n26837), .D(index_i[4]), .Z(n573)) /* synthesis lut_function=(!(A (B (D)+!B ((D)+!C))+!A (B (D)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_4_i573_3_lut_4_lut_4_lut_4_lut.init = 16'h11fc;
    LUT4 mux_198_Mux_10_i125_3_lut_4_lut_4_lut (.A(n27050), .B(index_i[3]), 
         .C(index_i[4]), .D(n26839), .Z(n125)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B (C (D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_10_i125_3_lut_4_lut_4_lut.init = 16'h3efe;
    L6MUX21 i20074 (.D0(n22515), .D1(n22516), .SD(index_i[6]), .Z(n22530));
    L6MUX21 i20075 (.D0(n22517), .D1(n22518), .SD(index_i[6]), .Z(n22531));
    LUT4 i20417_3_lut_4_lut (.A(n27050), .B(index_i[3]), .C(index_i[4]), 
         .D(n285_adj_2816), .Z(n22873)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20417_3_lut_4_lut.init = 16'hfe0e;
    L6MUX21 i20076 (.D0(n22519), .D1(n22520), .SD(index_i[6]), .Z(n22532));
    L6MUX21 i20077 (.D0(n22521), .D1(n22522), .SD(index_i[6]), .Z(n22533));
    L6MUX21 i20078 (.D0(n22523), .D1(n22524), .SD(index_i[6]), .Z(n22534));
    LUT4 mux_198_Mux_3_i573_3_lut_3_lut_4_lut (.A(n27050), .B(index_i[3]), 
         .C(n460_adj_2817), .D(index_i[4]), .Z(n573_adj_2818)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_3_i573_3_lut_3_lut_4_lut.init = 16'h11f0;
    L6MUX21 i21003 (.D0(n23451), .D1(n23452), .SD(index_i[6]), .Z(n23459));
    L6MUX21 i21004 (.D0(n23453), .D1(n23454), .SD(index_i[6]), .Z(n23460));
    L6MUX21 i21005 (.D0(n23455), .D1(n23456), .SD(index_i[6]), .Z(n23461));
    LUT4 mux_198_Mux_2_i573_3_lut_3_lut_4_lut (.A(n27050), .B(index_i[3]), 
         .C(n557_adj_2819), .D(index_i[4]), .Z(n573_adj_2820)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_2_i573_3_lut_3_lut_4_lut.init = 16'h11f0;
    LUT4 i22033_3_lut (.A(n109), .B(n124_adj_2821), .C(index_i[4]), .Z(n21611)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22033_3_lut.init = 16'hcaca;
    LUT4 i20770_3_lut_4_lut (.A(n26839), .B(index_i[3]), .C(index_i[4]), 
         .D(n220), .Z(n23226)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20770_3_lut_4_lut.init = 16'hf808;
    LUT4 i20765_3_lut_4_lut (.A(n26839), .B(index_i[3]), .C(index_i[4]), 
         .D(n46), .Z(n23221)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20765_3_lut_4_lut.init = 16'h8f80;
    PFUMX i20990 (.BLUT(n875), .ALUT(n890_adj_2792), .C0(index_i[4]), 
          .Z(n23446));
    L6MUX21 i21006 (.D0(n23457), .D1(n23458), .SD(index_i[6]), .Z(n23462));
    LUT4 i20717_3_lut (.A(n23170), .B(n23171), .C(index_i[8]), .Z(n23173)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20717_3_lut.init = 16'hcaca;
    LUT4 i20716_3_lut (.A(n23168), .B(n23169), .C(index_i[8]), .Z(n23172)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20716_3_lut.init = 16'hcaca;
    PFUMX i20991 (.BLUT(n908), .ALUT(n923), .C0(index_i[4]), .Z(n23447));
    LUT4 i22526_3_lut (.A(n574_adj_2822), .B(n637), .C(index_i[6]), .Z(n21559)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22526_3_lut.init = 16'hcaca;
    PFUMX i20992 (.BLUT(n939), .ALUT(n954), .C0(index_i[4]), .Z(n23448));
    LUT4 i20595_3_lut (.A(n23047), .B(n23048), .C(index_i[8]), .Z(n23051)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20595_3_lut.init = 16'hcaca;
    LUT4 i20946_3_lut (.A(n23399), .B(n23400), .C(index_i[8]), .Z(n23402)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20946_3_lut.init = 16'hcaca;
    LUT4 i20945_3_lut (.A(n23397), .B(n23398), .C(index_i[8]), .Z(n23401)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20945_3_lut.init = 16'hcaca;
    PFUMX i19445 (.BLUT(n21880), .ALUT(n21881), .C0(index_i[4]), .Z(n21882));
    LUT4 i19468_3_lut_4_lut (.A(n26969), .B(index_i[2]), .C(index_i[3]), 
         .D(n27013), .Z(n21905)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19468_3_lut_4_lut.init = 16'hdfd0;
    L6MUX21 i20129 (.D0(n21636), .D1(n21639), .SD(index_i[6]), .Z(n22585));
    PFUMX i20993 (.BLUT(n971), .ALUT(n986), .C0(index_i[4]), .Z(n23449));
    LUT4 i20046_3_lut_4_lut_4_lut (.A(n26824), .B(index_i[4]), .C(index_i[5]), 
         .D(n26800), .Z(n22502)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C)+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20046_3_lut_4_lut_4_lut.init = 16'h0434;
    LUT4 mux_198_Mux_8_i892_3_lut_4_lut (.A(n26824), .B(index_i[4]), .C(index_i[5]), 
         .D(n860), .Z(n892)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_8_i892_3_lut_4_lut.init = 16'h4f40;
    L6MUX21 i20673 (.D0(n23113), .D1(n23114), .SD(index_i[6]), .Z(n23129));
    L6MUX21 i20674 (.D0(n23115), .D1(n23116), .SD(index_i[6]), .Z(n23130));
    L6MUX21 i20130 (.D0(n21642), .D1(n21645), .SD(index_i[6]), .Z(n22586));
    PFUMX i20994 (.BLUT(n1002), .ALUT(n1017), .C0(index_i[4]), .Z(n23450));
    L6MUX21 i20131 (.D0(n21648), .D1(n21651), .SD(index_i[6]), .Z(n22587));
    PFUMX i20132 (.BLUT(n21654), .ALUT(n892_adj_2823), .C0(index_i[6]), 
          .Z(n22588));
    LUT4 i19438_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n21875)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(D))+!A (B (D)+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19438_3_lut_4_lut_4_lut_4_lut.init = 16'hd52b;
    PFUMX i19448 (.BLUT(n21883), .ALUT(n21884), .C0(index_i[4]), .Z(n21885));
    PFUMX i19451 (.BLUT(n21886), .ALUT(n21887), .C0(index_i[4]), .Z(n21888));
    LUT4 mux_198_Mux_2_i270_3_lut (.A(n27012), .B(n26951), .C(index_i[3]), 
         .Z(n270)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_2_i270_3_lut.init = 16'hcaca;
    LUT4 i22067_3_lut (.A(n94), .B(n27223), .C(index_i[5]), .Z(n21581)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22067_3_lut.init = 16'hcaca;
    PFUMX i19457 (.BLUT(n21892), .ALUT(n21893), .C0(index_i[4]), .Z(n21894));
    L6MUX21 i20675 (.D0(n23117), .D1(n23118), .SD(index_i[6]), .Z(n23131));
    LUT4 index_i_2__bdd_4_lut_25583 (.A(index_i[2]), .B(index_i[6]), .C(index_i[5]), 
         .D(index_i[0]), .Z(n28288)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C (D)))+!A (B+(C+(D)))) */ ;
    defparam index_i_2__bdd_4_lut_25583.init = 16'hd7fe;
    LUT4 index_i_2__bdd_3_lut_25598 (.A(index_i[2]), .B(n28288), .C(index_i[1]), 
         .Z(n28289)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam index_i_2__bdd_3_lut_25598.init = 16'hcaca;
    LUT4 index_i_2__bdd_4_lut_25597 (.A(index_i[2]), .B(n26837), .C(index_i[6]), 
         .D(index_i[5]), .Z(n28290)) /* synthesis lut_function=(!(A (B+!((D)+!C))+!A (B ((D)+!C)))) */ ;
    defparam index_i_2__bdd_4_lut_25597.init = 16'h3353;
    PFUMX i19463 (.BLUT(n21898), .ALUT(n21899), .C0(index_i[4]), .Z(n21900));
    LUT4 mux_198_Mux_9_i763_3_lut_4_lut (.A(n27037), .B(n26966), .C(index_i[4]), 
         .D(n26845), .Z(n763)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;
    defparam mux_198_Mux_9_i763_3_lut_4_lut.init = 16'hf101;
    LUT4 i15575_4_lut (.A(index_i[0]), .B(index_i[4]), .C(index_i[1]), 
         .D(n26966), .Z(n286)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i15575_4_lut.init = 16'hccc8;
    PFUMX i19119 (.BLUT(n318), .ALUT(n381), .C0(index_i[6]), .Z(n21556));
    PFUMX i19466 (.BLUT(n21901), .ALUT(n21902), .C0(index_i[4]), .Z(n21903));
    LUT4 mux_198_Mux_8_i763_3_lut_4_lut (.A(n27037), .B(n26966), .C(index_i[4]), 
         .D(n26845), .Z(n15052)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam mux_198_Mux_8_i763_3_lut_4_lut.init = 16'hfe0e;
    LUT4 i9445_3_lut_4_lut (.A(n26959), .B(index_i[2]), .C(n27049), .D(n27018), 
         .Z(n444)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9445_3_lut_4_lut.init = 16'h6f60;
    PFUMX i19469 (.BLUT(n21904), .ALUT(n21905), .C0(index_i[4]), .Z(n21906));
    LUT4 n24548_bdd_3_lut_26181 (.A(n24548), .B(n24541), .C(index_i[7]), 
         .Z(n24549)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n24548_bdd_3_lut_26181.init = 16'hcaca;
    LUT4 mux_198_Mux_4_i747_3_lut_4_lut (.A(n26959), .B(index_i[2]), .C(index_i[3]), 
         .D(n29479), .Z(n747_adj_2824)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_4_i747_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_198_Mux_6_i251_3_lut_4_lut (.A(n26959), .B(index_i[2]), .C(index_i[3]), 
         .D(n27018), .Z(n251_adj_2825)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_6_i251_3_lut_4_lut.init = 16'hf606;
    LUT4 n262_bdd_2_lut_24219_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[3]), 
         .Z(n26042)) /* synthesis lut_function=(A (B+(C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n262_bdd_2_lut_24219_3_lut.init = 16'hf9f9;
    LUT4 n773_bdd_3_lut_23285_4_lut (.A(n26953), .B(index_i[2]), .C(n27008), 
         .D(index_i[3]), .Z(n25022)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n773_bdd_3_lut_23285_4_lut.init = 16'hf066;
    PFUMX i20677 (.BLUT(n23121), .ALUT(n23122), .C0(index_i[6]), .Z(n23133));
    LUT4 mux_198_Mux_0_i93_3_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .Z(n93_adj_2805)) /* synthesis lut_function=(A (B)+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i93_3_lut_3_lut.init = 16'h9c9c;
    LUT4 mux_198_Mux_3_i668_3_lut_4_lut (.A(n26953), .B(index_i[2]), .C(index_i[3]), 
         .D(n27015), .Z(n668_adj_2826)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_3_i668_3_lut_4_lut.init = 16'h6f60;
    L6MUX21 i20678 (.D0(n23123), .D1(n23124), .SD(index_i[6]), .Z(n23134));
    L6MUX21 i20679 (.D0(n23125), .D1(n23126), .SD(index_i[6]), .Z(n23135));
    PFUMX i20680 (.BLUT(n23127), .ALUT(n23128), .C0(index_i[6]), .Z(n23136));
    L6MUX21 i20126 (.D0(n22949), .D1(n22956), .SD(index_i[6]), .Z(n22582));
    LUT4 mux_198_Mux_4_i763_3_lut_4_lut (.A(n26953), .B(index_i[2]), .C(index_i[4]), 
         .D(n747_adj_2824), .Z(n763_adj_2827)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_4_i763_3_lut_4_lut.init = 16'h6f60;
    LUT4 i19389_3_lut_3_lut_4_lut (.A(index_i[2]), .B(n27037), .C(n645), 
         .D(index_i[3]), .Z(n21826)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (B (C (D))+!B (C+!(D)))) */ ;
    defparam i19389_3_lut_3_lut_4_lut.init = 16'hf099;
    LUT4 n476_bdd_3_lut_23594_3_lut_4_lut (.A(index_i[2]), .B(n27037), .C(n491_adj_2828), 
         .D(index_i[4]), .Z(n25356)) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))+!A !(B ((D)+!C)+!B !(C+(D)))) */ ;
    defparam n476_bdd_3_lut_23594_3_lut_4_lut.init = 16'h99f0;
    LUT4 i19071_3_lut_3_lut_4_lut (.A(index_i[2]), .B(n27037), .C(n26948), 
         .D(index_i[3]), .Z(n21508)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (B (C (D))+!B (C+!(D)))) */ ;
    defparam i19071_3_lut_3_lut_4_lut.init = 16'hf099;
    PFUMX i20700 (.BLUT(n797), .ALUT(n828), .C0(index_i[5]), .Z(n23156));
    LUT4 mux_198_Mux_7_i443_3_lut_4_lut (.A(index_i[2]), .B(n27037), .C(index_i[3]), 
         .D(n26948), .Z(n443_adj_2829)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;
    defparam mux_198_Mux_7_i443_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_198_Mux_3_i860_3_lut_4_lut (.A(index_i[2]), .B(n27037), .C(index_i[4]), 
         .D(n859), .Z(n860_adj_2830)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam mux_198_Mux_3_i860_3_lut_4_lut.init = 16'hf606;
    L6MUX21 i20704 (.D0(n23144), .D1(n23145), .SD(index_i[6]), .Z(n23160));
    L6MUX21 i20705 (.D0(n23146), .D1(n23147), .SD(index_i[6]), .Z(n23161));
    L6MUX21 i20706 (.D0(n23148), .D1(n23149), .SD(index_i[6]), .Z(n23162));
    L6MUX21 i20707 (.D0(n23150), .D1(n23151), .SD(index_i[6]), .Z(n23163));
    L6MUX21 i20708 (.D0(n23152), .D1(n23153), .SD(index_i[6]), .Z(n23164));
    L6MUX21 i20711 (.D0(n23158), .D1(n23159), .SD(index_i[6]), .Z(n23167));
    LUT4 mux_198_Mux_0_i971_3_lut (.A(n29482), .B(n27038), .C(index_i[3]), 
         .Z(n971)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i971_3_lut.init = 16'hcaca;
    LUT4 i21553_3_lut (.A(n21835), .B(n27142), .C(index_i[4]), .Z(n21837)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21553_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_3_i924_3_lut (.A(n908_adj_2831), .B(index_i[0]), .C(index_i[4]), 
         .Z(n924_adj_2832)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_3_i924_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_3_i891_3_lut (.A(n541_adj_2833), .B(n890_adj_2814), 
         .C(index_i[4]), .Z(n891_adj_2834)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_3_i891_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_3_i669_3_lut (.A(n653_adj_2835), .B(n668_adj_2826), 
         .C(index_i[4]), .Z(n669)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_3_i669_3_lut.init = 16'hcaca;
    LUT4 i11149_3_lut_4_lut (.A(n26712), .B(index_i[7]), .C(index_i[8]), 
         .D(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2126[14])) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11149_3_lut_4_lut.init = 16'hffe0;
    LUT4 i9465_4_lut (.A(n27050), .B(n26839), .C(index_i[3]), .D(index_i[4]), 
         .Z(n12026)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B ((D)+!C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9465_4_lut.init = 16'h3afa;
    LUT4 i21570_3_lut (.A(n21823), .B(n21824), .C(index_i[4]), .Z(n21825)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21570_3_lut.init = 16'hcaca;
    PFUMX mux_198_Mux_1_i636 (.BLUT(n620_adj_2836), .ALUT(n635_adj_2837), 
          .C0(index_i[4]), .Z(n636)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 mux_198_Mux_3_i476_3_lut (.A(n460_adj_2813), .B(n285), .C(index_i[4]), 
         .Z(n476_adj_2838)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_3_i476_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_3_i413_3_lut (.A(n397_adj_2839), .B(n26944), .C(index_i[4]), 
         .Z(n413)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_3_i413_3_lut.init = 16'hcaca;
    LUT4 i22568_2_lut_rep_686 (.A(index_i[0]), .B(index_i[1]), .Z(n27009)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i22568_2_lut_rep_686.init = 16'h9999;
    LUT4 i19078_3_lut_4_lut (.A(n27053), .B(index_i[1]), .C(index_i[3]), 
         .D(n404), .Z(n21515)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19078_3_lut_4_lut.init = 16'hdfd0;
    LUT4 i12123_3_lut (.A(index_i[2]), .B(index_i[1]), .C(index_i[0]), 
         .Z(n1001)) /* synthesis lut_function=(A (B)+!A (B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i12123_3_lut.init = 16'hdcdc;
    LUT4 mux_198_Mux_3_i286_4_lut (.A(n93_adj_2840), .B(index_i[2]), .C(index_i[4]), 
         .D(n14831), .Z(n286_adj_2841)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_3_i286_4_lut.init = 16'h3aca;
    LUT4 mux_198_Mux_1_i620_3_lut_4_lut (.A(n27053), .B(index_i[1]), .C(index_i[3]), 
         .D(n27017), .Z(n620_adj_2836)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_1_i620_3_lut_4_lut.init = 16'hdfd0;
    LUT4 mux_198_Mux_0_i173_3_lut_4_lut (.A(n27053), .B(index_i[1]), .C(index_i[3]), 
         .D(n27015), .Z(n173_adj_2842)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i173_3_lut_4_lut.init = 16'hdfd0;
    LUT4 mux_198_Mux_8_i732_3_lut (.A(index_i[3]), .B(n15052), .C(index_i[5]), 
         .Z(n732_adj_2843)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_8_i732_3_lut.init = 16'h3a3a;
    LUT4 i20052_4_lut_4_lut (.A(n26760), .B(n26881), .C(index_i[5]), .D(index_i[4]), 
         .Z(n22508)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C+(D))+!B !(C (D)+!C !(D)))) */ ;
    defparam i20052_4_lut_4_lut.init = 16'hcf50;
    PFUMX mux_198_Mux_2_i891 (.BLUT(n875_adj_2844), .ALUT(n890_adj_2845), 
          .C0(index_i[4]), .Z(n891_adj_2846)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    PFUMX mux_198_Mux_2_i860 (.BLUT(n844_adj_2785), .ALUT(n859_adj_2847), 
          .C0(index_i[4]), .Z(n860_adj_2848)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 mux_198_Mux_2_i955_then_4_lut (.A(index_i[4]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n27163)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B (C+!(D))+!B !(C (D)))) */ ;
    defparam mux_198_Mux_2_i955_then_4_lut.init = 16'he95d;
    LUT4 i9477_3_lut_4_lut (.A(index_i[0]), .B(n27052), .C(index_i[4]), 
         .D(n588), .Z(n12038)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9477_3_lut_4_lut.init = 16'h4f40;
    LUT4 mux_198_Mux_2_i859_3_lut_4_lut (.A(index_i[0]), .B(n27052), .C(index_i[3]), 
         .D(n26954), .Z(n859_adj_2847)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_2_i859_3_lut_4_lut.init = 16'h4f40;
    LUT4 i19395_3_lut_4_lut (.A(index_i[0]), .B(n27052), .C(index_i[3]), 
         .D(n26964), .Z(n21832)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19395_3_lut_4_lut.init = 16'hf404;
    PFUMX i19079 (.BLUT(n21514), .ALUT(n21515), .C0(index_i[4]), .Z(n21516));
    LUT4 mux_198_Mux_3_i158_3_lut (.A(n142), .B(n26761), .C(index_i[4]), 
         .Z(n158)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_3_i158_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_3_i125_3_lut (.A(n46_adj_2849), .B(n526_adj_2850), 
         .C(index_i[4]), .Z(n125_adj_2851)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_3_i125_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_2_i316_3_lut (.A(n27016), .B(n26958), .C(index_i[3]), 
         .Z(n316_adj_2852)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_2_i316_3_lut.init = 16'hcaca;
    LUT4 i21596_3_lut (.A(n21403), .B(n21404), .C(index_i[4]), .Z(n21405)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i21596_3_lut.init = 16'hcaca;
    PFUMX mux_198_Mux_3_i763 (.BLUT(n747_adj_2853), .ALUT(n762_adj_2854), 
          .C0(index_i[4]), .Z(n763_adj_2855)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 n62_bdd_3_lut_25943 (.A(n62_adj_2787), .B(n125), .C(index_i[6]), 
         .Z(n28615)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n62_bdd_3_lut_25943.init = 16'hcaca;
    LUT4 n22508_bdd_4_lut_25940 (.A(n252_adj_2856), .B(n26868), .C(index_i[4]), 
         .D(index_i[5]), .Z(n28613)) /* synthesis lut_function=(A (B (D)+!B ((D)+!C))+!A !(B+(C+(D)))) */ ;
    defparam n22508_bdd_4_lut_25940.init = 16'haa03;
    LUT4 mux_198_Mux_2_i397_3_lut (.A(n29496), .B(n26948), .C(index_i[3]), 
         .Z(n397_adj_2857)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_2_i397_3_lut.init = 16'hcaca;
    LUT4 n62_bdd_4_lut_25944 (.A(n26966), .B(n26838), .C(index_i[6]), 
         .D(index_i[4]), .Z(n28616)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C+(D)))+!A (B ((D)+!C)+!B !(C)))) */ ;
    defparam n62_bdd_4_lut_25944.init = 16'h3af0;
    LUT4 n627_bdd_3_lut_24208 (.A(n27005), .B(n29482), .C(index_i[3]), 
         .Z(n26034)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n627_bdd_3_lut_24208.init = 16'hcaca;
    PFUMX i19172 (.BLUT(n21607), .ALUT(n21608), .C0(index_i[5]), .Z(n21609));
    LUT4 mux_198_Mux_2_i955_else_4_lut (.A(index_i[4]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n27162)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+(D)))+!A !(B (C+!(D))+!B !(C+!(D))))) */ ;
    defparam mux_198_Mux_2_i955_else_4_lut.init = 16'h49c6;
    PFUMX i19175 (.BLUT(n21610), .ALUT(n21611), .C0(index_i[5]), .Z(n21612));
    LUT4 n262_bdd_3_lut_24220 (.A(n26957), .B(n29496), .C(index_i[3]), 
         .Z(n26043)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n262_bdd_3_lut_24220.init = 16'hcaca;
    LUT4 i20672_4_lut (.A(n21816), .B(n1002_adj_2858), .C(index_i[5]), 
         .D(index_i[4]), .Z(n23128)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;
    defparam i20672_4_lut.init = 16'hfaca;
    LUT4 mux_198_Mux_4_i860_3_lut (.A(n506_adj_2859), .B(n15), .C(index_i[4]), 
         .Z(n860_adj_2860)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_4_i860_3_lut.init = 16'hcaca;
    LUT4 i21628_3_lut (.A(n21805), .B(n21806), .C(index_i[4]), .Z(n21807)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21628_3_lut.init = 16'hcaca;
    LUT4 n627_bdd_3_lut_24246 (.A(n27005), .B(n588), .C(index_i[3]), .Z(n26045)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n627_bdd_3_lut_24246.init = 16'hacac;
    LUT4 i21630_3_lut (.A(n21802), .B(n21803), .C(index_i[4]), .Z(n21804)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21630_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_3_i653_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n653_adj_2835)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A !(B (D)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_3_i653_3_lut_4_lut_4_lut.init = 16'h4d99;
    LUT4 n28754_bdd_3_lut (.A(n28754), .B(index_i[1]), .C(index_i[4]), 
         .Z(n28755)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n28754_bdd_3_lut.init = 16'hcaca;
    LUT4 index_i_1__bdd_4_lut_25935 (.A(index_i[1]), .B(index_i[3]), .C(index_i[0]), 
         .D(index_i[2]), .Z(n28754)) /* synthesis lut_function=(A (B (C+(D))+!B (C (D)))+!A !(B (C)+!B !(C+(D)))) */ ;
    defparam index_i_1__bdd_4_lut_25935.init = 16'hbd94;
    LUT4 mux_198_Mux_4_i700_3_lut (.A(n684_adj_2861), .B(index_i[1]), .C(index_i[4]), 
         .Z(n700_adj_2862)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_4_i700_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_4_i669_3_lut (.A(n781_adj_2863), .B(n668_adj_2864), 
         .C(index_i[4]), .Z(n669_adj_2865)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_4_i669_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_4_i542_3_lut (.A(n526_adj_2850), .B(n506_adj_2866), 
         .C(index_i[4]), .Z(n542_adj_2867)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_4_i542_3_lut.init = 16'hcaca;
    LUT4 i11208_3_lut_4_lut (.A(index_i[4]), .B(n27036), .C(index_i[5]), 
         .D(n26969), .Z(n892_adj_2868)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11208_3_lut_4_lut.init = 16'hf8f0;
    LUT4 i20666_4_lut (.A(n26814), .B(n27134), .C(index_i[5]), .D(index_i[4]), 
         .Z(n23122)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam i20666_4_lut.init = 16'hc5ca;
    LUT4 mux_198_Mux_6_i844_3_lut_4_lut (.A(n26969), .B(index_i[2]), .C(index_i[3]), 
         .D(n26970), .Z(n844_adj_2869)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_6_i844_3_lut_4_lut.init = 16'hf808;
    LUT4 index_i_6__bdd_3_lut_23065_4_lut_4_lut (.A(n26969), .B(index_i[2]), 
         .C(index_i[5]), .D(index_i[3]), .Z(n24773)) /* synthesis lut_function=(!(A (B (C)+!B ((D)+!C))+!A (B (C (D))+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam index_i_6__bdd_3_lut_23065_4_lut_4_lut.init = 16'h0c7c;
    LUT4 mux_198_Mux_4_i286_3_lut (.A(n270_adj_2870), .B(n15_adj_2871), 
         .C(index_i[4]), .Z(n286_adj_2872)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_4_i286_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_8_i157_3_lut_4_lut (.A(n26969), .B(index_i[2]), .C(index_i[3]), 
         .D(n26949), .Z(n15_adj_2873)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_8_i157_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_198_Mux_4_i94_3_lut (.A(n61), .B(n26945), .C(index_i[4]), 
         .Z(n94_adj_2874)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_4_i94_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_8_i301_3_lut_4_lut (.A(n26969), .B(index_i[2]), .C(index_i[3]), 
         .D(n70), .Z(n301)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_8_i301_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_198_Mux_2_i890_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n890_adj_2845)) /* synthesis lut_function=(A (B (C)+!B !(C+!(D)))+!A !(B (C+(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_2_i890_3_lut_4_lut_4_lut.init = 16'h9394;
    LUT4 mux_198_Mux_8_i173_3_lut_3_lut_4_lut (.A(n26969), .B(index_i[2]), 
         .C(n954_adj_2875), .D(index_i[4]), .Z(n173)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_8_i173_3_lut_3_lut_4_lut.init = 16'hf077;
    LUT4 mux_198_Mux_3_i251_3_lut_4_lut (.A(n26969), .B(index_i[2]), .C(index_i[3]), 
         .D(n26880), .Z(n15054)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_3_i251_3_lut_4_lut.init = 16'h8f80;
    PFUMX i19082 (.BLUT(n21517), .ALUT(n21518), .C0(index_i[4]), .Z(n21519));
    LUT4 mux_198_Mux_8_i653_3_lut_rep_400_3_lut_4_lut (.A(n26969), .B(index_i[2]), 
         .C(index_i[3]), .D(n26879), .Z(n26723)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_8_i653_3_lut_rep_400_3_lut_4_lut.init = 16'h08f8;
    LUT4 i19458_3_lut_3_lut_4_lut (.A(n26969), .B(index_i[2]), .C(n1001), 
         .D(index_i[3]), .Z(n21895)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19458_3_lut_3_lut_4_lut.init = 16'hf077;
    LUT4 index_i_6__bdd_3_lut_23410_4_lut_3_lut_4_lut (.A(n26969), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[5]), .Z(n24774)) /* synthesis lut_function=(!(A (B (D)+!B !(C+(D)))+!A !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam index_i_6__bdd_3_lut_23410_4_lut_3_lut_4_lut.init = 16'h77f8;
    LUT4 mux_198_Mux_9_i364_3_lut_3_lut_4_lut (.A(n26969), .B(index_i[2]), 
         .C(n26880), .D(index_i[3]), .Z(n364)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_9_i364_3_lut_3_lut_4_lut.init = 16'h77f0;
    LUT4 n21407_bdd_3_lut (.A(n27012), .B(n26948), .C(index_i[3]), .Z(n26089)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n21407_bdd_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_3_i828_3_lut_3_lut_4_lut_4_lut_4_lut (.A(n26969), .B(index_i[2]), 
         .C(index_i[4]), .D(index_i[3]), .Z(n828)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C (D)+!C !(D)))+!A !(B (C+!(D))+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_3_i828_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h70c7;
    LUT4 i22643_2_lut_rep_412_3_lut_4_lut (.A(n26969), .B(index_i[2]), .C(index_i[5]), 
         .D(n26968), .Z(n26735)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i22643_2_lut_rep_412_3_lut_4_lut.init = 16'h0f7f;
    LUT4 mux_198_Mux_3_i1018_3_lut_4_lut (.A(index_i[1]), .B(n26966), .C(index_i[4]), 
         .D(n19863), .Z(n1018)) /* synthesis lut_function=(A (C+!(D))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_3_i1018_3_lut_4_lut.init = 16'he0ef;
    LUT4 mux_198_Mux_2_i700_3_lut_4_lut (.A(index_i[1]), .B(n26966), .C(index_i[4]), 
         .D(n684_adj_2809), .Z(n700_adj_2876)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_2_i700_3_lut_4_lut.init = 16'hefe0;
    PFUMX i19184 (.BLUT(n21619), .ALUT(n21620), .C0(index_i[5]), .Z(n21621));
    LUT4 mux_198_Mux_4_i62_4_lut (.A(n27051), .B(n61), .C(index_i[4]), 
         .D(index_i[3]), .Z(n62_adj_2877)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_4_i62_4_lut.init = 16'hc5ca;
    LUT4 mux_198_Mux_4_i31_4_lut (.A(n15_adj_2871), .B(n26802), .C(index_i[4]), 
         .D(index_i[3]), .Z(n31)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_4_i31_4_lut.init = 16'h3aca;
    LUT4 mux_198_Mux_3_i31_3_lut (.A(n781_adj_2863), .B(n30), .C(index_i[4]), 
         .Z(n31_adj_2878)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_3_i31_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_8_i124_3_lut_3_lut_4_lut (.A(n27037), .B(index_i[2]), 
         .C(n26970), .D(index_i[3]), .Z(n124_adj_2821)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_8_i124_3_lut_3_lut_4_lut.init = 16'h11f0;
    LUT4 mux_198_Mux_6_i890_3_lut_3_lut_4_lut (.A(n27037), .B(index_i[2]), 
         .C(n27038), .D(index_i[3]), .Z(n890_adj_2879)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_6_i890_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 mux_198_Mux_0_i1002_3_lut_3_lut_4_lut (.A(n27037), .B(index_i[2]), 
         .C(n1001), .D(index_i[3]), .Z(n1002)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i1002_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 mux_198_Mux_8_i475_3_lut_3_lut_4_lut (.A(n27037), .B(index_i[2]), 
         .C(n26880), .D(index_i[3]), .Z(n475_adj_2880)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_8_i475_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 mux_198_Mux_9_i31_3_lut_4_lut_then_4_lut (.A(index_i[4]), .B(index_i[0]), 
         .C(index_i[2]), .D(index_i[1]), .Z(n27169)) /* synthesis lut_function=(A (B (C (D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_9_i31_3_lut_4_lut_then_4_lut.init = 16'hd550;
    LUT4 mux_198_Mux_9_i31_3_lut_4_lut_else_4_lut (.A(index_i[4]), .B(index_i[2]), 
         .Z(n27168)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_9_i31_3_lut_4_lut_else_4_lut.init = 16'h2222;
    PFUMX i19085 (.BLUT(n21520), .ALUT(n21521), .C0(index_i[4]), .Z(n21522));
    LUT4 mux_198_Mux_3_i93_3_lut_4_lut (.A(n27037), .B(index_i[2]), .C(index_i[3]), 
         .D(n70), .Z(n93_adj_2840)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_3_i93_3_lut_4_lut.init = 16'hefe0;
    LUT4 mux_198_Mux_7_i890_3_lut_3_lut_4_lut (.A(n27037), .B(index_i[2]), 
         .C(n26879), .D(index_i[3]), .Z(n890)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_7_i890_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 index_i_4__bdd_4_lut_25331 (.A(index_i[4]), .B(n26778), .C(n24542), 
         .D(index_i[5]), .Z(n26705)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (B (C (D))+!B (C+!(D)))) */ ;
    defparam index_i_4__bdd_4_lut_25331.init = 16'hf099;
    LUT4 mux_198_Mux_0_i795_3_lut_3_lut_rep_793 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29466)) /* synthesis lut_function=(A (B+(C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i795_3_lut_3_lut_rep_793.init = 16'hadad;
    LUT4 i21682_3_lut (.A(n716_adj_2881), .B(n731), .C(index_i[4]), .Z(n732_adj_2882)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21682_3_lut.init = 16'hcaca;
    LUT4 i20426_3_lut_4_lut (.A(n26837), .B(index_i[3]), .C(index_i[4]), 
         .D(n26824), .Z(n22882)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20426_3_lut_4_lut.init = 16'hfe0e;
    LUT4 mux_198_Mux_2_i669_3_lut (.A(n653_adj_2883), .B(n25049), .C(index_i[4]), 
         .Z(n669_adj_2884)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_2_i669_3_lut.init = 16'hcaca;
    PFUMX i19187 (.BLUT(n21622), .ALUT(n21623), .C0(index_i[5]), .Z(n21624));
    LUT4 mux_198_Mux_2_i605_3_lut (.A(n142), .B(n604_adj_2885), .C(index_i[4]), 
         .Z(n605)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_2_i605_3_lut.init = 16'hcaca;
    LUT4 i12264_1_lut_2_lut_3_lut_4_lut (.A(n26837), .B(index_i[3]), .C(index_i[5]), 
         .D(index_i[4]), .Z(n381)) /* synthesis lut_function=(!(A (C+(D))+!A (B (C+(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i12264_1_lut_2_lut_3_lut_4_lut.init = 16'h010f;
    LUT4 mux_198_Mux_10_i413_3_lut_3_lut_4_lut (.A(n26837), .B(index_i[3]), 
         .C(n26800), .D(index_i[4]), .Z(n413_adj_2886)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_10_i413_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 i21687_3_lut (.A(n29499), .B(n21854), .C(index_i[4]), .Z(n21855)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21687_3_lut.init = 16'hcaca;
    LUT4 index_i_7__bdd_4_lut_24932 (.A(index_i[7]), .B(n14956), .C(n24714), 
         .D(index_i[5]), .Z(n26708)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(B (C+(D))+!B !((D)+!C)))) */ ;
    defparam index_i_7__bdd_4_lut_24932.init = 16'h66f0;
    PFUMX i19190 (.BLUT(n21625), .ALUT(n21626), .C0(index_i[5]), .Z(n21627));
    LUT4 i20424_3_lut_3_lut_4_lut (.A(n26837), .B(index_i[3]), .C(n412_adj_2887), 
         .D(index_i[4]), .Z(n22880)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20424_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 i21694_3_lut (.A(n21850), .B(n21851), .C(index_i[4]), .Z(n21852)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21694_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_10_i252_3_lut_4_lut_4_lut (.A(n26837), .B(index_i[3]), 
         .C(index_i[4]), .D(n26839), .Z(n252_adj_2856)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B (C (D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_10_i252_3_lut_4_lut_4_lut.init = 16'h3efe;
    LUT4 mux_198_Mux_2_i413_3_lut (.A(n397_adj_2857), .B(n954_adj_2875), 
         .C(index_i[4]), .Z(n413_adj_2888)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_2_i413_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_2_i317_3_lut (.A(n668_adj_2826), .B(n316_adj_2852), 
         .C(index_i[4]), .Z(n317_adj_2889)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_2_i317_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_2_i286_3_lut (.A(n270), .B(n653_adj_2835), .C(index_i[4]), 
         .Z(n286_adj_2890)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_2_i286_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_0_i796_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n796)) /* synthesis lut_function=(A (B (C+(D))+!B (C (D)))+!A !(B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i796_3_lut_4_lut_4_lut.init = 16'hadc0;
    LUT4 i21707_3_lut (.A(n142_adj_2891), .B(n14052), .C(index_i[4]), 
         .Z(n158_adj_2892)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21707_3_lut.init = 16'hcaca;
    PFUMX i20659 (.BLUT(n158_adj_2893), .ALUT(n189_adj_2894), .C0(index_i[5]), 
          .Z(n23115));
    LUT4 mux_198_Mux_0_i939_4_lut (.A(n588), .B(n26959), .C(index_i[3]), 
         .D(index_i[2]), .Z(n939)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i939_4_lut.init = 16'hfaca;
    PFUMX i20780 (.BLUT(n23220), .ALUT(n23221), .C0(index_i[5]), .Z(n23236));
    PFUMX i20781 (.BLUT(n23222), .ALUT(n23223), .C0(index_i[5]), .Z(n23237));
    L6MUX21 i20782 (.D0(n23224), .D1(n23225), .SD(index_i[5]), .Z(n23238));
    LUT4 i19687_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n22124)) /* synthesis lut_function=(A (B (C)+!B !(C (D)+!C !(D)))+!A (B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19687_3_lut_4_lut_4_lut.init = 16'hd6a5;
    PFUMX i20783 (.BLUT(n23226), .ALUT(n23227), .C0(index_i[5]), .Z(n23239));
    PFUMX i19088 (.BLUT(n21523), .ALUT(n21524), .C0(index_i[4]), .Z(n21525));
    LUT4 n21317_bdd_3_lut_23288 (.A(n29483), .B(n27010), .C(index_i[3]), 
         .Z(n25025)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n21317_bdd_3_lut_23288.init = 16'hcaca;
    L6MUX21 i20785 (.D0(n23230), .D1(n23231), .SD(index_i[5]), .Z(n23241));
    PFUMX mux_198_Mux_5_i732 (.BLUT(n12012), .ALUT(n731_adj_2895), .C0(index_i[4]), 
          .Z(n732_adj_2896)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 n21559_bdd_3_lut (.A(n26715), .B(n701), .C(index_i[6]), .Z(n26236)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n21559_bdd_3_lut.init = 16'hacac;
    L6MUX21 i20786 (.D0(n23232), .D1(n23233), .SD(index_i[5]), .Z(n23242));
    L6MUX21 i20787 (.D0(n23234), .D1(n23235), .SD(index_i[5]), .Z(n23243));
    PFUMX i19193 (.BLUT(n21628), .ALUT(n21629), .C0(index_i[5]), .Z(n21630));
    LUT4 n953_bdd_3_lut_23293 (.A(n26954), .B(index_i[3]), .C(n27018), 
         .Z(n25029)) /* synthesis lut_function=(A (B+(C))+!A !(B+!(C))) */ ;
    defparam n953_bdd_3_lut_23293.init = 16'hb8b8;
    LUT4 n26239_bdd_3_lut (.A(n28618), .B(n22505), .C(index_i[8]), .Z(n26240)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n26239_bdd_3_lut.init = 16'hcaca;
    LUT4 n285_bdd_3_lut (.A(n26954), .B(n29479), .C(index_i[3]), .Z(n25032)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n285_bdd_3_lut.init = 16'hacac;
    PFUMX i19196 (.BLUT(n21631), .ALUT(n21632), .C0(index_i[5]), .Z(n21633));
    LUT4 mux_198_Mux_5_i891_3_lut (.A(n875_adj_2897), .B(n379_adj_2898), 
         .C(index_i[4]), .Z(n891_adj_2899)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_5_i891_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_5_i860_3_lut (.A(n15_adj_2900), .B(n859_adj_2901), 
         .C(index_i[4]), .Z(n860_adj_2902)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_5_i860_3_lut.init = 16'hcaca;
    LUT4 i21744_3_lut (.A(n22123), .B(n22124), .C(index_i[4]), .Z(n22125)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21744_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_5_i636_4_lut (.A(n157_adj_2903), .B(n26829), .C(index_i[4]), 
         .D(index_i[3]), .Z(n636_adj_2904)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_5_i636_4_lut.init = 16'h3aca;
    LUT4 n21506_bdd_3_lut_24029 (.A(n29481), .B(n29482), .C(index_i[3]), 
         .Z(n25047)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n21506_bdd_3_lut_24029.init = 16'hcaca;
    LUT4 i21747_3_lut (.A(n17792), .B(n17793), .C(index_i[4]), .Z(n17794)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21747_3_lut.init = 16'hcaca;
    LUT4 n308_bdd_3_lut_24032 (.A(n29467), .B(n27011), .C(index_i[3]), 
         .Z(n25050)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n308_bdd_3_lut_24032.init = 16'hacac;
    LUT4 mux_198_Mux_5_i507_3_lut (.A(n491), .B(n506_adj_2859), .C(index_i[4]), 
         .Z(n507)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_5_i507_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_5_i476_3_lut (.A(n460_adj_2905), .B(n475), .C(index_i[4]), 
         .Z(n476_adj_2906)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_5_i476_3_lut.init = 16'hcaca;
    PFUMX i23395 (.BLUT(n26837), .ALUT(n25132), .C0(index_i[3]), .Z(n25133));
    LUT4 mux_198_Mux_5_i413_3_lut (.A(n397_adj_2907), .B(n251_adj_2825), 
         .C(index_i[4]), .Z(n413_adj_2908)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_5_i413_3_lut.init = 16'hcaca;
    LUT4 n25054_bdd_3_lut (.A(n25054), .B(n157_adj_2909), .C(index_i[4]), 
         .Z(n25055)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n25054_bdd_3_lut.init = 16'hcaca;
    LUT4 i15563_3_lut (.A(n17825), .B(n17826), .C(index_i[4]), .Z(n17827)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15563_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_5_i125_3_lut (.A(n109_adj_2910), .B(n124_adj_2911), 
         .C(index_i[4]), .Z(n125_adj_2912)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_5_i125_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_5_i94_3_lut (.A(n653_adj_2913), .B(n635_adj_2914), 
         .C(index_i[4]), .Z(n94_adj_2915)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_5_i94_3_lut.init = 16'hcaca;
    LUT4 i20004_3_lut_4_lut (.A(n26765), .B(n26771), .C(index_i[5]), .D(index_i[6]), 
         .Z(n22460)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (B+((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20004_3_lut_4_lut.init = 16'hffc5;
    LUT4 n254_bdd_4_lut (.A(index_i[5]), .B(index_i[3]), .C(index_i[6]), 
         .D(index_i[4]), .Z(n26271)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;
    defparam n254_bdd_4_lut.init = 16'hf8f0;
    LUT4 mux_198_Mux_5_i31_3_lut (.A(n15_adj_2900), .B(n30_adj_2916), .C(index_i[4]), 
         .Z(n31_adj_2917)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_5_i31_3_lut.init = 16'hcaca;
    LUT4 i12141_3_lut (.A(index_i[3]), .B(index_i[1]), .C(index_i[0]), 
         .Z(n14825)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i12141_3_lut.init = 16'hecec;
    PFUMX i19199 (.BLUT(n21634), .ALUT(n21635), .C0(index_i[5]), .Z(n21636));
    LUT4 n26276_bdd_3_lut (.A(n27196), .B(n26272), .C(index_i[7]), .Z(n26277)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n26276_bdd_3_lut.init = 16'hcaca;
    LUT4 i9478_3_lut (.A(n12038), .B(n27017), .C(index_i[3]), .Z(n12039)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9478_3_lut.init = 16'hcaca;
    PFUMX i19202 (.BLUT(n21637), .ALUT(n21638), .C0(index_i[5]), .Z(n21639));
    PFUMX i19205 (.BLUT(n21640), .ALUT(n21641), .C0(index_i[5]), .Z(n21642));
    LUT4 mux_198_Mux_5_i124_3_lut (.A(n645), .B(n26971), .C(index_i[3]), 
         .Z(n124_adj_2911)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_5_i124_3_lut.init = 16'hcaca;
    L6MUX21 i23385 (.D0(n25122), .D1(n25120), .SD(index_i[7]), .Z(n25123));
    L6MUX21 i24569 (.D0(n26519), .D1(n26516), .SD(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2126[4]));
    PFUMX i24567 (.BLUT(n26518), .ALUT(n26517), .C0(index_i[8]), .Z(n26519));
    PFUMX i24564 (.BLUT(n26515), .ALUT(n23140), .C0(index_i[8]), .Z(n26516));
    LUT4 n25034_bdd_3_lut_25709 (.A(n25034), .B(n23347), .C(index_i[6]), 
         .Z(n26324)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n25034_bdd_3_lut_25709.init = 16'hcaca;
    LUT4 mux_198_Mux_1_i924_3_lut (.A(n316_adj_2790), .B(n412_adj_2887), 
         .C(index_i[4]), .Z(n924_adj_2918)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_1_i924_3_lut.init = 16'hcaca;
    LUT4 i19692_3_lut (.A(n26957), .B(n27007), .C(index_i[3]), .Z(n22129)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19692_3_lut.init = 16'hcaca;
    PFUMX i19208 (.BLUT(n21643), .ALUT(n21644), .C0(index_i[5]), .Z(n21645));
    LUT4 i21807_3_lut (.A(n21895), .B(n21896), .C(index_i[4]), .Z(n21897)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21807_3_lut.init = 16'hcaca;
    PFUMX i19211 (.BLUT(n21646), .ALUT(n21647), .C0(index_i[5]), .Z(n21648));
    PFUMX i23383 (.BLUT(n25121), .ALUT(n21581), .C0(index_i[6]), .Z(n25122));
    LUT4 mux_198_Mux_5_i700_3_lut (.A(n460_adj_2905), .B(n27010), .C(index_i[4]), 
         .Z(n700_adj_2919)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_5_i700_3_lut.init = 16'hcaca;
    PFUMX i19214 (.BLUT(n21649), .ALUT(n21650), .C0(index_i[5]), .Z(n21651));
    PFUMX i23381 (.BLUT(n25119), .ALUT(n24771), .C0(index_i[4]), .Z(n25120));
    LUT4 n25034_bdd_3_lut_24425 (.A(n23348), .B(n25052), .C(index_i[6]), 
         .Z(n26323)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n25034_bdd_3_lut_24425.init = 16'hcaca;
    LUT4 n25028_bdd_3_lut (.A(n25028), .B(n23343), .C(index_i[6]), .Z(n26326)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n25028_bdd_3_lut.init = 16'hcaca;
    LUT4 i9364_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n11925)) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B ((D)+!C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9364_3_lut_4_lut_4_lut.init = 16'hcdad;
    LUT4 mux_198_Mux_6_i731_3_lut (.A(n26948), .B(n26950), .C(index_i[3]), 
         .Z(n731_adj_2920)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_6_i731_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_1_i349_3_lut (.A(n506_adj_2866), .B(n348_adj_2921), 
         .C(index_i[4]), .Z(n349)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_1_i349_3_lut.init = 16'hcaca;
    LUT4 i21824_3_lut (.A(n21871), .B(n21872), .C(index_i[4]), .Z(n21873)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21824_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_1_i94_3_lut (.A(index_i[0]), .B(n93_adj_2922), .C(index_i[4]), 
         .Z(n94_adj_2923)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_1_i94_3_lut.init = 16'hcaca;
    LUT4 i20901_3_lut_4_lut_4_lut (.A(n26814), .B(index_i[5]), .C(index_i[4]), 
         .D(n26780), .Z(n23357)) /* synthesis lut_function=(A (B+(C (D)))+!A (B+((D)+!C))) */ ;
    defparam i20901_3_lut_4_lut_4_lut.init = 16'hfdcd;
    LUT4 mux_198_Mux_6_i891_3_lut (.A(n301), .B(n890_adj_2879), .C(index_i[4]), 
         .Z(n891_adj_2924)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_6_i891_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_6_i828_4_lut (.A(n812_adj_2925), .B(n13955), .C(index_i[4]), 
         .D(index_i[2]), .Z(n828_adj_2926)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_6_i828_4_lut.init = 16'hfaca;
    LUT4 mux_198_Mux_6_i797_3_lut (.A(n781_adj_2863), .B(n26722), .C(index_i[4]), 
         .Z(n797_adj_2927)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_6_i797_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_4_i15_3_lut (.A(n29466), .B(n588), .C(index_i[3]), 
         .Z(n15_adj_2871)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_4_i15_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_6_i669_3_lut (.A(n653_adj_2913), .B(n668_adj_2928), 
         .C(index_i[4]), .Z(n669_adj_2929)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_6_i669_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_6_i542_3_lut (.A(n26956), .B(n541_adj_2833), .C(index_i[4]), 
         .Z(n542_adj_2930)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_6_i542_3_lut.init = 16'hcaca;
    PFUMX i20421 (.BLUT(n22873), .ALUT(n22874), .C0(index_i[5]), .Z(n22877));
    LUT4 mux_198_Mux_6_i252_4_lut (.A(index_i[2]), .B(n251_adj_2825), .C(index_i[4]), 
         .D(n11191), .Z(n252_adj_2931)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_6_i252_4_lut.init = 16'hc5ca;
    LUT4 i22220_3_lut (.A(n25714), .B(n252_adj_2931), .C(index_i[5]), 
         .Z(n23345)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22220_3_lut.init = 16'hcaca;
    PFUMX i20422 (.BLUT(n22875), .ALUT(n22876), .C0(index_i[5]), .Z(n22878));
    PFUMX i20428 (.BLUT(n22880), .ALUT(n22881), .C0(index_i[5]), .Z(n22884));
    PFUMX i20429 (.BLUT(n22882), .ALUT(n22883), .C0(index_i[5]), .Z(n22885));
    LUT4 i12341_2_lut_3_lut_4_lut (.A(n26778), .B(index_i[4]), .C(index_i[6]), 
         .D(index_i[5]), .Z(n15034)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i12341_2_lut_3_lut_4_lut.init = 16'hfef0;
    LUT4 mux_198_Mux_10_i574_4_lut_4_lut (.A(n26778), .B(index_i[4]), .C(index_i[5]), 
         .D(n26755), .Z(n574_adj_2822)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_10_i574_4_lut_4_lut.init = 16'h1f1c;
    LUT4 mux_198_Mux_2_i284_rep_794 (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .Z(n29467)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_2_i284_rep_794.init = 16'h4d4d;
    LUT4 mux_198_Mux_4_i61_3_lut (.A(n26958), .B(n26942), .C(index_i[3]), 
         .Z(n61)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_4_i61_3_lut.init = 16'hcaca;
    LUT4 n24775_bdd_3_lut (.A(n24775), .B(n24772), .C(index_i[3]), .Z(n25119)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n24775_bdd_3_lut.init = 16'hcaca;
    LUT4 i22490_3_lut_4_lut (.A(n26878), .B(n19786), .C(index_i[8]), .D(n766), 
         .Z(n21527)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i22490_3_lut_4_lut.init = 16'hefe0;
    LUT4 mux_198_Mux_7_i892_3_lut (.A(n62), .B(n891), .C(index_i[5]), 
         .Z(n892_adj_2823)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_7_i892_3_lut.init = 16'hcaca;
    LUT4 n21581_bdd_3_lut_25627 (.A(n62), .B(n27170), .C(index_i[5]), 
         .Z(n25121)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n21581_bdd_3_lut_25627.init = 16'hacac;
    LUT4 i19213_3_lut (.A(n747), .B(n762), .C(index_i[4]), .Z(n21650)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19213_3_lut.init = 16'hcaca;
    LUT4 i19212_3_lut (.A(n716_adj_2932), .B(n14798), .C(index_i[4]), 
         .Z(n21649)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19212_3_lut.init = 16'hcaca;
    LUT4 i19210_3_lut (.A(n93_adj_2933), .B(n699), .C(index_i[4]), .Z(n21647)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19210_3_lut.init = 16'hcaca;
    LUT4 i19209_3_lut (.A(n653_adj_2808), .B(n26750), .C(index_i[4]), 
         .Z(n21646)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19209_3_lut.init = 16'hcaca;
    LUT4 i8612_4_lut_4_lut (.A(index_i[3]), .B(index_i[0]), .C(index_i[1]), 
         .D(index_i[2]), .Z(n11109)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (D)+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i8612_4_lut_4_lut.init = 16'h0bf4;
    LUT4 mux_198_Mux_0_i30_3_lut (.A(n26970), .B(n26949), .C(index_i[3]), 
         .Z(n30_adj_2934)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i30_3_lut.init = 16'hcaca;
    LUT4 n23140_bdd_3_lut (.A(n23133), .B(n23134), .C(index_i[7]), .Z(n26515)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n23140_bdd_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_0_i220_3_lut (.A(n26950), .B(n27011), .C(index_i[3]), 
         .Z(n220)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i220_3_lut.init = 16'hcaca;
    LUT4 n25361_bdd_3_lut_24566 (.A(n25361), .B(n23131), .C(index_i[7]), 
         .Z(n26517)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n25361_bdd_3_lut_24566.init = 16'hacac;
    LUT4 n25361_bdd_3_lut_25635 (.A(n23129), .B(n23130), .C(index_i[7]), 
         .Z(n26518)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n25361_bdd_3_lut_25635.init = 16'hcaca;
    LUT4 i19203_3_lut (.A(n526_adj_2935), .B(n15_adj_2936), .C(index_i[4]), 
         .Z(n21640)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19203_3_lut.init = 16'hcaca;
    LUT4 i19200_3_lut (.A(n397_adj_2937), .B(n475_adj_2807), .C(index_i[4]), 
         .Z(n21637)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19200_3_lut.init = 16'hcaca;
    L6MUX21 i20887 (.D0(n21492), .D1(n21495), .SD(index_i[5]), .Z(n23343));
    LUT4 i19198_3_lut (.A(n348_adj_2938), .B(n443_adj_2829), .C(index_i[4]), 
         .Z(n21635)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19198_3_lut.init = 16'hcaca;
    LUT4 i19197_3_lut (.A(n397_adj_2937), .B(n731_adj_2920), .C(index_i[4]), 
         .Z(n21634)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19197_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_7_i333_3_lut (.A(n27039), .B(n645), .C(index_i[3]), 
         .Z(n333)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_7_i333_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_7_i348_3_lut (.A(n26972), .B(n27042), .C(index_i[3]), 
         .Z(n348_adj_2938)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_7_i348_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_7_i397_3_lut (.A(n26972), .B(n27039), .C(index_i[3]), 
         .Z(n397_adj_2937)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_7_i397_3_lut.init = 16'hcaca;
    L6MUX21 i20891 (.D0(n21501), .D1(n17791), .SD(index_i[5]), .Z(n23347));
    LUT4 i19195_3_lut (.A(n364_adj_2939), .B(n379_adj_2898), .C(index_i[4]), 
         .Z(n21632)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19195_3_lut.init = 16'hcaca;
    LUT4 i19194_3_lut (.A(n333), .B(n348_adj_2938), .C(index_i[4]), .Z(n21631)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19194_3_lut.init = 16'hcaca;
    L6MUX21 i20892 (.D0(n21504), .D1(n11988), .SD(index_i[5]), .Z(n23348));
    LUT4 i1_4_lut (.A(index_i[6]), .B(n26845), .C(index_i[5]), .D(index_i[4]), 
         .Z(n20356)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i1_4_lut.init = 16'hfffe;
    L6MUX21 i20486 (.D0(n22940), .D1(n22941), .SD(index_i[5]), .Z(n22942));
    PFUMX i20894 (.BLUT(n542_adj_2930), .ALUT(n573_adj_2940), .C0(index_i[5]), 
          .Z(n23350));
    PFUMX i20895 (.BLUT(n605_adj_2941), .ALUT(n636_adj_2942), .C0(index_i[5]), 
          .Z(n23351));
    PFUMX i20896 (.BLUT(n669_adj_2929), .ALUT(n700_adj_2943), .C0(index_i[5]), 
          .Z(n23352));
    PFUMX i20897 (.BLUT(n732_adj_2944), .ALUT(n21510), .C0(index_i[5]), 
          .Z(n23353));
    PFUMX i20898 (.BLUT(n797_adj_2927), .ALUT(n828_adj_2926), .C0(index_i[5]), 
          .Z(n23354));
    LUT4 mux_198_Mux_5_i731_3_lut (.A(n27007), .B(n29479), .C(index_i[3]), 
         .Z(n731_adj_2895)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_5_i731_3_lut.init = 16'hcaca;
    PFUMX i20899 (.BLUT(n860_adj_2945), .ALUT(n891_adj_2924), .C0(index_i[5]), 
          .Z(n23355));
    L6MUX21 i20493 (.D0(n22947), .D1(n22948), .SD(index_i[5]), .Z(n22949));
    LUT4 i19086_3_lut (.A(n325), .B(n27007), .C(index_i[3]), .Z(n21523)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19086_3_lut.init = 16'hcaca;
    LUT4 i20771_3_lut (.A(n26965), .B(n251), .C(index_i[4]), .Z(n23227)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20771_3_lut.init = 16'hcaca;
    L6MUX21 i20500 (.D0(n22954), .D1(n22955), .SD(index_i[5]), .Z(n22956));
    PFUMX i20918 (.BLUT(n94_adj_2923), .ALUT(n21864), .C0(index_i[5]), 
          .Z(n23374));
    LUT4 i20764_3_lut (.A(n15_adj_2936), .B(n30_adj_2934), .C(index_i[4]), 
         .Z(n23220)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20764_3_lut.init = 16'hcaca;
    L6MUX21 i20919 (.D0(n21867), .D1(n21870), .SD(index_i[5]), .Z(n23375));
    LUT4 n25138_bdd_3_lut (.A(n28291), .B(n25133), .C(index_i[4]), .Z(n25139)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n25138_bdd_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_4_i158_3_lut (.A(n142_adj_2946), .B(n157_adj_2903), 
         .C(index_i[4]), .Z(n158_adj_2893)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_4_i158_3_lut.init = 16'hcaca;
    LUT4 i19191_3_lut_4_lut_4_lut (.A(n26879), .B(index_i[4]), .C(index_i[3]), 
         .D(n26837), .Z(n21628)) /* synthesis lut_function=(A (B (C)+!B !(C+!(D)))+!A (B (C)+!B (C+(D)))) */ ;
    defparam i19191_3_lut_4_lut_4_lut.init = 16'hd3d0;
    L6MUX21 i20507 (.D0(n22961), .D1(n22962), .SD(index_i[5]), .Z(n22963));
    LUT4 i20488_3_lut_3_lut (.A(n27039), .B(index_i[3]), .C(n29496), .Z(n22944)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam i20488_3_lut_3_lut.init = 16'h7474;
    PFUMX i20921 (.BLUT(n21873), .ALUT(n317_adj_2947), .C0(index_i[5]), 
          .Z(n23377));
    PFUMX i20922 (.BLUT(n349), .ALUT(n21876), .C0(index_i[5]), .Z(n23378));
    LUT4 n26237_bdd_3_lut_3_lut (.A(n1021), .B(index_i[8]), .C(n26237), 
         .Z(n26238)) /* synthesis lut_function=(A (B+(C))+!A !(B+!(C))) */ ;
    defparam n26237_bdd_3_lut_3_lut.init = 16'hb8b8;
    L6MUX21 i20923 (.D0(n21879), .D1(n21882), .SD(index_i[5]), .Z(n23379));
    LUT4 mux_198_Mux_7_i364_3_lut_3_lut (.A(n27039), .B(index_i[3]), .C(n26972), 
         .Z(n364_adj_2939)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;
    defparam mux_198_Mux_7_i364_3_lut_3_lut.init = 16'hd1d1;
    LUT4 mux_198_Mux_4_i668_3_lut_3_lut (.A(n27039), .B(index_i[3]), .C(n29496), 
         .Z(n668_adj_2864)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;
    defparam mux_198_Mux_4_i668_3_lut_3_lut.init = 16'hd1d1;
    L6MUX21 i20924 (.D0(n21885), .D1(n21888), .SD(index_i[5]), .Z(n23380));
    LUT4 mux_198_Mux_7_i379_3_lut_3_lut (.A(n27039), .B(index_i[3]), .C(n27042), 
         .Z(n379_adj_2898)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam mux_198_Mux_7_i379_3_lut_3_lut.init = 16'h7474;
    LUT4 i19186_3_lut (.A(n491_adj_2948), .B(n506_adj_2866), .C(index_i[4]), 
         .Z(n21623)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19186_3_lut.init = 16'hcaca;
    LUT4 i19360_3_lut_3_lut (.A(n27039), .B(index_i[3]), .C(n1001), .Z(n21797)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam i19360_3_lut_3_lut.init = 16'h7474;
    LUT4 i19185_3_lut (.A(n460_adj_2817), .B(n475_adj_2880), .C(index_i[4]), 
         .Z(n21622)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19185_3_lut.init = 16'hcaca;
    PFUMX i24438 (.BLUT(n26339), .ALUT(n29496), .C0(index_i[3]), .Z(n26340));
    LUT4 i19084_3_lut (.A(n27019), .B(n29479), .C(index_i[3]), .Z(n21521)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19084_3_lut.init = 16'hcaca;
    LUT4 i19083_3_lut (.A(n27013), .B(n29482), .C(index_i[3]), .Z(n21520)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19083_3_lut.init = 16'hcaca;
    L6MUX21 i24430 (.D0(n26327), .D1(n26325), .SD(index_i[8]), .Z(n26328));
    LUT4 i11619_3_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .Z(n11191)) /* synthesis lut_function=(!((B (C))+!A)) */ ;
    defparam i11619_3_lut.init = 16'h2a2a;
    PFUMX i24428 (.BLUT(n26326), .ALUT(n23359), .C0(index_i[7]), .Z(n26327));
    L6MUX21 i20926 (.D0(n21894), .D1(n636), .SD(index_i[5]), .Z(n23382));
    LUT4 i19183_3_lut (.A(n251_adj_2789), .B(n443_adj_2788), .C(index_i[4]), 
         .Z(n21620)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19183_3_lut.init = 16'hcaca;
    LUT4 i19182_3_lut (.A(n460_adj_2817), .B(n14798), .C(index_i[4]), 
         .Z(n21619)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;
    defparam i19182_3_lut.init = 16'h3a3a;
    LUT4 mux_198_Mux_6_i653_3_lut (.A(n27014), .B(n85), .C(index_i[3]), 
         .Z(n653_adj_2913)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_6_i653_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_6_i668_3_lut (.A(n108), .B(n27041), .C(index_i[3]), 
         .Z(n668_adj_2928)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_6_i668_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_6_i684_3_lut (.A(n645), .B(n29496), .C(index_i[3]), 
         .Z(n684_adj_2949)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_6_i684_3_lut.init = 16'hcaca;
    LUT4 i19443_3_lut_3_lut_4_lut (.A(index_i[0]), .B(n27050), .C(index_i[3]), 
         .D(n26880), .Z(n21880)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A !(C+(D))) */ ;
    defparam i19443_3_lut_3_lut_4_lut.init = 16'h808f;
    PFUMX i24426 (.BLUT(n26324), .ALUT(n26323), .C0(index_i[7]), .Z(n26325));
    PFUMX i20927 (.BLUT(n21897), .ALUT(n700_adj_2796), .C0(index_i[5]), 
          .Z(n23383));
    LUT4 i11099_2_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n844)) /* synthesis lut_function=(A (B+!(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11099_2_lut_3_lut_4_lut.init = 16'h9ff9;
    LUT4 i19081_3_lut (.A(n29467), .B(n29482), .C(index_i[3]), .Z(n21518)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19081_3_lut.init = 16'hcaca;
    LUT4 i19410_3_lut_3_lut_4_lut (.A(index_i[0]), .B(n27050), .C(n26880), 
         .D(index_i[3]), .Z(n21847)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(C+(D)))) */ ;
    defparam i19410_3_lut_3_lut_4_lut.init = 16'h77f0;
    LUT4 i22430_3_lut_rep_392_4_lut (.A(n26844), .B(index_i[5]), .C(index_i[8]), 
         .D(n1021), .Z(n26715)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i22430_3_lut_rep_392_4_lut.init = 16'hf808;
    LUT4 i11181_3_lut_4_lut (.A(index_i[0]), .B(n27050), .C(n26968), .D(index_i[5]), 
         .Z(n318)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (C (D))) */ ;
    defparam i11181_3_lut_4_lut.init = 16'hf800;
    LUT4 i17561_4_lut (.A(n27049), .B(n892_adj_2868), .C(index_i[6]), 
         .D(index_i[5]), .Z(n19848)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D))))) */ ;
    defparam i17561_4_lut.init = 16'h3a35;
    LUT4 n699_bdd_4_lut_4_lut_4_lut (.A(index_i[0]), .B(n27050), .C(index_i[4]), 
         .D(index_i[3]), .Z(n24684)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (D))+!A (B (C (D)+!C !(D))+!B (D)))) */ ;
    defparam n699_bdd_4_lut_4_lut_4_lut.init = 16'h0c73;
    PFUMX i19694 (.BLUT(n22129), .ALUT(n22130), .C0(index_i[4]), .Z(n22131));
    L6MUX21 i20929 (.D0(n21900), .D1(n21903), .SD(index_i[5]), .Z(n23385));
    LUT4 mux_198_Mux_1_i986_3_lut (.A(n26972), .B(n27011), .C(index_i[3]), 
         .Z(n986_adj_2950)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_1_i986_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_6_i15_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n15)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C))+!A !(B (C+!(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_6_i15_3_lut_4_lut_4_lut.init = 16'h5ad6;
    LUT4 i9379_4_lut_4_lut (.A(n27053), .B(index_i[1]), .C(index_i[3]), 
         .D(n20685), .Z(n11940)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A (B (C)+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9379_4_lut_4_lut.init = 16'h0e3e;
    PFUMX i20931 (.BLUT(n924_adj_2918), .ALUT(n21909), .C0(index_i[5]), 
          .Z(n23387));
    LUT4 i19173_3_lut (.A(n301), .B(n93_adj_2933), .C(index_i[4]), .Z(n21610)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19173_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_0_i572_3_lut_4_lut (.A(n27053), .B(index_i[1]), .C(index_i[3]), 
         .D(n29482), .Z(n572)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i572_3_lut_4_lut.init = 16'hefe0;
    LUT4 index_i_3__bdd_3_lut_22891_3_lut_4_lut (.A(n27053), .B(index_i[1]), 
         .C(index_i[4]), .D(index_i[3]), .Z(n24545)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam index_i_3__bdd_3_lut_22891_3_lut_4_lut.init = 16'hf10f;
    LUT4 i11161_2_lut_rep_416_3_lut_4_lut (.A(n27053), .B(index_i[1]), .C(index_i[4]), 
         .D(index_i[3]), .Z(n26739)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11161_2_lut_rep_416_3_lut_4_lut.init = 16'hfef0;
    LUT4 i19170_3_lut (.A(n15_adj_2873), .B(n526_adj_2850), .C(index_i[4]), 
         .Z(n21607)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19170_3_lut.init = 16'hcaca;
    PFUMX i20932 (.BLUT(n987), .ALUT(n21921), .C0(index_i[5]), .Z(n23388));
    LUT4 i19188_4_lut_4_lut_3_lut_4_lut (.A(n27053), .B(index_i[1]), .C(index_i[4]), 
         .D(index_i[3]), .Z(n21625)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19188_4_lut_4_lut_3_lut_4_lut.init = 16'h11ef;
    LUT4 i9380_3_lut_4_lut_4_lut (.A(n27052), .B(index_i[3]), .C(index_i[5]), 
         .D(n26879), .Z(n11941)) /* synthesis lut_function=(A (B+(C (D)))+!A (B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9380_3_lut_4_lut_4_lut.init = 16'hf8c8;
    LUT4 i20419_3_lut_3_lut_4_lut_4_lut (.A(n27052), .B(index_i[3]), .C(index_i[4]), 
         .D(n26837), .Z(n22875)) /* synthesis lut_function=(!(A (B (C)+!B ((D)+!C))+!A (B+((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20419_3_lut_3_lut_4_lut_4_lut.init = 16'h0838;
    LUT4 mux_198_Mux_3_i747_3_lut (.A(n26957), .B(n404), .C(index_i[3]), 
         .Z(n747_adj_2853)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_3_i747_3_lut.init = 16'hcaca;
    LUT4 index_i_3__bdd_3_lut_22918_4_lut_4_lut (.A(n27052), .B(index_i[3]), 
         .C(index_i[4]), .D(n26839), .Z(n24546)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C))+!A !(B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam index_i_3__bdd_3_lut_22918_4_lut_4_lut.init = 16'h838f;
    LUT4 mux_198_Mux_5_i15_3_lut (.A(n27012), .B(n29484), .C(index_i[3]), 
         .Z(n15_adj_2900)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_5_i15_3_lut.init = 16'hcaca;
    LUT4 i11152_2_lut_3_lut_4_lut (.A(n26837), .B(n26968), .C(index_i[6]), 
         .D(index_i[5]), .Z(n254)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i11152_2_lut_3_lut_4_lut.init = 16'hfef0;
    PFUMX i20917 (.BLUT(n12039), .ALUT(n62_adj_2951), .C0(index_i[5]), 
          .Z(n23373));
    LUT4 i19077_3_lut (.A(n26957), .B(n29482), .C(index_i[3]), .Z(n21514)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19077_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_5_i397_3_lut (.A(n27019), .B(n332), .C(index_i[3]), 
         .Z(n397_adj_2907)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_5_i397_3_lut.init = 16'hcaca;
    PFUMX i24391 (.BLUT(n26277), .ALUT(n1022), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2126[12]));
    LUT4 mux_198_Mux_5_i506_3_lut (.A(n29480), .B(n29466), .C(index_i[3]), 
         .Z(n506_adj_2859)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_5_i506_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_5_i859_3_lut (.A(n141), .B(n27012), .C(index_i[3]), 
         .Z(n859_adj_2901)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_5_i859_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_5_i875_3_lut (.A(n645), .B(n26972), .C(index_i[3]), 
         .Z(n875_adj_2897)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_5_i875_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_0_i923_3_lut (.A(n26948), .B(n27042), .C(index_i[3]), 
         .Z(n923)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i923_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_6_i732_3_lut_4_lut (.A(n27039), .B(index_i[3]), .C(index_i[4]), 
         .D(n731_adj_2920), .Z(n732_adj_2944)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_6_i732_3_lut_4_lut.init = 16'hf909;
    LUT4 mux_198_Mux_13_i511_4_lut_4_lut (.A(n26712), .B(index_i[7]), .C(index_i[8]), 
         .D(n254), .Z(n511)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (B (C+!(D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_13_i511_4_lut_4_lut.init = 16'h1c10;
    PFUMX i23320 (.BLUT(n25055), .ALUT(n26941), .C0(index_i[5]), .Z(n25056));
    LUT4 index_i_8__bdd_3_lut_then_4_lut (.A(index_i[4]), .B(index_i[6]), 
         .C(index_i[5]), .D(n26760), .Z(n27195)) /* synthesis lut_function=(!(A (B (C+(D)))+!A (B (C)))) */ ;
    defparam index_i_8__bdd_3_lut_then_4_lut.init = 16'h373f;
    PFUMX i20567 (.BLUT(n31_adj_2917), .ALUT(n21513), .C0(index_i[5]), 
          .Z(n23023));
    LUT4 i20425_3_lut_4_lut_3_lut (.A(index_i[3]), .B(index_i[4]), .C(n26839), 
         .Z(n22881)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20425_3_lut_4_lut_3_lut.init = 16'h6464;
    PFUMX i20568 (.BLUT(n94_adj_2915), .ALUT(n125_adj_2912), .C0(index_i[5]), 
          .Z(n23024));
    PFUMX i24387 (.BLUT(n254_adj_2952), .ALUT(n26271), .C0(index_i[8]), 
          .Z(n26272));
    LUT4 mux_198_Mux_6_i700_3_lut_4_lut (.A(n27039), .B(index_i[3]), .C(index_i[4]), 
         .D(n684_adj_2949), .Z(n700_adj_2943)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_6_i700_3_lut_4_lut.init = 16'h9f90;
    PFUMX i20569 (.BLUT(n17827), .ALUT(n14449), .C0(index_i[5]), .Z(n23025));
    LUT4 i20044_3_lut_4_lut_4_lut (.A(n26845), .B(index_i[4]), .C(index_i[5]), 
         .D(n26760), .Z(n22500)) /* synthesis lut_function=(A ((C+!(D))+!B)+!A (B (C+!(D))+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20044_3_lut_4_lut_4_lut.init = 16'he3ef;
    L6MUX21 i20571 (.D0(n21516), .D1(n21519), .SD(index_i[5]), .Z(n23027));
    PFUMX i23318 (.BLUT(n26955), .ALUT(n25053), .C0(index_i[2]), .Z(n25054));
    L6MUX21 i20572 (.D0(n21522), .D1(n21525), .SD(index_i[5]), .Z(n23028));
    PFUMX i20573 (.BLUT(n413_adj_2908), .ALUT(n444), .C0(index_i[5]), 
          .Z(n23029));
    L6MUX21 i23316 (.D0(n25051), .D1(n25048), .SD(index_i[5]), .Z(n25052));
    PFUMX i20574 (.BLUT(n476_adj_2906), .ALUT(n507), .C0(index_i[5]), 
          .Z(n23030));
    LUT4 index_i_8__bdd_3_lut_else_4_lut (.A(n26838), .B(index_i[4]), .C(index_i[6]), 
         .D(index_i[5]), .Z(n27194)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;
    defparam index_i_8__bdd_3_lut_else_4_lut.init = 16'hf080;
    PFUMX i23314 (.BLUT(n25050), .ALUT(n25049), .C0(index_i[4]), .Z(n25051));
    PFUMX i20575 (.BLUT(n17794), .ALUT(n573_adj_2953), .C0(index_i[5]), 
          .Z(n23031));
    LUT4 i19482_3_lut (.A(n29480), .B(n26964), .C(index_i[3]), .Z(n21919)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19482_3_lut.init = 16'hcaca;
    LUT4 i21786_3_lut (.A(n21919), .B(n21920), .C(index_i[4]), .Z(n21921)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21786_3_lut.init = 16'hcaca;
    PFUMX i20576 (.BLUT(n605_adj_2954), .ALUT(n636_adj_2904), .C0(index_i[5]), 
          .Z(n23032));
    PFUMX i20577 (.BLUT(n22125), .ALUT(n700_adj_2919), .C0(index_i[5]), 
          .Z(n23033));
    PFUMX i23311 (.BLUT(n25047), .ALUT(n21506), .C0(index_i[4]), .Z(n25048));
    L6MUX21 i20578 (.D0(n732_adj_2896), .D1(n22131), .SD(index_i[5]), 
            .Z(n23034));
    PFUMX i20579 (.BLUT(n797_adj_2955), .ALUT(n828_adj_2956), .C0(index_i[5]), 
          .Z(n23035));
    LUT4 i22109_3_lut (.A(n28755), .B(n27226), .C(index_i[5]), .Z(n23127)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22109_3_lut.init = 16'hcaca;
    PFUMX i20580 (.BLUT(n860_adj_2902), .ALUT(n891_adj_2899), .C0(index_i[5]), 
          .Z(n23036));
    LUT4 i22114_3_lut (.A(n542_adj_2867), .B(n573), .C(index_i[5]), .Z(n23121)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22114_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_12_i254_4_lut (.A(n26735), .B(n20563), .C(index_i[6]), 
         .D(n26839), .Z(n254_adj_2952)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_12_i254_4_lut.init = 16'hca0a;
    LUT4 i19470_3_lut (.A(n1001), .B(n588), .C(index_i[3]), .Z(n21907)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19470_3_lut.init = 16'hcaca;
    LUT4 i21793_3_lut (.A(n21907), .B(n21908), .C(index_i[4]), .Z(n21909)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21793_3_lut.init = 16'hcaca;
    LUT4 i22443_3_lut (.A(n19848), .B(n20356), .C(index_i[7]), .Z(n22547)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22443_3_lut.init = 16'hcaca;
    PFUMX i24363 (.BLUT(n26240), .ALUT(n26238), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2126[10]));
    L6MUX21 i23298 (.D0(n25033), .D1(n25031), .SD(index_i[5]), .Z(n25034));
    LUT4 i11100_4_lut_4_lut (.A(index_i[3]), .B(index_i[2]), .C(index_i[0]), 
         .D(index_i[1]), .Z(n875)) /* synthesis lut_function=((B (C)+!B (D))+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11100_4_lut_4_lut.init = 16'hf7d5;
    PFUMX i23296 (.BLUT(n25032), .ALUT(n285), .C0(index_i[4]), .Z(n25033));
    LUT4 mux_198_Mux_4_i270_3_lut (.A(n27017), .B(n29480), .C(index_i[3]), 
         .Z(n270_adj_2870)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_4_i270_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_1_i987_3_lut_4_lut_4_lut (.A(index_i[3]), .B(n986_adj_2950), 
         .C(index_i[4]), .D(n26950), .Z(n987)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_1_i987_3_lut_4_lut_4_lut.init = 16'hc5c0;
    PFUMX i23294 (.BLUT(n25030), .ALUT(n25029), .C0(index_i[4]), .Z(n25031));
    LUT4 mux_198_Mux_4_i348_3_lut (.A(n27005), .B(n27015), .C(index_i[3]), 
         .Z(n348_adj_2957)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_4_i348_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_2_i221_4_lut_4_lut (.A(index_i[3]), .B(index_i[4]), 
         .C(n26879), .D(n26755), .Z(n221_adj_2958)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (B+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_2_i221_4_lut_4_lut.init = 16'hf7c4;
    LUT4 i19216_4_lut_3_lut (.A(index_i[3]), .B(index_i[4]), .C(n26879), 
         .Z(n21653)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19216_4_lut_3_lut.init = 16'h6565;
    LUT4 i9381_3_lut_3_lut (.A(index_i[3]), .B(index_i[4]), .C(n11941), 
         .Z(n11942)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9381_3_lut_3_lut.init = 16'h7474;
    LUT4 mux_198_Mux_4_i684_3_lut (.A(n85), .B(n108), .C(index_i[3]), 
         .Z(n684_adj_2861)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_4_i684_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_3_i796_3_lut_3_lut (.A(index_i[4]), .B(n731_adj_2920), 
         .C(index_i[2]), .Z(n796_adj_2959)) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam mux_198_Mux_3_i796_3_lut_3_lut.init = 16'he4e4;
    LUT4 i20071_4_lut_4_lut (.A(index_i[4]), .B(index_i[5]), .C(n27164), 
         .D(n908_adj_2960), .Z(n22527)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam i20071_4_lut_4_lut.init = 16'hd1c0;
    L6MUX21 i23291 (.D0(n25027), .D1(n25024), .SD(index_i[5]), .Z(n25028));
    PFUMX i23289 (.BLUT(n15), .ALUT(n25025), .C0(index_i[4]), .Z(n25027));
    PFUMX i24361 (.BLUT(n21559), .ALUT(n26236), .C0(index_i[7]), .Z(n26237));
    PFUMX i23286 (.BLUT(n25023), .ALUT(n25022), .C0(index_i[4]), .Z(n25024));
    LUT4 i22365_3_lut (.A(n22527), .B(n26047), .C(index_i[6]), .Z(n22536)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22365_3_lut.init = 16'hcaca;
    LUT4 i22718_2_lut (.A(index_i[5]), .B(index_i[4]), .Z(n22297)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i22718_2_lut.init = 16'heeee;
    LUT4 i1_3_lut (.A(index_i[0]), .B(index_i[4]), .C(index_i[2]), .Z(n20685)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i1_3_lut.init = 16'hfefe;
    LUT4 i12147_3_lut (.A(index_i[3]), .B(index_i[1]), .C(index_i[0]), 
         .Z(n14831)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i12147_3_lut.init = 16'hc8c8;
    LUT4 mux_198_Mux_3_i348_3_lut (.A(n27011), .B(n27013), .C(index_i[3]), 
         .Z(n348_adj_2961)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_3_i348_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_3_i908_3_lut (.A(n26964), .B(n26942), .C(index_i[3]), 
         .Z(n908_adj_2831)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_3_i908_3_lut.init = 16'hcaca;
    LUT4 i22168_3_lut (.A(n286), .B(n317), .C(index_i[5]), .Z(n22499)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22168_3_lut.init = 16'hcaca;
    LUT4 i19693_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n22130)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A (B (C (D)+!C !(D))+!B (D))) */ ;
    defparam i19693_3_lut_4_lut.init = 16'hd926;
    L6MUX21 i20995 (.D0(n23435), .D1(n23436), .SD(index_i[5]), .Z(n23451));
    L6MUX21 i20996 (.D0(n23437), .D1(n23438), .SD(index_i[5]), .Z(n23452));
    L6MUX21 i20997 (.D0(n23439), .D1(n23440), .SD(index_i[5]), .Z(n23453));
    LUT4 i12081_2_lut_rep_596 (.A(index_i[2]), .B(index_i[0]), .Z(n26919)) /* synthesis lut_function=(A (B)) */ ;
    defparam i12081_2_lut_rep_596.init = 16'h8888;
    LUT4 mux_198_Mux_3_i700_3_lut_4_lut (.A(index_i[4]), .B(index_i[3]), 
         .C(n684_adj_2962), .D(n29483), .Z(n700_adj_2963)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_3_i700_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i22686_2_lut_rep_597 (.A(index_i[4]), .B(index_i[3]), .Z(n26920)) /* synthesis lut_function=((B)+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i22686_2_lut_rep_597.init = 16'hdddd;
    L6MUX21 i20998 (.D0(n23441), .D1(n23442), .SD(index_i[5]), .Z(n23454));
    LUT4 mux_198_Mux_0_i716_3_lut (.A(n26962), .B(n26942), .C(index_i[3]), 
         .Z(n716_adj_2812)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i716_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_3_i797_3_lut_4_lut (.A(index_i[4]), .B(index_i[3]), 
         .C(n796_adj_2959), .D(n70), .Z(n797)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_3_i797_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i20941_3_lut (.A(n23389), .B(n23390), .C(index_i[7]), .Z(n23397)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20941_3_lut.init = 16'hcaca;
    LUT4 i20934_3_lut (.A(n23375), .B(n25755), .C(index_i[6]), .Z(n23390)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20934_3_lut.init = 16'hcaca;
    LUT4 i20943_3_lut (.A(n23393), .B(n23394), .C(index_i[7]), .Z(n23399)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20943_3_lut.init = 16'hcaca;
    LUT4 i20937_3_lut (.A(n25767), .B(n23382), .C(index_i[6]), .Z(n23393)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20937_3_lut.init = 16'hcaca;
    PFUMX i20059 (.BLUT(n158_adj_2892), .ALUT(n189_adj_2798), .C0(index_i[5]), 
          .Z(n22515));
    LUT4 i20714_3_lut (.A(n23164), .B(n23165), .C(index_i[7]), .Z(n23170)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20714_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_0_i653_3_lut (.A(n645), .B(n29480), .C(index_i[3]), 
         .Z(n653)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i653_3_lut.init = 16'hcaca;
    LUT4 i20709_3_lut (.A(n23154), .B(n23155), .C(index_i[6]), .Z(n23165)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20709_3_lut.init = 16'hcaca;
    PFUMX i20060 (.BLUT(n221_adj_2958), .ALUT(n21843), .C0(index_i[5]), 
          .Z(n22516));
    PFUMX i20061 (.BLUT(n286_adj_2890), .ALUT(n317_adj_2889), .C0(index_i[5]), 
          .Z(n22517));
    PFUMX i20062 (.BLUT(n349_adj_2964), .ALUT(n21846), .C0(index_i[5]), 
          .Z(n22518));
    LUT4 mux_198_Mux_0_i620_3_lut (.A(n26972), .B(n27017), .C(index_i[3]), 
         .Z(n620_adj_2806)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i620_3_lut.init = 16'hcaca;
    LUT4 i20588_3_lut (.A(n23033), .B(n23034), .C(index_i[6]), .Z(n23044)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20588_3_lut.init = 16'hcaca;
    LUT4 i20081_3_lut (.A(n25291), .B(n22530), .C(index_i[7]), .Z(n22537)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20081_3_lut.init = 16'hcaca;
    PFUMX i20063 (.BLUT(n413_adj_2888), .ALUT(n21849), .C0(index_i[5]), 
          .Z(n22519));
    LUT4 mux_198_Mux_0_i589_3_lut (.A(n27042), .B(n588), .C(index_i[3]), 
         .Z(n589)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i589_3_lut.init = 16'hcaca;
    L6MUX21 i20999 (.D0(n23443), .D1(n23444), .SD(index_i[5]), .Z(n23455));
    PFUMX i20064 (.BLUT(n21852), .ALUT(n507_adj_2965), .C0(index_i[5]), 
          .Z(n22520));
    LUT4 i20005_3_lut (.A(n22453), .B(n25139), .C(index_i[7]), .Z(n22461)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20005_3_lut.init = 16'hcaca;
    L6MUX21 i21000 (.D0(n23445), .D1(n23446), .SD(index_i[5]), .Z(n23456));
    PFUMX i20065 (.BLUT(n21855), .ALUT(n573_adj_2820), .C0(index_i[5]), 
          .Z(n22521));
    PFUMX i20066 (.BLUT(n605), .ALUT(n21858), .C0(index_i[5]), .Z(n22522));
    PFUMX i20067 (.BLUT(n669_adj_2884), .ALUT(n700_adj_2876), .C0(index_i[5]), 
          .Z(n22523));
    PFUMX i20068 (.BLUT(n732_adj_2882), .ALUT(n763_adj_2966), .C0(index_i[5]), 
          .Z(n22524));
    LUT4 mux_198_Mux_1_i732_3_lut (.A(n716), .B(n491), .C(index_i[4]), 
         .Z(n732)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_1_i732_3_lut.init = 16'hcaca;
    PFUMX i24759 (.BLUT(n27168), .ALUT(n27169), .C0(index_i[3]), .Z(n27170));
    LUT4 mux_198_Mux_0_i684_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n684_adj_2810)) /* synthesis lut_function=(!(A ((D)+!B)+!A !(B (D)+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i684_3_lut_4_lut_4_lut.init = 16'h5498;
    L6MUX21 i21001 (.D0(n23447), .D1(n23448), .SD(index_i[5]), .Z(n23457));
    LUT4 i22215_3_lut (.A(n924), .B(n955), .C(index_i[5]), .Z(n23356)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22215_3_lut.init = 16'hcaca;
    L6MUX21 i20070 (.D0(n860_adj_2848), .D1(n891_adj_2846), .SD(index_i[5]), 
            .Z(n22526));
    L6MUX21 i21002 (.D0(n23449), .D1(n23450), .SD(index_i[5]), .Z(n23458));
    LUT4 i19440_3_lut (.A(n26958), .B(n27007), .C(index_i[3]), .Z(n21877)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19440_3_lut.init = 16'hcaca;
    PFUMX mux_198_Mux_1_i891 (.BLUT(n882), .ALUT(n890_adj_2967), .C0(n26920), 
          .Z(n891_adj_2804)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 n627_bdd_3_lut_24196_4_lut_4_lut (.A(index_i[2]), .B(n85), .C(index_i[3]), 
         .D(n26969), .Z(n26033)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B ((D)+!C)+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n627_bdd_3_lut_24196_4_lut_4_lut.init = 16'h5c0c;
    LUT4 i21822_3_lut (.A(n21874), .B(n21875), .C(index_i[4]), .Z(n21876)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21822_3_lut.init = 16'hcaca;
    PFUMX i20688 (.BLUT(n31_adj_2878), .ALUT(n62_adj_2968), .C0(index_i[5]), 
          .Z(n23144));
    LUT4 mux_198_Mux_1_i317_3_lut (.A(n301_adj_2969), .B(n908_adj_2960), 
         .C(index_i[4]), .Z(n317_adj_2947)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_1_i317_3_lut.init = 16'hcaca;
    PFUMX i20657 (.BLUT(n31), .ALUT(n62_adj_2877), .C0(index_i[5]), .Z(n23113));
    LUT4 i22452_3_lut (.A(n25056), .B(n23345), .C(index_i[6]), .Z(n23359)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22452_3_lut.init = 16'hcaca;
    LUT4 i20140_3_lut (.A(n22594), .B(n22595), .C(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2126[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20140_3_lut.init = 16'hcaca;
    LUT4 i20916_3_lut (.A(n26328), .B(n23371), .C(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2126[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20916_3_lut.init = 16'hcaca;
    LUT4 i20915_3_lut (.A(n23368), .B(n23369), .C(index_i[8]), .Z(n23371)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20915_3_lut.init = 16'hcaca;
    LUT4 mux_195_i16_3_lut (.A(\quarter_wave_sample_register_q[15] ), .B(o_val_pipeline_i_0__15__N_2157[15]), 
         .C(phase_negation_i[1]), .Z(n1212[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam mux_195_i16_3_lut.init = 16'hcaca;
    LUT4 mux_195_i15_3_lut (.A(quarter_wave_sample_register_i[14]), .B(o_val_pipeline_i_0__15__N_2157[14]), 
         .C(phase_negation_i[1]), .Z(n1212[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam mux_195_i15_3_lut.init = 16'hcaca;
    LUT4 mux_195_i14_3_lut (.A(quarter_wave_sample_register_i[13]), .B(o_val_pipeline_i_0__15__N_2157[13]), 
         .C(phase_negation_i[1]), .Z(n1212[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam mux_195_i14_3_lut.init = 16'hcaca;
    LUT4 mux_195_i13_3_lut (.A(quarter_wave_sample_register_i[12]), .B(o_val_pipeline_i_0__15__N_2157[12]), 
         .C(phase_negation_i[1]), .Z(n1212[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam mux_195_i13_3_lut.init = 16'hcaca;
    LUT4 mux_195_i12_3_lut (.A(quarter_wave_sample_register_i[11]), .B(o_val_pipeline_i_0__15__N_2157[11]), 
         .C(phase_negation_i[1]), .Z(n1212[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam mux_195_i12_3_lut.init = 16'hcaca;
    LUT4 mux_195_i11_3_lut (.A(quarter_wave_sample_register_i[10]), .B(o_val_pipeline_i_0__15__N_2157[10]), 
         .C(phase_negation_i[1]), .Z(n1212[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam mux_195_i11_3_lut.init = 16'hcaca;
    LUT4 mux_195_i10_3_lut (.A(quarter_wave_sample_register_i[9]), .B(o_val_pipeline_i_0__15__N_2157[9]), 
         .C(phase_negation_i[1]), .Z(n1212[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam mux_195_i10_3_lut.init = 16'hcaca;
    LUT4 mux_195_i9_3_lut (.A(quarter_wave_sample_register_i[8]), .B(o_val_pipeline_i_0__15__N_2157[8]), 
         .C(phase_negation_i[1]), .Z(n1212[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam mux_195_i9_3_lut.init = 16'hcaca;
    LUT4 mux_195_i8_3_lut (.A(quarter_wave_sample_register_i[7]), .B(o_val_pipeline_i_0__15__N_2157[7]), 
         .C(phase_negation_i[1]), .Z(n1212[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam mux_195_i8_3_lut.init = 16'hcaca;
    L6MUX21 i24257 (.D0(n26092), .D1(n26090), .SD(index_i[5]), .Z(n26093));
    LUT4 mux_195_i7_3_lut (.A(quarter_wave_sample_register_i[6]), .B(o_val_pipeline_i_0__15__N_2157[6]), 
         .C(phase_negation_i[1]), .Z(n1212[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam mux_195_i7_3_lut.init = 16'hcaca;
    LUT4 n25285_bdd_3_lut (.A(n25285), .B(n476), .C(index_i[5]), .Z(n25286)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n25285_bdd_3_lut.init = 16'hcaca;
    LUT4 mux_195_i6_3_lut (.A(quarter_wave_sample_register_i[5]), .B(o_val_pipeline_i_0__15__N_2157[5]), 
         .C(phase_negation_i[1]), .Z(n1212[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam mux_195_i6_3_lut.init = 16'hcaca;
    LUT4 mux_195_i5_3_lut (.A(quarter_wave_sample_register_i[4]), .B(o_val_pipeline_i_0__15__N_2157[4]), 
         .C(phase_negation_i[1]), .Z(n1212[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam mux_195_i5_3_lut.init = 16'hcaca;
    PFUMX i24255 (.BLUT(n26091), .ALUT(n645), .C0(index_i[3]), .Z(n26092));
    LUT4 mux_195_i4_3_lut (.A(quarter_wave_sample_register_i[3]), .B(o_val_pipeline_i_0__15__N_2157[3]), 
         .C(phase_negation_i[1]), .Z(n1212[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam mux_195_i4_3_lut.init = 16'hcaca;
    LUT4 i19405_3_lut_4_lut_4_lut (.A(index_i[2]), .B(n141), .C(index_i[3]), 
         .D(n26969), .Z(n21842)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19405_3_lut_4_lut_4_lut.init = 16'hc5c0;
    LUT4 mux_195_i3_3_lut (.A(quarter_wave_sample_register_i[2]), .B(o_val_pipeline_i_0__15__N_2157[2]), 
         .C(phase_negation_i[1]), .Z(n1212[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam mux_195_i3_3_lut.init = 16'hcaca;
    LUT4 mux_195_i2_3_lut (.A(quarter_wave_sample_register_i[1]), .B(o_val_pipeline_i_0__15__N_2157[1]), 
         .C(phase_negation_i[1]), .Z(n1212[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam mux_195_i2_3_lut.init = 16'hcaca;
    LUT4 mux_195_i1_3_lut (.A(quarter_wave_sample_register_i[0]), .B(o_val_pipeline_i_0__15__N_2157[0]), 
         .C(phase_negation_i[1]), .Z(n1212[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam mux_195_i1_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_4_i491_3_lut_4_lut_4_lut (.A(index_i[2]), .B(n26972), 
         .C(index_i[3]), .D(n27037), .Z(n491_adj_2828)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_4_i491_3_lut_4_lut_4_lut.init = 16'hfc5c;
    LUT4 n25289_bdd_3_lut (.A(n27152), .B(n25287), .C(index_i[5]), .Z(n25290)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n25289_bdd_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_7_i506_3_lut_4_lut_4_lut (.A(index_i[2]), .B(n26972), 
         .C(index_i[3]), .D(n26969), .Z(n506)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B ((D)+!C)+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_7_i506_3_lut_4_lut_4_lut.init = 16'h5c0c;
    LUT4 i19075_3_lut (.A(n26971), .B(n29496), .C(index_i[3]), .Z(n21512)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19075_3_lut.init = 16'hcaca;
    LUT4 n133_bdd_3_lut_24139_4_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .Z(n25053)) /* synthesis lut_function=(A (B)+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n133_bdd_3_lut_24139_4_lut_3_lut.init = 16'hd9d9;
    LUT4 mux_198_Mux_0_i715_3_lut_3_lut_rep_619_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26942)) /* synthesis lut_function=(A (B (C))+!A !(B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i715_3_lut_3_lut_rep_619_3_lut.init = 16'h9595;
    LUT4 i11095_2_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n668)) /* synthesis lut_function=(!(A ((D)+!B)+!A (B ((D)+!C)+!B (C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11095_2_lut_4_lut_4_lut_4_lut.init = 16'h00c9;
    PFUMX i24253 (.BLUT(n26089), .ALUT(n21407), .C0(index_i[4]), .Z(n26090));
    LUT4 mux_198_Mux_6_i573_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[4]), .D(n572_adj_2970), .Z(n573_adj_2940)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_6_i573_3_lut_4_lut.init = 16'hf909;
    LUT4 mux_198_Mux_0_i908_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n908)) /* synthesis lut_function=(!(A (B (C (D))+!B !(D))+!A (B+((D)+!C)))) */ ;
    defparam mux_198_Mux_0_i908_3_lut_4_lut_4_lut.init = 16'h2a98;
    LUT4 mux_198_Mux_7_i45_3_lut_3_lut_rep_628_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26951)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_7_i45_3_lut_3_lut_rep_628_3_lut.init = 16'h3939;
    PFUMX i24755 (.BLUT(n27162), .ALUT(n27163), .C0(index_i[0]), .Z(n27164));
    LUT4 i9461_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[4]), .D(n27036), .Z(n189_adj_2894)) /* synthesis lut_function=(A (B (C (D)))+!A !(B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9461_3_lut_4_lut_4_lut_4_lut.init = 16'h9555;
    LUT4 i23595_then_4_lut (.A(index_i[2]), .B(index_i[4]), .C(index_i[1]), 
         .D(index_i[3]), .Z(n27127)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B (C)+!B !(C (D)+!C !(D))))) */ ;
    defparam i23595_then_4_lut.init = 16'h3c2d;
    LUT4 mux_198_Mux_5_i924_4_lut_3_lut (.A(index_i[2]), .B(n14825), .C(index_i[4]), 
         .Z(n924_adj_2971)) /* synthesis lut_function=(!(A (B+(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_5_i924_4_lut_3_lut.init = 16'h5656;
    LUT4 i19446_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n21883)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !(B (C+!(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19446_3_lut_4_lut_4_lut.init = 16'ha5a9;
    LUT4 i21756_3_lut (.A(n21511), .B(n21512), .C(index_i[4]), .Z(n21513)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21756_3_lut.init = 16'hcaca;
    LUT4 i18970_3_lut (.A(n26972), .B(n141), .C(index_i[3]), .Z(n21407)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18970_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_6_i498_3_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n404)) /* synthesis lut_function=(A (B+!(C))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_6_i498_3_lut_4_lut_3_lut.init = 16'h9b9b;
    LUT4 mux_198_Mux_2_i604_3_lut_4_lut_4_lut_4_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n604_adj_2885)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)+!C !(D)))+!A (B (C)+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_2_i604_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'h3c9f;
    LUT4 i19417_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21854)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D))+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19417_3_lut_4_lut.init = 16'hccdb;
    LUT4 mux_198_Mux_1_i93_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n93_adj_2922)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C+(D)))+!A !(B (C (D)+!C !(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_1_i93_3_lut_4_lut_4_lut_4_lut.init = 16'h955a;
    LUT4 i21839_3_lut (.A(n21508), .B(n21509), .C(index_i[4]), .Z(n21510)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21839_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_0_i134_3_lut_4_lut_3_lut_rep_687 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27010)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i134_3_lut_4_lut_3_lut_rep_687.init = 16'h6969;
    LUT4 mux_198_Mux_0_i219_3_lut_3_lut_3_lut_rep_688 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27011)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i219_3_lut_3_lut_3_lut_rep_688.init = 16'h9393;
    PFUMX i20658 (.BLUT(n94_adj_2874), .ALUT(n21786), .C0(index_i[5]), 
          .Z(n23114));
    LUT4 mux_198_Mux_7_i77_3_lut_3_lut_rep_689 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27012)) /* synthesis lut_function=(A (B)+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_7_i77_3_lut_3_lut_rep_689.init = 16'h9c9c;
    LUT4 mux_198_Mux_0_i660_3_lut_rep_690 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27013)) /* synthesis lut_function=(A (B)+!A (B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i660_3_lut_rep_690.init = 16'hc9c9;
    LUT4 mux_198_Mux_6_i645_3_lut_4_lut_3_lut_rep_691 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27014)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_6_i645_3_lut_4_lut_3_lut_rep_691.init = 16'h1919;
    LUT4 mux_198_Mux_0_i165_3_lut_4_lut_3_lut_rep_692 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27015)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i165_3_lut_4_lut_3_lut_rep_692.init = 16'h9292;
    LUT4 mux_198_Mux_3_i676_3_lut_4_lut_3_lut_rep_693 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27016)) /* synthesis lut_function=(A (B (C))+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_3_i676_3_lut_4_lut_3_lut_rep_693.init = 16'h9494;
    LUT4 i19069_3_lut (.A(n404), .B(n27013), .C(index_i[3]), .Z(n21506)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19069_3_lut.init = 16'hcaca;
    PFUMX i20660 (.BLUT(n221_adj_2972), .ALUT(n252_adj_2973), .C0(index_i[5]), 
          .Z(n23116));
    PFUMX i20661 (.BLUT(n286_adj_2872), .ALUT(n21789), .C0(index_i[5]), 
          .Z(n23117));
    LUT4 mux_198_Mux_4_i262_3_lut_3_lut_rep_694 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27017)) /* synthesis lut_function=(A (B+(C))+!A !(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_4_i262_3_lut_3_lut_rep_694.init = 16'ha9a9;
    LUT4 mux_198_Mux_6_i134_3_lut_4_lut_3_lut_rep_695 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27018)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_6_i134_3_lut_4_lut_3_lut_rep_695.init = 16'h9696;
    LUT4 mux_198_Mux_6_i356_3_lut_4_lut_3_lut_rep_696 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27019)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_6_i356_3_lut_4_lut_3_lut_rep_696.init = 16'h4949;
    PFUMX i20662 (.BLUT(n349_adj_2974), .ALUT(n21792), .C0(index_i[5]), 
          .Z(n23118));
    LUT4 mux_198_Mux_6_i564_3_lut_4_lut_3_lut_rep_697 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27020)) /* synthesis lut_function=(A (B)+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_6_i564_3_lut_4_lut_3_lut_rep_697.init = 16'hd9d9;
    LUT4 mux_198_Mux_6_i572_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n572_adj_2970)) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_6_i572_3_lut_4_lut.init = 16'hccd9;
    LUT4 i19437_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21874)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (D))+!A !(B (C (D))+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19437_3_lut_3_lut_4_lut.init = 16'h4933;
    LUT4 n284_bdd_3_lut_23967_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n25764)) /* synthesis lut_function=(A (B (C+(D))+!B ((D)+!C))+!A !(B (C+(D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n284_bdd_3_lut_23967_4_lut.init = 16'haa96;
    LUT4 i23595_else_4_lut (.A(index_i[2]), .B(index_i[4]), .C(index_i[1]), 
         .D(index_i[3]), .Z(n27126)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A (B ((D)+!C)+!B !((D)+!C)))) */ ;
    defparam i23595_else_4_lut.init = 16'h39c3;
    LUT4 i19428_3_lut (.A(n900), .B(n27013), .C(index_i[3]), .Z(n21865)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19428_3_lut.init = 16'hcaca;
    LUT4 i19392_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21829)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A !(B (D)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19392_3_lut_3_lut_4_lut.init = 16'ha955;
    LUT4 mux_198_Mux_3_i397_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n397_adj_2839)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !(B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_3_i397_3_lut_4_lut_4_lut.init = 16'ha95a;
    LUT4 n572_bdd_3_lut_24509_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n25762)) /* synthesis lut_function=(A (B (C+(D)))+!A (B ((D)+!C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n572_bdd_3_lut_24509_4_lut.init = 16'hcc94;
    LUT4 mux_198_Mux_3_i684_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[4]), .Z(n684_adj_2962)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A !(B ((D)+!C)+!B (C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_3_i684_3_lut_3_lut_4_lut.init = 16'h5594;
    LUT4 mux_198_Mux_2_i653_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n653_adj_2883)) /* synthesis lut_function=(A (B (C+!(D))+!B !(D))+!A !(B (C+!(D))+!B !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_2_i653_3_lut_4_lut.init = 16'h94aa;
    LUT4 i19407_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21844)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C))+!A !(B ((D)+!C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19407_3_lut_4_lut_4_lut.init = 16'h925a;
    LUT4 i20010_3_lut (.A(n22463), .B(n22464), .C(index_i[8]), .Z(n22466)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20010_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_0_i812_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n812)) /* synthesis lut_function=(A (B (C+(D))+!B !(C))+!A (B (D)+!B !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i812_3_lut_4_lut_4_lut_4_lut.init = 16'hcf92;
    LUT4 i19074_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21511)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(D))+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19074_3_lut_3_lut_4_lut.init = 16'h3319;
    PFUMX i20667 (.BLUT(n669_adj_2865), .ALUT(n700_adj_2862), .C0(index_i[5]), 
          .Z(n23123));
    LUT4 i19471_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21908)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C+(D)))+!A (B (C)+!B !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19471_3_lut_4_lut_4_lut.init = 16'hc95a;
    LUT4 mux_198_Mux_3_i859_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n859)) /* synthesis lut_function=(!(A (B (D)+!B !(D))+!A (B (C+(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_3_i859_3_lut_3_lut_4_lut.init = 16'h339c;
    LUT4 i19080_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21517)) /* synthesis lut_function=(A (B (C (D))+!B !(C (D)))+!A !(B (D)+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19080_3_lut_4_lut_4_lut.init = 16'h9366;
    L6MUX21 i24211 (.D0(n26046), .D1(n26044), .SD(index_i[5]), .Z(n26047));
    PFUMX i20668 (.BLUT(n21804), .ALUT(n763_adj_2827), .C0(index_i[5]), 
          .Z(n23124));
    LUT4 i19461_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21898)) /* synthesis lut_function=(A (B (C)+!B (C (D)+!C !(D)))+!A !(B (C+!(D))+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19461_3_lut_4_lut_4_lut.init = 16'ha593;
    LUT4 mux_198_Mux_0_i142_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n142_adj_2975)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C))+!A !(B (C (D)+!C !(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i142_3_lut_4_lut_4_lut.init = 16'ha569;
    PFUMX i24209 (.BLUT(n572_adj_2976), .ALUT(n26045), .C0(index_i[4]), 
          .Z(n26046));
    PFUMX i20669 (.BLUT(n21807), .ALUT(n828_adj_2977), .C0(index_i[5]), 
          .Z(n23125));
    PFUMX i20670 (.BLUT(n860_adj_2860), .ALUT(n21810), .C0(index_i[5]), 
          .Z(n23126));
    LUT4 i21830_3_lut (.A(n27149), .B(n21863), .C(index_i[4]), .Z(n21864)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21830_3_lut.init = 16'hcaca;
    PFUMX i24206 (.BLUT(n26043), .ALUT(n26042), .C0(index_i[4]), .Z(n26044));
    LUT4 i18967_3_lut (.A(n26972), .B(n645), .C(index_i[3]), .Z(n21404)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18967_3_lut.init = 16'hcaca;
    LUT4 i18966_3_lut (.A(n27041), .B(n141), .C(index_i[3]), .Z(n21403)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18966_3_lut.init = 16'hcaca;
    PFUMX i20133 (.BLUT(n956), .ALUT(n20328), .C0(index_i[6]), .Z(n22589));
    L6MUX21 i24199 (.D0(n26035), .D1(n26032), .SD(index_i[5]), .Z(n26036));
    LUT4 mux_198_Mux_7_i173_3_lut (.A(n27012), .B(n645), .C(index_i[3]), 
         .Z(n173_adj_2978)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_7_i173_3_lut.init = 16'hcaca;
    PFUMX i24197 (.BLUT(n26034), .ALUT(n26033), .C0(index_i[4]), .Z(n26035));
    LUT4 i19419_3_lut (.A(n404), .B(n26954), .C(index_i[3]), .Z(n21856)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19419_3_lut.init = 16'hcaca;
    LUT4 i21685_3_lut (.A(n21856), .B(n21857), .C(index_i[4]), .Z(n21858)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21685_3_lut.init = 16'hcaca;
    L6MUX21 i25831 (.D0(n28617), .D1(n28614), .SD(index_i[7]), .Z(n28618));
    PFUMX i25829 (.BLUT(n28616), .ALUT(n28615), .C0(index_i[5]), .Z(n28617));
    LUT4 mux_198_Mux_11_i638_4_lut_4_lut (.A(n26739), .B(index_i[5]), .C(index_i[6]), 
         .D(n26779), .Z(n638)) /* synthesis lut_function=(A (B (C (D))+!B !(C))+!A (B ((D)+!C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_11_i638_4_lut_4_lut.init = 16'hc707;
    PFUMX i24194 (.BLUT(n26729), .ALUT(n26031), .C0(index_i[4]), .Z(n26032));
    PFUMX i25827 (.BLUT(n22508), .ALUT(n28613), .C0(index_i[6]), .Z(n28614));
    LUT4 i9590_3_lut_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n12155)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A !(B (C+(D))+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9590_3_lut_3_lut_4_lut_4_lut.init = 16'h44db;
    LUT4 i20684_3_lut (.A(n23135), .B(n23136), .C(index_i[7]), .Z(n23140)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20684_3_lut.init = 16'hcaca;
    LUT4 i19414_3_lut (.A(n404), .B(n29467), .C(index_i[3]), .Z(n21851)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19414_3_lut.init = 16'hcaca;
    PFUMX mux_198_Mux_7_i190 (.BLUT(n21405), .ALUT(n173_adj_2978), .C0(index_i[5]), 
          .Z(n190)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    PFUMX i19120 (.BLUT(n445), .ALUT(n508), .C0(index_i[6]), .Z(n21557));
    LUT4 i19066_3_lut (.A(n404), .B(n26961), .C(index_i[3]), .Z(n21503)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19066_3_lut.init = 16'hcaca;
    LUT4 i19065_3_lut (.A(n27015), .B(n325), .C(index_i[3]), .Z(n21502)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19065_3_lut.init = 16'hcaca;
    PFUMX i20689 (.BLUT(n94_adj_2979), .ALUT(n125_adj_2851), .C0(index_i[5]), 
          .Z(n23145));
    LUT4 i1_2_lut_rep_713 (.A(index_i[3]), .B(index_i[2]), .Z(n27036)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i1_2_lut_rep_713.init = 16'h8888;
    PFUMX i20690 (.BLUT(n158), .ALUT(n189), .C0(index_i[5]), .Z(n23146));
    LUT4 mux_198_Mux_5_i572_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n572_adj_2976)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A !(B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_5_i572_3_lut_4_lut_4_lut.init = 16'ha9a5;
    LUT4 i19063_3_lut (.A(n27015), .B(n26961), .C(index_i[3]), .Z(n21500)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19063_3_lut.init = 16'hcaca;
    LUT4 i15562_3_lut_3_lut_3_lut_4_lut (.A(index_i[3]), .B(index_i[2]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n17826)) /* synthesis lut_function=(!(A (B (C)+!B !(C (D)+!C !(D)))+!A !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i15562_3_lut_3_lut_3_lut_4_lut.init = 16'h780f;
    LUT4 mux_198_Mux_0_i364_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n364_adj_2980)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A ((C+!(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i364_3_lut_3_lut_4_lut.init = 16'hdb55;
    LUT4 i20427_3_lut_3_lut_3_lut_4_lut (.A(index_i[3]), .B(index_i[2]), 
         .C(index_i[4]), .D(index_i[1]), .Z(n22883)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20427_3_lut_3_lut_3_lut_4_lut.init = 16'h878f;
    LUT4 i12228_2_lut_rep_477_3_lut (.A(index_i[3]), .B(index_i[2]), .C(index_i[1]), 
         .Z(n26800)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i12228_2_lut_rep_477_3_lut.init = 16'h8080;
    LUT4 i19062_3_lut (.A(n325), .B(n332), .C(index_i[3]), .Z(n21499)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19062_3_lut.init = 16'hcaca;
    LUT4 i12253_2_lut_rep_522_3_lut_4_lut (.A(index_i[3]), .B(index_i[2]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n26845)) /* synthesis lut_function=(A (B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i12253_2_lut_rep_522_3_lut_4_lut.init = 16'h8880;
    LUT4 i11775_2_lut_2_lut_3_lut (.A(index_i[3]), .B(index_i[2]), .C(index_i[0]), 
         .Z(n14450)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11775_2_lut_2_lut_3_lut.init = 16'h0808;
    LUT4 mux_198_Mux_3_i62_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[4]), .D(n812_adj_2925), .Z(n62_adj_2968)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_3_i62_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_198_Mux_3_i94_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[4]), .D(n93_adj_2840), .Z(n94_adj_2979)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_3_i94_3_lut_4_lut.init = 16'hf606;
    LUT4 i7335_3_lut_3_lut_4_lut (.A(index_i[3]), .B(index_i[2]), .C(index_i[1]), 
         .D(index_i[0]), .Z(n157_adj_2903)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(D))+!A !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i7335_3_lut_3_lut_4_lut.init = 16'h7780;
    LUT4 i9431_3_lut_3_lut_3_lut_4_lut (.A(index_i[3]), .B(index_i[2]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n541_adj_2833)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9431_3_lut_3_lut_3_lut_4_lut.init = 16'h870f;
    LUT4 i15561_3_lut_3_lut_4_lut (.A(index_i[3]), .B(index_i[2]), .C(index_i[1]), 
         .D(index_i[0]), .Z(n17825)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i15561_3_lut_3_lut_4_lut.init = 16'hf078;
    LUT4 i9474_3_lut_3_lut_3_lut_4_lut (.A(index_i[3]), .B(index_i[2]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n875_adj_2844)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(D))+!A !(D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9474_3_lut_3_lut_3_lut_4_lut.init = 16'h887f;
    LUT4 i19956_1_lut_2_lut (.A(index_i[3]), .B(index_i[2]), .Z(n22412)) /* synthesis lut_function=(!(A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19956_1_lut_2_lut.init = 16'h7777;
    LUT4 i9467_3_lut_3_lut_4_lut_3_lut_4_lut (.A(index_i[3]), .B(index_i[2]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n762_adj_2854)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C (D)+!C !(D)))+!A !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9467_3_lut_3_lut_4_lut_3_lut_4_lut.init = 16'h700f;
    PFUMX mux_198_Mux_8_i764 (.BLUT(n716_adj_2981), .ALUT(n732_adj_2843), 
          .C0(n22297), .Z(n764)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 i11180_2_lut_rep_448_3_lut_4_lut (.A(index_i[3]), .B(index_i[2]), 
         .C(index_i[4]), .D(n27037), .Z(n26771)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11180_2_lut_rep_448_3_lut_4_lut.init = 16'hf8f0;
    LUT4 mux_198_Mux_4_i828_3_lut_4_lut (.A(index_i[4]), .B(index_i[3]), 
         .C(n812_adj_2982), .D(n29483), .Z(n828_adj_2977)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_4_i828_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i20691 (.BLUT(n221_adj_2815), .ALUT(n252_adj_2786), .C0(index_i[5]), 
          .Z(n23147));
    LUT4 i11402_2_lut_rep_714 (.A(index_i[0]), .B(index_i[1]), .Z(n27037)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11402_2_lut_rep_714.init = 16'h8888;
    LUT4 mux_198_Mux_6_i781_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n781_adj_2863)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A (B (C (D)+!C !(D))+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_6_i781_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hc837;
    LUT4 mux_198_Mux_7_i262_3_lut_rep_627_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26950)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_7_i262_3_lut_rep_627_3_lut.init = 16'h3838;
    LUT4 mux_198_Mux_5_i797_3_lut_4_lut (.A(index_i[4]), .B(index_i[3]), 
         .C(n27140), .D(n26957), .Z(n797_adj_2955)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_5_i797_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_198_Mux_7_i526_3_lut_3_lut_4_lut_4_lut_3_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n526_adj_2935)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(D))+!A !(D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_7_i526_3_lut_3_lut_4_lut_4_lut_3_lut_4_lut.init = 16'h887f;
    PFUMX mux_198_Mux_8_i574 (.BLUT(n542), .ALUT(n11940), .C0(index_i[5]), 
          .Z(n574)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 i20480_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n22936)) /* synthesis lut_function=(A (B (C)+!B !(C (D)+!C !(D)))+!A !(B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20480_3_lut_4_lut_4_lut_4_lut.init = 16'h83f0;
    LUT4 mux_198_Mux_1_i763_3_lut_4_lut (.A(index_i[4]), .B(index_i[3]), 
         .C(n27148), .D(n26957), .Z(n763_adj_2800)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_1_i763_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i20692 (.BLUT(n286_adj_2841), .ALUT(n21819), .C0(index_i[5]), 
          .Z(n23148));
    LUT4 mux_198_Mux_8_i635_3_lut_4_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n635_adj_2794)) /* synthesis lut_function=(!(A (B (C (D))+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_8_i635_3_lut_4_lut_3_lut_4_lut.init = 16'h0ff8;
    LUT4 i4404_2_lut_rep_618 (.A(index_i[0]), .B(index_i[2]), .Z(n26941)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i4404_2_lut_rep_618.init = 16'h6666;
    LUT4 i11088_2_lut_rep_432_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n26755)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11088_2_lut_rep_432_3_lut_4_lut.init = 16'hf080;
    LUT4 mux_198_Mux_4_i1002_3_lut_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n1002_adj_2858)) /* synthesis lut_function=(A (B (C (D))+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_4_i1002_3_lut_3_lut_3_lut_4_lut.init = 16'hf007;
    LUT4 mux_198_Mux_8_i526_3_lut_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n526_adj_2793)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_8_i526_3_lut_3_lut_3_lut_4_lut.init = 16'h0f70;
    LUT4 i19444_3_lut_4_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n21881)) /* synthesis lut_function=(!(A (B (D)+!B !((D)+!C))+!A (B (C+(D))+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19444_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'h338f;
    LUT4 mux_198_Mux_4_i349_3_lut_4_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[4]), .D(n348_adj_2957), .Z(n349_adj_2974)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_4_i349_3_lut_4_lut.init = 16'hf606;
    PFUMX i20693 (.BLUT(n349_adj_2983), .ALUT(n21822), .C0(index_i[5]), 
          .Z(n23149));
    PFUMX i20694 (.BLUT(n413), .ALUT(n444_adj_2984), .C0(index_i[5]), 
          .Z(n23150));
    PFUMX i20695 (.BLUT(n476_adj_2838), .ALUT(n507_adj_2985), .C0(index_i[5]), 
          .Z(n23151));
    PFUMX i20696 (.BLUT(n21825), .ALUT(n573_adj_2818), .C0(index_i[5]), 
          .Z(n23152));
    LUT4 mux_198_Mux_1_i348_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n348_adj_2921)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A (B ((D)+!C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_1_i348_3_lut_4_lut_4_lut_4_lut.init = 16'h38f0;
    PFUMX i20697 (.BLUT(n12026), .ALUT(n21828), .C0(index_i[5]), .Z(n23153));
    LUT4 mux_198_Mux_7_i491_3_lut_4_lut_4_lut_4_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[2]), .D(index_i[3]), .Z(n491_adj_2803)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A (B ((D)+!C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_7_i491_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'h3870;
    LUT4 i12267_2_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(n27049), 
         .D(index_i[2]), .Z(n14956)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i12267_2_lut_3_lut_4_lut.init = 16'hf080;
    LUT4 i22764_2_lut_rep_501_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n26824)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i22764_2_lut_rep_501_3_lut_4_lut.init = 16'h0007;
    PFUMX i20698 (.BLUT(n669), .ALUT(n700_adj_2963), .C0(index_i[5]), 
          .Z(n23154));
    LUT4 mux_198_Mux_7_i141_3_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n141)) /* synthesis lut_function=(A ((C)+!B)+!A (B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_7_i141_3_lut_4_lut_3_lut.init = 16'he7e7;
    L6MUX21 i20699 (.D0(n21831), .D1(n763_adj_2855), .SD(index_i[5]), 
            .Z(n23155));
    LUT4 i21699_3_lut (.A(n21847), .B(n21848), .C(index_i[4]), .Z(n21849)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21699_3_lut.init = 16'hcaca;
    LUT4 n77_bdd_3_lut_24325_3_lut_4_lut_4_lut_3_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n25751)) /* synthesis lut_function=(A (B (C)+!B !(D))+!A !(D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n77_bdd_3_lut_24325_3_lut_4_lut_4_lut_3_lut_4_lut.init = 16'h80f7;
    LUT4 mux_198_Mux_6_i812_3_lut_4_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n812_adj_2925)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(D))+!A !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_6_i812_3_lut_4_lut_3_lut_4_lut.init = 16'h7780;
    LUT4 i11087_2_lut_rep_516_3_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .Z(n26839)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11087_2_lut_rep_516_3_lut.init = 16'hf8f8;
    LUT4 mux_198_Mux_3_i1002_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n19863)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (D))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_3_i1002_3_lut_3_lut_4_lut.init = 16'hf708;
    LUT4 i11280_2_lut_2_lut_3_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .Z(n13955)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11280_2_lut_2_lut_3_lut.init = 16'h0808;
    LUT4 i15529_3_lut_3_lut (.A(index_i[0]), .B(index_i[2]), .C(index_i[3]), 
         .Z(n17793)) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i15529_3_lut_3_lut.init = 16'h6a6a;
    LUT4 i11254_3_lut_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n13928)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (D))+!A (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11254_3_lut_3_lut_3_lut_4_lut.init = 16'h00f7;
    PFUMX i20701 (.BLUT(n860_adj_2830), .ALUT(n891_adj_2834), .C0(index_i[5]), 
          .Z(n23157));
    LUT4 i19408_3_lut (.A(n29467), .B(n26971), .C(index_i[3]), .Z(n21845)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19408_3_lut.init = 16'hcaca;
    LUT4 i11395_2_lut_rep_431_4_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n26754)) /* synthesis lut_function=(!(A (B (C+(D))+!B (C+!(D)))+!A (B+(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11395_2_lut_rep_431_4_lut_4_lut_4_lut_4_lut.init = 16'h0308;
    LUT4 mux_198_Mux_1_i890_4_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[3]), 
         .C(n645), .D(index_i[4]), .Z(n890_adj_2967)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (D))+!A !((C+(D))+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_1_i890_4_lut_4_lut_4_lut_4_lut.init = 16'h55f3;
    LUT4 i21701_3_lut (.A(n21844), .B(n21845), .C(index_i[4]), .Z(n21846)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21701_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_8_i172_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n70)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_8_i172_3_lut_3_lut.init = 16'h7c7c;
    LUT4 mux_198_Mux_0_i29_3_lut_rep_626_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26949)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i29_3_lut_rep_626_3_lut.init = 16'h8383;
    LUT4 mux_198_Mux_5_i573_3_lut_3_lut (.A(index_i[0]), .B(index_i[4]), 
         .C(n572_adj_2976), .Z(n573_adj_2953)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_5_i573_3_lut_3_lut.init = 16'hd1d1;
    LUT4 mux_198_Mux_2_i763_4_lut_4_lut (.A(index_i[0]), .B(n12030), .C(index_i[4]), 
         .D(n157_adj_2909), .Z(n763_adj_2966)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_2_i763_4_lut_4_lut.init = 16'hdfd0;
    PFUMX i20702 (.BLUT(n924_adj_2832), .ALUT(n21834), .C0(index_i[5]), 
          .Z(n23158));
    PFUMX i20703 (.BLUT(n21837), .ALUT(n1018), .C0(index_i[5]), .Z(n23159));
    LUT4 i1_2_lut_rep_545_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n26868)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i1_2_lut_rep_545_3_lut_4_lut.init = 16'h8000;
    LUT4 i19377_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n21814)) /* synthesis lut_function=(!(A (B (D)+!B !(D))+!A (B ((D)+!C)+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19377_3_lut_4_lut_4_lut_4_lut.init = 16'h33c8;
    LUT4 i19449_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n21886)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A (B (C)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19449_3_lut_4_lut_4_lut.init = 16'h3c8c;
    LUT4 mux_198_Mux_7_i620_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n620)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A !(B (C+!(D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_7_i620_3_lut_4_lut_4_lut_4_lut.init = 16'h8c33;
    LUT4 mux_198_Mux_8_i93_3_lut_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n93_adj_2933)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (D))+!A (B ((D)+!C)+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_8_i93_3_lut_3_lut_4_lut_4_lut.init = 16'h08f3;
    LUT4 mux_198_Mux_8_i29_3_lut_rep_715 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27038)) /* synthesis lut_function=(!(A (B (C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_8_i29_3_lut_rep_715.init = 16'h7e7e;
    LUT4 mux_198_Mux_7_i92_3_lut_rep_716 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27039)) /* synthesis lut_function=(A (B+!(C))+!A !((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_7_i92_3_lut_rep_716.init = 16'h8e8e;
    LUT4 mux_198_Mux_7_i60_3_lut_4_lut_3_lut_rep_718 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27041)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_7_i60_3_lut_4_lut_3_lut_rep_718.init = 16'h1818;
    LUT4 mux_198_Mux_0_i581_3_lut_3_lut_rep_719 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27042)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i581_3_lut_3_lut_rep_719.init = 16'hc7c7;
    LUT4 mux_198_Mux_5_i30_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n30_adj_2916)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A (B+!(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_5_i30_3_lut_4_lut.init = 16'hcc67;
    LUT4 i21705_3_lut (.A(n21841), .B(n21842), .C(index_i[4]), .Z(n21843)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21705_3_lut.init = 16'hcaca;
    LUT4 i19413_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21850)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+(D)))+!A !(B (D)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19413_3_lut_4_lut_4_lut.init = 16'h99c7;
    LUT4 n262_bdd_3_lut_24525_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n25554)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C))+!A (B (C (D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n262_bdd_3_lut_24525_3_lut_4_lut.init = 16'h0fc7;
    LUT4 n12151_bdd_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[4]), 
         .D(index_i[2]), .Z(n26091)) /* synthesis lut_function=(A (B)+!A !(B (D)+!B !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n12151_bdd_3_lut_4_lut.init = 16'h98cc;
    LUT4 i19429_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21866)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A (B (D)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19429_3_lut_4_lut.init = 16'h18cc;
    LUT4 mux_198_Mux_2_i557_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n557_adj_2819)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C+!(D))+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_2_i557_3_lut_3_lut_4_lut.init = 16'h0f18;
    LUT4 mux_198_Mux_7_i716_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n716_adj_2932)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C+!(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_7_i716_3_lut_3_lut_4_lut.init = 16'h0f81;
    LUT4 mux_198_Mux_4_i221_3_lut_3_lut (.A(index_i[0]), .B(index_i[4]), 
         .C(n205), .Z(n221_adj_2972)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_4_i221_3_lut_3_lut.init = 16'h7474;
    LUT4 i19386_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21823)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)))+!A !(B (C+!(D))+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19386_3_lut_3_lut_4_lut.init = 16'h71cc;
    LUT4 mux_198_Mux_4_i526_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n526_adj_2850)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A !(B ((D)+!C)+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_4_i526_3_lut_3_lut_4_lut.init = 16'h7e0f;
    LUT4 i19350_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21787)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A !(B (C+!(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19350_3_lut_4_lut_4_lut.init = 16'ha52b;
    LUT4 mux_198_Mux_2_i349_3_lut_3_lut (.A(index_i[0]), .B(index_i[4]), 
         .C(n348_adj_2986), .Z(n349_adj_2964)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_2_i349_3_lut_3_lut.init = 16'hd1d1;
    LUT4 i19396_3_lut (.A(n325), .B(n27013), .C(index_i[3]), .Z(n21833)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19396_3_lut.init = 16'hcaca;
    LUT4 i21555_3_lut (.A(n21832), .B(n21833), .C(index_i[4]), .Z(n21834)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21555_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_2_i507_3_lut_3_lut (.A(index_i[0]), .B(index_i[4]), 
         .C(n491_adj_2987), .Z(n507_adj_2965)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_2_i507_3_lut_3_lut.init = 16'h7474;
    LUT4 i19686_3_lut_4_lut_4_lut (.A(index_i[0]), .B(n26958), .C(index_i[3]), 
         .D(n27050), .Z(n22123)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19686_3_lut_4_lut_4_lut.init = 16'hcfc5;
    LUT4 mux_198_Mux_3_i444_3_lut_4_lut (.A(index_i[0]), .B(index_i[3]), 
         .C(n27050), .D(index_i[4]), .Z(n444_adj_2984)) /* synthesis lut_function=(!(A (B (D)+!B (C (D)))+!A !(B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_3_i444_3_lut_4_lut.init = 16'h46aa;
    L6MUX21 i22894 (.D0(n24547), .D1(n26705), .SD(index_i[6]), .Z(n24548));
    LUT4 mux_198_Mux_4_i252_4_lut_4_lut (.A(index_i[0]), .B(index_i[3]), 
         .C(n27052), .D(index_i[4]), .Z(n252_adj_2973)) /* synthesis lut_function=(!(A (B (D)+!B !(D))+!A !(B ((D)+!C)+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_4_i252_4_lut_4_lut.init = 16'h669d;
    PFUMX i25584 (.BLUT(n28290), .ALUT(n28289), .C0(index_i[3]), .Z(n28291));
    LUT4 i19393_3_lut (.A(n27016), .B(n29479), .C(index_i[3]), .Z(n21830)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19393_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_4_lut (.A(n26739), .B(index_i[5]), .C(index_i[8]), .D(n19786), 
         .Z(n20196)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i1_3_lut_4_lut.init = 16'hfff8;
    LUT4 i21568_3_lut (.A(n21826), .B(n21827), .C(index_i[4]), .Z(n21828)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21568_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_1_i62_3_lut_4_lut (.A(index_i[0]), .B(index_i[3]), 
         .C(index_i[2]), .D(index_i[4]), .Z(n62_adj_2951)) /* synthesis lut_function=(A (B (D)+!B ((D)+!C))+!A !(B (D)+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_1_i62_3_lut_4_lut.init = 16'haa56;
    PFUMX i22892 (.BLUT(n24546), .ALUT(n24545), .C0(index_i[5]), .Z(n24547));
    LUT4 i19384_3_lut (.A(n27007), .B(n29480), .C(index_i[3]), .Z(n21821)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19384_3_lut.init = 16'hcaca;
    LUT4 i20135_3_lut (.A(n22584), .B(n22585), .C(index_i[7]), .Z(n22591)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20135_3_lut.init = 16'hcaca;
    LUT4 i19383_3_lut (.A(n29482), .B(n27019), .C(index_i[3]), .Z(n21820)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19383_3_lut.init = 16'hcaca;
    LUT4 i21575_3_lut (.A(n21820), .B(n21821), .C(index_i[4]), .Z(n21822)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21575_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_2_i348_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n348_adj_2986)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_2_i348_3_lut_4_lut_4_lut.init = 16'h52a5;
    LUT4 i20134_3_lut (.A(n22582), .B(n22583), .C(index_i[7]), .Z(n22590)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20134_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_3_i349_3_lut_3_lut (.A(index_i[1]), .B(index_i[4]), 
         .C(n348_adj_2961), .Z(n349_adj_2983)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_3_i349_3_lut_3_lut.init = 16'hd1d1;
    LUT4 i19364_then_4_lut (.A(index_i[0]), .B(index_i[4]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n27133)) /* synthesis lut_function=(A (B (C)+!B (C (D)+!C !(D)))+!A !(B (C+!(D))+!B !(C+!(D)))) */ ;
    defparam i19364_then_4_lut.init = 16'hb493;
    PFUMX i20947 (.BLUT(n23401), .ALUT(n23402), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2126[1]));
    LUT4 i19381_3_lut (.A(n29496), .B(n27014), .C(index_i[3]), .Z(n21818)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19381_3_lut.init = 16'hcaca;
    PFUMX i20597 (.BLUT(n23051), .ALUT(n23052), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2126[5]));
    LUT4 i9462_2_lut_rep_726 (.A(index_i[3]), .B(index_i[4]), .Z(n27049)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9462_2_lut_rep_726.init = 16'h8888;
    LUT4 i11279_3_lut_3_lut_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[0]), 
         .Z(n85)) /* synthesis lut_function=(!(A ((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11279_3_lut_3_lut_3_lut.init = 16'h5d5d;
    LUT4 i1_2_lut_rep_555_3_lut (.A(index_i[3]), .B(index_i[4]), .C(index_i[5]), 
         .Z(n26878)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i1_2_lut_rep_555_3_lut.init = 16'hf8f8;
    LUT4 i19380_3_lut (.A(n27039), .B(n85), .C(index_i[3]), .Z(n21817)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19380_3_lut.init = 16'hcaca;
    LUT4 i9463_3_lut_3_lut_3_lut_4_lut (.A(index_i[3]), .B(index_i[4]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n444_adj_2988)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C))+!A (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9463_3_lut_3_lut_3_lut_4_lut.init = 16'h0f87;
    LUT4 i21578_3_lut (.A(n21817), .B(n21818), .C(index_i[4]), .Z(n21819)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21578_3_lut.init = 16'hcaca;
    LUT4 i20045_3_lut_3_lut_4_lut (.A(index_i[3]), .B(index_i[4]), .C(n413_adj_2886), 
         .D(index_i[5]), .Z(n22501)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20045_3_lut_3_lut_4_lut.init = 16'h77f0;
    LUT4 i1_2_lut_3_lut (.A(index_i[3]), .B(index_i[4]), .C(index_i[5]), 
         .Z(n20563)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i1_2_lut_3_lut.init = 16'h8080;
    LUT4 i11396_2_lut_rep_727 (.A(index_i[1]), .B(index_i[2]), .Z(n27050)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11396_2_lut_rep_727.init = 16'h8888;
    LUT4 i9469_2_lut_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[3]), 
         .Z(n12030)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9469_2_lut_3_lut.init = 16'h8080;
    LUT4 n476_bdd_3_lut_23593_3_lut (.A(index_i[1]), .B(index_i[4]), .C(n124_adj_2911), 
         .Z(n25285)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n476_bdd_3_lut_23593_3_lut.init = 16'hd1d1;
    LUT4 i19411_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .D(index_i[3]), .Z(n21848)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(D))+!A (B+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19411_3_lut_4_lut_4_lut_4_lut.init = 16'h3380;
    LUT4 i11193_2_lut_rep_491_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[3]), 
         .Z(n26814)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11193_2_lut_rep_491_3_lut.init = 16'hf8f8;
    LUT4 mux_198_Mux_0_i396_3_lut_4_lut_3_lut_rep_806 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29479)) /* synthesis lut_function=(A ((C)+!B)+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i396_3_lut_4_lut_3_lut_rep_806.init = 16'hb6b6;
    LUT4 i19369_3_lut_4_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n21806)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19369_3_lut_4_lut_3_lut_4_lut.init = 16'hf80f;
    LUT4 mux_198_Mux_4_i93_3_lut_4_lut_3_lut_rep_622_4_lut (.A(index_i[1]), 
         .B(index_i[2]), .C(index_i[3]), .D(index_i[0]), .Z(n26945)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_4_i93_3_lut_4_lut_3_lut_rep_622_4_lut.init = 16'h07f0;
    LUT4 i11717_2_lut_rep_556_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[0]), 
         .Z(n26879)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11717_2_lut_rep_556_3_lut.init = 16'h8080;
    LUT4 mux_198_Mux_6_i636_4_lut_4_lut (.A(index_i[1]), .B(index_i[4]), 
         .C(n635_adj_2914), .D(n14450), .Z(n636_adj_2942)) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_6_i636_4_lut_4_lut.init = 16'hf3d1;
    LUT4 mux_198_Mux_3_i142_3_lut_3_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .Z(n142)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_3_i142_3_lut_3_lut_3_lut.init = 16'h3838;
    LUT4 i11176_2_lut_rep_457_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n26780)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11176_2_lut_rep_457_3_lut_4_lut.init = 16'hf8f0;
    LUT4 mux_198_Mux_1_i301_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n301_adj_2969)) /* synthesis lut_function=(A (B (C+(D))+!B !(D))+!A !(B (C+(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_1_i301_3_lut_4_lut_4_lut.init = 16'h99b6;
    LUT4 i11772_2_lut_rep_506_2_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .Z(n26829)) /* synthesis lut_function=(A (B+!(C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11772_2_lut_rep_506_2_lut_3_lut.init = 16'h8f8f;
    LUT4 i11774_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[4]), 
         .C(n27036), .D(index_i[0]), .Z(n14449)) /* synthesis lut_function=(!(A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11774_3_lut_4_lut_4_lut_4_lut.init = 16'h55d5;
    PFUMX i20718 (.BLUT(n23172), .ALUT(n23173), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2126[3]));
    LUT4 mux_198_Mux_8_i491_3_lut_3_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n491_adj_2948)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_8_i491_3_lut_3_lut_3_lut_4_lut.init = 16'h7870;
    LUT4 i19348_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n21785)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C (D)+!C !(D)))+!A !(B (D)+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19348_3_lut_4_lut_4_lut_4_lut.init = 16'h7c03;
    LUT4 mux_198_Mux_2_i908_3_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .D(index_i[3]), .Z(n908_adj_2960)) /* synthesis lut_function=(!(A (B+!(D))+!A !(B+!(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_2_i908_3_lut_4_lut_4_lut.init = 16'h6645;
    LUT4 i11083_2_lut_rep_630 (.A(index_i[0]), .B(index_i[1]), .Z(n26953)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11083_2_lut_rep_630.init = 16'h4444;
    LUT4 mux_198_Mux_0_i954_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n954)) /* synthesis lut_function=(A (D)+!A !(B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i954_3_lut_4_lut_4_lut.init = 16'haf40;
    LUT4 i11714_2_lut_rep_728 (.A(index_i[1]), .B(index_i[2]), .C(index_i[0]), 
         .Z(n27051)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11714_2_lut_rep_728.init = 16'h7070;
    LUT4 mux_198_Mux_0_i1017_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .D(index_i[3]), .Z(n1017)) /* synthesis lut_function=(A (B (D)+!B !((D)+!C))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i1017_4_lut_4_lut_4_lut.init = 16'hdd70;
    LUT4 i20913_3_lut (.A(n23364), .B(n23365), .C(index_i[7]), .Z(n23369)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20913_3_lut.init = 16'hcaca;
    LUT4 i11405_2_lut_rep_729 (.A(index_i[1]), .B(index_i[2]), .Z(n27052)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11405_2_lut_rep_729.init = 16'heeee;
    LUT4 i19372_3_lut (.A(n29479), .B(n325), .C(index_i[3]), .Z(n21809)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19372_3_lut.init = 16'hcaca;
    LUT4 i19364_else_4_lut (.A(index_i[0]), .B(index_i[4]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n27132)) /* synthesis lut_function=(!(A (B (C)+!B !(C+!(D)))+!A (B (C)+!B (D)))) */ ;
    defparam i19364_else_4_lut.init = 16'h2c3f;
    LUT4 i21626_3_lut (.A(n21808), .B(n21809), .C(index_i[4]), .Z(n21810)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21626_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_0_i953_rep_631 (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .Z(n26954)) /* synthesis lut_function=(A (C)+!A !((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i953_rep_631.init = 16'ha4a4;
    LUT4 i11716_2_lut_rep_479_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[0]), 
         .Z(n26802)) /* synthesis lut_function=(A (C)+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11716_2_lut_rep_479_3_lut.init = 16'hf1f1;
    LUT4 mux_198_Mux_9_i93_3_lut_3_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .Z(n93)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_9_i93_3_lut_3_lut_3_lut.init = 16'hc1c1;
    LUT4 i19459_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21896)) /* synthesis lut_function=(!(A ((D)+!C)+!A !(B ((D)+!C)+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19459_3_lut_3_lut_4_lut.init = 16'h55a4;
    LUT4 mux_198_Mux_0_i781_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n781)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A (B (C)+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i781_4_lut_4_lut_4_lut.init = 16'h0cb4;
    LUT4 i4415_2_lut_rep_632 (.A(index_i[0]), .B(index_i[1]), .Z(n26955)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i4415_2_lut_rep_632.init = 16'h6666;
    LUT4 mux_198_Mux_4_i236_3_lut_4_lut_3_lut_rep_621_4_lut (.A(index_i[1]), 
         .B(index_i[2]), .C(index_i[3]), .D(index_i[0]), .Z(n26944)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_4_i236_3_lut_4_lut_3_lut_rep_621_4_lut.init = 16'hf01f;
    LUT4 mux_198_Mux_0_i588_3_lut_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n588)) /* synthesis lut_function=(!(A (B+(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i588_3_lut_3_lut_3_lut.init = 16'h5656;
    LUT4 i9443_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(n27036), .D(index_i[4]), .Z(n221)) /* synthesis lut_function=(!(A (B)+!A (B (C+(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9443_3_lut_4_lut_4_lut_4_lut.init = 16'h3336;
    LUT4 i19368_3_lut (.A(n588), .B(n26958), .C(index_i[3]), .Z(n21805)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19368_3_lut.init = 16'hcaca;
    LUT4 i19366_3_lut (.A(n900), .B(n325), .C(index_i[3]), .Z(n21803)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19366_3_lut.init = 16'hcaca;
    LUT4 n9791_bdd_3_lut_24306_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[4]), .D(index_i[3]), .Z(n24542)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C+(D)))+!A (B (C (D)+!C !(D))+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n9791_bdd_3_lut_24306_4_lut_4_lut_4_lut.init = 16'hc10f;
    LUT4 mux_198_Mux_9_i412_3_lut_3_lut_4_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .Z(n412_adj_2887)) /* synthesis lut_function=(!(A (B (C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_9_i412_3_lut_3_lut_4_lut_3_lut.init = 16'h7e7e;
    LUT4 i11185_2_lut_rep_558_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[3]), 
         .Z(n26881)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11185_2_lut_rep_558_3_lut.init = 16'he0e0;
    LUT4 i19347_3_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[3]), 
         .D(index_i[0]), .Z(n21784)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19347_3_lut_3_lut_4_lut.init = 16'h0fe0;
    LUT4 mux_198_Mux_7_i108_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n108)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_7_i108_3_lut_3_lut.init = 16'hc6c6;
    LUT4 mux_198_Mux_8_i412_3_lut_4_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .Z(n14798)) /* synthesis lut_function=(A (B+!(C))+!A !((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_8_i412_3_lut_4_lut_3_lut.init = 16'h8e8e;
    LUT4 i11186_2_lut_rep_456_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[4]), .D(index_i[3]), .Z(n26779)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11186_2_lut_rep_456_3_lut_4_lut.init = 16'hfef0;
    LUT4 mux_198_Mux_5_i828_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[4]), .D(n26966), .Z(n828_adj_2956)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_5_i828_4_lut_4_lut.init = 16'hc66c;
    LUT4 i19483_3_lut_3_lut_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[3]), 
         .Z(n21920)) /* synthesis lut_function=(A (C)+!A (B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19483_3_lut_3_lut_3_lut.init = 16'he5e5;
    LUT4 mux_198_Mux_0_i645_3_lut_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n645)) /* synthesis lut_function=(!(A (B)+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i645_3_lut_3_lut_3_lut.init = 16'h6363;
    LUT4 i19359_3_lut (.A(n29496), .B(n29484), .C(index_i[3]), .Z(n21796)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19359_3_lut.init = 16'hcaca;
    PFUMX i9427 (.BLUT(n12154), .ALUT(n12155), .C0(n22412), .Z(n11988));
    LUT4 i12144_2_lut_rep_730 (.A(index_i[2]), .B(index_i[0]), .Z(n27053)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i12144_2_lut_rep_730.init = 16'heeee;
    LUT4 mux_198_Mux_1_i882_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n882)) /* synthesis lut_function=(A ((C)+!B)+!A !((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_1_i882_3_lut_3_lut.init = 16'ha6a6;
    LUT4 mux_198_Mux_9_i125_3_lut_3_lut_4_lut_then_4_lut (.A(index_i[2]), 
         .B(index_i[4]), .C(index_i[1]), .D(index_i[0]), .Z(n27222)) /* synthesis lut_function=(!(A+((C (D))+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_9_i125_3_lut_3_lut_4_lut_then_4_lut.init = 16'h0444;
    LUT4 mux_198_Mux_2_i173_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[2]), 
         .B(index_i[0]), .C(index_i[3]), .D(index_i[1]), .Z(n173_adj_2797)) /* synthesis lut_function=(!(A (C)+!A (B (C+!(D))+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_2_i173_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h0f1a;
    LUT4 i1_2_lut_rep_557_3_lut (.A(index_i[2]), .B(index_i[0]), .C(index_i[1]), 
         .Z(n26880)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i1_2_lut_rep_557_3_lut.init = 16'hfefe;
    PFUMX i20011 (.BLUT(n22465), .ALUT(n22466), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2126[8]));
    LUT4 mux_198_Mux_8_i716_3_lut_4_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[1]), .D(index_i[3]), .Z(n716_adj_2981)) /* synthesis lut_function=(!(A (D)+!A !(B+(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_8_i716_3_lut_4_lut_4_lut_4_lut.init = 16'h55fe;
    LUT4 mux_198_Mux_5_i954_3_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[1]), .Z(n954_adj_2875)) /* synthesis lut_function=(!(A (C)+!A (B+((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_5_i954_3_lut_4_lut_4_lut.init = 16'h0a1a;
    LUT4 i11160_2_lut_rep_455_3_lut_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[1]), .Z(n26778)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11160_2_lut_rep_455_3_lut_4_lut.init = 16'hf0e0;
    LUT4 mux_198_Mux_9_i285_3_lut_3_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[1]), .Z(n285_adj_2816)) /* synthesis lut_function=(A (C)+!A !(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_9_i285_3_lut_3_lut_4_lut_4_lut.init = 16'ha0a1;
    LUT4 mux_198_Mux_0_i46_3_lut_4_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[1]), .D(index_i[3]), .Z(n46)) /* synthesis lut_function=(A (D)+!A (B+(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i46_3_lut_4_lut_4_lut_4_lut.init = 16'hfe55;
    LUT4 n172_bdd_2_lut_3_lut_3_lut_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[1]), .D(index_i[3]), .Z(n25654)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n172_bdd_2_lut_3_lut_3_lut_4_lut.init = 16'h00fe;
    LUT4 mux_198_Mux_3_i507_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[4]), .D(n491_adj_2802), .Z(n507_adj_2985)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_3_i507_3_lut_4_lut.init = 16'h6f60;
    PFUMX i20768 (.BLUT(n142_adj_2975), .ALUT(n157), .C0(index_i[4]), 
          .Z(n23224));
    PFUMX i20769 (.BLUT(n173_adj_2842), .ALUT(n188), .C0(index_i[4]), 
          .Z(n23225));
    LUT4 i20789_3_lut (.A(n23238), .B(n23239), .C(index_i[6]), .Z(n23245)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20789_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_9_i125_3_lut_3_lut_4_lut_else_4_lut (.A(index_i[2]), 
         .B(index_i[4]), .C(index_i[1]), .D(index_i[0]), .Z(n27221)) /* synthesis lut_function=(A (B+!(C))+!A ((C+(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_9_i125_3_lut_3_lut_4_lut_else_4_lut.init = 16'hdfdb;
    LUT4 n476_bdd_3_lut_24919 (.A(n476), .B(n25356), .C(index_i[5]), .Z(n25357)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n476_bdd_3_lut_24919.init = 16'hcaca;
    LUT4 mux_198_Mux_6_i442_rep_634 (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .Z(n26957)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_6_i442_rep_634.init = 16'h6464;
    LUT4 mux_198_Mux_0_i525_3_lut_3_lut_rep_635 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26958)) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i525_3_lut_3_lut_rep_635.init = 16'h6a6a;
    LUT4 mux_198_Mux_2_i491_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n491_adj_2987)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A !(B (C)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_2_i491_3_lut_4_lut_4_lut.init = 16'h6a5a;
    LUT4 i9449_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(n26968), .Z(n605_adj_2954)) /* synthesis lut_function=(!(A (B (C+(D))+!B (D))+!A !(B (C+(D))+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9449_3_lut_3_lut_4_lut.init = 16'h556a;
    LUT4 i19365_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21802)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19365_3_lut_4_lut.init = 16'h64cc;
    LUT4 n21839_bdd_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(n26966), 
         .D(index_i[4]), .Z(n25287)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+(D)))+!A (B (D)+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n21839_bdd_3_lut_3_lut_4_lut.init = 16'h336c;
    LUT4 i11403_2_lut_rep_636 (.A(index_i[0]), .B(index_i[1]), .Z(n26959)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11403_2_lut_rep_636.init = 16'h2222;
    PFUMX i20774 (.BLUT(n333_adj_2989), .ALUT(n348), .C0(index_i[4]), 
          .Z(n23230));
    LUT4 i19354_3_lut (.A(n27015), .B(n26957), .C(index_i[3]), .Z(n21791)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19354_3_lut.init = 16'hcaca;
    LUT4 i19353_3_lut (.A(n26954), .B(n325), .C(index_i[3]), .Z(n21790)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19353_3_lut.init = 16'hcaca;
    LUT4 i21636_3_lut (.A(n21790), .B(n21791), .C(index_i[4]), .Z(n21792)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21636_3_lut.init = 16'hcaca;
    LUT4 i19351_3_lut (.A(n27008), .B(n29480), .C(index_i[3]), .Z(n21788)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19351_3_lut.init = 16'hcaca;
    LUT4 i21638_3_lut (.A(n21787), .B(n21788), .C(index_i[4]), .Z(n21789)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21638_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_6_i157_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n157_adj_2909)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (D))+!A !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_6_i157_3_lut_4_lut_4_lut_4_lut.init = 16'h5d22;
    LUT4 mux_198_Mux_4_i205_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n205)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_4_i205_3_lut_4_lut_4_lut.init = 16'h5a2a;
    LUT4 i21641_3_lut (.A(n21784), .B(n21785), .C(index_i[4]), .Z(n21786)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21641_3_lut.init = 16'hcaca;
    LUT4 mux_198_Mux_0_i985_3_lut_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n985)) /* synthesis lut_function=(!(A (B+!(C))+!A (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i985_3_lut_3_lut_3_lut.init = 16'h2525;
    LUT4 i9589_3_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[4]), 
         .Z(n12154)) /* synthesis lut_function=(!(A (B)+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9589_3_lut_4_lut_3_lut.init = 16'h6262;
    LUT4 mux_198_Mux_0_i490_3_lut_4_lut_3_lut_rep_638 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26961)) /* synthesis lut_function=(!(A (B+!(C))+!A ((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i490_3_lut_4_lut_3_lut_rep_638.init = 16'h2424;
    LUT4 mux_198_Mux_5_i754_3_lut_4_lut_3_lut_rep_639 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26962)) /* synthesis lut_function=(!(A (B)+!A ((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_5_i754_3_lut_4_lut_3_lut_rep_639.init = 16'h2626;
    PFUMX i20775 (.BLUT(n364_adj_2980), .ALUT(n379), .C0(index_i[4]), 
          .Z(n23231));
    L6MUX21 i12906359_i1 (.D0(n23250), .D1(n23465), .SD(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2126[0]));
    LUT4 i19398_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21835)) /* synthesis lut_function=(!(A (B)+!A (B (C+(D))+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19398_3_lut_3_lut_4_lut.init = 16'h3326;
    LUT4 mux_198_Mux_0_i491_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n491_adj_2990)) /* synthesis lut_function=(!(A (B (D)+!B !(C+!(D)))+!A ((C+!(D))+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i491_3_lut_4_lut.init = 16'h24aa;
    LUT4 n316_bdd_3_lut_24662_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n25551)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A !(B ((D)+!C)+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n316_bdd_3_lut_24662_3_lut_4_lut.init = 16'h552c;
    LUT4 i19053_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21490)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C))+!A !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19053_3_lut_4_lut_4_lut.init = 16'h5a52;
    LUT4 i11404_2_lut_rep_640 (.A(index_i[0]), .B(index_i[1]), .Z(n26963)) /* synthesis lut_function=(A+!(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11404_2_lut_rep_640.init = 16'hbbbb;
    LUT4 i19420_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n21857)) /* synthesis lut_function=(A (C+(D))+!A !(B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19420_3_lut_4_lut_4_lut.init = 16'haba5;
    LUT4 mux_198_Mux_5_i781_3_lut_4_lut_4_lut_then_4_lut (.A(index_i[3]), 
         .B(index_i[0]), .C(index_i[4]), .D(index_i[2]), .Z(n27139)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_5_i781_3_lut_4_lut_4_lut_then_4_lut.init = 16'hece0;
    LUT4 mux_198_Mux_4_i900_3_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n900)) /* synthesis lut_function=(A ((C)+!B)+!A !(B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_4_i900_3_lut_4_lut_3_lut.init = 16'hb2b2;
    LUT4 n72_bdd_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n25713)) /* synthesis lut_function=(!(A (D)+!A !(B (D)+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n72_bdd_4_lut_4_lut_4_lut.init = 16'h54bb;
    LUT4 i23085_then_4_lut (.A(index_i[0]), .B(index_i[4]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n27225)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)+!C !(D))+!B (C (D)))) */ ;
    defparam i23085_then_4_lut.init = 16'hda0e;
    LUT4 i23085_else_4_lut (.A(index_i[0]), .B(index_i[4]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n27224)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C))+!A (B (C)+!B (C+(D)))) */ ;
    defparam i23085_else_4_lut.init = 16'hf178;
    LUT4 mux_198_Mux_6_i70_3_lut_rep_807 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29480)) /* synthesis lut_function=(!(A (B+(C))+!A !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_6_i70_3_lut_rep_807.init = 16'h5252;
    LUT4 mux_198_Mux_6_i332_3_lut_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n332)) /* synthesis lut_function=(!(A (C)+!A !((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_6_i332_3_lut_3_lut_3_lut.init = 16'h5b5b;
    LUT4 mux_198_Mux_5_i459_3_lut_4_lut_3_lut_rep_641 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26964)) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_5_i459_3_lut_4_lut_3_lut_rep_641.init = 16'h6b6b;
    LUT4 mux_198_Mux_5_i460_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n460_adj_2905)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A !(B (C)+!B !(C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_5_i460_3_lut_4_lut_4_lut.init = 16'h6b5a;
    LUT4 mux_198_Mux_4_i142_3_lut_3_lut_3_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[3]), .Z(n142_adj_2946)) /* synthesis lut_function=(A (B (C))+!A !(B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_4_i142_3_lut_3_lut_3_lut.init = 16'h9595;
    PFUMX i20776 (.BLUT(n397), .ALUT(n412), .C0(index_i[4]), .Z(n23232));
    PFUMX i20087 (.BLUT(n22541), .ALUT(n22542), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2126[2]));
    LUT4 n17999_bdd_4_lut_then_4_lut (.A(index_i[3]), .B(index_i[4]), .C(index_i[1]), 
         .D(index_i[2]), .Z(n27147)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B+(C (D)+!C !(D)))) */ ;
    defparam n17999_bdd_4_lut_then_4_lut.init = 16'hf44f;
    LUT4 i11209_4_lut (.A(n26878), .B(index_i[7]), .C(n892_adj_2868), 
         .D(index_i[6]), .Z(n1021)) /* synthesis lut_function=(A (B+(C (D)))+!A (B+(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11209_4_lut.init = 16'hfcdd;
    PFUMX i20777 (.BLUT(n428), .ALUT(n443), .C0(index_i[4]), .Z(n23233));
    LUT4 mux_198_Mux_0_i236_3_lut_3_lut_rep_642 (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[3]), .Z(n26965)) /* synthesis lut_function=(A (B+(C))+!A !(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i236_3_lut_3_lut_rep_642.init = 16'ha9a9;
    PFUMX i20094 (.BLUT(n22548), .ALUT(n22549), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2126[9]));
    PFUMX i20778 (.BLUT(n460), .ALUT(n475_adj_2801), .C0(index_i[4]), 
          .Z(n23234));
    LUT4 mux_198_Mux_4_i812_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[4]), .Z(n812_adj_2982)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A !(B (D)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_4_i812_3_lut_3_lut_4_lut.init = 16'ha955;
    LUT4 i11191_2_lut_rep_643 (.A(index_i[2]), .B(index_i[3]), .Z(n26966)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11191_2_lut_rep_643.init = 16'heeee;
    LUT4 n61_bdd_3_lut_24365_3_lut_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n25753)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n61_bdd_3_lut_24365_3_lut_3_lut_4_lut.init = 16'h0fe1;
    PFUMX i20779 (.BLUT(n491_adj_2990), .ALUT(n11109), .C0(index_i[4]), 
          .Z(n23235));
    LUT4 i9429_3_lut_3_lut_rep_633_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n26956)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9429_3_lut_3_lut_rep_633_4_lut.init = 16'h1ef0;
    LUT4 i11725_2_lut_rep_515_3_lut (.A(index_i[2]), .B(index_i[3]), .C(index_i[1]), 
         .Z(n26838)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11725_2_lut_rep_515_3_lut.init = 16'hfefe;
    PFUMX i19091 (.BLUT(n21526), .ALUT(n21527), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2126[11]));
    LUT4 i20790_3_lut (.A(n25556), .B(n23241), .C(index_i[6]), .Z(n23246)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20790_3_lut.init = 16'hcaca;
    LUT4 i9448_2_lut_rep_645 (.A(index_i[3]), .B(index_i[4]), .Z(n26968)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9448_2_lut_rep_645.init = 16'heeee;
    LUT4 i1_3_lut_rep_521_4_lut (.A(index_i[3]), .B(index_i[4]), .C(index_i[2]), 
         .D(n27037), .Z(n26844)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i1_3_lut_rep_521_4_lut.init = 16'hfffe;
    LUT4 i1_3_lut_4_lut_adj_91 (.A(index_i[3]), .B(index_i[4]), .C(index_i[5]), 
         .D(n27050), .Z(n20328)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i1_3_lut_4_lut_adj_91.init = 16'hfffe;
    LUT4 i9433_3_lut_4_lut (.A(index_i[3]), .B(index_i[4]), .C(n27009), 
         .D(n29496), .Z(n605_adj_2941)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9433_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i20079_3_lut (.A(n26036), .B(n22526), .C(index_i[6]), .Z(n22535)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20079_3_lut.init = 16'hcaca;
    LUT4 i11401_2_lut_rep_646 (.A(index_i[0]), .B(index_i[1]), .Z(n26969)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11401_2_lut_rep_646.init = 16'heeee;
    LUT4 mux_198_Mux_8_i506_3_lut_4_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n506_adj_2866)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_8_i506_3_lut_4_lut_3_lut_4_lut.init = 16'h0ef0;
    LUT4 mux_198_Mux_3_i157_3_lut_3_lut_rep_438_3_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n26761)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_3_i157_3_lut_3_lut_rep_438_3_lut_4_lut.init = 16'h1ff0;
    LUT4 mux_198_Mux_2_i142_3_lut_4_lut_4_lut_4_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n142_adj_2891)) /* synthesis lut_function=(!(A (B (D)+!B (C (D)+!C !(D)))+!A (B (D)+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_2_i142_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'h03ec;
    PFUMX i22887 (.BLUT(n21586), .ALUT(n24540), .C0(index_i[6]), .Z(n24541));
    L6MUX21 i23970 (.D0(n25766), .D1(n25763), .SD(index_i[5]), .Z(n25767));
    LUT4 mux_198_Mux_6_i860_3_lut_3_lut (.A(n26750), .B(index_i[4]), .C(n844_adj_2869), 
         .Z(n860_adj_2945)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam mux_198_Mux_6_i860_3_lut_3_lut.init = 16'h7474;
    PFUMX i23968 (.BLUT(n25765), .ALUT(n25764), .C0(index_i[4]), .Z(n25766));
    LUT4 n348_bdd_3_lut_24243_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n26031)) /* synthesis lut_function=(A (B (C)+!B (C+(D)))+!A (B (C)+!B !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n348_bdd_3_lut_24243_4_lut_4_lut_4_lut.init = 16'he3f0;
    LUT4 i12094_1_lut_rep_406_2_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n26729)) /* synthesis lut_function=(!(A (C+(D))+!A (B (C+(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i12094_1_lut_rep_406_2_lut_3_lut_4_lut.init = 16'h010f;
    LUT4 i22376_3_lut (.A(n11942), .B(n892), .C(index_i[6]), .Z(n22459)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22376_3_lut.init = 16'hcaca;
    LUT4 i11150_2_lut_rep_514_3_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .Z(n26837)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11150_2_lut_rep_514_3_lut.init = 16'he0e0;
    LUT4 i19404_3_lut_3_lut_4_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n21841)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19404_3_lut_3_lut_4_lut_3_lut_4_lut.init = 16'h11ef;
    LUT4 i11195_2_lut_rep_437_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n26760)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11195_2_lut_rep_437_3_lut_4_lut.init = 16'hfef0;
    PFUMX i23965 (.BLUT(n25762), .ALUT(n26754), .C0(index_i[4]), .Z(n25763));
    LUT4 mux_198_Mux_8_i460_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n460_adj_2817)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_8_i460_3_lut_3_lut_4_lut.init = 16'hf10f;
    L6MUX21 i23956 (.D0(n25754), .D1(n25752), .SD(index_i[4]), .Z(n25755));
    LUT4 mux_198_Mux_8_i46_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n46_adj_2849)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (B (C)+!B !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_8_i46_3_lut_4_lut_4_lut_4_lut.init = 16'hc1f0;
    PFUMX i23954 (.BLUT(n26755), .ALUT(n25753), .C0(index_i[5]), .Z(n25754));
    LUT4 i11377_3_lut_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n14052)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11377_3_lut_3_lut_3_lut_4_lut.init = 16'h10ff;
    LUT4 mux_198_Mux_5_i781_3_lut_4_lut_4_lut_else_4_lut (.A(index_i[3]), 
         .B(index_i[0]), .C(index_i[4]), .Z(n27138)) /* synthesis lut_function=(!(A (C)+!A (B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_5_i781_3_lut_4_lut_4_lut_else_4_lut.init = 16'h1f1f;
    LUT4 mux_198_Mux_11_i766_3_lut (.A(n638), .B(n765), .C(index_i[7]), 
         .Z(n766)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_11_i766_3_lut.init = 16'h3a3a;
    LUT4 mux_198_Mux_3_i30_3_lut_3_lut_4_lut_3_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n30)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_3_i30_3_lut_3_lut_4_lut_3_lut_4_lut.init = 16'hfe11;
    LUT4 i11397_2_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n635_adj_2837)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A (B (C+!(D))+!B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11397_2_lut_4_lut_4_lut.init = 16'hf1fc;
    LUT4 mux_198_Mux_0_i333_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n333_adj_2989)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i333_3_lut_3_lut_4_lut.init = 16'hf10e;
    LUT4 mux_198_Mux_7_i572_3_lut_rep_399_3_lut_3_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n26722)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_7_i572_3_lut_rep_399_3_lut_3_lut_4_lut.init = 16'hfe01;
    LUT4 i19441_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n21878)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B ((D)+!C)+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19441_3_lut_4_lut_4_lut.init = 16'hfc1c;
    PFUMX i23952 (.BLUT(n25751), .ALUT(n25750), .C0(index_i[5]), .Z(n25752));
    LUT4 mux_198_Mux_0_i915_3_lut_rep_625_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26948)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i915_3_lut_rep_625_3_lut.init = 16'he3e3;
    LUT4 i19171_3_lut_3_lut (.A(n26750), .B(index_i[4]), .C(n46_adj_2849), 
         .Z(n21608)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam i19171_3_lut_3_lut.init = 16'h7474;
    LUT4 mux_198_Mux_2_i716_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n716_adj_2881)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)+!C !(D)))+!A (B (D)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_2_i716_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h31cf;
    LUT4 n273_bdd_3_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .Z(n26339)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n273_bdd_3_lut_4_lut_3_lut.init = 16'h6161;
    LUT4 mux_198_Mux_8_i101_3_lut_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n101)) /* synthesis lut_function=(!(A (B (C))+!A (B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_8_i101_3_lut_3_lut_3_lut.init = 16'h3e3e;
    LUT4 mux_198_Mux_9_i62_3_lut_4_lut_then_4_lut (.A(index_i[4]), .B(index_i[2]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n27234)) /* synthesis lut_function=(!(A (B (C+(D)))+!A (B+(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_9_i62_3_lut_4_lut_then_4_lut.init = 16'h222b;
    LUT4 i11198_2_lut_rep_442_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[4]), .D(n27036), .Z(n26765)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11198_2_lut_rep_442_3_lut_4_lut.init = 16'hfef0;
    LUT4 mux_198_Mux_7_i924_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[4]), .D(n27036), .Z(n924_adj_2991)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_7_i924_3_lut_3_lut_4_lut.init = 16'hf10f;
    LUT4 mux_198_Mux_0_i15_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n15_adj_2936)) /* synthesis lut_function=(A (B (D)+!B (C+!(D)))+!A (B (D)+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i15_3_lut_4_lut_4_lut_4_lut.init = 16'hec33;
    LUT4 i19431_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n21868)) /* synthesis lut_function=(A (B (D)+!B ((D)+!C))+!A (B (D)+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19431_3_lut_4_lut_4_lut_4_lut.init = 16'hfe13;
    LUT4 mux_198_Mux_8_i45_3_lut_rep_647 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26970)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_8_i45_3_lut_rep_647.init = 16'hc1c1;
    LUT4 mux_198_Mux_5_i53_3_lut_4_lut_3_lut_rep_648 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26971)) /* synthesis lut_function=(A ((C)+!B)+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_5_i53_3_lut_4_lut_3_lut_rep_648.init = 16'he6e6;
    LUT4 mux_198_Mux_0_i698_3_lut_rep_649 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26972)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i698_3_lut_rep_649.init = 16'h1c1c;
    LUT4 i19464_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21901)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C (D)))+!A (B (C+(D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19464_4_lut_4_lut_4_lut.init = 16'h301c;
    LUT4 i19387_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21824)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19387_3_lut_3_lut_4_lut.init = 16'h0f1c;
    LUT4 mux_198_Mux_0_i699_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n699_adj_2811)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (D))+!A (B (C+!(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i699_3_lut_3_lut_4_lut.init = 16'h1c33;
    LUT4 mux_198_Mux_0_i557_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n557)) /* synthesis lut_function=(A ((D)+!C)+!A !((D)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_0_i557_3_lut_4_lut.init = 16'haa4e;
    PFUMX i15527 (.BLUT(n17789), .ALUT(n17790), .C0(index_i[4]), .Z(n17791));
    LUT4 mux_198_Mux_6_i635_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n635_adj_2914)) /* synthesis lut_function=(A (B (C+(D))+!B !(D))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_6_i635_3_lut_4_lut.init = 16'hcce6;
    LUT4 n22_bdd_3_lut_23720_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n25514)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C (D)+!C !(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n22_bdd_3_lut_23720_3_lut_4_lut.init = 16'h0fc1;
    PFUMX i23066 (.BLUT(n24774), .ALUT(n24773), .C0(index_i[6]), .Z(n24775));
    LUT4 mux_198_Mux_9_i62_3_lut_4_lut_else_4_lut (.A(index_i[4]), .B(index_i[2]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n27233)) /* synthesis lut_function=((B+(C (D)))+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_9_i62_3_lut_4_lut_else_4_lut.init = 16'hfddd;
    PFUMX i24747 (.BLUT(n27150), .ALUT(n27151), .C0(index_i[1]), .Z(n27152));
    LUT4 n25359_bdd_3_lut (.A(n27128), .B(n444_adj_2988), .C(index_i[5]), 
         .Z(n25360)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n25359_bdd_3_lut.init = 16'hcaca;
    PFUMX i23913 (.BLUT(n25713), .ALUT(n26941), .C0(index_i[4]), .Z(n25714));
    LUT4 i21008_3_lut (.A(n23461), .B(n23462), .C(index_i[7]), .Z(n23464)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21008_3_lut.init = 16'hcaca;
    PFUMX i20484 (.BLUT(n22936), .ALUT(n22937), .C0(index_i[4]), .Z(n22940));
    LUT4 i21007_3_lut (.A(n23459), .B(n23460), .C(index_i[7]), .Z(n23463)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21007_3_lut.init = 16'hcaca;
    LUT4 index_i_0__bdd_4_lut_25198 (.A(index_i[0]), .B(index_i[3]), .C(index_i[1]), 
         .D(index_i[2]), .Z(n27142)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C))+!A (B (C (D)+!C !(D))+!B !(C+!(D))))) */ ;
    defparam index_i_0__bdd_4_lut_25198.init = 16'h16d3;
    LUT4 i22492_3_lut (.A(n24549), .B(n22547), .C(index_i[8]), .Z(n22549)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22492_3_lut.init = 16'hcaca;
    PFUMX i20485 (.BLUT(n22938), .ALUT(n22939), .C0(index_i[4]), .Z(n22941));
    LUT4 mux_198_Mux_5_i109_3_lut_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .Z(n109_adj_2910)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_5_i109_3_lut_3_lut_3_lut.init = 16'h3939;
    PFUMX i20491 (.BLUT(n22943), .ALUT(n22944), .C0(index_i[4]), .Z(n22947));
    PFUMX i23871 (.BLUT(n25655), .ALUT(n25654), .C0(index_i[4]), .Z(n25656));
    PFUMX i20492 (.BLUT(n22945), .ALUT(n22946), .C0(index_i[4]), .Z(n22948));
    PFUMX i24745 (.BLUT(n27146), .ALUT(n27147), .C0(index_i[0]), .Z(n27148));
    LUT4 i19149_3_lut_3_lut_4_lut (.A(n26868), .B(index_i[4]), .C(n700), 
         .D(index_i[5]), .Z(n21586)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19149_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 n773_bdd_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n25023)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n773_bdd_3_lut_4_lut_4_lut.init = 16'ha5ad;
    PFUMX i20498 (.BLUT(n22950), .ALUT(n22951), .C0(index_i[4]), .Z(n22954));
    PFUMX i20979 (.BLUT(n526), .ALUT(n541), .C0(index_i[4]), .Z(n23435));
    PFUMX mux_198_Mux_13_i1023 (.BLUT(n511), .ALUT(n20196), .C0(index_i[9]), 
          .Z(quarter_wave_sample_register_i_15__N_2126[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    PFUMX i20499 (.BLUT(n22952), .ALUT(n22953), .C0(index_i[4]), .Z(n22955));
    PFUMX i20505 (.BLUT(n22957), .ALUT(n22958), .C0(index_i[4]), .Z(n22961));
    PFUMX i20506 (.BLUT(n22959), .ALUT(n22960), .C0(index_i[4]), .Z(n22962));
    L6MUX21 i23017 (.D0(n24718), .D1(n26708), .SD(index_i[6]), .Z(n24719));
    PFUMX i23015 (.BLUT(n24717), .ALUT(n26735), .C0(index_i[7]), .Z(n24718));
    LUT4 mux_198_Mux_10_i701_4_lut_4_lut (.A(n26868), .B(index_i[4]), .C(index_i[5]), 
         .D(n26780), .Z(n701)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B (C (D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_10_i701_4_lut_4_lut.init = 16'h3efe;
    L6MUX21 i23762 (.D0(n25555), .D1(n25552), .SD(index_i[5]), .Z(n25556));
    PFUMX i23760 (.BLUT(n25554), .ALUT(n25553), .C0(index_i[4]), .Z(n25555));
    PFUMX i23757 (.BLUT(n25551), .ALUT(n316_adj_2790), .C0(index_i[4]), 
          .Z(n25552));
    L6MUX21 i23723 (.D0(n25516), .D1(n25513), .SD(index_i[5]), .Z(n25517));
    PFUMX i23721 (.BLUT(n25515), .ALUT(n25514), .C0(index_i[4]), .Z(n25516));
    LUT4 i20006_3_lut (.A(n22455), .B(n22456), .C(index_i[7]), .Z(n22462)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20006_3_lut.init = 16'hcaca;
    FD1S3BX quarter_wave_sample_register_i_i14 (.D(quarter_wave_sample_register_i_15__N_2126[14]), 
            .CK(dac_clk_p_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_i[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i14.GSR = "DISABLED";
    PFUMX i23718 (.BLUT(n301), .ALUT(n25512), .C0(index_i[4]), .Z(n25513));
    LUT4 i19434_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21871)) /* synthesis lut_function=(!(A (B (C (D))+!B (C (D)+!C !(D)))+!A !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19434_3_lut_4_lut_4_lut.init = 16'h5aad;
    LUT4 mux_198_Mux_7_i956_3_lut_3_lut_4_lut (.A(n26868), .B(index_i[4]), 
         .C(n924_adj_2991), .D(index_i[5]), .Z(n956)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_198_Mux_7_i956_3_lut_3_lut_4_lut.init = 16'h11f0;
    L6MUX21 i22988 (.D0(n24687), .D1(n24685), .SD(index_i[6]), .Z(n24688));
    PFUMX i22986 (.BLUT(n924_adj_2971), .ALUT(n24686), .C0(index_i[5]), 
          .Z(n24687));
    FD1S3BX quarter_wave_sample_register_i_i13 (.D(quarter_wave_sample_register_i_15__N_2126[13]), 
            .CK(dac_clk_p_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_i[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i13.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i12 (.D(quarter_wave_sample_register_i_15__N_2126[12]), 
            .CK(dac_clk_p_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_i[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i12.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i11 (.D(quarter_wave_sample_register_i_15__N_2126[11]), 
            .CK(dac_clk_p_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_i[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i11.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i10 (.D(quarter_wave_sample_register_i_15__N_2126[10]), 
            .CK(dac_clk_p_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_i[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i10.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i9 (.D(quarter_wave_sample_register_i_15__N_2126[9]), 
            .CK(dac_clk_p_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_i[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i9.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i8 (.D(quarter_wave_sample_register_i_15__N_2126[8]), 
            .CK(dac_clk_p_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_i[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i8.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i7 (.D(quarter_wave_sample_register_i_15__N_2126[7]), 
            .CK(dac_clk_p_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_i[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i7.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i6 (.D(quarter_wave_sample_register_i_15__N_2126[6]), 
            .CK(dac_clk_p_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_i[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i6.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i5 (.D(quarter_wave_sample_register_i_15__N_2126[5]), 
            .CK(dac_clk_p_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_i[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i5.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i4 (.D(quarter_wave_sample_register_i_15__N_2126[4]), 
            .CK(dac_clk_p_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_i[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i4.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i3 (.D(quarter_wave_sample_register_i_15__N_2126[3]), 
            .CK(dac_clk_p_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_i[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i3.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i2 (.D(quarter_wave_sample_register_i_15__N_2126[2]), 
            .CK(dac_clk_p_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_i[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i2.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i1 (.D(quarter_wave_sample_register_i_15__N_2126[1]), 
            .CK(dac_clk_p_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_i[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i1.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i32 (.D(n1212[15]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(\o_val_pipeline_i[0] [15])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i32.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i31 (.D(n1212[14]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(\o_val_pipeline_i[0] [14])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i31.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i30 (.D(n1212[13]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(\o_val_pipeline_i[0] [13])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i30.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i29 (.D(n1212[12]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(\o_val_pipeline_i[0] [12])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i29.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i28 (.D(n1212[11]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(\o_val_pipeline_i[0] [11])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i28.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i27 (.D(n1212[10]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(\o_val_pipeline_i[0] [10])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i27.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i26 (.D(n1212[9]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(\o_val_pipeline_i[0] [9])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i26.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i25 (.D(n1212[8]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(\o_val_pipeline_i[0] [8])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i25.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i24 (.D(n1212[7]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(\o_val_pipeline_i[0] [7])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i24.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i23 (.D(n1212[6]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(\o_val_pipeline_i[0] [6])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i23.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i22 (.D(n1212[5]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(\o_val_pipeline_i[0] [5])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i22.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i21 (.D(n1212[4]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(\o_val_pipeline_i[0] [4])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i21.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i20 (.D(n1212[3]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(\o_val_pipeline_i[0] [3])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i20.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i19 (.D(n1212[2]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(\o_val_pipeline_i[0] [2])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i19.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i18 (.D(n1212[1]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(\o_val_pipeline_i[0] [1])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i18.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i17 (.D(n1212[0]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(\o_val_pipeline_i[0] [0])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i17.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i16 (.D(\o_val_pipeline_i[0] [15]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(modulation_output[15])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i16.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i15 (.D(\o_val_pipeline_i[0] [14]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(modulation_output[14])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i15.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i14 (.D(\o_val_pipeline_i[0] [13]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(modulation_output[13])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i14.GSR = "DISABLED";
    PFUMX i22984 (.BLUT(n24684), .ALUT(n26844), .C0(index_i[5]), .Z(n24685));
    
endmodule
//
// Verilog Description of module \nco(OW=12) 
//

module \nco(OW=12)  (dac_clk_p_c, i_resetb_N_301, increment, o_phase, 
            GND_net) /* synthesis syn_module_defined=1 */ ;
    input dac_clk_p_c;
    input i_resetb_N_301;
    input [30:0]increment;
    output [11:0]o_phase;
    input GND_net;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(28[49:58])
    wire [31:0]n233;
    wire [31:0]n133;
    
    wire n17690, n17689, n17688, n17687, n17686, n17685, n17684, 
        n17683, n17682, n17681, n17680, n17679, n17678, n17677, 
        n17676;
    
    FD1S3DX phase_register_549__i0 (.D(n133[0]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(n233[0])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_549__i0.GSR = "DISABLED";
    LUT4 i15479_2_lut (.A(increment[0]), .B(n233[0]), .Z(n133[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i15479_2_lut.init = 16'h6666;
    CCU2D phase_register_549_add_4_32 (.A0(increment[30]), .B0(o_phase[10]), 
          .C0(GND_net), .D0(GND_net), .A1(o_phase[11]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n17690), .S0(n133[30]), .S1(n133[31]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_549_add_4_32.INIT0 = 16'h5666;
    defparam phase_register_549_add_4_32.INIT1 = 16'hfaaa;
    defparam phase_register_549_add_4_32.INJECT1_0 = "NO";
    defparam phase_register_549_add_4_32.INJECT1_1 = "NO";
    CCU2D phase_register_549_add_4_30 (.A0(increment[28]), .B0(o_phase[8]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[29]), .B1(o_phase[9]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17689), .COUT(n17690), .S0(n133[28]), 
          .S1(n133[29]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_549_add_4_30.INIT0 = 16'h5666;
    defparam phase_register_549_add_4_30.INIT1 = 16'h5666;
    defparam phase_register_549_add_4_30.INJECT1_0 = "NO";
    defparam phase_register_549_add_4_30.INJECT1_1 = "NO";
    CCU2D phase_register_549_add_4_28 (.A0(increment[26]), .B0(o_phase[6]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[27]), .B1(o_phase[7]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17688), .COUT(n17689), .S0(n133[26]), 
          .S1(n133[27]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_549_add_4_28.INIT0 = 16'h5666;
    defparam phase_register_549_add_4_28.INIT1 = 16'h5666;
    defparam phase_register_549_add_4_28.INJECT1_0 = "NO";
    defparam phase_register_549_add_4_28.INJECT1_1 = "NO";
    CCU2D phase_register_549_add_4_26 (.A0(increment[24]), .B0(o_phase[4]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[25]), .B1(o_phase[5]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17687), .COUT(n17688), .S0(n133[24]), 
          .S1(n133[25]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_549_add_4_26.INIT0 = 16'h5666;
    defparam phase_register_549_add_4_26.INIT1 = 16'h5666;
    defparam phase_register_549_add_4_26.INJECT1_0 = "NO";
    defparam phase_register_549_add_4_26.INJECT1_1 = "NO";
    CCU2D phase_register_549_add_4_24 (.A0(increment[22]), .B0(o_phase[2]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[23]), .B1(o_phase[3]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17686), .COUT(n17687), .S0(n133[22]), 
          .S1(n133[23]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_549_add_4_24.INIT0 = 16'h5666;
    defparam phase_register_549_add_4_24.INIT1 = 16'h5666;
    defparam phase_register_549_add_4_24.INJECT1_0 = "NO";
    defparam phase_register_549_add_4_24.INJECT1_1 = "NO";
    CCU2D phase_register_549_add_4_22 (.A0(increment[20]), .B0(o_phase[0]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[21]), .B1(o_phase[1]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17685), .COUT(n17686), .S0(n133[20]), 
          .S1(n133[21]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_549_add_4_22.INIT0 = 16'h5666;
    defparam phase_register_549_add_4_22.INIT1 = 16'h5666;
    defparam phase_register_549_add_4_22.INJECT1_0 = "NO";
    defparam phase_register_549_add_4_22.INJECT1_1 = "NO";
    CCU2D phase_register_549_add_4_20 (.A0(increment[18]), .B0(n233[18]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[19]), .B1(n233[19]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17684), .COUT(n17685), .S0(n133[18]), 
          .S1(n133[19]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_549_add_4_20.INIT0 = 16'h5666;
    defparam phase_register_549_add_4_20.INIT1 = 16'h5666;
    defparam phase_register_549_add_4_20.INJECT1_0 = "NO";
    defparam phase_register_549_add_4_20.INJECT1_1 = "NO";
    CCU2D phase_register_549_add_4_18 (.A0(increment[16]), .B0(n233[16]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[17]), .B1(n233[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17683), .COUT(n17684), .S0(n133[16]), 
          .S1(n133[17]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_549_add_4_18.INIT0 = 16'h5666;
    defparam phase_register_549_add_4_18.INIT1 = 16'h5666;
    defparam phase_register_549_add_4_18.INJECT1_0 = "NO";
    defparam phase_register_549_add_4_18.INJECT1_1 = "NO";
    CCU2D phase_register_549_add_4_16 (.A0(increment[14]), .B0(n233[14]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[15]), .B1(n233[15]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17682), .COUT(n17683), .S0(n133[14]), 
          .S1(n133[15]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_549_add_4_16.INIT0 = 16'h5666;
    defparam phase_register_549_add_4_16.INIT1 = 16'h5666;
    defparam phase_register_549_add_4_16.INJECT1_0 = "NO";
    defparam phase_register_549_add_4_16.INJECT1_1 = "NO";
    CCU2D phase_register_549_add_4_14 (.A0(increment[12]), .B0(n233[12]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[13]), .B1(n233[13]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17681), .COUT(n17682), .S0(n133[12]), 
          .S1(n133[13]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_549_add_4_14.INIT0 = 16'h5666;
    defparam phase_register_549_add_4_14.INIT1 = 16'h5666;
    defparam phase_register_549_add_4_14.INJECT1_0 = "NO";
    defparam phase_register_549_add_4_14.INJECT1_1 = "NO";
    CCU2D phase_register_549_add_4_12 (.A0(increment[10]), .B0(n233[10]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[11]), .B1(n233[11]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17680), .COUT(n17681), .S0(n133[10]), 
          .S1(n133[11]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_549_add_4_12.INIT0 = 16'h5666;
    defparam phase_register_549_add_4_12.INIT1 = 16'h5666;
    defparam phase_register_549_add_4_12.INJECT1_0 = "NO";
    defparam phase_register_549_add_4_12.INJECT1_1 = "NO";
    CCU2D phase_register_549_add_4_10 (.A0(increment[8]), .B0(n233[8]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[9]), .B1(n233[9]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17679), .COUT(n17680), .S0(n133[8]), 
          .S1(n133[9]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_549_add_4_10.INIT0 = 16'h5666;
    defparam phase_register_549_add_4_10.INIT1 = 16'h5666;
    defparam phase_register_549_add_4_10.INJECT1_0 = "NO";
    defparam phase_register_549_add_4_10.INJECT1_1 = "NO";
    CCU2D phase_register_549_add_4_8 (.A0(increment[6]), .B0(n233[6]), .C0(GND_net), 
          .D0(GND_net), .A1(increment[7]), .B1(n233[7]), .C1(GND_net), 
          .D1(GND_net), .CIN(n17678), .COUT(n17679), .S0(n133[6]), .S1(n133[7]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_549_add_4_8.INIT0 = 16'h5666;
    defparam phase_register_549_add_4_8.INIT1 = 16'h5666;
    defparam phase_register_549_add_4_8.INJECT1_0 = "NO";
    defparam phase_register_549_add_4_8.INJECT1_1 = "NO";
    CCU2D phase_register_549_add_4_6 (.A0(increment[4]), .B0(n233[4]), .C0(GND_net), 
          .D0(GND_net), .A1(increment[5]), .B1(n233[5]), .C1(GND_net), 
          .D1(GND_net), .CIN(n17677), .COUT(n17678), .S0(n133[4]), .S1(n133[5]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_549_add_4_6.INIT0 = 16'h5666;
    defparam phase_register_549_add_4_6.INIT1 = 16'h5666;
    defparam phase_register_549_add_4_6.INJECT1_0 = "NO";
    defparam phase_register_549_add_4_6.INJECT1_1 = "NO";
    CCU2D phase_register_549_add_4_4 (.A0(increment[2]), .B0(n233[2]), .C0(GND_net), 
          .D0(GND_net), .A1(increment[3]), .B1(n233[3]), .C1(GND_net), 
          .D1(GND_net), .CIN(n17676), .COUT(n17677), .S0(n133[2]), .S1(n133[3]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_549_add_4_4.INIT0 = 16'h5666;
    defparam phase_register_549_add_4_4.INIT1 = 16'h5666;
    defparam phase_register_549_add_4_4.INJECT1_0 = "NO";
    defparam phase_register_549_add_4_4.INJECT1_1 = "NO";
    CCU2D phase_register_549_add_4_2 (.A0(increment[0]), .B0(n233[0]), .C0(GND_net), 
          .D0(GND_net), .A1(increment[1]), .B1(n233[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n17676), .S1(n133[1]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_549_add_4_2.INIT0 = 16'h7000;
    defparam phase_register_549_add_4_2.INIT1 = 16'h5666;
    defparam phase_register_549_add_4_2.INJECT1_0 = "NO";
    defparam phase_register_549_add_4_2.INJECT1_1 = "NO";
    FD1S3DX phase_register_549__i31 (.D(n133[31]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(o_phase[11])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_549__i31.GSR = "DISABLED";
    FD1S3DX phase_register_549__i30 (.D(n133[30]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(o_phase[10])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_549__i30.GSR = "DISABLED";
    FD1S3DX phase_register_549__i29 (.D(n133[29]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(o_phase[9])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_549__i29.GSR = "DISABLED";
    FD1S3DX phase_register_549__i28 (.D(n133[28]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(o_phase[8])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_549__i28.GSR = "DISABLED";
    FD1S3DX phase_register_549__i27 (.D(n133[27]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(o_phase[7])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_549__i27.GSR = "DISABLED";
    FD1S3DX phase_register_549__i26 (.D(n133[26]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(o_phase[6])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_549__i26.GSR = "DISABLED";
    FD1S3DX phase_register_549__i25 (.D(n133[25]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(o_phase[5])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_549__i25.GSR = "DISABLED";
    FD1S3DX phase_register_549__i24 (.D(n133[24]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(o_phase[4])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_549__i24.GSR = "DISABLED";
    FD1S3DX phase_register_549__i23 (.D(n133[23]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(o_phase[3])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_549__i23.GSR = "DISABLED";
    FD1S3DX phase_register_549__i22 (.D(n133[22]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(o_phase[2])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_549__i22.GSR = "DISABLED";
    FD1S3DX phase_register_549__i21 (.D(n133[21]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(o_phase[1])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_549__i21.GSR = "DISABLED";
    FD1S3DX phase_register_549__i20 (.D(n133[20]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(o_phase[0])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_549__i20.GSR = "DISABLED";
    FD1S3DX phase_register_549__i19 (.D(n133[19]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(n233[19])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_549__i19.GSR = "DISABLED";
    FD1S3DX phase_register_549__i18 (.D(n133[18]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(n233[18])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_549__i18.GSR = "DISABLED";
    FD1S3DX phase_register_549__i17 (.D(n133[17]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(n233[17])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_549__i17.GSR = "DISABLED";
    FD1S3DX phase_register_549__i16 (.D(n133[16]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(n233[16])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_549__i16.GSR = "DISABLED";
    FD1S3DX phase_register_549__i15 (.D(n133[15]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(n233[15])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_549__i15.GSR = "DISABLED";
    FD1S3DX phase_register_549__i14 (.D(n133[14]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(n233[14])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_549__i14.GSR = "DISABLED";
    FD1S3DX phase_register_549__i13 (.D(n133[13]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(n233[13])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_549__i13.GSR = "DISABLED";
    FD1S3DX phase_register_549__i12 (.D(n133[12]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(n233[12])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_549__i12.GSR = "DISABLED";
    FD1S3DX phase_register_549__i11 (.D(n133[11]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(n233[11])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_549__i11.GSR = "DISABLED";
    FD1S3DX phase_register_549__i10 (.D(n133[10]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(n233[10])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_549__i10.GSR = "DISABLED";
    FD1S3DX phase_register_549__i9 (.D(n133[9]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(n233[9])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_549__i9.GSR = "DISABLED";
    FD1S3DX phase_register_549__i8 (.D(n133[8]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(n233[8])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_549__i8.GSR = "DISABLED";
    FD1S3DX phase_register_549__i7 (.D(n133[7]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(n233[7])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_549__i7.GSR = "DISABLED";
    FD1S3DX phase_register_549__i6 (.D(n133[6]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(n233[6])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_549__i6.GSR = "DISABLED";
    FD1S3DX phase_register_549__i5 (.D(n133[5]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(n233[5])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_549__i5.GSR = "DISABLED";
    FD1S3DX phase_register_549__i4 (.D(n133[4]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(n233[4])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_549__i4.GSR = "DISABLED";
    FD1S3DX phase_register_549__i3 (.D(n133[3]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(n233[3])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_549__i3.GSR = "DISABLED";
    FD1S3DX phase_register_549__i2 (.D(n133[2]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(n233[2])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_549__i2.GSR = "DISABLED";
    FD1S3DX phase_register_549__i1 (.D(n133[1]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(n233[1])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_549__i1.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module dds_U2
//

module dds_U2 (dac_clk_p_c, i_resetb_N_301, carrier_increment, i_resetb_c, 
            o_baseband_q_c_7, o_baseband_i_c_7, o_baseband_i_c_15, o_baseband_i_c_14, 
            o_baseband_i_c_13, o_baseband_i_c_12, o_baseband_i_c_11, o_baseband_i_c_10, 
            n3655, o_baseband_i_c_8, \quarter_wave_sample_register_q[15] , 
            n29501, o_baseband_q_c_15, o_baseband_q_c_14, o_baseband_q_c_13, 
            o_baseband_q_c_12, o_baseband_q_c_11, o_baseband_q_c_10, n3656, 
            o_baseband_q_c_8, GND_net) /* synthesis syn_module_defined=1 */ ;
    input dac_clk_p_c;
    input i_resetb_N_301;
    input [30:0]carrier_increment;
    input i_resetb_c;
    output o_baseband_q_c_7;
    output o_baseband_i_c_7;
    output o_baseband_i_c_15;
    output o_baseband_i_c_14;
    output o_baseband_i_c_13;
    output o_baseband_i_c_12;
    output o_baseband_i_c_11;
    output o_baseband_i_c_10;
    output n3655;
    output o_baseband_i_c_8;
    output \quarter_wave_sample_register_q[15] ;
    input n29501;
    output o_baseband_q_c_15;
    output o_baseband_q_c_14;
    output o_baseband_q_c_13;
    output o_baseband_q_c_12;
    output o_baseband_q_c_11;
    output o_baseband_q_c_10;
    output n3656;
    output o_baseband_q_c_8;
    input GND_net;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(28[49:58])
    wire o_baseband_q_c_7 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[49:59])
    wire o_baseband_i_c_7 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[37:47])
    wire o_baseband_i_c_15 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[37:47])
    wire o_baseband_i_c_14 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[37:47])
    wire o_baseband_i_c_13 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[37:47])
    wire o_baseband_i_c_12 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[37:47])
    wire o_baseband_i_c_11 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[37:47])
    wire o_baseband_i_c_10 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[37:47])
    wire n3655 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[37:47])
    wire o_baseband_i_c_8 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[37:47])
    wire o_baseband_q_c_15 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[49:59])
    wire o_baseband_q_c_14 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[49:59])
    wire o_baseband_q_c_13 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[49:59])
    wire o_baseband_q_c_12 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[49:59])
    wire o_baseband_q_c_11 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[49:59])
    wire o_baseband_q_c_10 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[49:59])
    wire n3656 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[49:59])
    wire o_baseband_q_c_8 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[49:59])
    wire [30:0]increment;   // d:/documents/git_local/fm_modulator/rtl/dds.v(14[31:40])
    wire [11:0]o_phase;   // d:/documents/git_local/fm_modulator/rtl/dds.v(18[26:33])
    
    FD1S3DX increment_i0 (.D(carrier_increment[0]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(increment[0])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=67, LSE_RLINE=67 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i0.GSR = "DISABLED";
    FD1S3DX increment_i30 (.D(carrier_increment[30]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(increment[30])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=67, LSE_RLINE=67 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i30.GSR = "DISABLED";
    FD1S3DX increment_i29 (.D(carrier_increment[29]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(increment[29])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=67, LSE_RLINE=67 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i29.GSR = "DISABLED";
    FD1S3DX increment_i28 (.D(carrier_increment[28]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(increment[28])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=67, LSE_RLINE=67 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i28.GSR = "DISABLED";
    FD1S3DX increment_i27 (.D(carrier_increment[27]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(increment[27])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=67, LSE_RLINE=67 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i27.GSR = "DISABLED";
    FD1S3DX increment_i26 (.D(carrier_increment[26]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(increment[26])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=67, LSE_RLINE=67 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i26.GSR = "DISABLED";
    FD1S3DX increment_i25 (.D(carrier_increment[25]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(increment[25])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=67, LSE_RLINE=67 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i25.GSR = "DISABLED";
    FD1S3DX increment_i24 (.D(carrier_increment[24]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(increment[24])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=67, LSE_RLINE=67 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i24.GSR = "DISABLED";
    FD1S3DX increment_i23 (.D(carrier_increment[23]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(increment[23])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=67, LSE_RLINE=67 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i23.GSR = "DISABLED";
    FD1S3DX increment_i22 (.D(carrier_increment[22]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(increment[22])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=67, LSE_RLINE=67 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i22.GSR = "DISABLED";
    FD1S3DX increment_i21 (.D(carrier_increment[21]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(increment[21])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=67, LSE_RLINE=67 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i21.GSR = "DISABLED";
    FD1S3DX increment_i20 (.D(carrier_increment[20]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(increment[20])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=67, LSE_RLINE=67 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i20.GSR = "DISABLED";
    FD1S3DX increment_i19 (.D(carrier_increment[19]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(increment[19])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=67, LSE_RLINE=67 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i19.GSR = "DISABLED";
    FD1S3DX increment_i18 (.D(carrier_increment[18]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(increment[18])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=67, LSE_RLINE=67 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i18.GSR = "DISABLED";
    FD1S3DX increment_i17 (.D(carrier_increment[17]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(increment[17])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=67, LSE_RLINE=67 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i17.GSR = "DISABLED";
    FD1S3DX increment_i16 (.D(carrier_increment[16]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(increment[16])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=67, LSE_RLINE=67 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i16.GSR = "DISABLED";
    FD1S3DX increment_i15 (.D(carrier_increment[15]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(increment[15])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=67, LSE_RLINE=67 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i15.GSR = "DISABLED";
    FD1S3DX increment_i14 (.D(carrier_increment[14]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(increment[14])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=67, LSE_RLINE=67 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i14.GSR = "DISABLED";
    FD1S3DX increment_i13 (.D(carrier_increment[13]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(increment[13])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=67, LSE_RLINE=67 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i13.GSR = "DISABLED";
    FD1S3DX increment_i12 (.D(carrier_increment[12]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(increment[12])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=67, LSE_RLINE=67 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i12.GSR = "DISABLED";
    FD1S3DX increment_i11 (.D(carrier_increment[11]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(increment[11])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=67, LSE_RLINE=67 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i11.GSR = "DISABLED";
    FD1S3DX increment_i10 (.D(carrier_increment[10]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(increment[10])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=67, LSE_RLINE=67 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i10.GSR = "DISABLED";
    FD1S3DX increment_i9 (.D(carrier_increment[9]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(increment[9])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=67, LSE_RLINE=67 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i9.GSR = "DISABLED";
    FD1S3DX increment_i8 (.D(carrier_increment[8]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(increment[8])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=67, LSE_RLINE=67 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i8.GSR = "DISABLED";
    FD1S3DX increment_i7 (.D(carrier_increment[7]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(increment[7])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=67, LSE_RLINE=67 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i7.GSR = "DISABLED";
    FD1S3DX increment_i6 (.D(carrier_increment[6]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(increment[6])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=67, LSE_RLINE=67 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i6.GSR = "DISABLED";
    FD1S3DX increment_i5 (.D(carrier_increment[5]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(increment[5])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=67, LSE_RLINE=67 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i5.GSR = "DISABLED";
    FD1S3DX increment_i4 (.D(carrier_increment[4]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(increment[4])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=67, LSE_RLINE=67 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i4.GSR = "DISABLED";
    FD1S3DX increment_i3 (.D(carrier_increment[3]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(increment[3])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=67, LSE_RLINE=67 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i3.GSR = "DISABLED";
    FD1S3DX increment_i2 (.D(carrier_increment[2]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(increment[2])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=67, LSE_RLINE=67 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i2.GSR = "DISABLED";
    FD1S3DX increment_i1 (.D(carrier_increment[1]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(increment[1])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=4, LSE_RCOL=158, LSE_LLINE=67, LSE_RLINE=67 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(26[11] 30[5])
    defparam increment_i1.GSR = "DISABLED";
    quarter_wave_sine_lookup_U0 qtr_inst (.dac_clk_p_c(dac_clk_p_c), .i_resetb_c(i_resetb_c), 
            .o_phase({o_phase}), .i_resetb_N_301(i_resetb_N_301), .o_baseband_q_c_7(o_baseband_q_c_7), 
            .o_baseband_i_c_7(o_baseband_i_c_7), .o_baseband_i_c_15(o_baseband_i_c_15), 
            .o_baseband_i_c_14(o_baseband_i_c_14), .o_baseband_i_c_13(o_baseband_i_c_13), 
            .o_baseband_i_c_12(o_baseband_i_c_12), .o_baseband_i_c_11(o_baseband_i_c_11), 
            .o_baseband_i_c_10(o_baseband_i_c_10), .n3655(n3655), .o_baseband_i_c_8(o_baseband_i_c_8), 
            .\quarter_wave_sample_register_q[15] (\quarter_wave_sample_register_q[15] ), 
            .n29501(n29501), .o_baseband_q_c_15(o_baseband_q_c_15), .o_baseband_q_c_14(o_baseband_q_c_14), 
            .o_baseband_q_c_13(o_baseband_q_c_13), .o_baseband_q_c_12(o_baseband_q_c_12), 
            .o_baseband_q_c_11(o_baseband_q_c_11), .o_baseband_q_c_10(o_baseband_q_c_10), 
            .n3656(n3656), .o_baseband_q_c_8(o_baseband_q_c_8), .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(21[70:134])
    \nco(OW=12)_U1  nco_inst (.increment({increment}), .o_phase({o_phase}), 
            .GND_net(GND_net), .dac_clk_p_c(dac_clk_p_c), .i_resetb_N_301(i_resetb_N_301)) /* synthesis syn_module_defined=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/dds.v(20[49:100])
    
endmodule
//
// Verilog Description of module quarter_wave_sine_lookup_U0
//

module quarter_wave_sine_lookup_U0 (dac_clk_p_c, i_resetb_c, o_phase, 
            i_resetb_N_301, o_baseband_q_c_7, o_baseband_i_c_7, o_baseband_i_c_15, 
            o_baseband_i_c_14, o_baseband_i_c_13, o_baseband_i_c_12, o_baseband_i_c_11, 
            o_baseband_i_c_10, n3655, o_baseband_i_c_8, \quarter_wave_sample_register_q[15] , 
            n29501, o_baseband_q_c_15, o_baseband_q_c_14, o_baseband_q_c_13, 
            o_baseband_q_c_12, o_baseband_q_c_11, o_baseband_q_c_10, n3656, 
            o_baseband_q_c_8, GND_net) /* synthesis syn_module_defined=1 */ ;
    input dac_clk_p_c;
    input i_resetb_c;
    input [11:0]o_phase;
    input i_resetb_N_301;
    output o_baseband_q_c_7;
    output o_baseband_i_c_7;
    output o_baseband_i_c_15;
    output o_baseband_i_c_14;
    output o_baseband_i_c_13;
    output o_baseband_i_c_12;
    output o_baseband_i_c_11;
    output o_baseband_i_c_10;
    output n3655;
    output o_baseband_i_c_8;
    output \quarter_wave_sample_register_q[15] ;
    input n29501;
    output o_baseband_q_c_15;
    output o_baseband_q_c_14;
    output o_baseband_q_c_13;
    output o_baseband_q_c_12;
    output o_baseband_q_c_11;
    output o_baseband_q_c_10;
    output n3656;
    output o_baseband_q_c_8;
    input GND_net;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(28[49:58])
    wire o_baseband_q_c_7 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[49:59])
    wire [15:0]\o_val_pipeline_q[0]  /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(16[24:40])
    wire o_baseband_i_c_7 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[37:47])
    wire [15:0]\o_val_pipeline_i[0]  /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(15[24:40])
    wire o_baseband_i_c_15 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[37:47])
    wire o_baseband_i_c_14 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[37:47])
    wire o_baseband_i_c_13 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[37:47])
    wire o_baseband_i_c_12 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[37:47])
    wire o_baseband_i_c_11 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[37:47])
    wire o_baseband_i_c_10 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[37:47])
    wire n3655 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[37:47])
    wire o_baseband_i_c_8 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[37:47])
    wire o_baseband_q_c_15 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[49:59])
    wire o_baseband_q_c_14 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[49:59])
    wire o_baseband_q_c_13 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[49:59])
    wire o_baseband_q_c_12 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[49:59])
    wire o_baseband_q_c_11 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[49:59])
    wire o_baseband_q_c_10 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[49:59])
    wire n3656 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[49:59])
    wire o_baseband_q_c_8 /* synthesis syn_pipeline=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(111[49:59])
    
    wire n26893;
    wire [9:0]index_q;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(31[26:33])
    
    wire n14814, n252, n24733, n20555;
    wire [9:0]index_i;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(31[17:24])
    
    wire n26836, n254, n620, n635, n636, n23217, n23218, n23219, 
        n25444, n25443, n25445, n22780, n22781, n22785, n620_adj_2250, 
        n22842, n22843, n22847, n23279, n23280, n23281, n22866, 
        n22867, n22870, n22868, n22869, n22871, n23298, n23299, 
        n23306, n23300, n23301, n23307, n557, n572, n23405, n589, 
        n604, n23406, n22138, n22139, n22140, n620_adj_2251, n635_adj_2252, 
        n23407, n23002, n23003, n23006, n25412, n25409, n25413, 
        n653, n668, n23408, n684, n699, n23409, n23081, n21729, 
        n22860, n27143, n27144, n27145, n27106, n652, n653_adj_2253, 
        n716, n731, n23410, n23432, n23433, n23434, n660, n27105, 
        n668_adj_2254, n190, n253, n22859, n747, n762, n23411;
    wire [11:0]phase_q;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(12[17:24])
    wire [15:0]quarter_wave_sample_register_i;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(22[24:54])
    wire [14:0]quarter_wave_sample_register_i_15__N_2126;
    
    wire n541, n23104, n23105, n23109, n26733, n20559, n26861, 
        n254_adj_2255, n812, n781, n796, n23412, n26863, n11958, 
        n26887, n29485, n684_adj_2256, n812_adj_2257, n11914, n23413, 
        n557_adj_2258, n22064;
    wire [1:0]phase_negation_i;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(23[12:28])
    wire [11:0]phase_i;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(11[17:24])
    wire [1:0]phase_negation_q;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(23[30:46])
    wire [9:0]index_i_9__N_2106;
    wire [9:0]index_q_9__N_2116;
    wire [15:0]quarter_wave_sample_register_q;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(22[56:86])
    wire [14:0]quarter_wave_sample_register_q_15__N_2141;
    
    wire n22021, n30, n364, n22918, n844, n11917, n23414, o_val_pipeline_i_0__15__N_2156, 
        n875, n890, n23415, n26909, o_val_pipeline_i_0__15__N_2158, 
        o_val_pipeline_i_0__15__N_2160, o_val_pipeline_i_0__15__N_2162, 
        n26977, o_val_pipeline_i_0__15__N_2164, n23004, n23005, n23007, 
        n908, n923, n23416, o_val_pipeline_i_0__15__N_2166, n23494, 
        n23495, n23496, o_val_pipeline_i_0__15__N_2168, o_val_pipeline_i_0__15__N_2170, 
        o_val_pipeline_i_0__15__N_2172, n939, n954, n23417, n26748, 
        n844_adj_2259, n860, n22650, n22651, n22655, n22670, n22671, 
        n22676, n22672, n22673, n22677, n971, n986, n23418, n25583, 
        n27236, n27237, n62, n1002, n1017, n23419, n22697, n22698, 
        n22705, n22699, n22700, n22706, n22716, n22717, n22722, 
        n22718, n22719, n22723, n25493, n781_adj_2260, n22048, n22770, 
        n22771, n26856, n62_adj_2261, n22774, n22775, n22782, n22776, 
        n22777, n22783, n23315, n23316, n23322, n844_adj_2262, n12112, 
        n23476;
    wire [14:0]n1829;
    
    wire n26416, n22807, n22808, n22814, n851, n27058, n23078, 
        n22809, n22810, n22815, n22811, n22812, n22816, n22012, 
        n22830, n22831, n22841, n29495, n985, n875_adj_2263, n890_adj_2264, 
        n891, n22832, n22833, n22838, n22839, n22845, n382, n509, 
        n22852, n23009, n23010, n23013, n844_adj_2265, n859, n860_adj_2266, 
        n22862, n22863, n22864, n22865, n716_adj_2267, n23011, n23012, 
        n23014, n23302, n23303, n23308, n23317, n23318, n23323, 
        n17597;
    wire [15:0]o_val_pipeline_i_0__15__N_2157;
    
    wire n23319, n23320, n23324, n17596, n17595, n22142;
    wire [11:0]phase_q_11__N_2232;
    
    wire n27102, n23077, n27230, n27231, n27232, n23332, n23333, 
        n23334, n22989, n22990, n22996, n22991, n22992, n22997, 
        n27080, n27099, n21416, n22993, n22994, n22998, n21754, 
        n21755, n21756, n23016, n23017, n23020, n22488, n22489, 
        n22494, n23018, n23019, n23021, n23092, n23093, n23103, 
        n27095, n356, n21415, n21757, n21758, n21759, n23094, 
        n23095, n17594, n23100, n23101, n23107, n27085, n21773, 
        n23313, n25001, n23321, n653_adj_2268, n22567, n22568, n22575, 
        n23326, n26854, n21763, n21764, n21765, n22569, n22570, 
        n22576, n21417, n17593, n21769, n21770, n21771, n12164, 
        n397, n747_adj_2269, n762_adj_2270, n763, n21772, n21774, 
        n23304, n23305, n23309, n93, n21565, n21566, n21567, n23288, 
        n24971, n21775, n21776, n21777, n13947, n26978, n27135, 
        n27136, n27137, n23179, n23180, n23181, n475, n21574, 
        n21575, n21576, n22640, n22641, n22644, n22645, n22652, 
        n22646, n22647, n22653, n382_adj_2271, n509_adj_2272, n22660, 
        n21684, n21687, n22669, n21690, n21693, n21696, n21699, 
        n526, n24904, n17592, n17591, n21702, n892, n24964, n23287, 
        n27218, n27219, n27220, n157, n29477, n27104, n23076, 
        n27086, n23075, n25322, n23283, n22681, n22682, n22861, 
        n27215, n27216, n27217, n21427, n22683, n22684, n22858, 
        n27212, n27213, n27214, n22685, n22686, n22687, n22688, 
        n22689, n22690, n22701, n22693, n22694, n22703, n27209, 
        n27210, n27211, n12116, n21711, n22713, n27061, n23071, 
        n21717, n21720, n22715, n574, n21723, n21726, n764, n23205, 
        n23206, n23213, n23211, n23212, n23216, n22727, n22728, 
        n22743, n22729, n22730, n22744, n22731, n22732, n22745, 
        n21466, n316, n25734, n22735, n22736, n22747, n26796, 
        n189, n25731, n26872, n26772, n637, n12109, n27206, n27207, 
        n27208, n25652, n22737, n22738, n22748, n812_adj_2273, n17814, 
        n29494, n27107, n22739, n22740, n22749, n22741, n22742, 
        n22750, n26871, n93_adj_2274, n21725, n142, n22916, n716_adj_2275, 
        n797, n828, n10079, n765, n317, n22758, n22759, n26859, 
        n700, n24805, n428, n890_adj_2276, n891_adj_2277, n443, 
        n22760, n22761, n506, n26875, n24734, n22762, n22763, 
        n26849, n860_adj_2278, n46, n364_adj_2279, n22897, n716_adj_2280, 
        n25968, n62_adj_2281, n27034, n221, n26721, n955, n908_adj_2282, 
        n285, n25490, n12079, n731_adj_2283, n732, n444, n22764, 
        n22765, n251, n15108, n252_adj_2284, n812_adj_2285, n25492, 
        n25494, n22766, n22767, n22778, n22772, n22773, n26842, 
        n189_adj_2286, n26876, n316_adj_2287, n22895, n317_adj_2288, 
        n9918, n765_adj_2289, n93_adj_2290, n24783, n890_adj_2291, 
        n891_adj_2292, n21677, n26835, n700_adj_2293, n22791, n22792, 
        n22806, n22793, n22794, n26877, n26775, n637_adj_2294, n22085, 
        n221_adj_2295, n173, n27117, n22795, n22796, n22797, n22798, 
        n25707, n22799, n22800, n27088, n939_adj_2296, n24710, n747_adj_2297, 
        n25667, n27077, n21458, n22714, n22721, n762_adj_2298, n25670, 
        n732_adj_2299, n763_adj_2300, n220, n23257, n22067, n21457, 
        n21459, n27096, n29474, n21455, n22104, n891_adj_2301, n443_adj_2302, 
        n428_adj_2303, n22820, n22821, n22836, n46_adj_2304, n23252, 
        n762_adj_2305, n27129, n27130, n27131, n22824, n22825, n21391, 
        n21392, n21393, n22826, n22827, n22151, n22834, n22835, 
        n23267, n23268, n23275, n23273, n23274, n23278, n23067, 
        n23074, n21394, n21395, n21396, n22966, n22965, n25321, 
        n25318, n22013, n251_adj_2306, n25320, n25319, n21732, n21735, 
        n21738, n21741, n252_adj_2307, n443_adj_2308, n333, n379, 
        n21744, n21747, n23070, n443_adj_2309, n379_adj_2310, n890_adj_2311, 
        n21750, n892_adj_2312, n699_adj_2313, n23055, n460, n23057, 
        n26747, n251_adj_2314, n109, n21440, n23056, n15, n412, 
        n25672, n22970, n26882, n26821, n22903, n763_adj_2315, n24486, 
        n252_adj_2316, n604_adj_2317, n22967, n684_adj_2318, n157_adj_2319, 
        n413, n24494, n24487, n24495, n412_adj_2320, n22901, n381, 
        n23290, n23291, n460_adj_2321, n23292, n23293, n23294, n23295, 
        n619, n26927, n25578, n23277, n109_adj_2322, n24642, n24640, 
        n24643, n23296, n23297, n27001, n29491, n364_adj_2323, n21451, 
        n21452, n21453, n541_adj_2324, n21400, n21401, n21402, n29493, 
        n526_adj_2325, n29497, n668_adj_2326, n26999, n379_adj_2327, 
        n21669, n21672, n574_adj_2328, n21675, n22668, n22675, n22666, 
        n22667, n22674, n38, n21995, n252_adj_2329, n716_adj_2330, 
        n684_adj_2331, n445, n26983, n27028, n25580, n716_adj_2332, 
        n21935, n21678, n764_adj_2333, n445_adj_2334, n412_adj_2335, 
        n27024, n25584, n22102, n699_adj_2336, n773, n25586, n890_adj_2337, 
        n684_adj_2338, n27200, n27201, n27202, n27022, n25602, n22898, 
        n22899, n23276, n22905, n22906, n22372, n26720, n955_adj_2339, 
        n22659, n22663, n924, n24641, n23328, n23329, n26986, 
        n25611, n22854, n22856, n27048, n526_adj_2340, n542, n635_adj_2341, 
        n21674, n26864, n24731, n28252, n27063, n635_adj_2342, n21722, 
        n526_adj_2343, n542_adj_2344, n700_adj_2345, n26714, n26996, 
        n27027, n22100, n541_adj_2346, n29489, n27025, n526_adj_2347, 
        n731_adj_2348, n25634, n23069, n22073, n27031, n22070, n109_adj_2349, 
        n23330, n23331, n254_adj_2350, n511, n15088, n1022, n24748, 
        n29500, n22919, n22920, n348, n29487, n22055, n20693, 
        n24639, n26860, n21958, n29488, n762_adj_2351, n22027, n173_adj_2352, 
        n189_adj_2353, n508, n26987, n668_adj_2354, n25316, n747_adj_2355, 
        n763_adj_2356, n124, n21707, n29473, n27072, n21446, n27098, 
        n21445, n21447, n22926, n22927, n15064, n1022_adj_2357, 
        n21443, n26732, n21439, n21442, n21444, n908_adj_2358, n14171, 
        n21692, n23062, n491, n506_adj_2359, n21686, n25317, n26911, 
        n812_adj_2360, n29490, n604_adj_2361, n27123, n27124, n27125, 
        n364_adj_2362, n124_adj_2363, n21659, n21434, n26913, n475_adj_2364, 
        n21433, n21435, n27081, n491_adj_2365, n27035, n189_adj_2366, 
        n22022, n24753, n21538, n1001, n21422, n19801, n25270, 
        n26974, n25271, n29492, n27071, n747_adj_2367, n29470, n796_adj_2368, 
        n27044, n27079, n444_adj_2369, n26918, n25268, n25269, n24736, 
        n21532, n397_adj_2370, n251_adj_2371, n25669, n27116, n19798, 
        n27197, n27198, n27199, n22573, n24712, n22578, n22571, 
        n22572, n22577, n796_adj_2372, n797_adj_2373, n22580, n22678, 
        n22679, n22150, n23310, n23311, n491_adj_2374, n27078, n23068, 
        n22973, n22974, n22988, n22975, n22976, n668_adj_2375, n931, 
        n188, n890_adj_2376, n475_adj_2377, n24619, n26700, n26417, 
        n124_adj_2378, n23254, n22977, n22978, n29471, n22979, n22980, 
        n12161, n22981, n22982, n27101, n25802, n27066, n25804, 
        n26982, n27032, n21965, n23420, n23421, n23428, n460_adj_2379, 
        n26993, n22061, n25813, n23422, n23423, n23429, n285_adj_2380, 
        n23424, n23425, n23430, n29472, n588, n25815, n22090, 
        n26995, n605, n27120, n23426, n23427, n23431, n22025, 
        n26923, n475_adj_2381, n491_adj_2382, n684_adj_2383, n29468, 
        n21950, n21691, n475_adj_2384, n70, n653_adj_2385, n21657, 
        n21660, n21689, n26356, n22497, n22495, n22476, n22477, 
        n22478, n22479, n22480, n22481, n22490, n22482, n22483, 
        n22491, n23000, n22995, n22999, n27046, n573, n285_adj_2386, 
        n22894, n573_adj_2387, n27119;
    wire [15:0]o_val_pipeline_q_0__15__N_2189;
    
    wire n22168, n124_adj_2388, n24782, n23325, n444_adj_2389, n732_adj_2390, 
        n763_adj_2391, n397_adj_2392, n573_adj_2393, n125, n22851, 
        n22855, n25237, n25234, n25238, n476, n24864, n24865, 
        n12149, n23054, n23058, n891_adj_2394, n142_adj_2395, n157_adj_2396, 
        n158, n22818, n23082, n23083, n23098, n22813, n22817, 
        n23086, n23087, n25236, n23059, n22720, n22724, n22708, 
        n93_adj_2397, n22702, n22707, n22710, n22654, n22657, n23088, 
        n23089, n29475, n22166, n22656, n27090, n573_adj_2398, n285_adj_2399, 
        n22915, n23096, n23097, n23061, n23065, n22156, n125_adj_2400, 
        n574_adj_2401, n21577, n124_adj_2402, n24804, n22579, n574_adj_2403, 
        n21568, n22152, n23108, n23111, n557_adj_2404, n573_adj_2405, 
        n23063, n23064, n23066, n23106, n23110, n573_adj_2406, n26994, 
        n15132, n22712, n26937, n173_adj_2407, n404, n21956, n27160, 
        n17577, n22846, n22849, n301, n908_adj_2408, n317_adj_2409, 
        n22551, n22552, n22844, n22848, n22553, n22554, n22555, 
        n22556, n22784, n22787, n17576, n22557, n22558, n397_adj_2410, 
        n22559, n22560, n22563, n22564, n22786, n22709, n27000, 
        n716_adj_2411, n23072, n28248, n28249, n142_adj_2412, n12157, 
        n12158, n22374, n12050, n28251, n23073, n15_adj_2413, n26898, 
        n763_adj_2414, n22169, n15106, n27103, n23079, n28269, n28270, 
        n318, n381_adj_2415, n23080, n716_adj_2416, n25733, n526_adj_2417, 
        n25233, n21914, n21982, n318_adj_2418, n21448, n635_adj_2419, 
        n21449, n25212, n25210, n25213, n21460, n27122, n21462, 
        n908_adj_2420, n924_adj_2421, n25211, n285_adj_2422, n27159, 
        n21705, n21708, n21910, n21911, n21912, n21421, n476_adj_2423, 
        n22597, n22598, n22613, n22599, n22600, n22614, n541_adj_2424, 
        n890_adj_2425, n891_adj_2426, n22601, n22602, n22615, n17808, 
        n17809, n17810, n444_adj_2427, n24868, n22605, n22606, n22617, 
        n22607, n22608, n22618, n22609, n22610, n22619, n22611, 
        n22612, n22620, n668_adj_2428, n669, n23482, n23483, n23490, 
        n11973, n23484, n23485, n23491, n23486, n23487, n23492, 
        n21925, n21926, n21927, n23488, n23489, n23493, n828_adj_2429, 
        n21450, n22628, n22629, n460_adj_2430, n476_adj_2431, n23175, 
        n23176, n397_adj_2432, n27056, n413_adj_2433, n21931, n21932, 
        n21933, n23177, n23178, n27083, n25965, n21934, n21936, 
        n93_adj_2434, n13941, n286, n22630, n22631, n22632, n22633, 
        n21940, n21941, n21942, n27189, n27190, n27191, n22634, 
        n22635, n22636, n22637, n22648, n572_adj_2435, n142_adj_2436, 
        n157_adj_2437, n158_adj_2438, n491_adj_2439, n125_adj_2440, 
        n22642, n22643, n26713, n21971, n23008, n23015, n956, 
        n20334, n24902, n24903, n27065, n21413, n892_adj_2441, n21412, 
        n21414, n28534, n252_adj_2442, n28532, n21441, n1002_adj_2443, 
        n94, n125_adj_2444, n28535, n25209, n25208, n506_adj_2445, 
        n25447, n860_adj_2446, n17830, n14440, n21430, n21431, n21432, 
        n28556, n21957, n21960, n21963, n21966, n413_adj_2447, n444_adj_2448, 
        n26737, n26773, n638, n28554, n476_adj_2449, n507, n27084, 
        n26014, n17811, n17812, n17813, n17816, n573_adj_2450, n28557, 
        n892_adj_2451, n605_adj_2452, n636_adj_2453, n21969, n700_adj_2454, 
        n22691, n27091, n61, n62_adj_2455, n15_adj_2456, n26834, 
        n31, n27094, n828_adj_2457, n21972, n22692, n797_adj_2458, 
        n828_adj_2459, n21943, n21944, n21945, n26512, n23189, n23190, 
        n14871, n860_adj_2460, n891_adj_2461, n23191, n23192, n21428, 
        n21429, n23193, n23194, n23207, n684_adj_2462, n700_adj_2463, 
        n653_adj_2464, n669_adj_2465, n22148, n542_adj_2466, n26816, 
        n27161, n30_adj_2467, n31_adj_2468, n24907, n12015, n270, 
        n286_adj_2469, n700_adj_2470, n19881, n1018, n15_adj_2471, 
        n30_adj_2472, n31_adj_2473, n348_adj_2474, n27047, n61_adj_2475, 
        n62_adj_2476, n491_adj_2477, n15_adj_2478, n26792, n31_adj_2479, 
        n27057, n94_adj_2480, n30_adj_2481, n31_adj_2482, n23199, 
        n23200, n23210, n21955, n23201, n23202, n12103, n12104, 
        n23203, n23204, n26813, n26776, n26781, n23337, n94_adj_2483, 
        n21975, n1002_adj_2484, n221_adj_2485, n252_adj_2486, n93_adj_2487, 
        n12134, n22116, n286_adj_2488, n21978, n221_adj_2489, n21959, 
        n21961, n21962, n349, n21981, n890_adj_2490, n475_adj_2491, 
        n26973, n700_adj_2492, n22401, n28805, n28806, n26991, n24962, 
        n22113, n173_adj_2493, n875_adj_2494, n891_adj_2495, n15_adj_2496, 
        n859_adj_2497, n860_adj_2498, n21397, n21398, n21399, n157_adj_2499, 
        n26892, n636_adj_2500, n731_adj_2501, n796_adj_2502, n26928, 
        n24617, n669_adj_2503, n700_adj_2504, n17786, n17787, n17788, 
        n21964, n22002, n22005, n828_adj_2505, n26900, n27026, n124_adj_2506, 
        n491_adj_2507, n507_adj_2508, n460_adj_2509, n476_adj_2510, 
        n860_adj_2511, n22008, n397_adj_2512, n413_adj_2513, n21970, 
        n27023, n24959, n17822, n17823, n17824, n109_adj_2514, n124_adj_2515, 
        n125_adj_2516, n797_adj_2517, n94_adj_2518, n26934, n24965, 
        n24966, n30_adj_2519, n31_adj_2520, n26989, n24969, n557_adj_2521, 
        n572_adj_2522, n23467, n286_adj_2523, n29040, n29041, n29039, 
        n26767, n23184, n29038, n29042, n589_adj_2524, n23468, n29043, 
        n29044, n29045, n94_adj_2525, n125_adj_2526, n17575, n316_adj_2527, 
        n923_adj_2528, n924_adj_2529, n158_adj_2530, n27186, n27187, 
        n27188, n24973, n157_adj_2531, n24974, n21766, n21767, n21768, 
        n27064, n125_adj_2532, n26706, n15124, n26707, n29159, n22133, 
        n29158, n27003, n24994, n29160, n29161, n29162, n29163, 
        n29164, n29165, n286_adj_2533, n22017, n24998, n22103, n25000, 
        n349_adj_2534, n22020, n620_adj_2535, n635_adj_2536, n23469, 
        n24488, n26709, n349_adj_2537, n308, n22040, n413_adj_2538, 
        n22147, n22149, n189_adj_2539, n476_adj_2540, n507_adj_2541, 
        n22023, n508_adj_2542, n21985, n21986, n21987, n12091, n22026, 
        n892_adj_2543, n669_adj_2544, n700_adj_2545, n22768, n22029, 
        n22769, n860_adj_2546, n891_adj_2547, n27068, n620_adj_2548, 
        n635_adj_2549, n636_adj_2550, n924_adj_2551, n22032, n93_adj_2552, 
        n94_adj_2553, n348_adj_2554, n27082, n12016, n22035, n653_adj_2555, 
        n668_adj_2556, n23470, n716_adj_2557, n732_adj_2558, n22399, 
        n21917, n699_adj_2559, n23471, n21737, n684_adj_2560, n26215, 
        n732_adj_2561, n158_adj_2562, n26564, n26561, n21922, n21923, 
        n21924, n21988, n21989, n21990, n26216, n26221, n221_adj_2563, 
        n22041, n475_adj_2564, n26223, n286_adj_2565, n317_adj_2566, 
        n716_adj_2567, n23472, n78, n891_adj_2568, n26563, n26562, 
        n653_adj_2569, n349_adj_2570, n22044, n21739, n413_adj_2571, 
        n22047, n26224, n26229, n22050, n507_adj_2572, n13909, n828_adj_2573, 
        n26719, n797_adj_2574, n22053, n605_adj_2575, n22056, n669_adj_2576, 
        n669_adj_2577, n732_adj_2578, n763_adj_2579, n24624, n24625, 
        n747_adj_2580, n23473, n24623, n24622, n22802, n26560, n22624, 
        n21994, n17574, n812_adj_2581, n542_adj_2582, n12119, n11119, 
        n252_adj_2583, n25900, n22471, n20197, n94_adj_2584, n22062, 
        n22065, n22068, n22822, n22071, n317_adj_2585, n286_adj_2586, 
        n26716, n701, n26246, n349_adj_2587, n22074, n22077, n22080, 
        n22083, n22086, n28559, n26250, n17573, n22092, n22829, 
        n26717, n701_adj_2588, n26261, n22095, n28537, n26265, n27092, 
        n22098, n22101, n924_adj_2589, n22107, n498, n62_adj_2590, 
        n747_adj_2591, n908_adj_2592, n21746, n14928, n21745, n173_adj_2593, 
        n26766, n26770, n93_adj_2594, n21743, n987, n22110, n21742, 
        n526_adj_2595, n21736, n22014, n397_adj_2596, n21733, n781_adj_2597, 
        n23474, n348_adj_2598, n443_adj_2599, n21731, n781_adj_2600, 
        n21730, n24869, n26296, n21728, n23475, n333_adj_2601, n21727, 
        n26294, n23251, n17572, n27174, n26297, n27182, n27183, 
        n27184, n23253, n27002, n931_adj_2602, n188_adj_2603, n26513, 
        n26514, n731_adj_2604, n732_adj_2605, n26967, n13925, n653_adj_2606, 
        n669_adj_2607, n954_adj_2608, n23255, n23256, n23269, n604_adj_2609, 
        n605_adj_2610, n27141, n21479, n21480, n23258, n23270, n27193, 
        n22134, n21475, n21476, n21477, n22028, n397_adj_2611, n413_adj_2612, 
        n25736, n23060, n23261, n23262, n23272, n27192, n124_adj_2613, 
        n316_adj_2614, n317_adj_2615, n270_adj_2616, n286_adj_2617, 
        n23263, n23264, n26011, n158_adj_2618, n23265, n23266, n27176, 
        n986_adj_2619, n684_adj_2620, n700_adj_2621, n26768, n26769, 
        n22115, n875_adj_2622, n890_adj_2623, n891_adj_2624, n27062, 
        n22114, n22112, n22111, n844_adj_2625, n859_adj_2626, n860_adj_2627, 
        n21976, n28254, n23214, n25495, n23215, n27029, n22108, 
        n956_adj_2628, n20333, n22109, n491_adj_2629, n21719, n21655, 
        n21656, n475_adj_2630, n21718, n22474, n26351, n22105, n22106, 
        n21658, n21716, n21715, n12055, n22097, n542_adj_2631, n573_adj_2632, 
        n636_adj_2633, n22473, n26352, n669_adj_2634, n700_adj_2635, 
        n26753, n21949, n22082, n491_adj_2636, n22024, n22075, n732_adj_2637, 
        n21951, n25449, n22469, n26354, n797_adj_2638, n828_adj_2639, 
        n22072, n891_adj_2640, n731_adj_2641, n25096, n25097, n26933, 
        n653_adj_2642, n21706, n204, n397_adj_2643, n26759, n985_adj_2644, 
        n986_adj_2645, n971_adj_2646, n859_adj_2647, n27087, n21703, 
        n301_adj_2648, n506_adj_2649, n26848, n939_adj_2650, n923_adj_2651, 
        n21698, n14858, n21697, n93_adj_2652, n21695, n21694, n443_adj_2653, 
        n30_adj_2654, n142_adj_2655, n158_adj_2656, n26932, n27178, 
        n27179, n27180, n859_adj_2657, n21667, n21668, n17571, n875_adj_2658, 
        n21670, n21671, n723, n22063, n27185, n526_adj_2659, n541_adj_2660, 
        n21688, n21916, n26817, n27175, n397_adj_2661, n21685, n860_adj_2662, 
        n892_adj_2663, n491_adj_2664, n25408, n859_adj_2665, n860_adj_2666, 
        n844_adj_2667, n860_adj_2668, n21673, n22054, n348_adj_2669, 
        n21683, n21676, n21682, n19855, n1018_adj_2670, n21680, 
        n333_adj_2671, n21679, n700_adj_2672, n747_adj_2673, n22896, 
        n27177, n25098, n25101, n21704, n270_adj_2674, n348_adj_2675, 
        n22049, n22902, n26774, n491_adj_2676, n25102, n875_adj_2677, 
        n23477, n22045, n22046, n108, n684_adj_2678, n22043, n27181, 
        n22042, n22904, n22039, n301_adj_2679, n763_adj_2680, n812_adj_2681, 
        n14178, n26809, n26874, n766, n21533, n26870, n766_adj_2682, 
        n21539, n21681, n668_adj_2683, n541_adj_2684, n396, n22031, 
        n14875, n22030, n348_adj_2685, n15_adj_2686, n251_adj_2687, 
        n11274, n252_adj_2688, n25653, n23285, n26988, n908_adj_2689, 
        n236, n24708, n22019, n22018, n22066, n21595, n24618, 
        n21472, n22917, n22016, n22015, n22922, n22923, n270_adj_2690, 
        n316_adj_2691, n189_adj_2692, n397_adj_2693, n22924, n22925, 
        n908_adj_2694, n23478, n22159, n22754, n954_adj_2695, n23479, 
        n30_adj_2696, n24807, n22007, n20689, n22093, n22094, n21724, 
        n22006, n23480, n26355, n26353, n1017_adj_2697, n23481, 
        n22003, n22001, n348_adj_2698, n986_adj_2699, n22069, n12120, 
        n24492, n732_adj_2700, n27093, n22485, n24626, n22662, n22664, 
        n763_adj_2701, n22076, n731_adj_2702, n22078, n22079, n22081, 
        n22084, n653_adj_2703, n475_adj_2704, n142_adj_2705, n22052, 
        n954_adj_2706, n653_adj_2707, n27033, n27100, n14203, n684_adj_2708, 
        n12046, n22091, n22033, n26738, n890_adj_2709, n22096, n22099, 
        n26777, n638_adj_2710, n397_adj_2711, n26976, n21983, n21721, 
        n21984, n21980, n21979, n22968, n22969, n21977, n882, 
        n890_adj_2712, n26925, n30_adj_2713, n24785, n46_adj_2714, 
        n12047, n21973, n21974, n1002_adj_2715, n22004, n460_adj_2716, 
        n254_adj_2717, n22000, n542_adj_2718, n221_adj_2719, n21468, 
        n349_adj_2720, n21471, n900, n21474, n142_adj_2721, n157_adj_2722, 
        n507_adj_2723, n1021, n26979, n21483, n26298, n26295, n21953, 
        n763_adj_2724, n21952, n21954, n26840, n1021_adj_2725, n25446, 
        n732_adj_2726, n26990, n22984, n21967, n21968, n26794, n17815, 
        n491_adj_2727, n475_adj_2728, n17828, n17829, n109_adj_2729, 
        n635_adj_2730, n700_adj_2731, n204_adj_2732, n20362, n27045, 
        n19870, n23404, n20198, n21734, n21740, n511_adj_2733, n23022, 
        n173_adj_2734, n26263, n22177, n173_adj_2735, n26262, n26248, 
        n21918, n27097, n26247, n14441, n11929, n573_adj_2736, n605_adj_2737, 
        n636_adj_2738, n27076, n27070, n62_adj_2739, n94_adj_2740, 
        n348_adj_2741, n205, n882_adj_2742, n253_adj_2743, n190_adj_2744, 
        n21409, n21410, n21411, n348_adj_2745, n828_adj_2746, n924_adj_2747, 
        n12165, n507_adj_2748, n22779, n62_adj_2749, n22837, n25607, 
        n22840, n25613, n23099, n23084, n25970, n23102, n26016, 
        n23091, n22649, n22638, n22639, n24908, n11334, n24809, 
        n22143, n22413, n21701, n12048, n26922, n22985, n25817, 
        n22561, n22562, n21467, n24999, n26992, n506_adj_2750, n25635, 
        n24787, n22158, n22161, n22167, n22170, n22179, n22803, 
        n24975, n27021, n24972, n24970, n24967, n21780, n987_adj_2751, 
        n21783, n157_adj_2752, n24963, n24961, n14460, n62_adj_2753, 
        n890_adj_2754, n24491, n573_adj_2755, n24960, n25491, n605_adj_2756, 
        n700_adj_2757, n924_adj_2758, n25577, n25605, n26731, n333_adj_2759, 
        n221_adj_2760, n572_adj_2761, n22725, n12160, n62_adj_2762, 
        n413_adj_2763, n491_adj_2764, n221_adj_2765, n252_adj_2766, 
        n25610, n22420, n349_adj_2767, n924_adj_2768, n924_adj_2769, 
        n23466, n22406, n26015, n26012, n28558, n28555, n26013, 
        n25706, n26746, n28536, n28533, n684_adj_2770, n25801, n25830, 
        n21749, n25969, n25967, n26851, n11977, n25966, n20366, 
        n19907, n349_adj_2771, n444_adj_2772, n21456, n25588, n364_adj_2773, 
        n924_adj_2774, n93_adj_2775, n12095, n28253, n28250, n348_adj_2776, 
        n21481, n21482, n22141, n491_adj_2777, n22157, n22160, n22165, 
        n25899, n21473, n22178, n12148, n25708, n25828, n348_adj_2778, 
        n572_adj_2779, n14464, n205_adj_2780, n21604, n21781, n25608, 
        n21782, n21778, n25829, n21779, n24808, n24806, n25816, 
        n25814, n25812, n25805, n25803, n25806, n27075, n142_adj_2781, 
        n27118, n24786, n24784, n364_adj_2782, n620_adj_2783, n14525, 
        n21470, n11354, n25735, n25732, n21469, n12121, n24751, 
        n27073, n25582, n25632, n24752, n25671, n25668, n572_adj_2784, 
        n25603, n26975, n21454, n25636, n25633, n25637, n24735, 
        n22964, n25612, n25609, n26749, n25606, n25604, n25587, 
        n25585, n25581, n25579, n24493, n24711, n24709, n25448;
    
    LUT4 mux_197_Mux_3_i252_3_lut_4_lut (.A(n26893), .B(index_q[3]), .C(index_q[4]), 
         .D(n14814), .Z(n252)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_3_i252_3_lut_4_lut.init = 16'h08f8;
    LUT4 mux_196_Mux_12_i254_4_lut (.A(n24733), .B(n20555), .C(index_i[6]), 
         .D(n26836), .Z(n254)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_12_i254_4_lut.init = 16'hca0a;
    PFUMX mux_196_Mux_1_i636 (.BLUT(n620), .ALUT(n635), .C0(index_i[4]), 
          .Z(n636)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    PFUMX i20763 (.BLUT(n23217), .ALUT(n23218), .C0(index_i[8]), .Z(n23219));
    PFUMX i23672 (.BLUT(n25444), .ALUT(n25443), .C0(index_q[4]), .Z(n25445));
    L6MUX21 i20329 (.D0(n22780), .D1(n22781), .SD(index_i[7]), .Z(n22785));
    LUT4 mux_196_Mux_7_i620_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n620_adj_2250)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B ((D)+!C)+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_7_i620_3_lut_4_lut_4_lut.init = 16'h83c3;
    L6MUX21 i20391 (.D0(n22842), .D1(n22843), .SD(index_i[7]), .Z(n22847));
    PFUMX i20825 (.BLUT(n23279), .ALUT(n23280), .C0(index_q[8]), .Z(n23281));
    PFUMX i20414 (.BLUT(n22866), .ALUT(n22867), .C0(index_q[8]), .Z(n22870));
    L6MUX21 i20415 (.D0(n22868), .D1(n22869), .SD(index_q[8]), .Z(n22871));
    PFUMX i20850 (.BLUT(n23298), .ALUT(n23299), .C0(index_i[7]), .Z(n23306));
    PFUMX i20851 (.BLUT(n23300), .ALUT(n23301), .C0(index_i[7]), .Z(n23307));
    PFUMX i20949 (.BLUT(n557), .ALUT(n572), .C0(index_q[4]), .Z(n23405));
    PFUMX i20950 (.BLUT(n589), .ALUT(n604), .C0(index_q[4]), .Z(n23406));
    PFUMX i19703 (.BLUT(n22138), .ALUT(n22139), .C0(index_q[4]), .Z(n22140));
    PFUMX i20951 (.BLUT(n620_adj_2251), .ALUT(n635_adj_2252), .C0(index_q[4]), 
          .Z(n23407));
    PFUMX i20550 (.BLUT(n23002), .ALUT(n23003), .C0(index_i[4]), .Z(n23006));
    PFUMX i23645 (.BLUT(n25412), .ALUT(n25409), .C0(index_q[6]), .Z(n25413));
    PFUMX i20952 (.BLUT(n653), .ALUT(n668), .C0(index_q[4]), .Z(n23408));
    PFUMX i20953 (.BLUT(n684), .ALUT(n699), .C0(index_q[4]), .Z(n23409));
    LUT4 i20404_3_lut (.A(n23081), .B(n21729), .C(index_q[6]), .Z(n22860)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20404_3_lut.init = 16'hcaca;
    PFUMX i24743 (.BLUT(n27143), .ALUT(n27144), .C0(index_q[0]), .Z(n27145));
    LUT4 mux_197_Mux_6_i653_3_lut (.A(n27106), .B(n652), .C(index_q[3]), 
         .Z(n653_adj_2253)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_6_i653_3_lut.init = 16'hcaca;
    PFUMX i20954 (.BLUT(n716), .ALUT(n731), .C0(index_q[4]), .Z(n23410));
    PFUMX i20978 (.BLUT(n23432), .ALUT(n23433), .C0(index_q[8]), .Z(n23434));
    LUT4 mux_197_Mux_6_i668_3_lut (.A(n660), .B(n27105), .C(index_q[3]), 
         .Z(n668_adj_2254)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_6_i668_3_lut.init = 16'hcaca;
    LUT4 i20403_3_lut (.A(n190), .B(n253), .C(index_q[6]), .Z(n22859)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20403_3_lut.init = 16'hcaca;
    PFUMX i20955 (.BLUT(n747), .ALUT(n762), .C0(index_q[4]), .Z(n23411));
    FD1P3AX phase_q__i1 (.D(o_phase[0]), .SP(i_resetb_c), .CK(dac_clk_p_c), 
            .Q(phase_q[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_q__i1.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i14 (.D(quarter_wave_sample_register_i_15__N_2126[14]), 
            .CK(dac_clk_p_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_i[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i14.GSR = "DISABLED";
    LUT4 mux_197_Mux_4_i541_3_lut_4_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n541)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_4_i541_3_lut_4_lut_3_lut_4_lut.init = 16'h0ef0;
    L6MUX21 i20653 (.D0(n23104), .D1(n23105), .SD(index_q[7]), .Z(n23109));
    FD1S3BX quarter_wave_sample_register_i_i13 (.D(quarter_wave_sample_register_i_15__N_2126[13]), 
            .CK(dac_clk_p_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_i[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i13.GSR = "DISABLED";
    LUT4 mux_197_Mux_12_i254_4_lut (.A(n26733), .B(n20559), .C(index_q[6]), 
         .D(n26861), .Z(n254_adj_2255)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_12_i254_4_lut.init = 16'hca0a;
    LUT4 mux_197_Mux_6_i812_3_lut_4_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n812)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(D))+!A !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_6_i812_3_lut_4_lut_3_lut_4_lut.init = 16'h7780;
    FD1S3BX quarter_wave_sample_register_i_i12 (.D(quarter_wave_sample_register_i_15__N_2126[12]), 
            .CK(dac_clk_p_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_i[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i12.GSR = "DISABLED";
    PFUMX i20956 (.BLUT(n781), .ALUT(n796), .C0(index_q[4]), .Z(n23412));
    FD1S3BX quarter_wave_sample_register_i_i11 (.D(quarter_wave_sample_register_i_15__N_2126[11]), 
            .CK(dac_clk_p_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_i[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i11.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_540_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n26863)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_2_lut_rep_540_3_lut_4_lut.init = 16'h8000;
    LUT4 i9397_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n11958)) /* synthesis lut_function=(!(A (B (D)+!B (C+!(D)))+!A !(B (D)+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9397_3_lut_4_lut_4_lut.init = 16'h4699;
    LUT4 mux_197_Mux_6_i684_3_lut (.A(n26887), .B(n29485), .C(index_q[3]), 
         .Z(n684_adj_2256)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_6_i684_3_lut.init = 16'hcaca;
    FD1S3BX quarter_wave_sample_register_i_i10 (.D(quarter_wave_sample_register_i_15__N_2126[10]), 
            .CK(dac_clk_p_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_i[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i10.GSR = "DISABLED";
    PFUMX i20957 (.BLUT(n812_adj_2257), .ALUT(n11914), .C0(index_q[4]), 
          .Z(n23413));
    FD1S3BX quarter_wave_sample_register_i_i9 (.D(quarter_wave_sample_register_i_15__N_2126[9]), 
            .CK(dac_clk_p_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_i[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i9.GSR = "DISABLED";
    LUT4 mux_196_Mux_2_i557_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n557_adj_2258)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C+!(D))+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_2_i557_3_lut_3_lut_4_lut.init = 16'h0f18;
    LUT4 i19627_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n22064)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A (B (D)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19627_3_lut_4_lut.init = 16'h18cc;
    FD1S3BX quarter_wave_sample_register_i_i8 (.D(quarter_wave_sample_register_i_15__N_2126[8]), 
            .CK(dac_clk_p_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_i[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i8.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i7 (.D(quarter_wave_sample_register_i_15__N_2126[7]), 
            .CK(dac_clk_p_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_i[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i7.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i1 (.D(\o_val_pipeline_q[0] [7]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(o_baseband_q_c_7)) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_q_1__i1.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i6 (.D(quarter_wave_sample_register_i_15__N_2126[6]), 
            .CK(dac_clk_p_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_i[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i6.GSR = "DISABLED";
    FD1S3DX phase_negation_i_i0 (.D(phase_i[11]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(phase_negation_i[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_negation_i_i0.GSR = "DISABLED";
    FD1S3DX phase_negation_q_i0 (.D(phase_q[11]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(phase_negation_q[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_negation_q_i0.GSR = "DISABLED";
    FD1S3DX index_i_i0 (.D(index_i_9__N_2106[0]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(index_i[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_i_i0.GSR = "DISABLED";
    FD1S3DX index_q_i0 (.D(index_q_9__N_2116[0]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(index_q[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_q_i0.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i0 (.D(quarter_wave_sample_register_q_15__N_2141[0]), 
            .CK(dac_clk_p_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_q[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_q_i0.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i1 (.D(\o_val_pipeline_i[0] [7]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(o_baseband_i_c_7)) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i1.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i0 (.D(quarter_wave_sample_register_i_15__N_2126[0]), 
            .CK(dac_clk_p_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_i[0])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i0.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i5 (.D(quarter_wave_sample_register_i_15__N_2126[5]), 
            .CK(dac_clk_p_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_i[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i5.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i4 (.D(quarter_wave_sample_register_i_15__N_2126[4]), 
            .CK(dac_clk_p_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_i[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i4.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i3 (.D(quarter_wave_sample_register_i_15__N_2126[3]), 
            .CK(dac_clk_p_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_i[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i3.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_i_i2 (.D(quarter_wave_sample_register_i_15__N_2126[2]), 
            .CK(dac_clk_p_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_i[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i2.GSR = "DISABLED";
    LUT4 i19584_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n22021)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)))+!A !(B (C+!(D))+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19584_3_lut_3_lut_4_lut.init = 16'h71cc;
    LUT4 mux_196_Mux_8_i30_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n30)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A !(B ((D)+!C)+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_8_i30_3_lut_3_lut_4_lut.init = 16'h7e0f;
    LUT4 i20462_3_lut_4_lut (.A(n26893), .B(index_q[3]), .C(index_q[4]), 
         .D(n364), .Z(n22918)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20462_3_lut_4_lut.init = 16'h8f80;
    FD1S3BX quarter_wave_sample_register_i_i1 (.D(quarter_wave_sample_register_i_15__N_2126[1]), 
            .CK(dac_clk_p_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_i[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_i_i1.GSR = "DISABLED";
    PFUMX i20958 (.BLUT(n844), .ALUT(n11917), .C0(index_q[4]), .Z(n23414));
    FD1S3DX o_val_pipeline_i_1__i18 (.D(o_val_pipeline_i_0__15__N_2156), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(\o_val_pipeline_i[0] [15])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i18.GSR = "DISABLED";
    PFUMX i20959 (.BLUT(n875), .ALUT(n890), .C0(index_q[4]), .Z(n23415));
    LUT4 i22580_2_lut_rep_586 (.A(index_i[1]), .B(index_i[2]), .Z(n26909)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i22580_2_lut_rep_586.init = 16'h9999;
    FD1S3DX o_val_pipeline_i_1__i17 (.D(o_val_pipeline_i_0__15__N_2158), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(\o_val_pipeline_i[0] [14])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i17.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i16 (.D(o_val_pipeline_i_0__15__N_2160), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(\o_val_pipeline_i[0] [13])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i16.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i15 (.D(o_val_pipeline_i_0__15__N_2162), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(\o_val_pipeline_i[0] [12])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i15.GSR = "DISABLED";
    LUT4 mux_196_Mux_4_i204_3_lut_4_lut_4_lut_3_lut_rep_654 (.A(index_i[0]), 
         .B(index_i[2]), .C(index_i[1]), .Z(n26977)) /* synthesis lut_function=(!(A (B+(C))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_4_i204_3_lut_4_lut_4_lut_3_lut_rep_654.init = 16'h4646;
    FD1S3DX o_val_pipeline_i_1__i14 (.D(o_val_pipeline_i_0__15__N_2164), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(\o_val_pipeline_i[0] [11])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i14.GSR = "DISABLED";
    PFUMX i20551 (.BLUT(n23004), .ALUT(n23005), .C0(index_i[4]), .Z(n23007));
    PFUMX i20960 (.BLUT(n908), .ALUT(n923), .C0(index_q[4]), .Z(n23416));
    FD1S3DX o_val_pipeline_i_1__i13 (.D(o_val_pipeline_i_0__15__N_2166), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(\o_val_pipeline_i[0] [10])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i13.GSR = "DISABLED";
    PFUMX i21040 (.BLUT(n23494), .ALUT(n23495), .C0(index_i[8]), .Z(n23496));
    FD1S3DX o_val_pipeline_i_1__i12 (.D(o_val_pipeline_i_0__15__N_2168), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(\o_val_pipeline_i[0] [9])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i12.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i11 (.D(o_val_pipeline_i_0__15__N_2170), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(\o_val_pipeline_i[0] [8])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i11.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i10 (.D(o_val_pipeline_i_0__15__N_2172), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(\o_val_pipeline_i[0] [7])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i10.GSR = "DISABLED";
    PFUMX i20961 (.BLUT(n939), .ALUT(n954), .C0(index_q[4]), .Z(n23417));
    LUT4 mux_196_Mux_6_i860_3_lut_3_lut (.A(n26748), .B(index_i[4]), .C(n844_adj_2259), 
         .Z(n860)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam mux_196_Mux_6_i860_3_lut_3_lut.init = 16'h7474;
    FD1S3DX o_val_pipeline_i_1__i9 (.D(\o_val_pipeline_i[0] [15]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(o_baseband_i_c_15)) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i9.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i8 (.D(\o_val_pipeline_i[0] [14]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(o_baseband_i_c_14)) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i8.GSR = "DISABLED";
    L6MUX21 i20199 (.D0(n22650), .D1(n22651), .SD(index_q[7]), .Z(n22655));
    L6MUX21 i20220 (.D0(n22670), .D1(n22671), .SD(index_i[7]), .Z(n22676));
    L6MUX21 i20221 (.D0(n22672), .D1(n22673), .SD(index_i[7]), .Z(n22677));
    PFUMX i20962 (.BLUT(n971), .ALUT(n986), .C0(index_q[4]), .Z(n23418));
    LUT4 n442_bdd_2_lut_23803_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[3]), 
         .Z(n25583)) /* synthesis lut_function=(A (B+(C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n442_bdd_2_lut_23803_3_lut.init = 16'hf9f9;
    FD1S3DX o_val_pipeline_i_1__i7 (.D(\o_val_pipeline_i[0] [13]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(o_baseband_i_c_13)) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i7.GSR = "DISABLED";
    PFUMX i24803 (.BLUT(n27236), .ALUT(n27237), .C0(index_i[3]), .Z(n62));
    PFUMX i20963 (.BLUT(n1002), .ALUT(n1017), .C0(index_q[4]), .Z(n23419));
    FD1S3DX o_val_pipeline_i_1__i6 (.D(\o_val_pipeline_i[0] [12]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(o_baseband_i_c_12)) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i6.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i5 (.D(\o_val_pipeline_i[0] [11]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(o_baseband_i_c_11)) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i5.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i4 (.D(\o_val_pipeline_i[0] [10]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(o_baseband_i_c_10)) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i4.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i3 (.D(\o_val_pipeline_i[0] [9]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(n3655)) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i3.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_i_1__i2 (.D(\o_val_pipeline_i[0] [8]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(o_baseband_i_c_8)) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_i_1__i2.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i11 (.D(o_phase[11]), .SP(i_resetb_c), .CK(dac_clk_p_c), 
            .Q(phase_i[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i11.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i10 (.D(o_phase[10]), .SP(i_resetb_c), .CK(dac_clk_p_c), 
            .Q(phase_i[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i10.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i9 (.D(o_phase[9]), .SP(i_resetb_c), .CK(dac_clk_p_c), 
            .Q(phase_i[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i9.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i8 (.D(o_phase[8]), .SP(i_resetb_c), .CK(dac_clk_p_c), 
            .Q(phase_i[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i8.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i7 (.D(o_phase[7]), .SP(i_resetb_c), .CK(dac_clk_p_c), 
            .Q(phase_i[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i7.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i6 (.D(o_phase[6]), .SP(i_resetb_c), .CK(dac_clk_p_c), 
            .Q(phase_i[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i6.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i5 (.D(o_phase[5]), .SP(i_resetb_c), .CK(dac_clk_p_c), 
            .Q(phase_i[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i5.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i4 (.D(o_phase[4]), .SP(i_resetb_c), .CK(dac_clk_p_c), 
            .Q(phase_i[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i4.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i3 (.D(o_phase[3]), .SP(i_resetb_c), .CK(dac_clk_p_c), 
            .Q(phase_i[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i3.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i2 (.D(o_phase[2]), .SP(i_resetb_c), .CK(dac_clk_p_c), 
            .Q(phase_i[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i2.GSR = "DISABLED";
    FD1P3AX phase_i_i0_i1 (.D(o_phase[1]), .SP(i_resetb_c), .CK(dac_clk_p_c), 
            .Q(phase_i[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_i_i0_i1.GSR = "DISABLED";
    L6MUX21 i20249 (.D0(n22697), .D1(n22698), .SD(index_i[7]), .Z(n22705));
    L6MUX21 i20250 (.D0(n22699), .D1(n22700), .SD(index_i[7]), .Z(n22706));
    L6MUX21 i20266 (.D0(n22716), .D1(n22717), .SD(index_q[7]), .Z(n22722));
    PFUMX i20267 (.BLUT(n22718), .ALUT(n22719), .C0(index_q[7]), .Z(n22723));
    LUT4 index_i_5__bdd_3_lut_23790_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n25493)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C))+!A (B (C (D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam index_i_5__bdd_3_lut_23790_3_lut_4_lut.init = 16'h0fc7;
    FD1S3BX quarter_wave_sample_register_q_i15 (.D(n29501), .CK(dac_clk_p_c), 
            .PD(i_resetb_N_301), .Q(\quarter_wave_sample_register_q[15] )) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_q_i15.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i14 (.D(quarter_wave_sample_register_q_15__N_2141[14]), 
            .CK(dac_clk_p_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_q[14])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_q_i14.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i13 (.D(quarter_wave_sample_register_q_15__N_2141[13]), 
            .CK(dac_clk_p_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_q[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_q_i13.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i12 (.D(quarter_wave_sample_register_q_15__N_2141[12]), 
            .CK(dac_clk_p_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_q[12])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_q_i12.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i11 (.D(quarter_wave_sample_register_q_15__N_2141[11]), 
            .CK(dac_clk_p_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_q[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_q_i11.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i10 (.D(quarter_wave_sample_register_q_15__N_2141[10]), 
            .CK(dac_clk_p_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_q[10])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_q_i10.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i9 (.D(quarter_wave_sample_register_q_15__N_2141[9]), 
            .CK(dac_clk_p_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_q[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_q_i9.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i8 (.D(quarter_wave_sample_register_q_15__N_2141[8]), 
            .CK(dac_clk_p_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_q[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_q_i8.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i7 (.D(quarter_wave_sample_register_q_15__N_2141[7]), 
            .CK(dac_clk_p_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_q[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_q_i7.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i6 (.D(quarter_wave_sample_register_q_15__N_2141[6]), 
            .CK(dac_clk_p_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_q[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_q_i6.GSR = "DISABLED";
    LUT4 mux_196_Mux_6_i781_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n781_adj_2260)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A (B (C (D)+!C !(D))+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_6_i781_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hc837;
    FD1S3BX quarter_wave_sample_register_q_i5 (.D(quarter_wave_sample_register_q_15__N_2141[5]), 
            .CK(dac_clk_p_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_q[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_q_i5.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i4 (.D(quarter_wave_sample_register_q_15__N_2141[4]), 
            .CK(dac_clk_p_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_q[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_q_i4.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i3 (.D(quarter_wave_sample_register_q_15__N_2141[3]), 
            .CK(dac_clk_p_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_q[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_q_i3.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i2 (.D(quarter_wave_sample_register_q_15__N_2141[2]), 
            .CK(dac_clk_p_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_q[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_q_i2.GSR = "DISABLED";
    FD1S3BX quarter_wave_sample_register_q_i1 (.D(quarter_wave_sample_register_q_15__N_2141[1]), 
            .CK(dac_clk_p_c), .PD(i_resetb_N_301), .Q(quarter_wave_sample_register_q[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam quarter_wave_sample_register_q_i1.GSR = "DISABLED";
    FD1S3DX index_q_i9 (.D(index_q_9__N_2116[9]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(index_q[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_q_i9.GSR = "DISABLED";
    FD1S3DX index_q_i8 (.D(index_q_9__N_2116[8]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(index_q[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_q_i8.GSR = "DISABLED";
    FD1S3DX index_q_i7 (.D(index_q_9__N_2116[7]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(index_q[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_q_i7.GSR = "DISABLED";
    FD1S3DX index_q_i6 (.D(index_q_9__N_2116[6]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(index_q[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_q_i6.GSR = "DISABLED";
    LUT4 i19611_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n22048)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+(D)))+!A !(B (D)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19611_3_lut_4_lut_4_lut.init = 16'h99c7;
    FD1S3DX index_q_i5 (.D(index_q_9__N_2116[5]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(index_q[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_q_i5.GSR = "DISABLED";
    FD1S3DX index_q_i4 (.D(index_q_9__N_2116[4]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(index_q[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_q_i4.GSR = "DISABLED";
    FD1S3DX index_q_i3 (.D(index_q_9__N_2116[3]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(index_q[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_q_i3.GSR = "DISABLED";
    FD1S3DX index_q_i2 (.D(index_q_9__N_2116[2]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(index_q[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_q_i2.GSR = "DISABLED";
    FD1S3DX index_q_i1 (.D(index_q_9__N_2116[1]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(index_q[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_q_i1.GSR = "DISABLED";
    FD1S3DX index_i_i9 (.D(index_i_9__N_2106[9]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(index_i[9])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_i_i9.GSR = "DISABLED";
    L6MUX21 i20324 (.D0(n22770), .D1(n22771), .SD(index_i[6]), .Z(n22780));
    FD1S3DX index_i_i8 (.D(index_i_9__N_2106[8]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(index_i[8])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_i_i8.GSR = "DISABLED";
    LUT4 mux_197_Mux_10_i62_3_lut_3_lut_4_lut (.A(n26893), .B(index_q[3]), 
         .C(n26856), .D(index_q[4]), .Z(n62_adj_2261)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_10_i62_3_lut_3_lut_4_lut.init = 16'hf077;
    L6MUX21 i20326 (.D0(n22774), .D1(n22775), .SD(index_i[7]), .Z(n22782));
    L6MUX21 i20327 (.D0(n22776), .D1(n22777), .SD(index_i[7]), .Z(n22783));
    FD1S3DX index_i_i7 (.D(index_i_9__N_2106[7]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(index_i[7])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_i_i7.GSR = "DISABLED";
    FD1S3DX index_i_i6 (.D(index_i_9__N_2106[6]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(index_i[6])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_i_i6.GSR = "DISABLED";
    FD1S3DX index_i_i5 (.D(index_i_9__N_2106[5]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(index_i[5])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_i_i5.GSR = "DISABLED";
    FD1S3DX index_i_i4 (.D(index_i_9__N_2106[4]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(index_i[4])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_i_i4.GSR = "DISABLED";
    LUT4 i20866_3_lut (.A(n23315), .B(n23316), .C(index_i[7]), .Z(n23322)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20866_3_lut.init = 16'hcaca;
    FD1S3DX index_i_i3 (.D(index_i_9__N_2106[3]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(index_i[3])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_i_i3.GSR = "DISABLED";
    FD1S3DX index_i_i2 (.D(index_i_9__N_2106[2]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(index_i[2])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_i_i2.GSR = "DISABLED";
    FD1S3DX index_i_i1 (.D(index_i_9__N_2106[1]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(index_i[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam index_i_i1.GSR = "DISABLED";
    FD1S3DX phase_negation_q_i1 (.D(phase_negation_q[0]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(phase_negation_q[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_negation_q_i1.GSR = "DISABLED";
    FD1S3DX phase_negation_i_i1 (.D(phase_negation_i[0]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(phase_negation_i[1])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_negation_i_i1.GSR = "DISABLED";
    PFUMX i21020 (.BLUT(n844_adj_2262), .ALUT(n12112), .C0(index_i[4]), 
          .Z(n23476));
    FD1S3DX o_val_pipeline_q_1__i18 (.D(n1829[14]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(\o_val_pipeline_q[0] [15])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_q_1__i18.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i17 (.D(n1829[13]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(\o_val_pipeline_q[0] [14])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_q_1__i17.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i16 (.D(n1829[12]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(\o_val_pipeline_q[0] [13])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_q_1__i16.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i15 (.D(n1829[11]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(\o_val_pipeline_q[0] [12])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_q_1__i15.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i14 (.D(n1829[10]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(\o_val_pipeline_q[0] [11])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_q_1__i14.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i13 (.D(n1829[9]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(\o_val_pipeline_q[0] [10])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_q_1__i13.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i12 (.D(n1829[8]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(\o_val_pipeline_q[0] [9])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_q_1__i12.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i11 (.D(n1829[7]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(\o_val_pipeline_q[0] [8])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_q_1__i11.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i10 (.D(n1829[6]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(\o_val_pipeline_q[0] [7])) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_q_1__i10.GSR = "DISABLED";
    LUT4 n903_bdd_3_lut_4_lut_3_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .Z(n26416)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n903_bdd_3_lut_4_lut_3_lut.init = 16'h6161;
    L6MUX21 i20358 (.D0(n22807), .D1(n22808), .SD(index_i[7]), .Z(n22814));
    FD1S3DX o_val_pipeline_q_1__i9 (.D(\o_val_pipeline_q[0] [15]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(o_baseband_q_c_15)) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_q_1__i9.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i8 (.D(\o_val_pipeline_q[0] [14]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(o_baseband_q_c_14)) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_q_1__i8.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i7 (.D(\o_val_pipeline_q[0] [13]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(o_baseband_q_c_13)) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_q_1__i7.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i6 (.D(\o_val_pipeline_q[0] [12]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(o_baseband_q_c_12)) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_q_1__i6.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i5 (.D(\o_val_pipeline_q[0] [11]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(o_baseband_q_c_11)) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_q_1__i5.GSR = "DISABLED";
    LUT4 i20622_3_lut (.A(n851), .B(n27058), .C(index_q[3]), .Z(n23078)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20622_3_lut.init = 16'hcaca;
    L6MUX21 i20359 (.D0(n22809), .D1(n22810), .SD(index_i[7]), .Z(n22815));
    PFUMX i20360 (.BLUT(n22811), .ALUT(n22812), .C0(index_i[7]), .Z(n22816));
    LUT4 i19575_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n22012)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B (C+!(D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19575_3_lut_4_lut_4_lut.init = 16'h3c38;
    FD1S3DX o_val_pipeline_q_1__i4 (.D(\o_val_pipeline_q[0] [10]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(o_baseband_q_c_10)) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_q_1__i4.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i3 (.D(\o_val_pipeline_q[0] [9]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(n3656)) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_q_1__i3.GSR = "DISABLED";
    FD1S3DX o_val_pipeline_q_1__i2 (.D(\o_val_pipeline_q[0] [8]), .CK(dac_clk_p_c), 
            .CD(i_resetb_N_301), .Q(o_baseband_q_c_8)) /* synthesis syn_pipeline=1, LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam o_val_pipeline_q_1__i2.GSR = "DISABLED";
    L6MUX21 i20385 (.D0(n22830), .D1(n22831), .SD(index_i[6]), .Z(n22841));
    LUT4 mux_197_Mux_0_i986_3_lut (.A(n29495), .B(n985), .C(index_q[3]), 
         .Z(n986)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i986_3_lut.init = 16'hcaca;
    PFUMX mux_196_Mux_2_i891 (.BLUT(n875_adj_2263), .ALUT(n890_adj_2264), 
          .C0(index_i[4]), .Z(n891)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    L6MUX21 i20386 (.D0(n22832), .D1(n22833), .SD(index_i[6]), .Z(n22842));
    L6MUX21 i20389 (.D0(n22838), .D1(n22839), .SD(index_i[7]), .Z(n22845));
    L6MUX21 i20396 (.D0(n382), .D1(n509), .SD(index_q[7]), .Z(n22852));
    PFUMX i20557 (.BLUT(n23009), .ALUT(n23010), .C0(index_i[4]), .Z(n23013));
    PFUMX mux_196_Mux_2_i860 (.BLUT(n844_adj_2265), .ALUT(n859), .C0(index_i[4]), 
          .Z(n860_adj_2266)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    L6MUX21 i20412 (.D0(n22862), .D1(n22863), .SD(index_q[7]), .Z(n22868));
    L6MUX21 i20413 (.D0(n22864), .D1(n22865), .SD(index_q[7]), .Z(n22869));
    LUT4 mux_196_Mux_7_i716_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n716_adj_2267)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C+!(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_7_i716_3_lut_3_lut_4_lut.init = 16'h0f81;
    PFUMX i20558 (.BLUT(n23011), .ALUT(n23012), .C0(index_i[4]), .Z(n23014));
    L6MUX21 i20852 (.D0(n23302), .D1(n23303), .SD(index_i[7]), .Z(n23308));
    L6MUX21 i20867 (.D0(n23317), .D1(n23318), .SD(index_i[7]), .Z(n23323));
    CCU2D add_376_15 (.A0(quarter_wave_sample_register_i[14]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(\quarter_wave_sample_register_q[15] ), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17597), .S0(o_val_pipeline_i_0__15__N_2157[14]), 
          .S1(o_val_pipeline_i_0__15__N_2157[15]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam add_376_15.INIT0 = 16'hf555;
    defparam add_376_15.INIT1 = 16'hf555;
    defparam add_376_15.INJECT1_0 = "NO";
    defparam add_376_15.INJECT1_1 = "NO";
    PFUMX i20868 (.BLUT(n23319), .ALUT(n23320), .C0(index_i[7]), .Z(n23324));
    CCU2D add_376_13 (.A0(quarter_wave_sample_register_i[12]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[13]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17596), .COUT(n17597), 
          .S0(o_val_pipeline_i_0__15__N_2157[12]), .S1(o_val_pipeline_i_0__15__N_2157[13]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam add_376_13.INIT0 = 16'hf555;
    defparam add_376_13.INIT1 = 16'hf555;
    defparam add_376_13.INJECT1_0 = "NO";
    defparam add_376_13.INJECT1_1 = "NO";
    CCU2D add_376_11 (.A0(quarter_wave_sample_register_i[10]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[11]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17595), .COUT(n17596), 
          .S0(o_val_pipeline_i_0__15__N_2157[10]), .S1(o_val_pipeline_i_0__15__N_2157[11]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam add_376_11.INIT0 = 16'hf555;
    defparam add_376_11.INIT1 = 16'hf555;
    defparam add_376_11.INJECT1_0 = "NO";
    defparam add_376_11.INJECT1_1 = "NO";
    LUT4 i19705_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n22142)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C+(D)))+!A (B (C (D)+!C !(D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19705_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h3ef0;
    FD1P3AX phase_q__i11 (.D(phase_q_11__N_2232[11]), .SP(i_resetb_c), .CK(dac_clk_p_c), 
            .Q(phase_q[11])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam phase_q__i11.GSR = "DISABLED";
    LUT4 i20621_3_lut (.A(n652), .B(n27102), .C(index_q[3]), .Z(n23077)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20621_3_lut.init = 16'hcaca;
    PFUMX i24799 (.BLUT(n27230), .ALUT(n27231), .C0(index_i[1]), .Z(n27232));
    L6MUX21 i20878 (.D0(n23332), .D1(n23333), .SD(index_i[7]), .Z(n23334));
    L6MUX21 i20540 (.D0(n22989), .D1(n22990), .SD(index_q[7]), .Z(n22996));
    L6MUX21 i20541 (.D0(n22991), .D1(n22992), .SD(index_q[7]), .Z(n22997));
    LUT4 i18979_3_lut (.A(n27080), .B(n27099), .C(index_q[3]), .Z(n21416)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18979_3_lut.init = 16'hcaca;
    PFUMX i20542 (.BLUT(n22993), .ALUT(n22994), .C0(index_q[7]), .Z(n22998));
    PFUMX i19319 (.BLUT(n21754), .ALUT(n21755), .C0(index_q[4]), .Z(n21756));
    PFUMX i20564 (.BLUT(n23016), .ALUT(n23017), .C0(index_i[4]), .Z(n23020));
    L6MUX21 i20038 (.D0(n22488), .D1(n22489), .SD(index_q[7]), .Z(n22494));
    PFUMX i20565 (.BLUT(n23018), .ALUT(n23019), .C0(index_i[4]), .Z(n23021));
    L6MUX21 i20647 (.D0(n23092), .D1(n23093), .SD(index_q[6]), .Z(n23103));
    LUT4 i18978_3_lut (.A(n27095), .B(n356), .C(index_q[3]), .Z(n21415)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18978_3_lut.init = 16'hcaca;
    PFUMX i19322 (.BLUT(n21757), .ALUT(n21758), .C0(index_q[4]), .Z(n21759));
    L6MUX21 i20648 (.D0(n23094), .D1(n23095), .SD(index_q[6]), .Z(n23104));
    CCU2D add_376_9 (.A0(quarter_wave_sample_register_i[8]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[9]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17594), .COUT(n17595), 
          .S0(o_val_pipeline_i_0__15__N_2157[8]), .S1(o_val_pipeline_i_0__15__N_2157[9]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam add_376_9.INIT0 = 16'hf555;
    defparam add_376_9.INIT1 = 16'hf555;
    defparam add_376_9.INJECT1_0 = "NO";
    defparam add_376_9.INJECT1_1 = "NO";
    L6MUX21 i20651 (.D0(n23100), .D1(n23101), .SD(index_q[7]), .Z(n23107));
    LUT4 i19336_3_lut_4_lut (.A(n27085), .B(index_q[2]), .C(index_q[3]), 
         .D(n29495), .Z(n21773)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19336_3_lut_4_lut.init = 16'hf404;
    LUT4 i20865_3_lut (.A(n23313), .B(n25001), .C(index_i[7]), .Z(n23321)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20865_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_3_i653_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n653_adj_2268)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A !(B (D)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_3_i653_3_lut_4_lut_4_lut.init = 16'h4d99;
    L6MUX21 i20119 (.D0(n22567), .D1(n22568), .SD(index_q[7]), .Z(n22575));
    LUT4 i20870_3_lut (.A(n23323), .B(n23324), .C(index_i[8]), .Z(n23326)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20870_3_lut.init = 16'hcaca;
    LUT4 i11238_2_lut_rep_531_3_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .Z(n26854)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11238_2_lut_rep_531_3_lut.init = 16'he0e0;
    PFUMX i19328 (.BLUT(n21763), .ALUT(n21764), .C0(index_q[4]), .Z(n21765));
    L6MUX21 i20120 (.D0(n22569), .D1(n22570), .SD(index_q[7]), .Z(n22576));
    LUT4 i21605_3_lut (.A(n21415), .B(n21416), .C(index_q[4]), .Z(n21417)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21605_3_lut.init = 16'hcaca;
    CCU2D add_376_7 (.A0(quarter_wave_sample_register_i[6]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[7]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17593), .COUT(n17594), 
          .S1(o_val_pipeline_i_0__15__N_2157[7]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam add_376_7.INIT0 = 16'hf555;
    defparam add_376_7.INIT1 = 16'hf555;
    defparam add_376_7.INJECT1_0 = "NO";
    defparam add_376_7.INJECT1_1 = "NO";
    PFUMX i19334 (.BLUT(n21769), .ALUT(n21770), .C0(index_q[4]), .Z(n21771));
    LUT4 i9599_3_lut_4_lut_3_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[4]), 
         .Z(n12164)) /* synthesis lut_function=(A (B)+!A !(B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9599_3_lut_4_lut_3_lut.init = 16'h9898;
    LUT4 mux_197_Mux_8_i397_3_lut_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n397)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_8_i397_3_lut_3_lut_3_lut_4_lut.init = 16'hf10f;
    PFUMX mux_196_Mux_3_i763 (.BLUT(n747_adj_2269), .ALUT(n762_adj_2270), 
          .C0(index_i[4]), .Z(n763)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    PFUMX i19337 (.BLUT(n21772), .ALUT(n21773), .C0(index_q[4]), .Z(n21774));
    LUT4 i20853_3_lut (.A(n23304), .B(n23305), .C(index_i[7]), .Z(n23309)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20853_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_0_i93_3_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .Z(n93)) /* synthesis lut_function=(A (B)+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_0_i93_3_lut_3_lut.init = 16'h9c9c;
    L6MUX21 i19130 (.D0(n21565), .D1(n21566), .SD(index_i[7]), .Z(n21567));
    LUT4 i20845_3_lut (.A(n23288), .B(n24971), .C(index_i[6]), .Z(n23301)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20845_3_lut.init = 16'hcaca;
    PFUMX i19340 (.BLUT(n21775), .ALUT(n21776), .C0(index_q[4]), .Z(n21777));
    LUT4 i11272_3_lut_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n13947)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11272_3_lut_3_lut_3_lut_4_lut.init = 16'h10ff;
    LUT4 mux_196_Mux_4_i77_3_lut_4_lut_3_lut_rep_655 (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[1]), .Z(n26978)) /* synthesis lut_function=(A (B (C))+!A !(B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_4_i77_3_lut_4_lut_3_lut_rep_655.init = 16'h9595;
    PFUMX i24738 (.BLUT(n27135), .ALUT(n27136), .C0(index_i[1]), .Z(n27137));
    L6MUX21 i20725 (.D0(n23179), .D1(n23180), .SD(index_q[7]), .Z(n23181));
    LUT4 mux_197_Mux_5_i475_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n475)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_5_i475_3_lut_4_lut_4_lut.init = 16'hd4a5;
    L6MUX21 i19139 (.D0(n21574), .D1(n21575), .SD(index_q[7]), .Z(n21576));
    L6MUX21 i20194 (.D0(n22640), .D1(n22641), .SD(index_q[6]), .Z(n22650));
    L6MUX21 i20196 (.D0(n22644), .D1(n22645), .SD(index_q[7]), .Z(n22652));
    L6MUX21 i20197 (.D0(n22646), .D1(n22647), .SD(index_q[7]), .Z(n22653));
    L6MUX21 i20204 (.D0(n382_adj_2271), .D1(n509_adj_2272), .SD(index_i[7]), 
            .Z(n22660));
    L6MUX21 i20213 (.D0(n21684), .D1(n21687), .SD(index_i[6]), .Z(n22669));
    L6MUX21 i20214 (.D0(n21690), .D1(n21693), .SD(index_i[6]), .Z(n22670));
    L6MUX21 i20215 (.D0(n21696), .D1(n21699), .SD(index_i[6]), .Z(n22671));
    LUT4 n22037_bdd_3_lut_3_lut (.A(index_i[1]), .B(n526), .C(index_i[4]), 
         .Z(n24904)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n22037_bdd_3_lut_3_lut.init = 16'h5c5c;
    CCU2D add_376_5 (.A0(quarter_wave_sample_register_i[4]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[5]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17592), .COUT(n17593));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam add_376_5.INIT0 = 16'hf555;
    defparam add_376_5.INIT1 = 16'hf555;
    defparam add_376_5.INJECT1_0 = "NO";
    defparam add_376_5.INJECT1_1 = "NO";
    CCU2D add_376_3 (.A0(quarter_wave_sample_register_i[2]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_i[3]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17591), .COUT(n17592));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam add_376_3.INIT0 = 16'hf555;
    defparam add_376_3.INIT1 = 16'hf555;
    defparam add_376_3.INJECT1_0 = "NO";
    defparam add_376_3.INJECT1_1 = "NO";
    PFUMX i20216 (.BLUT(n21702), .ALUT(n892), .C0(index_i[6]), .Z(n22672));
    LUT4 i20844_3_lut (.A(n24964), .B(n23287), .C(index_i[6]), .Z(n23300)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20844_3_lut.init = 16'hcaca;
    LUT4 i11642_2_lut_rep_533_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n26856)) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11642_2_lut_rep_533_3_lut_4_lut.init = 16'he000;
    PFUMX i24791 (.BLUT(n27218), .ALUT(n27219), .C0(index_i[2]), .Z(n27220));
    LUT4 mux_197_Mux_0_i157_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n157)) /* synthesis lut_function=(A (B (C+!(D))+!B !(D))+!A (B (D)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i157_3_lut_4_lut.init = 16'hd4aa;
    LUT4 i20620_3_lut (.A(n29477), .B(n27104), .C(index_q[3]), .Z(n23076)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20620_3_lut.init = 16'hcaca;
    LUT4 i20619_3_lut (.A(n27058), .B(n27086), .C(index_q[3]), .Z(n23075)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20619_3_lut.init = 16'hcaca;
    LUT4 i20842_3_lut (.A(n25322), .B(n23283), .C(index_i[6]), .Z(n23298)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20842_3_lut.init = 16'hcaca;
    L6MUX21 i20241 (.D0(n22681), .D1(n22682), .SD(index_i[6]), .Z(n22697));
    LUT4 i20411_3_lut (.A(n22860), .B(n22861), .C(index_q[7]), .Z(n22867)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20411_3_lut.init = 16'hcaca;
    PFUMX i24789 (.BLUT(n27215), .ALUT(n27216), .C0(index_i[1]), .Z(n27217));
    LUT4 i18990_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21427)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18990_3_lut_4_lut.init = 16'h64cc;
    L6MUX21 i20242 (.D0(n22683), .D1(n22684), .SD(index_i[6]), .Z(n22698));
    LUT4 i20410_3_lut (.A(n22858), .B(n22859), .C(index_q[7]), .Z(n22866)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20410_3_lut.init = 16'hcaca;
    PFUMX i24787 (.BLUT(n27212), .ALUT(n27213), .C0(index_q[3]), .Z(n27214));
    CCU2D add_376_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(quarter_wave_sample_register_i[0]), .B1(quarter_wave_sample_register_i[1]), 
          .C1(GND_net), .D1(GND_net), .COUT(n17591));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(74[29:60])
    defparam add_376_1.INIT0 = 16'hF000;
    defparam add_376_1.INIT1 = 16'ha666;
    defparam add_376_1.INJECT1_0 = "NO";
    defparam add_376_1.INJECT1_1 = "NO";
    L6MUX21 i20243 (.D0(n22685), .D1(n22686), .SD(index_i[6]), .Z(n22699));
    L6MUX21 i20244 (.D0(n22687), .D1(n22688), .SD(index_i[6]), .Z(n22700));
    L6MUX21 i20245 (.D0(n22689), .D1(n22690), .SD(index_i[6]), .Z(n22701));
    L6MUX21 i20247 (.D0(n22693), .D1(n22694), .SD(index_i[6]), .Z(n22703));
    PFUMX i24785 (.BLUT(n27209), .ALUT(n27210), .C0(index_i[1]), .Z(n27211));
    PFUMX i20257 (.BLUT(n12116), .ALUT(n21711), .C0(index_q[6]), .Z(n22713));
    LUT4 i20615_3_lut (.A(n27061), .B(n27086), .C(index_q[3]), .Z(n23071)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20615_3_lut.init = 16'hcaca;
    L6MUX21 i20259 (.D0(n21717), .D1(n21720), .SD(index_q[6]), .Z(n22715));
    L6MUX21 i20260 (.D0(n574), .D1(n21723), .SD(index_q[6]), .Z(n22716));
    L6MUX21 i20261 (.D0(n21726), .D1(n764), .SD(index_q[6]), .Z(n22717));
    L6MUX21 i20757 (.D0(n23205), .D1(n23206), .SD(index_i[6]), .Z(n23213));
    L6MUX21 i20760 (.D0(n23211), .D1(n23212), .SD(index_i[6]), .Z(n23216));
    L6MUX21 i20287 (.D0(n22727), .D1(n22728), .SD(index_i[6]), .Z(n22743));
    L6MUX21 i20288 (.D0(n22729), .D1(n22730), .SD(index_i[6]), .Z(n22744));
    L6MUX21 i20289 (.D0(n22731), .D1(n22732), .SD(index_i[6]), .Z(n22745));
    LUT4 i19029_3_lut_3_lut_4_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n21466)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19029_3_lut_3_lut_4_lut_3_lut_4_lut.init = 16'h11ef;
    LUT4 mux_197_Mux_9_i316_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), 
         .B(index_q[2]), .C(index_q[3]), .D(index_q[0]), .Z(n316)) /* synthesis lut_function=(!(A (B (C)+!B !(C+(D)))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_9_i316_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h7e7c;
    LUT4 n11074_bdd_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .D(index_q[0]), .Z(n25734)) /* synthesis lut_function=(A (B (C)+!B ((D)+!C))+!A (B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n11074_bdd_3_lut_4_lut_4_lut_4_lut.init = 16'he7c7;
    PFUMX i20291 (.BLUT(n22735), .ALUT(n22736), .C0(index_i[6]), .Z(n22747));
    LUT4 i9551_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n12112)) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B ((D)+!C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9551_3_lut_4_lut_4_lut.init = 16'hcdad;
    LUT4 mux_197_Mux_3_i189_3_lut_3_lut_4_lut (.A(n26893), .B(index_q[3]), 
         .C(index_q[4]), .D(n26796), .Z(n189)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_3_i189_3_lut_3_lut_4_lut.init = 16'h08f8;
    LUT4 n78_bdd_3_lut_23991_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .D(index_q[0]), .Z(n25731)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A !((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n78_bdd_3_lut_23991_4_lut_4_lut_4_lut.init = 16'h7173;
    LUT4 mux_197_Mux_10_i637_3_lut_4_lut_4_lut (.A(n26872), .B(index_q[4]), 
         .C(index_q[5]), .D(n26772), .Z(n637)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_10_i637_3_lut_4_lut_4_lut.init = 16'h1f1c;
    LUT4 i9548_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n12109)) /* synthesis lut_function=(A (B (D)+!B !((D)+!C))+!A (((D)+!C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9548_3_lut_4_lut_4_lut_4_lut.init = 16'hdd35;
    PFUMX i24783 (.BLUT(n27206), .ALUT(n27207), .C0(index_i[0]), .Z(n27208));
    LUT4 n303_bdd_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[2]), .C(index_i[1]), 
         .D(index_i[3]), .Z(n25652)) /* synthesis lut_function=(!(A (B)+!A !(B (C+(D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n303_bdd_4_lut_4_lut_4_lut.init = 16'h6763;
    L6MUX21 i20292 (.D0(n22737), .D1(n22738), .SD(index_i[6]), .Z(n22748));
    LUT4 mux_196_Mux_4_i812_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[4]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n812_adj_2273)) /* synthesis lut_function=(A (B (C+(D)))+!A !(B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_4_i812_3_lut_3_lut_4_lut.init = 16'h9995;
    LUT4 i15550_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[1]), .Z(n17814)) /* synthesis lut_function=(A (B (C (D))+!B !(C))+!A (B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i15550_3_lut_4_lut_4_lut_4_lut.init = 16'hd656;
    LUT4 mux_197_Mux_0_i971_3_lut (.A(n29494), .B(n27107), .C(index_q[3]), 
         .Z(n971)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i971_3_lut.init = 16'hcaca;
    L6MUX21 i20293 (.D0(n22739), .D1(n22740), .SD(index_i[6]), .Z(n22749));
    PFUMX i20294 (.BLUT(n22741), .ALUT(n22742), .C0(index_i[6]), .Z(n22750));
    LUT4 i19288_3_lut_3_lut_4_lut (.A(n26871), .B(index_q[3]), .C(n93_adj_2274), 
         .D(index_q[4]), .Z(n21725)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19288_3_lut_3_lut_4_lut.init = 16'h11f0;
    LUT4 mux_196_Mux_2_i142_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n142)) /* synthesis lut_function=(!(A (B)+!A (B (C)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_2_i142_3_lut_4_lut_4_lut_4_lut.init = 16'h3626;
    LUT4 i20460_3_lut_3_lut_4_lut (.A(n26871), .B(index_q[3]), .C(n316), 
         .D(index_q[4]), .Z(n22916)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20460_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 mux_196_Mux_2_i716_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), 
         .B(index_i[2]), .C(index_i[3]), .D(index_i[0]), .Z(n716_adj_2275)) /* synthesis lut_function=(!(A (B)+!A !(B (C+!(D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_2_i716_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h6367;
    PFUMX i20314 (.BLUT(n797), .ALUT(n828), .C0(index_i[5]), .Z(n22770));
    LUT4 i9353_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n11914)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))+!A !(B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9353_3_lut_4_lut_4_lut.init = 16'hb5b3;
    LUT4 i11465_3_lut_4_lut (.A(n26871), .B(index_q[3]), .C(n10079), .D(index_q[6]), 
         .Z(n765)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11465_3_lut_4_lut.init = 16'hffe0;
    LUT4 i9356_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n11917)) /* synthesis lut_function=(A (B+!((D)+!C))+!A (B ((D)+!C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9356_3_lut_4_lut_4_lut.init = 16'hcdad;
    LUT4 mux_197_Mux_10_i317_3_lut_3_lut_4_lut (.A(n26871), .B(index_q[3]), 
         .C(n26796), .D(index_q[4]), .Z(n317)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_10_i317_3_lut_3_lut_4_lut.init = 16'hf011;
    L6MUX21 i20318 (.D0(n22758), .D1(n22759), .SD(index_i[6]), .Z(n22774));
    LUT4 mux_197_Mux_9_i700_3_lut_4_lut (.A(n26871), .B(index_q[3]), .C(index_q[4]), 
         .D(n26859), .Z(n700)) /* synthesis lut_function=(!(A (C+!(D))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_9_i700_3_lut_4_lut.init = 16'h1f10;
    LUT4 n124_bdd_3_lut_24479_4_lut (.A(n26871), .B(index_q[3]), .C(index_q[4]), 
         .D(n93_adj_2274), .Z(n24805)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n124_bdd_3_lut_24479_4_lut.init = 16'hfe0e;
    LUT4 mux_196_Mux_0_i428_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[2]), 
         .B(index_i[0]), .C(index_i[1]), .D(index_i[3]), .Z(n428)) /* synthesis lut_function=(A (B (C+!(D))+!B !((D)+!C))+!A (B (D)+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_0_i428_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hd5a9;
    LUT4 mux_197_Mux_7_i891_3_lut_4_lut (.A(n26871), .B(index_q[3]), .C(index_q[4]), 
         .D(n890_adj_2276), .Z(n891_adj_2277)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_7_i891_3_lut_4_lut.init = 16'hfe0e;
    LUT4 mux_197_Mux_0_i443_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[0]), .D(index_q[3]), .Z(n443)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C (D))+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i443_3_lut_4_lut_4_lut_4_lut.init = 16'h0ed5;
    L6MUX21 i20319 (.D0(n22760), .D1(n22761), .SD(index_i[6]), .Z(n22775));
    LUT4 mux_196_Mux_8_i506_3_lut_4_lut_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[0]), .D(index_i[1]), .Z(n506)) /* synthesis lut_function=(!(A (B+!(C+(D)))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_8_i506_3_lut_4_lut_3_lut_4_lut.init = 16'h6664;
    LUT4 index_i_4__bdd_3_lut_23033_4_lut (.A(n26875), .B(index_i[3]), .C(index_i[5]), 
         .D(index_i[4]), .Z(n24734)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam index_i_4__bdd_3_lut_23033_4_lut.init = 16'hf080;
    L6MUX21 i20320 (.D0(n22762), .D1(n22763), .SD(index_i[6]), .Z(n22776));
    LUT4 mux_196_Mux_8_i860_3_lut_4_lut (.A(n26875), .B(index_i[3]), .C(index_i[4]), 
         .D(n26849), .Z(n860_adj_2278)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_8_i860_3_lut_4_lut.init = 16'h08f8;
    LUT4 mux_196_Mux_0_i46_3_lut_4_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n46)) /* synthesis lut_function=(A (B)+!A ((C+(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_0_i46_3_lut_4_lut_4_lut_4_lut.init = 16'hddd9;
    LUT4 i20441_3_lut_4_lut (.A(n26875), .B(index_i[3]), .C(index_i[4]), 
         .D(n364_adj_2279), .Z(n22897)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20441_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_196_Mux_8_i716_3_lut_4_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n716_adj_2280)) /* synthesis lut_function=(!(A (B)+!A !(B+(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_8_i716_3_lut_4_lut_4_lut_4_lut.init = 16'h7776;
    LUT4 n61_bdd_3_lut_24287_4_lut_3_lut_4_lut (.A(index_q[1]), .B(index_q[3]), 
         .C(index_q[2]), .D(index_q[0]), .Z(n25968)) /* synthesis lut_function=(!(A (B (D)+!B ((D)+!C))+!A !(B (D)+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n61_bdd_3_lut_24287_4_lut_3_lut_4_lut.init = 16'h55a9;
    LUT4 mux_196_Mux_10_i62_3_lut_3_lut_4_lut (.A(n26875), .B(index_i[3]), 
         .C(n26849), .D(index_i[4]), .Z(n62_adj_2281)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_10_i62_3_lut_3_lut_4_lut.init = 16'hf077;
    LUT4 i9389_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[0]), 
         .C(index_q[4]), .D(n27034), .Z(n221)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A !(B+(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9389_3_lut_4_lut_4_lut_4_lut.init = 16'h5556;
    LUT4 mux_196_Mux_6_i955_3_lut_4_lut (.A(n26875), .B(index_i[3]), .C(index_i[4]), 
         .D(n26721), .Z(n955)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_6_i955_3_lut_4_lut.init = 16'h8f80;
    LUT4 n908_bdd_3_lut (.A(n908_adj_2282), .B(n285), .C(index_i[5]), 
         .Z(n25490)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n908_bdd_3_lut.init = 16'hacac;
    PFUMX mux_196_Mux_5_i732 (.BLUT(n12079), .ALUT(n731_adj_2283), .C0(index_i[4]), 
          .Z(n732)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 i9410_3_lut_4_lut_3_lut_4_lut (.A(index_q[1]), .B(index_q[3]), 
         .C(index_q[4]), .D(index_q[0]), .Z(n444)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A !(((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9410_3_lut_4_lut_3_lut_4_lut.init = 16'h5595;
    L6MUX21 i20321 (.D0(n22764), .D1(n22765), .SD(index_i[6]), .Z(n22777));
    LUT4 mux_197_Mux_0_i251_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[0]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n251)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A !(B ((D)+!C)+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i251_3_lut_4_lut_4_lut_4_lut.init = 16'h543c;
    LUT4 mux_196_Mux_3_i252_3_lut_4_lut (.A(n26875), .B(index_i[3]), .C(index_i[4]), 
         .D(n15108), .Z(n252_adj_2284)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_3_i252_3_lut_4_lut.init = 16'h08f8;
    LUT4 mux_197_Mux_4_i812_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[4]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n812_adj_2285)) /* synthesis lut_function=(A (B (C+(D)))+!A !(B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_4_i812_3_lut_3_lut_4_lut.init = 16'h9995;
    LUT4 n25493_bdd_3_lut (.A(n25493), .B(n25492), .C(index_i[5]), .Z(n25494)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n25493_bdd_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_0_i747_3_lut_4_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[2]), 
         .C(index_q[3]), .D(index_q[1]), .Z(n747)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C+(D)))+!A !(B ((D)+!C)+!B (C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i747_3_lut_4_lut_3_lut_4_lut.init = 16'h5596;
    L6MUX21 i20322 (.D0(n22766), .D1(n22767), .SD(index_i[6]), .Z(n22778));
    L6MUX21 i20325 (.D0(n22772), .D1(n22773), .SD(index_i[6]), .Z(n22781));
    LUT4 mux_196_Mux_3_i189_3_lut_3_lut_4_lut (.A(n26875), .B(index_i[3]), 
         .C(index_i[4]), .D(n26842), .Z(n189_adj_2286)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_3_i189_3_lut_3_lut_4_lut.init = 16'h08f8;
    LUT4 i20439_3_lut_3_lut_4_lut (.A(n26876), .B(index_i[3]), .C(n316_adj_2287), 
         .D(index_i[4]), .Z(n22895)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20439_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 mux_196_Mux_10_i317_3_lut_3_lut_4_lut (.A(n26876), .B(index_i[3]), 
         .C(n26842), .D(index_i[4]), .Z(n317_adj_2288)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_10_i317_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 i11392_3_lut_4_lut (.A(n26876), .B(index_i[3]), .C(n9918), .D(index_i[6]), 
         .Z(n765_adj_2289)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11392_3_lut_4_lut.init = 16'hffe0;
    LUT4 n699_bdd_3_lut_24516_4_lut (.A(n26876), .B(index_i[3]), .C(index_i[4]), 
         .D(n93_adj_2290), .Z(n24783)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n699_bdd_3_lut_24516_4_lut.init = 16'hfe0e;
    LUT4 mux_196_Mux_7_i891_3_lut_4_lut (.A(n26876), .B(index_i[3]), .C(index_i[4]), 
         .D(n890_adj_2291), .Z(n891_adj_2292)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_7_i891_3_lut_4_lut.init = 16'hfe0e;
    LUT4 i19240_3_lut_3_lut_4_lut (.A(n26876), .B(index_i[3]), .C(n93_adj_2290), 
         .D(index_i[4]), .Z(n21677)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19240_3_lut_3_lut_4_lut.init = 16'h11f0;
    LUT4 mux_196_Mux_9_i700_3_lut_4_lut (.A(n26876), .B(index_i[3]), .C(index_i[4]), 
         .D(n26835), .Z(n700_adj_2293)) /* synthesis lut_function=(!(A (C+!(D))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_9_i700_3_lut_4_lut.init = 16'h1f10;
    L6MUX21 i20350 (.D0(n22791), .D1(n22792), .SD(index_i[6]), .Z(n22806));
    L6MUX21 i20351 (.D0(n22793), .D1(n22794), .SD(index_i[6]), .Z(n22807));
    LUT4 mux_196_Mux_10_i637_3_lut_4_lut_4_lut (.A(n26877), .B(index_i[4]), 
         .C(index_i[5]), .D(n26775), .Z(n637_adj_2294)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_10_i637_3_lut_4_lut_4_lut.init = 16'h1f1c;
    LUT4 i19648_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n22085)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B (C+!(D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19648_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h1c18;
    LUT4 mux_197_Mux_3_i221_3_lut_4_lut (.A(n26861), .B(index_q[3]), .C(index_q[4]), 
         .D(n26863), .Z(n221_adj_2295)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;
    defparam mux_197_Mux_3_i221_3_lut_4_lut.init = 16'h08f8;
    LUT4 mux_196_Mux_2_i173_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n173)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_2_i173_3_lut_4_lut_4_lut_4_lut.init = 16'h0e1e;
    LUT4 i23643_then_4_lut (.A(index_q[0]), .B(index_q[4]), .C(index_q[1]), 
         .D(index_q[3]), .Z(n27117)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam i23643_then_4_lut.init = 16'h3c69;
    L6MUX21 i20352 (.D0(n22795), .D1(n22796), .SD(index_i[6]), .Z(n22808));
    L6MUX21 i20353 (.D0(n22797), .D1(n22798), .SD(index_i[6]), .Z(n22809));
    LUT4 n45_bdd_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n25707)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n45_bdd_3_lut_4_lut_4_lut_4_lut.init = 16'h1e1c;
    L6MUX21 i20354 (.D0(n22799), .D1(n22800), .SD(index_i[6]), .Z(n22810));
    LUT4 n867_bdd_4_lut (.A(n27088), .B(n939_adj_2296), .C(index_q[4]), 
         .D(index_q[3]), .Z(n24710)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D)))) */ ;
    defparam n867_bdd_4_lut.init = 16'hcacc;
    LUT4 mux_196_Mux_7_i747_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n747_adj_2297)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))+!A (B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_7_i747_3_lut_4_lut_4_lut_4_lut.init = 16'he1e3;
    LUT4 n301_bdd_3_lut_24599_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n25667)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A !((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n301_bdd_3_lut_24599_4_lut_4_lut_4_lut.init = 16'h7173;
    LUT4 i19021_3_lut (.A(n356), .B(n27077), .C(index_q[3]), .Z(n21458)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19021_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_9_i316_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), 
         .B(index_i[2]), .C(index_i[3]), .D(index_i[0]), .Z(n316_adj_2287)) /* synthesis lut_function=(!(A (B (C)+!B !(C+(D)))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_9_i316_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h7e7c;
    LUT4 i20265_3_lut (.A(n22714), .B(n22715), .C(index_q[7]), .Z(n22721)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20265_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_7_i762_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), 
         .B(index_i[2]), .C(index_i[3]), .D(index_i[0]), .Z(n762_adj_2298)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B ((D)+!C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_7_i762_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h3878;
    LUT4 n45_bdd_3_lut_24602_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n25670)) /* synthesis lut_function=(A (B (C)+!B ((D)+!C))+!A (B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n45_bdd_3_lut_24602_4_lut_4_lut_4_lut.init = 16'he7c7;
    PFUMX i20375 (.BLUT(n732_adj_2299), .ALUT(n763_adj_2300), .C0(index_i[5]), 
          .Z(n22831));
    LUT4 i20801_3_lut_4_lut (.A(n26861), .B(index_q[3]), .C(index_q[4]), 
         .D(n220), .Z(n23257)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;
    defparam i20801_3_lut_4_lut.init = 16'hf808;
    LUT4 i19630_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n22067)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B (C+(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19630_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h7c78;
    LUT4 i21539_3_lut (.A(n21457), .B(n21458), .C(index_q[4]), .Z(n21459)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21539_3_lut.init = 16'hcaca;
    LUT4 i19018_3_lut (.A(n27096), .B(n29474), .C(index_q[3]), .Z(n21455)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19018_3_lut.init = 16'hcaca;
    L6MUX21 i20377 (.D0(n22104), .D1(n891_adj_2301), .SD(index_i[5]), 
            .Z(n22833));
    LUT4 mux_196_Mux_0_i443_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .D(index_i[3]), .Z(n443_adj_2302)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C (D))+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_0_i443_3_lut_4_lut_4_lut_4_lut.init = 16'h0ed5;
    LUT4 mux_197_Mux_0_i428_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_q[2]), 
         .B(index_q[0]), .C(index_q[1]), .D(index_q[3]), .Z(n428_adj_2303)) /* synthesis lut_function=(A (B (C+!(D))+!B !((D)+!C))+!A (B (D)+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i428_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hd5a9;
    L6MUX21 i20380 (.D0(n22820), .D1(n22821), .SD(index_i[6]), .Z(n22836));
    LUT4 i9537_3_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[3]), .C(index_i[0]), 
         .D(index_i[1]), .Z(n844_adj_2265)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9537_3_lut_4_lut_4_lut.init = 16'hf00e;
    LUT4 mux_197_Mux_0_i731_3_lut_4_lut (.A(n27085), .B(index_q[2]), .C(index_q[3]), 
         .D(n27102), .Z(n731)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i731_3_lut_4_lut.init = 16'h4f40;
    LUT4 i20796_3_lut_4_lut (.A(n26861), .B(index_q[3]), .C(index_q[4]), 
         .D(n46_adj_2304), .Z(n23252)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam i20796_3_lut_4_lut.init = 16'h8f80;
    LUT4 i9414_3_lut_3_lut_4_lut_4_lut (.A(index_q[2]), .B(index_q[3]), 
         .C(index_q[0]), .D(index_q[1]), .Z(n762_adj_2305)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C (D)+!C !(D)))+!A !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9414_3_lut_3_lut_4_lut_4_lut.init = 16'h700f;
    PFUMX i24734 (.BLUT(n27129), .ALUT(n27130), .C0(index_q[1]), .Z(n27131));
    L6MUX21 i20382 (.D0(n22824), .D1(n22825), .SD(index_i[6]), .Z(n22838));
    PFUMX i18956 (.BLUT(n21391), .ALUT(n21392), .C0(index_q[4]), .Z(n21393));
    L6MUX21 i20383 (.D0(n22826), .D1(n22827), .SD(index_i[6]), .Z(n22839));
    LUT4 i19714_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n22151)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(D))+!A (B (D)+!B ((D)+!C))) */ ;
    defparam i19714_3_lut_4_lut_4_lut.init = 16'hd52b;
    L6MUX21 i20387 (.D0(n22834), .D1(n22835), .SD(index_i[6]), .Z(n22843));
    L6MUX21 i20819 (.D0(n23267), .D1(n23268), .SD(index_q[6]), .Z(n23275));
    L6MUX21 i20822 (.D0(n23273), .D1(n23274), .SD(index_q[6]), .Z(n23278));
    LUT4 mux_197_Mux_0_i604_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n604)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)+!C !(D)))+!A (B (C (D))+!B (C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i604_3_lut_4_lut_4_lut.init = 16'h0e65;
    LUT4 mux_197_Mux_0_i890_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n890)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)+!C !(D)))+!A !(B (C)+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i890_3_lut_4_lut_4_lut.init = 16'h70ca;
    L6MUX21 i20402 (.D0(n23067), .D1(n23074), .SD(index_q[6]), .Z(n22858));
    LUT4 mux_196_Mux_8_i61_3_lut_rep_425_4_lut_4_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[2]), .D(index_i[3]), .Z(n26748)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A (B (C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_8_i61_3_lut_rep_425_4_lut_4_lut_4_lut.init = 16'he0f8;
    PFUMX i18959 (.BLUT(n21394), .ALUT(n21395), .C0(index_q[4]), .Z(n21396));
    LUT4 i20510_3_lut_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n22966)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C+!(D))+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20510_3_lut_3_lut_4_lut_4_lut.init = 16'h1f81;
    LUT4 i20509_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n22965)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20509_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hf81f;
    L6MUX21 i23558 (.D0(n25321), .D1(n25318), .SD(index_i[5]), .Z(n25322));
    LUT4 i19576_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n22013)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C))+!A (B (C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19576_3_lut_4_lut_4_lut_4_lut.init = 16'he078;
    LUT4 mux_196_Mux_8_i251_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n251_adj_2306)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_8_i251_3_lut_4_lut_4_lut_4_lut.init = 16'h07e0;
    PFUMX i23556 (.BLUT(n25320), .ALUT(n25319), .C0(index_i[4]), .Z(n25321));
    L6MUX21 i20405 (.D0(n21732), .D1(n21735), .SD(index_q[6]), .Z(n22861));
    L6MUX21 i20406 (.D0(n21738), .D1(n21741), .SD(index_q[6]), .Z(n22862));
    LUT4 mux_197_Mux_5_i252_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[4]), .Z(n252_adj_2307)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+(D)))+!A (B (C (D))+!B !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_5_i252_3_lut_4_lut.init = 16'hc993;
    LUT4 mux_196_Mux_8_i443_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n443_adj_2308)) /* synthesis lut_function=(A (B (C+!(D))+!B !((D)+!C))+!A !(B (D)+!B ((D)+!C))) */ ;
    defparam mux_196_Mux_8_i443_3_lut_4_lut_4_lut.init = 16'h80fc;
    LUT4 mux_197_Mux_0_i333_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n333)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i333_3_lut_3_lut_4_lut.init = 16'hf10e;
    LUT4 mux_196_Mux_0_i379_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n379)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !((D)+!C))+!A !(B ((D)+!C)+!B (D))) */ ;
    defparam mux_196_Mux_0_i379_3_lut_4_lut_4_lut.init = 16'h8079;
    L6MUX21 i20407 (.D0(n21744), .D1(n21747), .SD(index_q[6]), .Z(n22863));
    LUT4 i20614_3_lut (.A(n29477), .B(n660), .C(index_q[3]), .Z(n23070)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20614_3_lut.init = 16'hcaca;
    LUT4 i19321_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21758)) /* synthesis lut_function=(A (C)+!A !(B (C)+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19321_3_lut_4_lut_4_lut.init = 16'hb4b5;
    LUT4 mux_197_Mux_8_i443_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n443_adj_2309)) /* synthesis lut_function=(A (B (C+!(D))+!B !((D)+!C))+!A !(B (D)+!B ((D)+!C))) */ ;
    defparam mux_197_Mux_8_i443_3_lut_4_lut_4_lut.init = 16'h80fc;
    LUT4 mux_197_Mux_0_i379_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n379_adj_2310)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !((D)+!C))+!A !(B ((D)+!C)+!B (D))) */ ;
    defparam mux_197_Mux_0_i379_3_lut_4_lut_4_lut.init = 16'h8079;
    LUT4 i19338_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n21775)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B+(C+(D))))) */ ;
    defparam i19338_3_lut_4_lut_4_lut_4_lut.init = 16'h2aab;
    LUT4 mux_197_Mux_6_i890_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), 
         .B(index_q[1]), .C(index_q[2]), .D(index_q[3]), .Z(n890_adj_2311)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !((D)+!C))+!A !(B ((D)+!C)+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_6_i890_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h7e07;
    PFUMX i20408 (.BLUT(n21750), .ALUT(n892_adj_2312), .C0(index_q[6]), 
          .Z(n22864));
    LUT4 mux_197_Mux_7_i699_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n699_adj_2313)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C+!(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_7_i699_3_lut_4_lut_4_lut.init = 16'hf07e;
    LUT4 i20599_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n23055)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20599_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hf81f;
    LUT4 mux_197_Mux_0_i460_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n460)) /* synthesis lut_function=(A (B+(C (D)+!C !(D)))+!A (B (C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i460_3_lut_4_lut_4_lut.init = 16'hf8cb;
    LUT4 i20601_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n23057)) /* synthesis lut_function=(A (B (C+!(D))+!B !((D)+!C))+!A !(B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20601_3_lut_4_lut_4_lut.init = 16'h81f8;
    LUT4 mux_197_Mux_6_i859_3_lut_rep_424_4_lut_4_lut_4_lut (.A(index_q[0]), 
         .B(index_q[1]), .C(index_q[2]), .D(index_q[3]), .Z(n26747)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A (B (C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_6_i859_3_lut_rep_424_4_lut_4_lut_4_lut.init = 16'he0f8;
    LUT4 mux_197_Mux_8_i251_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), 
         .B(index_q[1]), .C(index_q[2]), .D(index_q[3]), .Z(n251_adj_2314)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_8_i251_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h07e0;
    LUT4 mux_197_Mux_8_i109_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n109)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C+!(D)))+!A (B (C (D)+!C !(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_8_i109_3_lut_4_lut_4_lut.init = 16'hf83e;
    LUT4 i19003_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n21440)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C))+!A (B (C)+!B !((D)+!C))) */ ;
    defparam i19003_3_lut_4_lut_4_lut_4_lut.init = 16'he078;
    LUT4 i20600_3_lut_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n23056)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C+!(D))+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20600_3_lut_3_lut_4_lut_4_lut.init = 16'h1f81;
    LUT4 mux_197_Mux_8_i15_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n15)) /* synthesis lut_function=(A (B (C)+!B !(C (D)+!C !(D)))+!A !(B ((D)+!C)+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_8_i15_3_lut_4_lut_4_lut.init = 16'h83e0;
    LUT4 mux_197_Mux_0_i412_3_lut_4_lut_4_lut (.A(index_q[2]), .B(index_q[0]), 
         .C(index_q[1]), .D(index_q[3]), .Z(n412)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C (D)))+!A (B (C+!(D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i412_3_lut_4_lut_4_lut.init = 16'hf14c;
    LUT4 i20859_3_lut (.A(n25672), .B(n22970), .C(index_i[6]), .Z(n23315)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20859_3_lut.init = 16'hcaca;
    LUT4 i20447_3_lut_4_lut (.A(n26882), .B(index_i[3]), .C(index_i[4]), 
         .D(n26821), .Z(n22903)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20447_3_lut_4_lut.init = 16'hfe0e;
    LUT4 n21604_bdd_4_lut_24668 (.A(n27034), .B(n763_adj_2315), .C(index_q[5]), 
         .D(index_q[4]), .Z(n24486)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam n21604_bdd_4_lut_24668.init = 16'hcfca;
    LUT4 mux_196_Mux_10_i252_3_lut_4_lut_4_lut (.A(n26882), .B(index_i[3]), 
         .C(index_i[4]), .D(n26836), .Z(n252_adj_2316)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B (C (D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_10_i252_3_lut_4_lut_4_lut.init = 16'h3efe;
    LUT4 mux_196_Mux_0_i604_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n604_adj_2317)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)+!C !(D)))+!A (B (C (D))+!B (C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_0_i604_3_lut_4_lut_4_lut.init = 16'h0e65;
    LUT4 i20511_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n22967)) /* synthesis lut_function=(A (B (C+!(D))+!B !((D)+!C))+!A !(B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;
    defparam i20511_3_lut_4_lut_4_lut_4_lut.init = 16'h81f8;
    LUT4 mux_197_Mux_1_i684_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n684_adj_2318)) /* synthesis lut_function=(A (B ((D)+!C)+!B !((D)+!C))+!A !(B (C+(D))+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_1_i684_3_lut_4_lut_4_lut.init = 16'h992d;
    LUT4 mux_196_Mux_3_i828_3_lut_3_lut_4_lut (.A(n26882), .B(index_i[3]), 
         .C(n157_adj_2319), .D(index_i[4]), .Z(n828)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_3_i828_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 mux_196_Mux_10_i413_3_lut_3_lut_4_lut (.A(n26882), .B(index_i[3]), 
         .C(n26842), .D(index_i[4]), .Z(n413)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_10_i413_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 n24494_bdd_3_lut_26080 (.A(n24494), .B(n24487), .C(index_q[7]), 
         .Z(n24495)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n24494_bdd_3_lut_26080.init = 16'hcaca;
    LUT4 i20445_3_lut_3_lut_4_lut (.A(n26882), .B(index_i[3]), .C(n412_adj_2320), 
         .D(index_i[4]), .Z(n22901)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20445_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 i12468_1_lut_2_lut_3_lut_4_lut (.A(n26882), .B(index_i[3]), .C(index_i[5]), 
         .D(index_i[4]), .Z(n381)) /* synthesis lut_function=(!(A (C+(D))+!A (B (C+(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i12468_1_lut_2_lut_3_lut_4_lut.init = 16'h010f;
    L6MUX21 i20846 (.D0(n23290), .D1(n23291), .SD(index_i[6]), .Z(n23302));
    LUT4 mux_196_Mux_0_i460_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n460_adj_2321)) /* synthesis lut_function=(A (B+(C (D)+!C !(D)))+!A (B (C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_0_i460_3_lut_4_lut_4_lut.init = 16'hf8cb;
    L6MUX21 i20847 (.D0(n23292), .D1(n23293), .SD(index_i[6]), .Z(n23303));
    L6MUX21 i20848 (.D0(n23294), .D1(n23295), .SD(index_i[6]), .Z(n23304));
    LUT4 index_i_5__bdd_4_lut_23861 (.A(n619), .B(index_i[2]), .C(index_i[3]), 
         .D(n26927), .Z(n25578)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (B+!(C (D))))) */ ;
    defparam index_i_5__bdd_4_lut_23861.init = 16'h3a0a;
    LUT4 i20824_3_lut (.A(n23277), .B(n23278), .C(index_q[7]), .Z(n23280)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20824_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_8_i109_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n109_adj_2322)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C+!(D)))+!A (B (C (D)+!C !(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_8_i109_3_lut_4_lut_4_lut.init = 16'hf83e;
    L6MUX21 i22956 (.D0(n24642), .D1(n24640), .SD(index_i[6]), .Z(n24643));
    PFUMX i20849 (.BLUT(n23296), .ALUT(n23297), .C0(index_i[6]), .Z(n23305));
    LUT4 mux_196_Mux_7_i364_3_lut_3_lut (.A(n27001), .B(index_i[3]), .C(n29491), 
         .Z(n364_adj_2323)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;
    defparam mux_196_Mux_7_i364_3_lut_3_lut.init = 16'hd1d1;
    LUT4 i21544_3_lut (.A(n21451), .B(n21452), .C(index_q[4]), .Z(n21453)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21544_3_lut.init = 16'hcaca;
    LUT4 i11916_2_lut (.A(index_q[1]), .B(index_q[3]), .Z(n541_adj_2324)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i11916_2_lut.init = 16'h1111;
    PFUMX i18965 (.BLUT(n21400), .ALUT(n21401), .C0(index_q[4]), .Z(n21402));
    LUT4 mux_197_Mux_0_i526_3_lut (.A(n27080), .B(n29493), .C(index_q[3]), 
         .Z(n526_adj_2325)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i526_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_4_i668_3_lut_3_lut (.A(n27001), .B(index_i[3]), .C(n29497), 
         .Z(n668_adj_2326)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;
    defparam mux_196_Mux_4_i668_3_lut_3_lut.init = 16'hd1d1;
    LUT4 mux_196_Mux_7_i379_3_lut_3_lut (.A(n27001), .B(index_i[3]), .C(n26999), 
         .Z(n379_adj_2327)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam mux_196_Mux_7_i379_3_lut_3_lut.init = 16'h7474;
    L6MUX21 i20860 (.D0(n21669), .D1(n21672), .SD(index_i[6]), .Z(n23316));
    L6MUX21 i20861 (.D0(n574_adj_2328), .D1(n21675), .SD(index_i[6]), 
            .Z(n23317));
    LUT4 i20219_3_lut (.A(n22668), .B(n22669), .C(index_i[7]), .Z(n22675)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20219_3_lut.init = 16'hcaca;
    LUT4 i20218_3_lut (.A(n22666), .B(n22667), .C(index_i[7]), .Z(n22674)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20218_3_lut.init = 16'hcaca;
    LUT4 i19558_3_lut_3_lut (.A(n27001), .B(index_i[3]), .C(n38), .Z(n21995)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam i19558_3_lut_3_lut.init = 16'h7474;
    LUT4 mux_196_Mux_5_i252_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[4]), .Z(n252_adj_2329)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+(D)))+!A (B (C (D))+!B !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_5_i252_3_lut_4_lut.init = 16'hc993;
    LUT4 i20547_3_lut_3_lut (.A(n27001), .B(index_i[3]), .C(n29497), .Z(n23003)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam i20547_3_lut_3_lut.init = 16'h7474;
    LUT4 mux_196_Mux_1_i716_3_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[1]), .D(index_i[3]), .Z(n716_adj_2330)) /* synthesis lut_function=(!(A (B (D)+!B !(C))+!A !(B (C (D))+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_1_i716_3_lut_4_lut_4_lut.init = 16'h70a9;
    LUT4 mux_196_Mux_1_i684_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n684_adj_2331)) /* synthesis lut_function=(A (B ((D)+!C)+!B !((D)+!C))+!A !(B (C+(D))+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_1_i684_3_lut_4_lut_4_lut.init = 16'h992d;
    LUT4 mux_196_Mux_11_i445_3_lut_4_lut_4_lut_4_lut (.A(index_i[3]), .B(index_i[4]), 
         .C(index_i[5]), .D(n26882), .Z(n445)) /* synthesis lut_function=(!(A (B (C))+!A !(B+(C+(D))))) */ ;
    defparam mux_196_Mux_11_i445_3_lut_4_lut_4_lut_4_lut.init = 16'h7f7e;
    LUT4 n348_bdd_3_lut_24656 (.A(n26983), .B(n27028), .C(index_i[3]), 
         .Z(n25580)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n348_bdd_3_lut_24656.init = 16'hcaca;
    LUT4 mux_197_Mux_1_i716_3_lut_4_lut_4_lut (.A(index_q[2]), .B(index_q[0]), 
         .C(index_q[1]), .D(index_q[3]), .Z(n716_adj_2332)) /* synthesis lut_function=(!(A (B (D)+!B !(C))+!A !(B (C (D))+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_1_i716_3_lut_4_lut_4_lut.init = 16'h70a9;
    LUT4 i19498_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21935)) /* synthesis lut_function=(A (C)+!A !(B (C)+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19498_3_lut_4_lut_4_lut.init = 16'hb4b5;
    L6MUX21 i20862 (.D0(n21678), .D1(n764_adj_2333), .SD(index_i[6]), 
            .Z(n23318));
    LUT4 mux_197_Mux_11_i445_3_lut_4_lut_4_lut_4_lut (.A(index_q[3]), .B(index_q[4]), 
         .C(index_q[5]), .D(n26854), .Z(n445_adj_2334)) /* synthesis lut_function=(!(A (B (C))+!A !(B+(C+(D))))) */ ;
    defparam mux_197_Mux_11_i445_3_lut_4_lut_4_lut_4_lut.init = 16'h7f7e;
    LUT4 mux_196_Mux_0_i412_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n412_adj_2335)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(D))+!A (B (D)+!B !(C+!(D)))) */ ;
    defparam mux_196_Mux_0_i412_3_lut_4_lut_4_lut.init = 16'hcd2a;
    LUT4 n442_bdd_3_lut_23804 (.A(n27024), .B(n29497), .C(index_i[3]), 
         .Z(n25584)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n442_bdd_3_lut_23804.init = 16'hcaca;
    LUT4 i19665_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n22102)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B+(C+(D))))) */ ;
    defparam i19665_3_lut_4_lut_4_lut_4_lut.init = 16'h2aab;
    LUT4 mux_196_Mux_7_i699_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n699_adj_2336)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C+!(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_7_i699_3_lut_4_lut_4_lut.init = 16'hf07e;
    LUT4 n300_bdd_3_lut (.A(n26983), .B(n773), .C(index_i[3]), .Z(n25586)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n300_bdd_3_lut.init = 16'hacac;
    LUT4 mux_196_Mux_0_i890_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n890_adj_2337)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)+!C !(D)))+!A !(B (C)+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_0_i890_3_lut_4_lut_4_lut.init = 16'h70ca;
    LUT4 mux_196_Mux_0_i684_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n684_adj_2338)) /* synthesis lut_function=(!(A ((D)+!B)+!A !(B (D)+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_0_i684_3_lut_4_lut_4_lut_4_lut.init = 16'h5498;
    PFUMX i24779 (.BLUT(n27200), .ALUT(n27201), .C0(index_q[8]), .Z(n27202));
    LUT4 n518_bdd_3_lut_23817 (.A(n27028), .B(n27022), .C(index_i[3]), 
         .Z(n25602)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n518_bdd_3_lut_23817.init = 16'hcaca;
    L6MUX21 i20444 (.D0(n22898), .D1(n22899), .SD(index_i[6]), .Z(n382_adj_2271));
    LUT4 i20823_3_lut (.A(n23275), .B(n23276), .C(index_q[7]), .Z(n23279)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20823_3_lut.init = 16'hcaca;
    L6MUX21 i20451 (.D0(n22905), .D1(n22906), .SD(index_i[6]), .Z(n509_adj_2272));
    LUT4 i22679_2_lut (.A(index_i[5]), .B(index_i[4]), .Z(n22372)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i22679_2_lut.init = 16'heeee;
    LUT4 mux_197_Mux_6_i955_3_lut_4_lut (.A(n26893), .B(index_q[3]), .C(index_q[4]), 
         .D(n26720), .Z(n955_adj_2339)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_6_i955_3_lut_4_lut.init = 16'h8f80;
    LUT4 i20207_3_lut (.A(n22659), .B(n22660), .C(index_i[8]), .Z(n22663)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20207_3_lut.init = 16'hcaca;
    PFUMX i22954 (.BLUT(n924), .ALUT(n24641), .C0(index_i[5]), .Z(n24642));
    PFUMX i20876 (.BLUT(n23328), .ALUT(n23329), .C0(index_i[6]), .Z(n23332));
    LUT4 n92_bdd_3_lut_23897 (.A(n27001), .B(n26986), .C(index_i[3]), 
         .Z(n25611)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n92_bdd_3_lut_23897.init = 16'hcaca;
    LUT4 n17993_bdd_4_lut_else_4_lut (.A(index_q[3]), .B(index_q[4]), .C(index_q[1]), 
         .D(index_q[2]), .Z(n27143)) /* synthesis lut_function=(!(A (B (D)+!B ((D)+!C))+!A !(B+!((D)+!C)))) */ ;
    defparam n17993_bdd_4_lut_else_4_lut.init = 16'h44fc;
    LUT4 i22509_3_lut (.A(n24495), .B(n22854), .C(index_q[8]), .Z(n22856)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22509_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_8_i542_3_lut_4_lut (.A(n27048), .B(index_i[3]), .C(index_i[4]), 
         .D(n526_adj_2340), .Z(n542)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_8_i542_3_lut_4_lut.init = 16'h6f60;
    LUT4 i19237_3_lut_4_lut (.A(n27048), .B(index_i[3]), .C(index_i[4]), 
         .D(n635_adj_2341), .Z(n21674)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19237_3_lut_4_lut.init = 16'hf606;
    LUT4 index_i_4__bdd_4_lut_23130 (.A(index_i[4]), .B(n26864), .C(index_i[7]), 
         .D(n26835), .Z(n24731)) /* synthesis lut_function=(A (C+!(D))+!A (B+!(C))) */ ;
    defparam index_i_4__bdd_4_lut_23130.init = 16'he5ef;
    LUT4 n26998_bdd_2_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[4]), .Z(n28252)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C (D)))+!A (B+!(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n26998_bdd_2_lut_4_lut.init = 16'h3800;
    LUT4 i19285_3_lut_4_lut (.A(n27063), .B(index_q[3]), .C(index_q[4]), 
         .D(n635_adj_2342), .Z(n21722)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19285_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_197_Mux_8_i542_3_lut_4_lut (.A(n27063), .B(index_q[3]), .C(index_q[4]), 
         .D(n526_adj_2343), .Z(n542_adj_2344)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_8_i542_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_196_Mux_1_i700_3_lut_4_lut (.A(n26909), .B(index_i[3]), .C(index_i[4]), 
         .D(n684_adj_2331), .Z(n700_adj_2345)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_1_i700_3_lut_4_lut.init = 16'hefe0;
    LUT4 i11375_3_lut_4_lut (.A(n26714), .B(index_i[7]), .C(index_i[8]), 
         .D(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2126[14])) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11375_3_lut_4_lut.init = 16'hffe0;
    LUT4 i19663_3_lut_4_lut (.A(n26996), .B(index_i[2]), .C(index_i[3]), 
         .D(n27027), .Z(n22100)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19663_3_lut_4_lut.init = 16'hf404;
    LUT4 i12193_2_lut (.A(index_i[1]), .B(index_i[3]), .Z(n541_adj_2346)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i12193_2_lut.init = 16'h1111;
    LUT4 mux_196_Mux_0_i526_3_lut (.A(n29489), .B(n27025), .C(index_i[3]), 
         .Z(n526_adj_2347)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_0_i526_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_0_i731_3_lut_4_lut (.A(n26996), .B(index_i[2]), .C(index_i[3]), 
         .D(n29491), .Z(n731_adj_2348)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_0_i731_3_lut_4_lut.init = 16'h4f40;
    LUT4 n389_bdd_3_lut_23850 (.A(n27107), .B(n29485), .C(index_q[3]), 
         .Z(n25634)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n389_bdd_3_lut_23850.init = 16'hcaca;
    LUT4 i20613_3_lut (.A(n652), .B(n27104), .C(index_q[3]), .Z(n23069)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20613_3_lut.init = 16'hcaca;
    LUT4 i19636_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n22073)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(D))+!A (B (D)+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19636_3_lut_4_lut_4_lut_4_lut.init = 16'hd52b;
    LUT4 i19633_3_lut_4_lut (.A(index_i[0]), .B(n27048), .C(index_i[3]), 
         .D(n27031), .Z(n22070)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19633_3_lut_4_lut.init = 16'hfb0b;
    LUT4 mux_197_Mux_3_i109_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n109_adj_2349)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (D)+!B !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_3_i109_3_lut_4_lut_4_lut.init = 16'hcf10;
    PFUMX i20877 (.BLUT(n23330), .ALUT(n23331), .C0(index_i[6]), .Z(n23333));
    LUT4 mux_196_Mux_14_i511_4_lut_4_lut (.A(n26714), .B(index_i[7]), .C(index_i[8]), 
         .D(n254_adj_2350), .Z(n511)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (B (C+!(D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_14_i511_4_lut_4_lut.init = 16'h1c10;
    LUT4 i11466_4_lut (.A(n15088), .B(index_q[8]), .C(n765), .D(index_q[7]), 
         .Z(n1022)) /* synthesis lut_function=(A (B+(C (D)))+!A (B+(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11466_4_lut.init = 16'hfcdd;
    LUT4 i12060_3_lut_3_lut_rep_812 (.A(index_q[2]), .B(index_q[0]), .C(index_q[1]), 
         .Z(n29485)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12060_3_lut_3_lut_rep_812.init = 16'hd0d0;
    LUT4 i19015_3_lut_4_lut_4_lut (.A(index_q[2]), .B(index_q[0]), .C(index_q[1]), 
         .D(index_q[3]), .Z(n21452)) /* synthesis lut_function=(A (B (C)+!B !(C+!(D)))+!A (B (C)+!B !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19015_3_lut_4_lut_4_lut.init = 16'hc3d0;
    LUT4 index_q_4__bdd_4_lut_23209 (.A(index_q[4]), .B(n26863), .C(index_q[7]), 
         .D(n26859), .Z(n24748)) /* synthesis lut_function=(A (C+!(D))+!A (B+!(C))) */ ;
    defparam index_q_4__bdd_4_lut_23209.init = 16'he5ef;
    LUT4 index_i_1__bdd_4_lut (.A(index_i[1]), .B(index_i[3]), .C(index_i[2]), 
         .D(index_i[0]), .Z(n29500)) /* synthesis lut_function=(!(A (B (C (D))+!B (C+!(D)))+!A !(B (C (D)+!C !(D))+!B ((D)+!C)))) */ ;
    defparam index_i_1__bdd_4_lut.init = 16'h5b8d;
    L6MUX21 i20465 (.D0(n22919), .D1(n22920), .SD(index_q[6]), .Z(n382));
    LUT4 mux_197_Mux_1_i348_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n348)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A (B ((D)+!C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_1_i348_3_lut_4_lut_4_lut_4_lut.init = 16'h38f0;
    LUT4 mux_196_Mux_4_i389_3_lut_3_lut_3_lut_rep_814 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29487)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_4_i389_3_lut_3_lut_3_lut_rep_814.init = 16'h9393;
    LUT4 i19618_3_lut_4_lut (.A(index_i[0]), .B(index_i[2]), .C(index_i[1]), 
         .D(index_i[3]), .Z(n22055)) /* synthesis lut_function=(A (B+(D))+!A !(B (C+(D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19618_3_lut_4_lut.init = 16'haa9d;
    LUT4 i1_3_lut (.A(index_i[0]), .B(index_i[4]), .C(index_i[2]), .Z(n20693)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i1_3_lut.init = 16'hfefe;
    PFUMX i22952 (.BLUT(n24639), .ALUT(n26860), .C0(index_i[5]), .Z(n24640));
    LUT4 i19521_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21958)) /* synthesis lut_function=(A (B (C (D))+!B !(C (D)))+!A !(B (D)+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19521_3_lut_4_lut_4_lut.init = 16'h9366;
    LUT4 mux_196_Mux_4_i262_3_lut_3_lut_rep_815 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29488)) /* synthesis lut_function=(A (B+(C))+!A !(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_4_i262_3_lut_3_lut_rep_815.init = 16'ha9a9;
    LUT4 mux_196_Mux_0_i762_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n762_adj_2351)) /* synthesis lut_function=(A (B+!((D)+!C))+!A !(B (D)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_0_i762_3_lut_4_lut_4_lut.init = 16'h98fc;
    LUT4 i19590_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n22027)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A !(B (D)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19590_3_lut_3_lut_4_lut.init = 16'ha955;
    LUT4 mux_196_Mux_6_i389_3_lut_4_lut_4_lut_3_lut_rep_816 (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[2]), .Z(n29489)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_6_i389_3_lut_4_lut_4_lut_3_lut_rep_816.init = 16'h9292;
    LUT4 mux_197_Mux_2_i189_3_lut_3_lut_4_lut (.A(index_q[1]), .B(n27034), 
         .C(n173_adj_2352), .D(index_q[4]), .Z(n189_adj_2353)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(C+(D)))) */ ;
    defparam mux_197_Mux_2_i189_3_lut_3_lut_4_lut.init = 16'h77f0;
    LUT4 i11481_2_lut_3_lut_4_lut (.A(index_q[1]), .B(n27034), .C(index_q[5]), 
         .D(index_q[4]), .Z(n508)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;
    defparam i11481_2_lut_3_lut_4_lut.init = 16'hf080;
    LUT4 mux_196_Mux_3_i668_3_lut_4_lut (.A(n26987), .B(index_i[2]), .C(index_i[3]), 
         .D(n29489), .Z(n668_adj_2354)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_3_i668_3_lut_4_lut.init = 16'h6f60;
    LUT4 n53_bdd_3_lut_23552_4_lut (.A(n26987), .B(index_i[2]), .C(n27031), 
         .D(index_i[3]), .Z(n25316)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n53_bdd_3_lut_23552_4_lut.init = 16'hf066;
    LUT4 mux_196_Mux_4_i763_3_lut_4_lut (.A(n26987), .B(index_i[2]), .C(index_i[4]), 
         .D(n747_adj_2355), .Z(n763_adj_2356)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_4_i763_3_lut_4_lut.init = 16'h6f60;
    LUT4 i21847_3_lut (.A(n109), .B(n124), .C(index_q[4]), .Z(n21707)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21847_3_lut.init = 16'hcaca;
    LUT4 i19009_3_lut (.A(n29473), .B(n27072), .C(index_q[3]), .Z(n21446)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19009_3_lut.init = 16'hcaca;
    LUT4 i19008_3_lut (.A(n29494), .B(n27098), .C(index_q[3]), .Z(n21445)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19008_3_lut.init = 16'hcaca;
    LUT4 i21550_3_lut (.A(n21445), .B(n21446), .C(index_q[4]), .Z(n21447)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21550_3_lut.init = 16'hcaca;
    L6MUX21 i20472 (.D0(n22926), .D1(n22927), .SD(index_q[6]), .Z(n509));
    LUT4 i11393_4_lut (.A(n15064), .B(index_i[8]), .C(n765_adj_2289), 
         .D(index_i[7]), .Z(n1022_adj_2357)) /* synthesis lut_function=(A (B+(C (D)))+!A (B+(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11393_4_lut.init = 16'hfcdd;
    LUT4 i19006_3_lut (.A(n29485), .B(n27106), .C(index_q[3]), .Z(n21443)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19006_3_lut.init = 16'hcaca;
    LUT4 i12159_1_lut_rep_409_2_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n26732)) /* synthesis lut_function=(!(A (C+(D))+!A (B (C+(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12159_1_lut_rep_409_2_lut_3_lut_4_lut.init = 16'h010f;
    LUT4 i19002_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n21439)) /* synthesis lut_function=(!(A (B (D)+!B !(D))+!A (B ((D)+!C)+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19002_3_lut_4_lut_4_lut_4_lut.init = 16'h33c8;
    LUT4 i19005_3_lut (.A(n27104), .B(n652), .C(index_q[3]), .Z(n21442)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19005_3_lut.init = 16'hcaca;
    LUT4 i21557_3_lut (.A(n21442), .B(n21443), .C(index_q[4]), .Z(n21444)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21557_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_2_i908_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[1]), .D(index_i[3]), .Z(n908_adj_2358)) /* synthesis lut_function=(!(A (B (C)+!B !(C (D)))+!A (B (C)+!B !(C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_2_i908_3_lut_4_lut_4_lut.init = 16'h3c0d;
    LUT4 i21859_3_lut (.A(n620_adj_2250), .B(n14171), .C(index_i[4]), 
         .Z(n21692)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21859_3_lut.init = 16'hcaca;
    LUT4 i20606_3_lut_3_lut (.A(n27104), .B(index_q[3]), .C(n29485), .Z(n23062)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam i20606_3_lut_3_lut.init = 16'h7474;
    LUT4 i21869_3_lut (.A(n491), .B(n506_adj_2359), .C(index_i[4]), .Z(n21686)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21869_3_lut.init = 16'hcaca;
    PFUMX i23553 (.BLUT(n25317), .ALUT(n25316), .C0(index_i[4]), .Z(n25318));
    LUT4 i22709_2_lut_rep_588 (.A(index_q[4]), .B(index_q[3]), .Z(n26911)) /* synthesis lut_function=((B)+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i22709_2_lut_rep_588.init = 16'hdddd;
    LUT4 mux_196_Mux_0_i812_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n812_adj_2360)) /* synthesis lut_function=(A (B (C+(D))+!B !(C))+!A (B (D)+!B !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_0_i812_3_lut_4_lut_4_lut_4_lut.init = 16'hcf92;
    LUT4 mux_196_Mux_7_i45_3_lut_3_lut_3_lut_rep_817 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29490)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_7_i45_3_lut_3_lut_3_lut_rep_817.init = 16'h3939;
    LUT4 mux_196_Mux_2_i604_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n604_adj_2361)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)+!C !(D)))+!A (B (D)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_2_i604_3_lut_4_lut_4_lut_4_lut.init = 16'h39cf;
    PFUMX i24730 (.BLUT(n27123), .ALUT(n27124), .C0(index_i[0]), .Z(n27125));
    LUT4 mux_197_Mux_7_i364_3_lut_3_lut (.A(n27104), .B(index_q[3]), .C(n27102), 
         .Z(n364_adj_2362)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;
    defparam mux_197_Mux_7_i364_3_lut_3_lut.init = 16'hd1d1;
    LUT4 i21899_3_lut (.A(n109_adj_2322), .B(n124_adj_2363), .C(index_i[4]), 
         .Z(n21659)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21899_3_lut.init = 16'hcaca;
    LUT4 i18997_3_lut (.A(n29474), .B(n356), .C(index_q[3]), .Z(n21434)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18997_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_0_i475_3_lut_4_lut (.A(n26913), .B(index_q[1]), .C(index_q[3]), 
         .D(n26861), .Z(n475_adj_2364)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i475_3_lut_4_lut.init = 16'h4f40;
    LUT4 i21585_3_lut (.A(n21433), .B(n21434), .C(index_q[4]), .Z(n21435)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21585_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_3_i491_3_lut_4_lut (.A(n26913), .B(index_q[1]), .C(index_q[3]), 
         .D(n27081), .Z(n491_adj_2365)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_3_i491_3_lut_4_lut.init = 16'h4f40;
    LUT4 i9526_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[4]), .D(n27035), .Z(n189_adj_2366)) /* synthesis lut_function=(A (B (C (D)))+!A !(B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9526_3_lut_4_lut_4_lut_4_lut.init = 16'h9555;
    LUT4 mux_196_Mux_7_i340_3_lut_rep_818 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29491)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B (C)+!B !(C)))) */ ;
    defparam mux_196_Mux_7_i340_3_lut_rep_818.init = 16'h1c1c;
    LUT4 i19585_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n22022)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B (C (D)+!C !(D))))) */ ;
    defparam i19585_3_lut_3_lut_4_lut.init = 16'h0f1c;
    LUT4 i19101_3_lut (.A(n24753), .B(n21576), .C(index_q[8]), .Z(n21538)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19101_3_lut.init = 16'hcaca;
    LUT4 i18985_3_lut_3_lut (.A(n27104), .B(index_q[3]), .C(n1001), .Z(n21422)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam i18985_3_lut_3_lut.init = 16'h7474;
    LUT4 i7422_2_lut (.A(index_i[4]), .B(index_i[5]), .Z(n9918)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i7422_2_lut.init = 16'h8888;
    LUT4 i1_2_lut (.A(index_i[6]), .B(index_i[7]), .Z(n19801)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i1_2_lut.init = 16'heeee;
    PFUMX i23510 (.BLUT(n25270), .ALUT(n26974), .C0(index_q[5]), .Z(n25271));
    LUT4 mux_196_Mux_8_i116_3_lut_rep_819 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29492)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B !(C))) */ ;
    defparam mux_196_Mux_8_i116_3_lut_rep_819.init = 16'hc1c1;
    LUT4 mux_197_Mux_4_i747_3_lut_4_lut (.A(n27071), .B(index_q[2]), .C(index_q[3]), 
         .D(n29474), .Z(n747_adj_2367)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_4_i747_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_196_Mux_5_i505_3_lut_3_lut_rep_797 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29470)) /* synthesis lut_function=(A (B+(C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_5_i505_3_lut_3_lut_rep_797.init = 16'hadad;
    LUT4 mux_196_Mux_0_i796_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n796_adj_2368)) /* synthesis lut_function=(A (B (C+(D))+!B (C (D)))+!A !(B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_0_i796_3_lut_4_lut_4_lut.init = 16'hadc0;
    LUT4 i9391_3_lut_4_lut (.A(n27071), .B(index_q[2]), .C(n27044), .D(n27079), 
         .Z(n444_adj_2369)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9391_3_lut_4_lut.init = 16'h6f60;
    PFUMX i23508 (.BLUT(n26918), .ALUT(n25268), .C0(index_q[2]), .Z(n25269));
    LUT4 i19095_3_lut (.A(n24736), .B(n21567), .C(index_i[8]), .Z(n21532)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19095_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_0_i397_3_lut (.A(n27086), .B(n29474), .C(index_q[3]), 
         .Z(n397_adj_2370)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i397_3_lut.init = 16'hcaca;
    LUT4 i7583_2_lut (.A(index_q[4]), .B(index_q[5]), .Z(n10079)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i7583_2_lut.init = 16'h8888;
    LUT4 mux_197_Mux_6_i251_3_lut_4_lut (.A(n27071), .B(index_q[2]), .C(index_q[3]), 
         .D(n27079), .Z(n251_adj_2371)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_6_i251_3_lut_4_lut.init = 16'hf606;
    LUT4 n45_bdd_3_lut_23885_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n25669)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C (D)+!C !(D))+!B (C)))) */ ;
    defparam n45_bdd_3_lut_23885_3_lut_4_lut.init = 16'h0fc1;
    LUT4 i23643_else_4_lut (.A(index_q[0]), .B(index_q[4]), .C(index_q[1]), 
         .D(index_q[3]), .Z(n27116)) /* synthesis lut_function=(!(A (B (C)+!B !(C (D)+!C !(D)))+!A (B ((D)+!C)+!B !((D)+!C)))) */ ;
    defparam i23643_else_4_lut.init = 16'h394b;
    LUT4 i1_2_lut_adj_82 (.A(index_q[6]), .B(index_q[7]), .Z(n19798)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_2_lut_adj_82.init = 16'heeee;
    PFUMX i24777 (.BLUT(n27197), .ALUT(n27198), .C0(index_i[8]), .Z(n27199));
    LUT4 i20122_3_lut (.A(n22573), .B(n24712), .C(index_q[7]), .Z(n22578)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20122_3_lut.init = 16'hcaca;
    LUT4 i20121_3_lut (.A(n22571), .B(n22572), .C(index_q[7]), .Z(n22577)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20121_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_3_i797_3_lut_4_lut (.A(index_q[4]), .B(index_q[3]), 
         .C(n796_adj_2372), .D(n27088), .Z(n797_adj_2373)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_3_i797_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i22522_3_lut (.A(n22577), .B(n22578), .C(index_q[8]), .Z(n22580)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22522_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_0_i525_3_lut_3_lut_rep_820 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29493)) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i525_3_lut_3_lut_rep_820.init = 16'h6a6a;
    LUT4 i20224_3_lut (.A(n22678), .B(n22679), .C(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2126[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20224_3_lut.init = 16'hcaca;
    LUT4 i19713_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n22150)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (D))+!A !(B (C (D))+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19713_3_lut_3_lut_4_lut.init = 16'h4933;
    LUT4 i20856_3_lut (.A(n23310), .B(n23311), .C(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2126[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20856_3_lut.init = 16'hcaca;
    LUT4 i20855_3_lut (.A(n23308), .B(n23309), .C(index_i[8]), .Z(n23311)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20855_3_lut.init = 16'hcaca;
    LUT4 i6430_2_lut (.A(phase_q[0]), .B(phase_i[10]), .Z(index_i_9__N_2106[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i6430_2_lut.init = 16'h6666;
    LUT4 i22538_2_lut (.A(phase_q[0]), .B(phase_i[10]), .Z(index_q_9__N_2116[0])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i22538_2_lut.init = 16'h9999;
    LUT4 quarter_wave_sample_register_i_15__I_0_3_lut (.A(\quarter_wave_sample_register_q[15] ), 
         .B(o_val_pipeline_i_0__15__N_2157[15]), .C(phase_negation_i[1]), 
         .Z(o_val_pipeline_i_0__15__N_2156)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[14] 77[8])
    defparam quarter_wave_sample_register_i_15__I_0_3_lut.init = 16'hcaca;
    LUT4 quarter_wave_sample_register_i_14__I_0_3_lut (.A(quarter_wave_sample_register_i[14]), 
         .B(o_val_pipeline_i_0__15__N_2157[14]), .C(phase_negation_i[1]), 
         .Z(o_val_pipeline_i_0__15__N_2158)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[14] 77[8])
    defparam quarter_wave_sample_register_i_14__I_0_3_lut.init = 16'hcaca;
    LUT4 quarter_wave_sample_register_i_13__I_0_3_lut (.A(quarter_wave_sample_register_i[13]), 
         .B(o_val_pipeline_i_0__15__N_2157[13]), .C(phase_negation_i[1]), 
         .Z(o_val_pipeline_i_0__15__N_2160)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[14] 77[8])
    defparam quarter_wave_sample_register_i_13__I_0_3_lut.init = 16'hcaca;
    LUT4 quarter_wave_sample_register_i_12__I_0_3_lut (.A(quarter_wave_sample_register_i[12]), 
         .B(o_val_pipeline_i_0__15__N_2157[12]), .C(phase_negation_i[1]), 
         .Z(o_val_pipeline_i_0__15__N_2162)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[14] 77[8])
    defparam quarter_wave_sample_register_i_12__I_0_3_lut.init = 16'hcaca;
    LUT4 quarter_wave_sample_register_i_11__I_0_3_lut (.A(quarter_wave_sample_register_i[11]), 
         .B(o_val_pipeline_i_0__15__N_2157[11]), .C(phase_negation_i[1]), 
         .Z(o_val_pipeline_i_0__15__N_2164)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[14] 77[8])
    defparam quarter_wave_sample_register_i_11__I_0_3_lut.init = 16'hcaca;
    LUT4 i12177_3_lut (.A(index_i[2]), .B(index_i[1]), .C(index_i[0]), 
         .Z(n38)) /* synthesis lut_function=(A (B)+!A (B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i12177_3_lut.init = 16'hdcdc;
    LUT4 mux_197_Mux_2_i491_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n491_adj_2374)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A !(B (C)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_2_i491_3_lut_4_lut_4_lut.init = 16'h6a5a;
    LUT4 mux_197_Mux_0_i963_3_lut_3_lut_rep_821 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29494)) /* synthesis lut_function=(!(A (B)+!A (B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i963_3_lut_3_lut_rep_821.init = 16'h3636;
    LUT4 i20612_3_lut (.A(n26887), .B(n27078), .C(index_q[3]), .Z(n23068)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20612_3_lut.init = 16'hcaca;
    LUT4 quarter_wave_sample_register_i_10__I_0_3_lut (.A(quarter_wave_sample_register_i[10]), 
         .B(o_val_pipeline_i_0__15__N_2157[10]), .C(phase_negation_i[1]), 
         .Z(o_val_pipeline_i_0__15__N_2166)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[14] 77[8])
    defparam quarter_wave_sample_register_i_10__I_0_3_lut.init = 16'hcaca;
    LUT4 quarter_wave_sample_register_i_9__I_0_3_lut (.A(quarter_wave_sample_register_i[9]), 
         .B(o_val_pipeline_i_0__15__N_2157[9]), .C(phase_negation_i[1]), 
         .Z(o_val_pipeline_i_0__15__N_2168)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[14] 77[8])
    defparam quarter_wave_sample_register_i_9__I_0_3_lut.init = 16'hcaca;
    L6MUX21 i20532 (.D0(n22973), .D1(n22974), .SD(index_q[6]), .Z(n22988));
    L6MUX21 i20533 (.D0(n22975), .D1(n22976), .SD(index_q[6]), .Z(n22989));
    LUT4 mux_197_Mux_4_i668_3_lut_3_lut (.A(n27104), .B(index_q[3]), .C(n29485), 
         .Z(n668_adj_2375)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;
    defparam mux_197_Mux_4_i668_3_lut_3_lut.init = 16'hd1d1;
    LUT4 mux_197_Mux_0_i188_3_lut (.A(n27105), .B(n931), .C(index_q[3]), 
         .Z(n188)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i188_3_lut.init = 16'hcaca;
    LUT4 quarter_wave_sample_register_i_8__I_0_3_lut (.A(quarter_wave_sample_register_i[8]), 
         .B(o_val_pipeline_i_0__15__N_2157[8]), .C(phase_negation_i[1]), 
         .Z(o_val_pipeline_i_0__15__N_2170)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[14] 77[8])
    defparam quarter_wave_sample_register_i_8__I_0_3_lut.init = 16'hcaca;
    LUT4 quarter_wave_sample_register_i_7__I_0_3_lut (.A(quarter_wave_sample_register_i[7]), 
         .B(o_val_pipeline_i_0__15__N_2157[7]), .C(phase_negation_i[1]), 
         .Z(o_val_pipeline_i_0__15__N_2172)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(75[14] 77[8])
    defparam quarter_wave_sample_register_i_7__I_0_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_5_i890_3_lut_3_lut (.A(n27104), .B(index_q[3]), .C(n27086), 
         .Z(n890_adj_2376)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam mux_197_Mux_5_i890_3_lut_3_lut.init = 16'h7474;
    LUT4 mux_197_Mux_6_i475_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n475_adj_2377)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A !(B (C+(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_6_i475_3_lut_4_lut_4_lut.init = 16'h9936;
    LUT4 index_i_4__bdd_4_lut_25482 (.A(index_i[4]), .B(n26775), .C(n24619), 
         .D(index_i[5]), .Z(n26700)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (B (C (D))+!B (C+!(D)))) */ ;
    defparam index_i_4__bdd_4_lut_25482.init = 16'hf099;
    LUT4 i21919_3_lut (.A(n26417), .B(n124_adj_2378), .C(index_q[4]), 
         .Z(n23254)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21919_3_lut.init = 16'hcaca;
    L6MUX21 i20534 (.D0(n22977), .D1(n22978), .SD(index_q[6]), .Z(n22990));
    LUT4 mux_196_Mux_6_i435_3_lut_4_lut_4_lut_3_lut_rep_798 (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[2]), .Z(n29471)) /* synthesis lut_function=(A (B+!(C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_6_i435_3_lut_4_lut_4_lut_3_lut_rep_798.init = 16'hdbdb;
    LUT4 mux_197_Mux_0_i978_3_lut_3_lut_rep_822 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29495)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i978_3_lut_3_lut_rep_822.init = 16'h6c6c;
    LUT4 mux_197_Mux_0_i124_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n124_adj_2378)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A !(B (D)+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i124_3_lut_4_lut_4_lut.init = 16'h6c99;
    L6MUX21 i20535 (.D0(n22979), .D1(n22980), .SD(index_q[6]), .Z(n22991));
    LUT4 i9596_3_lut_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n12161)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A !(B (C+(D))+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9596_3_lut_3_lut_4_lut_4_lut.init = 16'h44db;
    L6MUX21 i20536 (.D0(n22981), .D1(n22982), .SD(index_q[6]), .Z(n22992));
    LUT4 index_q_5__bdd_4_lut_24347 (.A(n652), .B(index_q[2]), .C(index_q[3]), 
         .D(n27101), .Z(n25802)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (B+!(C (D))))) */ ;
    defparam index_q_5__bdd_4_lut_24347.init = 16'h3a0a;
    LUT4 n812_bdd_3_lut_24495 (.A(n27066), .B(n29494), .C(index_q[3]), 
         .Z(n25804)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n812_bdd_3_lut_24495.init = 16'hcaca;
    LUT4 i19528_3_lut_4_lut (.A(n26982), .B(index_i[2]), .C(index_i[3]), 
         .D(n27032), .Z(n21965)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19528_3_lut_4_lut.init = 16'h6f60;
    L6MUX21 i20972 (.D0(n23420), .D1(n23421), .SD(index_q[6]), .Z(n23428));
    LUT4 mux_196_Mux_3_i460_3_lut_4_lut (.A(n26982), .B(index_i[2]), .C(index_i[3]), 
         .D(n27025), .Z(n460_adj_2379)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_3_i460_3_lut_4_lut.init = 16'h6f60;
    LUT4 i19624_3_lut_4_lut (.A(n26982), .B(index_i[2]), .C(index_i[3]), 
         .D(n26993), .Z(n22061)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19624_3_lut_4_lut.init = 16'hf606;
    LUT4 n442_bdd_3_lut_24017 (.A(n27099), .B(n29485), .C(index_q[3]), 
         .Z(n25813)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n442_bdd_3_lut_24017.init = 16'hcaca;
    L6MUX21 i20973 (.D0(n23422), .D1(n23423), .SD(index_q[6]), .Z(n23429));
    LUT4 mux_196_Mux_6_i285_3_lut_4_lut (.A(n26982), .B(index_i[2]), .C(index_i[3]), 
         .D(n27022), .Z(n285_adj_2380)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_6_i285_3_lut_4_lut.init = 16'hf606;
    L6MUX21 i20974 (.D0(n23424), .D1(n23425), .SD(index_q[6]), .Z(n23430));
    LUT4 i11492_3_lut_3_lut_3_lut_rep_799 (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[1]), .Z(n29472)) /* synthesis lut_function=(!(A ((C)+!B)+!A (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11492_3_lut_3_lut_3_lut_rep_799.init = 16'h0d0d;
    LUT4 n627_bdd_3_lut_24559 (.A(n27066), .B(n588), .C(index_q[3]), .Z(n25815)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n627_bdd_3_lut_24559.init = 16'hacac;
    LUT4 i12179_3_lut_rep_824 (.A(index_i[2]), .B(index_i[1]), .C(index_i[0]), 
         .Z(n29497)) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i12179_3_lut_rep_824.init = 16'hc4c4;
    LUT4 i19653_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[2]), .C(index_i[1]), 
         .D(index_i[3]), .Z(n22090)) /* synthesis lut_function=(!(A ((C (D)+!C !(D))+!B)+!A (B (C (D)+!C !(D))+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19653_3_lut_4_lut_4_lut.init = 16'h0dc0;
    LUT4 mux_197_Mux_6_i420_3_lut_4_lut_3_lut_rep_800 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29473)) /* synthesis lut_function=(A (B+!(C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_6_i420_3_lut_4_lut_3_lut_rep_800.init = 16'hdbdb;
    LUT4 i9500_3_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[1]), .C(index_i[0]), 
         .D(n26995), .Z(n605)) /* synthesis lut_function=(A (B (C)+!B !(C+!(D)))+!A (B (C+!(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9500_3_lut_4_lut_4_lut.init = 16'hc3c4;
    LUT4 mux_197_Mux_9_i62_3_lut_4_lut_then_4_lut (.A(index_q[4]), .B(index_q[2]), 
         .C(index_q[1]), .D(index_q[0]), .Z(n27120)) /* synthesis lut_function=(!(A (B (C+(D)))+!A (B+(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_9_i62_3_lut_4_lut_then_4_lut.init = 16'h222b;
    L6MUX21 i20975 (.D0(n23426), .D1(n23427), .SD(index_q[6]), .Z(n23431));
    LUT4 i19588_3_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[1]), .C(index_i[0]), 
         .D(index_i[3]), .Z(n22025)) /* synthesis lut_function=(A (B (C)+!B !(C+!(D)))+!A (B (C+!(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19588_3_lut_4_lut_4_lut.init = 16'hc3c4;
    LUT4 mux_196_Mux_0_i475_3_lut_4_lut (.A(n26923), .B(index_i[1]), .C(index_i[3]), 
         .D(n26836), .Z(n475_adj_2381)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_0_i475_3_lut_4_lut.init = 16'h4f40;
    LUT4 mux_196_Mux_3_i491_3_lut_4_lut (.A(n26923), .B(index_i[1]), .C(index_i[3]), 
         .D(n29487), .Z(n491_adj_2382)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_3_i491_3_lut_4_lut.init = 16'h4f40;
    LUT4 mux_196_Mux_2_i684_3_lut_4_lut (.A(index_i[2]), .B(n26927), .C(index_i[3]), 
         .D(n29472), .Z(n684_adj_2383)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;
    defparam mux_196_Mux_2_i684_3_lut_4_lut.init = 16'h6f60;
    LUT4 i19513_3_lut_4_lut (.A(index_i[2]), .B(n26927), .C(index_i[3]), 
         .D(n29468), .Z(n21950)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;
    defparam i19513_3_lut_4_lut.init = 16'h6f60;
    LUT4 i19254_4_lut_4_lut_4_lut (.A(index_i[2]), .B(n26927), .C(index_i[4]), 
         .D(index_i[3]), .Z(n21691)) /* synthesis lut_function=(A (B+!(C+(D)))+!A !(B+!(C+(D)))) */ ;
    defparam i19254_4_lut_4_lut_4_lut.init = 16'h999a;
    LUT4 mux_196_Mux_7_i475_3_lut_4_lut (.A(index_i[2]), .B(n26927), .C(index_i[3]), 
         .D(n26999), .Z(n475_adj_2384)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+(D)))) */ ;
    defparam mux_196_Mux_7_i475_3_lut_4_lut.init = 16'h9f90;
    LUT4 mux_196_Mux_7_i653_3_lut_4_lut (.A(index_i[2]), .B(n26927), .C(index_i[3]), 
         .D(n70), .Z(n653_adj_2385)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam mux_196_Mux_7_i653_3_lut_4_lut.init = 16'hf606;
    L6MUX21 i20857 (.D0(n21657), .D1(n21660), .SD(index_i[6]), .Z(n23313));
    LUT4 i19252_3_lut_3_lut_4_lut_4_lut (.A(index_i[2]), .B(n26927), .C(index_i[3]), 
         .D(index_i[4]), .Z(n21689)) /* synthesis lut_function=(A (B+(C (D)))+!A !(B+(C (D)))) */ ;
    defparam i19252_3_lut_3_lut_4_lut_4_lut.init = 16'ha999;
    LUT4 i20416_3_lut (.A(n22870), .B(n22871), .C(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_2141[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20416_3_lut.init = 16'hcaca;
    LUT4 i20042_3_lut (.A(n26356), .B(n22497), .C(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_2141[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20042_3_lut.init = 16'hcaca;
    LUT4 i20041_3_lut (.A(n22494), .B(n22495), .C(index_q[8]), .Z(n22497)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20041_3_lut.init = 16'hcaca;
    LUT4 i22540_2_lut (.A(phase_i[9]), .B(phase_i[10]), .Z(index_q_9__N_2116[9])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i22540_2_lut.init = 16'h9999;
    LUT4 i22542_2_lut (.A(phase_i[8]), .B(phase_i[10]), .Z(index_q_9__N_2116[8])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i22542_2_lut.init = 16'h9999;
    L6MUX21 i20032 (.D0(n22476), .D1(n22477), .SD(index_q[6]), .Z(n22488));
    L6MUX21 i20033 (.D0(n22478), .D1(n22479), .SD(index_q[6]), .Z(n22489));
    LUT4 i22544_2_lut (.A(phase_i[7]), .B(phase_i[10]), .Z(index_q_9__N_2116[7])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i22544_2_lut.init = 16'h9999;
    L6MUX21 i20034 (.D0(n22480), .D1(n22481), .SD(index_q[6]), .Z(n22490));
    LUT4 i22546_2_lut (.A(phase_i[6]), .B(phase_i[10]), .Z(index_q_9__N_2116[6])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i22546_2_lut.init = 16'h9999;
    PFUMX i20035 (.BLUT(n22482), .ALUT(n22483), .C0(index_q[6]), .Z(n22491));
    LUT4 i22548_2_lut (.A(phase_i[5]), .B(phase_i[10]), .Z(index_q_9__N_2116[5])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i22548_2_lut.init = 16'h9999;
    LUT4 i22550_2_lut (.A(phase_i[4]), .B(phase_i[10]), .Z(index_q_9__N_2116[4])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i22550_2_lut.init = 16'h9999;
    LUT4 i22552_2_lut (.A(phase_i[3]), .B(phase_i[10]), .Z(index_q_9__N_2116[3])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i22552_2_lut.init = 16'h9999;
    LUT4 i22554_2_lut (.A(phase_i[2]), .B(phase_i[10]), .Z(index_q_9__N_2116[2])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i22554_2_lut.init = 16'h9999;
    LUT4 i22556_2_lut (.A(phase_i[1]), .B(phase_i[10]), .Z(index_q_9__N_2116[1])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i22556_2_lut.init = 16'h9999;
    LUT4 i6442_2_lut (.A(phase_i[9]), .B(phase_i[10]), .Z(index_i_9__N_2106[9])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i6442_2_lut.init = 16'h6666;
    LUT4 i6443_2_lut (.A(phase_i[8]), .B(phase_i[10]), .Z(index_i_9__N_2106[8])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i6443_2_lut.init = 16'h6666;
    LUT4 i6444_2_lut (.A(phase_i[7]), .B(phase_i[10]), .Z(index_i_9__N_2106[7])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i6444_2_lut.init = 16'h6666;
    LUT4 i6445_2_lut (.A(phase_i[6]), .B(phase_i[10]), .Z(index_i_9__N_2106[6])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i6445_2_lut.init = 16'h6666;
    LUT4 i6446_2_lut (.A(phase_i[5]), .B(phase_i[10]), .Z(index_i_9__N_2106[5])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i6446_2_lut.init = 16'h6666;
    LUT4 i6447_2_lut (.A(phase_i[4]), .B(phase_i[10]), .Z(index_i_9__N_2106[4])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i6447_2_lut.init = 16'h6666;
    LUT4 i6448_2_lut (.A(phase_i[3]), .B(phase_i[10]), .Z(index_i_9__N_2106[3])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i6448_2_lut.init = 16'h6666;
    LUT4 i6449_2_lut (.A(phase_i[2]), .B(phase_i[10]), .Z(index_i_9__N_2106[2])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i6449_2_lut.init = 16'h6666;
    LUT4 i6450_2_lut (.A(phase_i[1]), .B(phase_i[10]), .Z(index_i_9__N_2106[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(59[14] 62[8])
    defparam i6450_2_lut.init = 16'h6666;
    LUT4 i20544_3_lut (.A(n22997), .B(n22998), .C(index_q[8]), .Z(n23000)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20544_3_lut.init = 16'hcaca;
    LUT4 i20543_3_lut (.A(n22995), .B(n22996), .C(index_q[8]), .Z(n22999)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20543_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_2_i573_3_lut_3_lut_4_lut (.A(n27046), .B(index_i[3]), 
         .C(n557_adj_2258), .D(index_i[4]), .Z(n573)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_2_i573_3_lut_3_lut_4_lut.init = 16'h11f0;
    LUT4 i20438_3_lut_4_lut (.A(n27046), .B(index_i[3]), .C(index_i[4]), 
         .D(n285_adj_2386), .Z(n22894)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20438_3_lut_4_lut.init = 16'hfe0e;
    LUT4 mux_196_Mux_4_i573_3_lut_3_lut_4_lut_4_lut (.A(n27046), .B(index_i[3]), 
         .C(index_i[4]), .D(n26882), .Z(n573_adj_2387)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_4_i573_3_lut_3_lut_4_lut_4_lut.init = 16'h1f1c;
    LUT4 mux_197_Mux_9_i62_3_lut_4_lut_else_4_lut (.A(index_q[4]), .B(index_q[2]), 
         .C(index_q[1]), .D(index_q[0]), .Z(n27119)) /* synthesis lut_function=((B+(C (D)))+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_9_i62_3_lut_4_lut_else_4_lut.init = 16'hfddd;
    LUT4 mux_417_i9_3_lut (.A(\quarter_wave_sample_register_q[15] ), .B(o_val_pipeline_q_0__15__N_2189[15]), 
         .C(phase_negation_q[1]), .Z(n1829[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(80[29:60])
    defparam mux_417_i9_3_lut.init = 16'hcaca;
    LUT4 i19731_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n22168)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A (B (C)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19731_3_lut_4_lut_4_lut.init = 16'h3c8c;
    LUT4 n699_bdd_3_lut_23071_4_lut (.A(n27046), .B(index_i[3]), .C(index_i[4]), 
         .D(n124_adj_2388), .Z(n24782)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n699_bdd_3_lut_23071_4_lut.init = 16'hf101;
    LUT4 mux_417_i8_3_lut (.A(quarter_wave_sample_register_q[14]), .B(o_val_pipeline_q_0__15__N_2189[14]), 
         .C(phase_negation_q[1]), .Z(n1829[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(80[29:60])
    defparam mux_417_i8_3_lut.init = 16'hcaca;
    LUT4 mux_417_i7_3_lut (.A(quarter_wave_sample_register_q[13]), .B(o_val_pipeline_q_0__15__N_2189[13]), 
         .C(phase_negation_q[1]), .Z(n1829[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(80[29:60])
    defparam mux_417_i7_3_lut.init = 16'hcaca;
    LUT4 i22506_3_lut (.A(n23321), .B(n23322), .C(index_i[8]), .Z(n23325)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22506_3_lut.init = 16'hcaca;
    LUT4 mux_417_i6_3_lut (.A(quarter_wave_sample_register_q[12]), .B(o_val_pipeline_q_0__15__N_2189[12]), 
         .C(phase_negation_q[1]), .Z(n1829[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(80[29:60])
    defparam mux_417_i6_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_3_i444_3_lut_4_lut (.A(index_i[0]), .B(index_i[3]), 
         .C(n27046), .D(index_i[4]), .Z(n444_adj_2389)) /* synthesis lut_function=(!(A (B (D)+!B (C (D)))+!A !(B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_3_i444_3_lut_4_lut.init = 16'h46aa;
    LUT4 mux_417_i5_3_lut (.A(quarter_wave_sample_register_q[11]), .B(o_val_pipeline_q_0__15__N_2189[11]), 
         .C(phase_negation_q[1]), .Z(n1829[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(80[29:60])
    defparam mux_417_i5_3_lut.init = 16'hcaca;
    LUT4 mux_417_i4_3_lut (.A(quarter_wave_sample_register_q[10]), .B(o_val_pipeline_q_0__15__N_2189[10]), 
         .C(phase_negation_q[1]), .Z(n1829[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(80[29:60])
    defparam mux_417_i4_3_lut.init = 16'hcaca;
    PFUMX i20637 (.BLUT(n732_adj_2390), .ALUT(n763_adj_2391), .C0(index_q[5]), 
          .Z(n23093));
    LUT4 mux_417_i3_3_lut (.A(quarter_wave_sample_register_q[9]), .B(o_val_pipeline_q_0__15__N_2189[9]), 
         .C(phase_negation_q[1]), .Z(n1829[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(80[29:60])
    defparam mux_417_i3_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_3_i573_3_lut_3_lut_4_lut (.A(n27046), .B(index_i[3]), 
         .C(n397_adj_2392), .D(index_i[4]), .Z(n573_adj_2393)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_3_i573_3_lut_3_lut_4_lut.init = 16'h11f0;
    LUT4 mux_196_Mux_10_i125_3_lut_4_lut_4_lut (.A(n27046), .B(index_i[3]), 
         .C(index_i[4]), .D(n26836), .Z(n125)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B (C (D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_10_i125_3_lut_4_lut_4_lut.init = 16'h3efe;
    LUT4 mux_417_i2_3_lut (.A(quarter_wave_sample_register_q[8]), .B(o_val_pipeline_q_0__15__N_2189[8]), 
         .C(phase_negation_q[1]), .Z(n1829[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(80[29:60])
    defparam mux_417_i2_3_lut.init = 16'hcaca;
    LUT4 i20399_3_lut (.A(n22851), .B(n22852), .C(index_q[8]), .Z(n22855)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20399_3_lut.init = 16'hcaca;
    LUT4 mux_417_i1_3_lut (.A(quarter_wave_sample_register_q[7]), .B(o_val_pipeline_q_0__15__N_2189[7]), 
         .C(phase_negation_q[1]), .Z(n1829[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(80[29:60])
    defparam mux_417_i1_3_lut.init = 16'hcaca;
    L6MUX21 i23480 (.D0(n25237), .D1(n25234), .SD(index_q[5]), .Z(n25238));
    LUT4 n476_bdd_3_lut_23174 (.A(n476), .B(n24864), .C(index_i[5]), .Z(n24865)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n476_bdd_3_lut_23174.init = 16'hcaca;
    LUT4 i9584_3_lut_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n12149)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A !(B (C+(D))+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9584_3_lut_3_lut_4_lut_4_lut.init = 16'h44db;
    PFUMX i20602 (.BLUT(n23054), .ALUT(n23055), .C0(index_q[4]), .Z(n23058));
    L6MUX21 i20639 (.D0(n21777), .D1(n891_adj_2394), .SD(index_q[5]), 
            .Z(n23095));
    LUT4 mux_196_Mux_4_i158_3_lut (.A(n142_adj_2395), .B(n157_adj_2396), 
         .C(index_i[4]), .Z(n158)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_4_i158_3_lut.init = 16'hcaca;
    LUT4 i20362_3_lut (.A(n22815), .B(n22816), .C(index_i[8]), .Z(n22818)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20362_3_lut.init = 16'hcaca;
    L6MUX21 i20642 (.D0(n23082), .D1(n23083), .SD(index_q[6]), .Z(n23098));
    LUT4 i20361_3_lut (.A(n22813), .B(n22814), .C(index_i[8]), .Z(n22817)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20361_3_lut.init = 16'hcaca;
    L6MUX21 i20644 (.D0(n23086), .D1(n23087), .SD(index_q[6]), .Z(n23100));
    PFUMX i23478 (.BLUT(n25236), .ALUT(n475_adj_2377), .C0(index_q[4]), 
          .Z(n25237));
    LUT4 mux_197_Mux_0_i396_3_lut_4_lut_3_lut_rep_801 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29474)) /* synthesis lut_function=(A ((C)+!B)+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i396_3_lut_4_lut_3_lut_rep_801.init = 16'hb6b6;
    PFUMX i20603 (.BLUT(n23056), .ALUT(n23057), .C0(index_q[4]), .Z(n23059));
    LUT4 i22514_3_lut (.A(n22720), .B(n22721), .C(index_q[8]), .Z(n22724)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22514_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_83 (.A(o_phase[11]), .B(o_phase[10]), .Z(phase_q_11__N_2232[11])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i1_2_lut_adj_83.init = 16'h9999;
    LUT4 i20252_3_lut (.A(n22703), .B(n24643), .C(index_i[7]), .Z(n22708)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20252_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_1_i93_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[1]), .D(index_i[3]), .Z(n93_adj_2397)) /* synthesis lut_function=(A (B (C (D))+!B !(D))+!A !(B (C (D))+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_1_i93_3_lut_4_lut_4_lut.init = 16'h9566;
    LUT4 i20251_3_lut (.A(n22701), .B(n22702), .C(index_i[7]), .Z(n22707)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20251_3_lut.init = 16'hcaca;
    LUT4 i22536_3_lut (.A(n22707), .B(n22708), .C(index_i[8]), .Z(n22710)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22536_3_lut.init = 16'hcaca;
    LUT4 i20201_3_lut (.A(n22654), .B(n22655), .C(index_q[8]), .Z(n22657)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20201_3_lut.init = 16'hcaca;
    L6MUX21 i20645 (.D0(n23088), .D1(n23089), .SD(index_q[6]), .Z(n23101));
    LUT4 i19729_3_lut (.A(n29475), .B(n27079), .C(index_q[3]), .Z(n22166)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19729_3_lut.init = 16'hcaca;
    LUT4 i20200_3_lut (.A(n22652), .B(n22653), .C(index_q[8]), .Z(n22656)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20200_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_3_i573_3_lut_3_lut_4_lut (.A(n27090), .B(index_q[3]), 
         .C(n397), .D(index_q[4]), .Z(n573_adj_2398)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_3_i573_3_lut_3_lut_4_lut.init = 16'h11f0;
    LUT4 i20459_3_lut_4_lut (.A(n27090), .B(index_q[3]), .C(index_q[4]), 
         .D(n285_adj_2399), .Z(n22915)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20459_3_lut_4_lut.init = 16'hfe0e;
    L6MUX21 i20649 (.D0(n23096), .D1(n23097), .SD(index_q[6]), .Z(n23105));
    PFUMX i20609 (.BLUT(n23061), .ALUT(n23062), .C0(index_q[4]), .Z(n23065));
    LUT4 i19719_3_lut (.A(n29493), .B(n29473), .C(index_q[3]), .Z(n22156)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19719_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_10_i125_3_lut_4_lut_4_lut (.A(n27090), .B(index_q[3]), 
         .C(index_q[4]), .D(n26861), .Z(n125_adj_2400)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B (C (D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_10_i125_3_lut_4_lut_4_lut.init = 16'h3efe;
    LUT4 i22520_3_lut (.A(n574_adj_2401), .B(n637), .C(index_q[6]), .Z(n21577)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22520_3_lut.init = 16'hcaca;
    LUT4 n124_bdd_3_lut_23087_4_lut (.A(n27090), .B(index_q[3]), .C(index_q[4]), 
         .D(n124_adj_2402), .Z(n24804)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n124_bdd_3_lut_23087_4_lut.init = 16'hf101;
    LUT4 i20123_3_lut (.A(n22575), .B(n22576), .C(index_q[8]), .Z(n22579)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20123_3_lut.init = 16'hcaca;
    LUT4 i22524_3_lut (.A(n574_adj_2403), .B(n637_adj_2294), .C(index_i[6]), 
         .Z(n21568)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22524_3_lut.init = 16'hcaca;
    LUT4 i21690_3_lut (.A(n22150), .B(n22151), .C(index_q[4]), .Z(n22152)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21690_3_lut.init = 16'hcaca;
    LUT4 i20655_3_lut (.A(n23108), .B(n23109), .C(index_q[8]), .Z(n23111)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20655_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_2_i573_3_lut_3_lut_4_lut (.A(n27090), .B(index_q[3]), 
         .C(n557_adj_2404), .D(index_q[4]), .Z(n573_adj_2405)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_2_i573_3_lut_3_lut_4_lut.init = 16'h11f0;
    PFUMX i20610 (.BLUT(n23063), .ALUT(n23064), .C0(index_q[4]), .Z(n23066));
    LUT4 i20654_3_lut (.A(n23106), .B(n23107), .C(index_q[8]), .Z(n23110)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20654_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_4_i573_3_lut_3_lut_4_lut_4_lut (.A(n27090), .B(index_q[3]), 
         .C(index_q[4]), .D(n26854), .Z(n573_adj_2406)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_4_i573_3_lut_3_lut_4_lut_4_lut.init = 16'h1f1c;
    LUT4 mux_197_Mux_9_i763_3_lut_4_lut (.A(n27085), .B(n26994), .C(index_q[4]), 
         .D(n26856), .Z(n763_adj_2315)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;
    defparam mux_197_Mux_9_i763_3_lut_4_lut.init = 16'hf101;
    LUT4 mux_197_Mux_8_i763_3_lut_4_lut (.A(n27085), .B(n26994), .C(index_q[4]), 
         .D(n26856), .Z(n15132)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam mux_197_Mux_8_i763_3_lut_4_lut.init = 16'hfe0e;
    LUT4 i20264_3_lut (.A(n22712), .B(n22713), .C(index_q[7]), .Z(n22720)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20264_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_0_i173_3_lut_4_lut (.A(n26937), .B(index_i[1]), .C(index_i[3]), 
         .D(n29489), .Z(n173_adj_2407)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_0_i173_3_lut_4_lut.init = 16'hdfd0;
    LUT4 i19519_3_lut_4_lut (.A(n26937), .B(index_i[1]), .C(index_i[3]), 
         .D(n404), .Z(n21956)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19519_3_lut_4_lut.init = 16'hdfd0;
    LUT4 i18989_then_4_lut (.A(index_q[0]), .B(index_q[4]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n27160)) /* synthesis lut_function=(A (B (C)+!B (C (D)+!C !(D)))+!A !(B (C+!(D))+!B !(C+!(D)))) */ ;
    defparam i18989_then_4_lut.init = 16'hb493;
    LUT4 mux_196_Mux_1_i620_3_lut_4_lut (.A(n26937), .B(index_i[1]), .C(index_i[3]), 
         .D(n29488), .Z(n620)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_1_i620_3_lut_4_lut.init = 16'hdfd0;
    CCU2D add_377_15 (.A0(quarter_wave_sample_register_q[14]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(\quarter_wave_sample_register_q[15] ), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17577), .S0(o_val_pipeline_q_0__15__N_2189[14]), 
          .S1(o_val_pipeline_q_0__15__N_2189[15]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(80[29:60])
    defparam add_377_15.INIT0 = 16'hf555;
    defparam add_377_15.INIT1 = 16'hf555;
    defparam add_377_15.INJECT1_0 = "NO";
    defparam add_377_15.INJECT1_1 = "NO";
    LUT4 i20393_3_lut (.A(n22846), .B(n22847), .C(index_i[8]), .Z(n22849)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20393_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_1_i317_3_lut (.A(n301), .B(n908_adj_2408), .C(index_q[4]), 
         .Z(n317_adj_2409)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_1_i317_3_lut.init = 16'hcaca;
    L6MUX21 i20111 (.D0(n22551), .D1(n22552), .SD(index_q[6]), .Z(n22567));
    LUT4 i20392_3_lut (.A(n22844), .B(n22845), .C(index_i[8]), .Z(n22848)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20392_3_lut.init = 16'hcaca;
    L6MUX21 i20112 (.D0(n22553), .D1(n22554), .SD(index_q[6]), .Z(n22568));
    L6MUX21 i20113 (.D0(n22555), .D1(n22556), .SD(index_q[6]), .Z(n22569));
    LUT4 i20331_3_lut (.A(n22784), .B(n22785), .C(index_i[8]), .Z(n22787)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20331_3_lut.init = 16'hcaca;
    CCU2D add_377_13 (.A0(quarter_wave_sample_register_q[12]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_q[13]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17576), .COUT(n17577), 
          .S0(o_val_pipeline_q_0__15__N_2189[12]), .S1(o_val_pipeline_q_0__15__N_2189[13]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(80[29:60])
    defparam add_377_13.INIT0 = 16'hf555;
    defparam add_377_13.INIT1 = 16'hf555;
    defparam add_377_13.INJECT1_0 = "NO";
    defparam add_377_13.INJECT1_1 = "NO";
    L6MUX21 i20114 (.D0(n22557), .D1(n22558), .SD(index_q[6]), .Z(n22570));
    LUT4 mux_196_Mux_0_i397_3_lut (.A(n26999), .B(n27032), .C(index_i[3]), 
         .Z(n397_adj_2410)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_0_i397_3_lut.init = 16'hcaca;
    L6MUX21 i20115 (.D0(n22559), .D1(n22560), .SD(index_q[6]), .Z(n22571));
    L6MUX21 i20117 (.D0(n22563), .D1(n22564), .SD(index_q[6]), .Z(n22573));
    LUT4 i20330_3_lut (.A(n22782), .B(n22783), .C(index_i[8]), .Z(n22786)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20330_3_lut.init = 16'hcaca;
    LUT4 i20253_3_lut (.A(n22705), .B(n22706), .C(index_i[8]), .Z(n22709)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20253_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_0_i285_3_lut (.A(n27000), .B(n29497), .C(index_i[3]), 
         .Z(n285)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_0_i285_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_2_i716_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), 
         .B(index_q[1]), .C(index_q[3]), .D(index_q[2]), .Z(n716_adj_2411)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)+!C !(D)))+!A (B (D)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_2_i716_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h31cf;
    PFUMX i20616 (.BLUT(n23068), .ALUT(n23069), .C0(index_q[4]), .Z(n23072));
    LUT4 index_i_2__bdd_4_lut_25983 (.A(index_i[2]), .B(index_i[0]), .C(index_i[4]), 
         .D(index_i[1]), .Z(n28248)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((C (D))+!B))) */ ;
    defparam index_i_2__bdd_4_lut_25983.init = 16'h0cec;
    LUT4 index_i_2__bdd_3_lut_26320 (.A(index_i[2]), .B(index_i[0]), .C(index_i[4]), 
         .Z(n28249)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B (C)+!B !(C)))) */ ;
    defparam index_i_2__bdd_3_lut_26320.init = 16'h6969;
    LUT4 mux_197_Mux_2_i142_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n142_adj_2412)) /* synthesis lut_function=(!(A (B (D)+!B (C (D)+!C !(D)))+!A (B (D)+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_2_i142_3_lut_4_lut_4_lut_4_lut.init = 16'h03ec;
    PFUMX i9489 (.BLUT(n12157), .ALUT(n12158), .C0(n22374), .Z(n12050));
    LUT4 n26998_bdd_3_lut_25753 (.A(n26836), .B(n29487), .C(index_i[4]), 
         .Z(n28251)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n26998_bdd_3_lut_25753.init = 16'hcaca;
    PFUMX i20617 (.BLUT(n23070), .ALUT(n23071), .C0(index_q[4]), .Z(n23073));
    LUT4 mux_197_Mux_0_i15_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n15_adj_2413)) /* synthesis lut_function=(A (B (D)+!B (C+!(D)))+!A (B (D)+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i15_3_lut_4_lut_4_lut_4_lut.init = 16'hec33;
    LUT4 mux_196_Mux_9_i763_3_lut_4_lut (.A(n26996), .B(n26898), .C(index_i[4]), 
         .D(n26849), .Z(n763_adj_2414)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;
    defparam mux_196_Mux_9_i763_3_lut_4_lut.init = 16'hf101;
    LUT4 i19732_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n22169)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)+!C !(D)))+!A (B (C+!(D))+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19732_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h0e30;
    LUT4 mux_197_Mux_0_i723_3_lut_rep_779 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n27102)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i723_3_lut_rep_779.init = 16'h1c1c;
    LUT4 mux_196_Mux_8_i763_3_lut_4_lut (.A(n26996), .B(n26898), .C(index_i[4]), 
         .D(n26849), .Z(n15106)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam mux_196_Mux_8_i763_3_lut_4_lut.init = 16'hfe0e;
    LUT4 mux_197_Mux_5_i53_3_lut_4_lut_3_lut_rep_780 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n27103)) /* synthesis lut_function=(A ((C)+!B)+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_5_i53_3_lut_4_lut_3_lut_rep_780.init = 16'he6e6;
    PFUMX i20623 (.BLUT(n23075), .ALUT(n23076), .C0(index_q[4]), .Z(n23079));
    LUT4 mux_197_Mux_6_i691_3_lut_rep_781 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n27104)) /* synthesis lut_function=(A (B+!(C))+!A !((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_6_i691_3_lut_rep_781.init = 16'h8e8e;
    LUT4 index_i_1__bdd_4_lut_25685 (.A(index_i[1]), .B(index_i[3]), .C(index_i[2]), 
         .D(index_i[0]), .Z(n28269)) /* synthesis lut_function=(A (B (C+(D))+!B (C (D)))+!A !(B (D)+!B !(C+(D)))) */ ;
    defparam index_i_1__bdd_4_lut_25685.init = 16'hb9d4;
    LUT4 n28269_bdd_3_lut (.A(n28269), .B(index_i[1]), .C(index_i[4]), 
         .Z(n28270)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n28269_bdd_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_0_i180_3_lut_4_lut_3_lut_rep_782 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n27105)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i180_3_lut_4_lut_3_lut_rep_782.init = 16'h1818;
    LUT4 mux_197_Mux_5_i70_3_lut_4_lut_3_lut_rep_783 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n27106)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_5_i70_3_lut_4_lut_3_lut_rep_783.init = 16'h1919;
    LUT4 mux_197_Mux_0_i277_3_lut_rep_784 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n27107)) /* synthesis lut_function=(!(A (B (C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i277_3_lut_rep_784.init = 16'h7e7e;
    PFUMX i19137 (.BLUT(n318), .ALUT(n381_adj_2415), .C0(index_q[6]), 
          .Z(n21574));
    PFUMX i20624 (.BLUT(n23077), .ALUT(n23078), .C0(index_q[4]), .Z(n23080));
    LUT4 mux_197_Mux_7_i716_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n716_adj_2416)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C+!(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_7_i716_3_lut_3_lut_4_lut.init = 16'h0f81;
    LUT4 n11074_bdd_3_lut_23934_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n25733)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A (B (C (D)+!C !(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n11074_bdd_3_lut_23934_3_lut_4_lut.init = 16'h0fc1;
    LUT4 mux_197_Mux_4_i526_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n526_adj_2417)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A !(B ((D)+!C)+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_4_i526_3_lut_3_lut_4_lut.init = 16'h7e0f;
    PFUMX i23475 (.BLUT(n25233), .ALUT(n21914), .C0(index_q[4]), .Z(n25234));
    LUT4 i19545_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21982)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(D))+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19545_3_lut_3_lut_4_lut.init = 16'h3319;
    LUT4 i19702_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n22139)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A (B (D)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19702_3_lut_4_lut.init = 16'h18cc;
    PFUMX i19128 (.BLUT(n318_adj_2418), .ALUT(n381), .C0(index_i[6]), 
          .Z(n21565));
    LUT4 mux_197_Mux_2_i557_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n557_adj_2404)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C+!(D))+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_2_i557_3_lut_3_lut_4_lut.init = 16'h0f18;
    LUT4 i19011_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21448)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)))+!A !(B (C+!(D))+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19011_3_lut_3_lut_4_lut.init = 16'h71cc;
    LUT4 mux_197_Mux_6_i635_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n635_adj_2419)) /* synthesis lut_function=(A (B (C+(D))+!B !(D))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_6_i635_3_lut_4_lut.init = 16'hcce6;
    LUT4 i19012_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21449)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19012_3_lut_3_lut_4_lut.init = 16'h0f1c;
    LUT4 i19335_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21772)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C (D)))+!A (B (C+(D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19335_4_lut_4_lut_4_lut.init = 16'h301c;
    LUT4 mux_197_Mux_0_i699_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n699)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (D))+!A (B (C+!(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i699_3_lut_3_lut_4_lut.init = 16'h1c33;
    LUT4 mux_197_Mux_0_i557_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n557)) /* synthesis lut_function=(A ((D)+!C)+!A !((D)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i557_3_lut_4_lut.init = 16'haa4e;
    L6MUX21 i23458 (.D0(n25212), .D1(n25210), .SD(index_q[5]), .Z(n25213));
    LUT4 i21537_3_lut (.A(n21460), .B(n27122), .C(index_q[4]), .Z(n21462)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21537_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_3_i924_3_lut (.A(n908_adj_2420), .B(index_q[0]), .C(index_q[4]), 
         .Z(n924_adj_2421)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_3_i924_3_lut.init = 16'hcaca;
    PFUMX i23456 (.BLUT(n25211), .ALUT(n285_adj_2422), .C0(index_q[4]), 
          .Z(n25212));
    LUT4 i18989_else_4_lut (.A(index_q[0]), .B(index_q[4]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n27159)) /* synthesis lut_function=(!(A (B (C)+!B !(C+!(D)))+!A (B (C)+!B (D)))) */ ;
    defparam i18989_else_4_lut.init = 16'h2c3f;
    L6MUX21 i20256 (.D0(n21705), .D1(n21708), .SD(index_q[6]), .Z(n22712));
    PFUMX i19475 (.BLUT(n21910), .ALUT(n21911), .C0(index_q[4]), .Z(n21912));
    PFUMX i18986 (.BLUT(n21421), .ALUT(n21422), .C0(index_q[4]), .Z(n476_adj_2423));
    L6MUX21 i20157 (.D0(n22597), .D1(n22598), .SD(index_q[6]), .Z(n22613));
    L6MUX21 i20158 (.D0(n22599), .D1(n22600), .SD(index_q[6]), .Z(n22614));
    LUT4 mux_197_Mux_3_i891_3_lut (.A(n541_adj_2424), .B(n890_adj_2425), 
         .C(index_q[4]), .Z(n891_adj_2426)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_3_i891_3_lut.init = 16'hcaca;
    L6MUX21 i20159 (.D0(n22601), .D1(n22602), .SD(index_q[6]), .Z(n22615));
    PFUMX i15546 (.BLUT(n17808), .ALUT(n17809), .C0(index_q[4]), .Z(n17810));
    LUT4 n24867_bdd_3_lut (.A(n27220), .B(n444_adj_2427), .C(index_i[5]), 
         .Z(n24868)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n24867_bdd_3_lut.init = 16'hcaca;
    PFUMX i20161 (.BLUT(n22605), .ALUT(n22606), .C0(index_q[6]), .Z(n22617));
    L6MUX21 i20162 (.D0(n22607), .D1(n22608), .SD(index_q[6]), .Z(n22618));
    L6MUX21 i20163 (.D0(n22609), .D1(n22610), .SD(index_q[6]), .Z(n22619));
    PFUMX i20164 (.BLUT(n22611), .ALUT(n22612), .C0(index_q[6]), .Z(n22620));
    LUT4 mux_197_Mux_3_i669_3_lut (.A(n653_adj_2268), .B(n668_adj_2428), 
         .C(index_q[4]), .Z(n669)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_3_i669_3_lut.init = 16'hcaca;
    L6MUX21 i21034 (.D0(n23482), .D1(n23483), .SD(index_i[6]), .Z(n23490));
    LUT4 i9412_4_lut (.A(n27090), .B(n26861), .C(index_q[3]), .D(index_q[4]), 
         .Z(n11973)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B ((D)+!C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9412_4_lut.init = 16'h3afa;
    L6MUX21 i21035 (.D0(n23484), .D1(n23485), .SD(index_i[6]), .Z(n23491));
    L6MUX21 i21036 (.D0(n23486), .D1(n23487), .SD(index_i[6]), .Z(n23492));
    PFUMX i19490 (.BLUT(n21925), .ALUT(n21926), .C0(index_i[4]), .Z(n21927));
    L6MUX21 i21037 (.D0(n23488), .D1(n23489), .SD(index_i[6]), .Z(n23493));
    PFUMX i20184 (.BLUT(n797_adj_2373), .ALUT(n828_adj_2429), .C0(index_q[5]), 
          .Z(n22640));
    LUT4 i18964_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21401)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A (B (C (D)+!C !(D))+!B (D))) */ ;
    defparam i18964_3_lut_4_lut.init = 16'hd926;
    LUT4 i21546_3_lut (.A(n21448), .B(n21449), .C(index_q[4]), .Z(n21450)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21546_3_lut.init = 16'hcaca;
    L6MUX21 i20188 (.D0(n22628), .D1(n22629), .SD(index_q[6]), .Z(n22644));
    LUT4 mux_197_Mux_3_i476_3_lut (.A(n460_adj_2430), .B(n285_adj_2422), 
         .C(index_q[4]), .Z(n476_adj_2431)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_3_i476_3_lut.init = 16'hcaca;
    PFUMX i20723 (.BLUT(n23175), .ALUT(n23176), .C0(index_q[6]), .Z(n23179));
    LUT4 mux_197_Mux_3_i413_3_lut (.A(n397_adj_2432), .B(n27056), .C(index_q[4]), 
         .Z(n413_adj_2433)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_3_i413_3_lut.init = 16'hcaca;
    PFUMX i19496 (.BLUT(n21931), .ALUT(n21932), .C0(index_i[4]), .Z(n21933));
    PFUMX i20724 (.BLUT(n23177), .ALUT(n23178), .C0(index_q[6]), .Z(n23180));
    LUT4 n77_bdd_3_lut_24147 (.A(n27083), .B(n29494), .C(index_q[3]), 
         .Z(n25965)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n77_bdd_3_lut_24147.init = 16'hacac;
    PFUMX i19499 (.BLUT(n21934), .ALUT(n21935), .C0(index_i[4]), .Z(n21936));
    LUT4 mux_197_Mux_3_i286_4_lut (.A(n93_adj_2434), .B(index_q[2]), .C(index_q[4]), 
         .D(n13941), .Z(n286)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_3_i286_4_lut.init = 16'h3aca;
    L6MUX21 i20189 (.D0(n22630), .D1(n22631), .SD(index_q[6]), .Z(n22645));
    L6MUX21 i20190 (.D0(n22632), .D1(n22633), .SD(index_q[6]), .Z(n22646));
    PFUMX i19505 (.BLUT(n21940), .ALUT(n21941), .C0(index_i[4]), .Z(n21942));
    PFUMX i24771 (.BLUT(n27189), .ALUT(n27190), .C0(index_q[0]), .Z(n27191));
    L6MUX21 i20191 (.D0(n22634), .D1(n22635), .SD(index_q[6]), .Z(n22647));
    L6MUX21 i20192 (.D0(n22636), .D1(n22637), .SD(index_q[6]), .Z(n22648));
    LUT4 mux_196_Mux_5_i572_3_lut_4_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[1]), .D(index_i[3]), .Z(n572_adj_2435)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A !(B (C+(D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_5_i572_3_lut_4_lut.init = 16'haa95;
    LUT4 mux_197_Mux_3_i158_3_lut (.A(n142_adj_2436), .B(n157_adj_2437), 
         .C(index_q[4]), .Z(n158_adj_2438)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_3_i158_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_7_i491_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n491_adj_2439)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(D))+!A (B (C+!(D))+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_7_i491_3_lut_4_lut_4_lut_4_lut.init = 16'h3780;
    LUT4 mux_197_Mux_3_i125_3_lut (.A(n109_adj_2349), .B(n526_adj_2417), 
         .C(index_q[4]), .Z(n125_adj_2440)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_3_i125_3_lut.init = 16'hcaca;
    L6MUX21 i20195 (.D0(n22642), .D1(n22643), .SD(index_q[6]), .Z(n22651));
    LUT4 i11452_3_lut_4_lut (.A(n26713), .B(index_q[7]), .C(index_q[8]), 
         .D(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_2141[14])) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11452_3_lut_4_lut.init = 16'hffe0;
    LUT4 i19534_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21971)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A (B (C (D)+!C !(D))+!B (D))) */ ;
    defparam i19534_3_lut_4_lut.init = 16'hd926;
    L6MUX21 i20210 (.D0(n23008), .D1(n23015), .SD(index_i[6]), .Z(n22666));
    PFUMX i20217 (.BLUT(n956), .ALUT(n20334), .C0(index_i[6]), .Z(n22673));
    LUT4 n24902_bdd_3_lut (.A(n24902), .B(n476), .C(index_i[5]), .Z(n24903)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n24902_bdd_3_lut.init = 16'hcaca;
    LUT4 i18976_3_lut (.A(n27065), .B(n27072), .C(index_q[3]), .Z(n21413)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18976_3_lut.init = 16'hcaca;
    LUT4 i11607_3_lut_4_lut (.A(n27034), .B(index_q[4]), .C(index_q[5]), 
         .D(n27101), .Z(n892_adj_2441)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11607_3_lut_4_lut.init = 16'hf8f0;
    LUT4 i21608_3_lut (.A(n21412), .B(n21413), .C(index_q[4]), .Z(n21414)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21608_3_lut.init = 16'hcaca;
    LUT4 n62_bdd_3_lut_25962 (.A(n62_adj_2261), .B(n125_adj_2400), .C(index_q[6]), 
         .Z(n28534)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n62_bdd_3_lut_25962.init = 16'hcaca;
    LUT4 n23184_bdd_4_lut_25959 (.A(n252_adj_2442), .B(n26863), .C(index_q[4]), 
         .D(index_q[5]), .Z(n28532)) /* synthesis lut_function=(A (B (D)+!B ((D)+!C))+!A !(B+(C+(D)))) */ ;
    defparam n23184_bdd_4_lut_25959.init = 16'haa03;
    LUT4 i20156_4_lut (.A(n21441), .B(n1002_adj_2443), .C(index_q[5]), 
         .D(index_q[4]), .Z(n22612)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;
    defparam i20156_4_lut.init = 16'hfaca;
    PFUMX i20226 (.BLUT(n94), .ALUT(n125_adj_2444), .C0(index_i[5]), .Z(n22682));
    LUT4 n62_bdd_4_lut_25963 (.A(n26994), .B(n26859), .C(index_q[6]), 
         .D(index_q[4]), .Z(n28535)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C+(D)))+!A (B ((D)+!C)+!B !(C)))) */ ;
    defparam n62_bdd_4_lut_25963.init = 16'h3af0;
    PFUMX i23454 (.BLUT(n25209), .ALUT(n25208), .C0(index_q[4]), .Z(n25210));
    LUT4 mux_197_Mux_4_i860_3_lut (.A(n506_adj_2445), .B(n25447), .C(index_q[4]), 
         .Z(n860_adj_2446)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_4_i860_3_lut.init = 16'hcaca;
    PFUMX i20227 (.BLUT(n17830), .ALUT(n14440), .C0(index_i[5]), .Z(n22683));
    LUT4 i21587_3_lut (.A(n21430), .B(n21431), .C(index_q[4]), .Z(n21432)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21587_3_lut.init = 16'hcaca;
    LUT4 n62_bdd_3_lut_25953 (.A(n62_adj_2281), .B(n125), .C(index_i[6]), 
         .Z(n28556)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n62_bdd_3_lut_25953.init = 16'hcaca;
    L6MUX21 i20229 (.D0(n21957), .D1(n21960), .SD(index_i[5]), .Z(n22685));
    L6MUX21 i20230 (.D0(n21963), .D1(n21966), .SD(index_i[5]), .Z(n22686));
    PFUMX i20231 (.BLUT(n413_adj_2447), .ALUT(n444_adj_2448), .C0(index_i[5]), 
          .Z(n22687));
    LUT4 mux_197_Mux_11_i638_4_lut_4_lut (.A(n26737), .B(index_q[5]), .C(index_q[6]), 
         .D(n26773), .Z(n638)) /* synthesis lut_function=(A (B (C (D))+!B !(C))+!A (B ((D)+!C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_11_i638_4_lut_4_lut.init = 16'hc707;
    LUT4 n23337_bdd_4_lut_25950 (.A(n252_adj_2316), .B(n26864), .C(index_i[4]), 
         .D(index_i[5]), .Z(n28554)) /* synthesis lut_function=(A (B (D)+!B ((D)+!C))+!A !(B+(C+(D)))) */ ;
    defparam n23337_bdd_4_lut_25950.init = 16'haa03;
    PFUMX i20232 (.BLUT(n476_adj_2449), .ALUT(n507), .C0(index_i[5]), 
          .Z(n22688));
    LUT4 n715_bdd_3_lut_24265 (.A(n27104), .B(n27084), .C(index_q[3]), 
         .Z(n26014)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n715_bdd_3_lut_24265.init = 16'hcaca;
    PFUMX i15549 (.BLUT(n17811), .ALUT(n17812), .C0(index_i[4]), .Z(n17813));
    PFUMX i20233 (.BLUT(n17816), .ALUT(n573_adj_2450), .C0(index_i[5]), 
          .Z(n22689));
    LUT4 n62_bdd_4_lut_25954 (.A(n26898), .B(n26835), .C(index_i[6]), 
         .D(index_i[4]), .Z(n28557)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C+(D)))+!A (B ((D)+!C)+!B !(C)))) */ ;
    defparam n62_bdd_4_lut_25954.init = 16'h3af0;
    LUT4 i11445_3_lut_4_lut (.A(index_i[4]), .B(n27035), .C(index_i[5]), 
         .D(n26927), .Z(n892_adj_2451)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11445_3_lut_4_lut.init = 16'hf8f0;
    PFUMX i20234 (.BLUT(n605_adj_2452), .ALUT(n636_adj_2453), .C0(index_i[5]), 
          .Z(n22690));
    PFUMX i20235 (.BLUT(n21969), .ALUT(n700_adj_2454), .C0(index_i[5]), 
          .Z(n22691));
    LUT4 mux_197_Mux_4_i62_4_lut (.A(n27091), .B(n61), .C(index_q[4]), 
         .D(index_q[3]), .Z(n62_adj_2455)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_4_i62_4_lut.init = 16'hc5ca;
    LUT4 mux_197_Mux_4_i31_4_lut (.A(n15_adj_2456), .B(n26834), .C(index_q[4]), 
         .D(index_q[3]), .Z(n31)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_4_i31_4_lut.init = 16'h3aca;
    LUT4 mux_197_Mux_4_i828_3_lut_4_lut (.A(index_q[4]), .B(index_q[3]), 
         .C(n812_adj_2285), .D(n27094), .Z(n828_adj_2457)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_4_i828_3_lut_4_lut.init = 16'hf1e0;
    L6MUX21 i20236 (.D0(n732), .D1(n21972), .SD(index_i[5]), .Z(n22692));
    PFUMX i20237 (.BLUT(n797_adj_2458), .ALUT(n828_adj_2459), .C0(index_i[5]), 
          .Z(n22693));
    PFUMX i19508 (.BLUT(n21943), .ALUT(n21944), .C0(index_i[4]), .Z(n21945));
    LUT4 n715_bdd_3_lut_24561_4_lut (.A(n27101), .B(index_q[2]), .C(index_q[3]), 
         .D(n27104), .Z(n26512)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n715_bdd_3_lut_24561_4_lut.init = 16'hdfd0;
    PFUMX i20749 (.BLUT(n23189), .ALUT(n23190), .C0(index_i[5]), .Z(n23205));
    LUT4 i12185_3_lut (.A(index_i[3]), .B(index_i[1]), .C(index_i[0]), 
         .Z(n14871)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i12185_3_lut.init = 16'hecec;
    LUT4 i19339_3_lut_4_lut (.A(n27101), .B(index_q[2]), .C(index_q[3]), 
         .D(n27077), .Z(n21776)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19339_3_lut_4_lut.init = 16'hdfd0;
    PFUMX i20238 (.BLUT(n860_adj_2460), .ALUT(n891_adj_2461), .C0(index_i[5]), 
          .Z(n22694));
    PFUMX i20750 (.BLUT(n23191), .ALUT(n23192), .C0(index_i[5]), .Z(n23206));
    LUT4 i21599_3_lut (.A(n21427), .B(n21428), .C(index_q[4]), .Z(n21429)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21599_3_lut.init = 16'hcaca;
    L6MUX21 i20751 (.D0(n23193), .D1(n23194), .SD(index_i[5]), .Z(n23207));
    LUT4 mux_197_Mux_4_i700_3_lut (.A(n684_adj_2462), .B(index_q[1]), .C(index_q[4]), 
         .Z(n700_adj_2463)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_4_i700_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_4_i669_3_lut (.A(n653_adj_2464), .B(n668_adj_2375), 
         .C(index_q[4]), .Z(n669_adj_2465)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_4_i669_3_lut.init = 16'hcaca;
    LUT4 i19711_3_lut_4_lut (.A(index_q[0]), .B(n27063), .C(index_q[3]), 
         .D(n27065), .Z(n22148)) /* synthesis lut_function=(A ((D)+!C)+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19711_3_lut_4_lut.init = 16'hfb0b;
    LUT4 mux_197_Mux_4_i542_3_lut (.A(n526_adj_2417), .B(n541), .C(index_q[4]), 
         .Z(n542_adj_2466)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_4_i542_3_lut.init = 16'hcaca;
    LUT4 i20150_4_lut (.A(n26816), .B(n27161), .C(index_q[5]), .D(index_q[4]), 
         .Z(n22606)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam i20150_4_lut.init = 16'hc5ca;
    LUT4 mux_197_Mux_3_i31_3_lut (.A(n653_adj_2464), .B(n30_adj_2467), .C(index_q[4]), 
         .Z(n31_adj_2468)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_3_i31_3_lut.init = 16'hcaca;
    LUT4 n24906_bdd_3_lut_23422 (.A(n27217), .B(n24904), .C(index_i[5]), 
         .Z(n24907)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n24906_bdd_3_lut_23422.init = 16'hcaca;
    LUT4 i9454_3_lut_4_lut (.A(index_q[0]), .B(n27063), .C(index_q[4]), 
         .D(n588), .Z(n12015)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9454_3_lut_4_lut.init = 16'h4f40;
    LUT4 mux_197_Mux_4_i286_3_lut (.A(n270), .B(n15_adj_2456), .C(index_q[4]), 
         .Z(n286_adj_2469)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_4_i286_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_2_i700_3_lut_4_lut (.A(index_i[1]), .B(n26898), .C(index_i[4]), 
         .D(n684_adj_2383), .Z(n700_adj_2470)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_2_i700_3_lut_4_lut.init = 16'hefe0;
    LUT4 mux_196_Mux_3_i1018_3_lut_4_lut (.A(index_i[1]), .B(n26898), .C(index_i[4]), 
         .D(n19881), .Z(n1018)) /* synthesis lut_function=(A (C+!(D))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_3_i1018_3_lut_4_lut.init = 16'he0ef;
    LUT4 mux_196_Mux_5_i31_3_lut (.A(n15_adj_2471), .B(n30_adj_2472), .C(index_i[4]), 
         .Z(n31_adj_2473)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_5_i31_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_2_i348_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[1]), .D(index_i[3]), .Z(n348_adj_2474)) /* synthesis lut_function=(!(A (B (D)+!B (C+!(D)))+!A !(B (D)+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_2_i348_3_lut_4_lut_4_lut.init = 16'h4699;
    LUT4 mux_196_Mux_4_i62_4_lut (.A(n27047), .B(n61_adj_2475), .C(index_i[4]), 
         .D(index_i[3]), .Z(n62_adj_2476)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_4_i62_4_lut.init = 16'hc5ca;
    LUT4 mux_197_Mux_0_i491_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n491_adj_2477)) /* synthesis lut_function=(!(A (B (D)+!B !(C+!(D)))+!A ((C+!(D))+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i491_3_lut_4_lut.init = 16'h24aa;
    LUT4 mux_196_Mux_4_i31_4_lut (.A(n15_adj_2478), .B(n26792), .C(index_i[4]), 
         .D(index_i[3]), .Z(n31_adj_2479)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_4_i31_4_lut.init = 16'h3aca;
    LUT4 mux_197_Mux_4_i94_3_lut (.A(n61), .B(n27057), .C(index_q[4]), 
         .Z(n94_adj_2480)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_4_i94_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_3_i31_3_lut (.A(n781_adj_2260), .B(n30_adj_2481), .C(index_i[4]), 
         .Z(n31_adj_2482)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_3_i31_3_lut.init = 16'hcaca;
    L6MUX21 i20754 (.D0(n23199), .D1(n23200), .SD(index_i[5]), .Z(n23210));
    PFUMX i19520 (.BLUT(n21955), .ALUT(n21956), .C0(index_i[4]), .Z(n21957));
    L6MUX21 i20755 (.D0(n23201), .D1(n23202), .SD(index_i[5]), .Z(n23211));
    LUT4 i9543_3_lut (.A(n12103), .B(n29488), .C(index_i[3]), .Z(n12104)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9543_3_lut.init = 16'hcaca;
    L6MUX21 i20756 (.D0(n23203), .D1(n23204), .SD(index_i[5]), .Z(n23212));
    LUT4 i20841_3_lut_4_lut (.A(n26813), .B(n26776), .C(index_i[4]), .D(index_i[5]), 
         .Z(n23297)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (B+((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20841_3_lut_4_lut.init = 16'hffc5;
    LUT4 i20735_3_lut_3_lut_4_lut (.A(n26836), .B(index_i[3]), .C(n93), 
         .D(index_i[4]), .Z(n23191)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20735_3_lut_3_lut_4_lut.init = 16'hf077;
    LUT4 i20881_4_lut_4_lut (.A(n26781), .B(n26877), .C(index_i[5]), .D(index_i[4]), 
         .Z(n23337)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C+(D))+!B !(C (D)+!C !(D)))) */ ;
    defparam i20881_4_lut_4_lut.init = 16'hcf50;
    PFUMX i20272 (.BLUT(n94_adj_2483), .ALUT(n21975), .C0(index_i[5]), 
          .Z(n22728));
    LUT4 mux_196_Mux_7_i890_3_lut_4_lut (.A(n26996), .B(index_i[2]), .C(index_i[3]), 
         .D(n26876), .Z(n890_adj_2291)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_7_i890_3_lut_4_lut.init = 16'hf101;
    LUT4 mux_196_Mux_0_i1002_3_lut_3_lut_4_lut (.A(n26996), .B(index_i[2]), 
         .C(n38), .D(index_i[3]), .Z(n1002_adj_2484)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_0_i1002_3_lut_3_lut_4_lut.init = 16'hf011;
    PFUMX i20274 (.BLUT(n221_adj_2485), .ALUT(n252_adj_2486), .C0(index_i[5]), 
          .Z(n22730));
    LUT4 mux_196_Mux_9_i124_3_lut_4_lut (.A(n26996), .B(index_i[2]), .C(index_i[3]), 
         .D(n26875), .Z(n124_adj_2388)) /* synthesis lut_function=(!(A (C+!(D))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_9_i124_3_lut_4_lut.init = 16'h1f10;
    LUT4 mux_196_Mux_3_i93_3_lut_4_lut (.A(n26996), .B(index_i[2]), .C(index_i[3]), 
         .D(n70), .Z(n93_adj_2487)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_3_i93_3_lut_4_lut.init = 16'hefe0;
    L6MUX21 mux_197_Mux_7_i253 (.D0(n12134), .D1(n22116), .SD(index_q[5]), 
            .Z(n253)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    PFUMX i20275 (.BLUT(n286_adj_2488), .ALUT(n21978), .C0(index_i[5]), 
          .Z(n22731));
    LUT4 mux_196_Mux_3_i221_3_lut_4_lut (.A(n26836), .B(index_i[3]), .C(index_i[4]), 
         .D(n26864), .Z(n221_adj_2489)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_3_i221_3_lut_4_lut.init = 16'h08f8;
    PFUMX i19523 (.BLUT(n21958), .ALUT(n21959), .C0(index_i[4]), .Z(n21960));
    LUT4 mux_196_Mux_8_i124_3_lut_3_lut_4_lut (.A(n26996), .B(index_i[2]), 
         .C(n29492), .D(index_i[3]), .Z(n124_adj_2363)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_8_i124_3_lut_3_lut_4_lut.init = 16'h11f0;
    PFUMX i19526 (.BLUT(n21961), .ALUT(n21962), .C0(index_i[4]), .Z(n21963));
    PFUMX i20276 (.BLUT(n349), .ALUT(n21981), .C0(index_i[5]), .Z(n22732));
    LUT4 mux_196_Mux_6_i890_3_lut_4_lut (.A(n26996), .B(index_i[2]), .C(index_i[3]), 
         .D(n27000), .Z(n890_adj_2490)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_6_i890_3_lut_4_lut.init = 16'hf101;
    LUT4 mux_196_Mux_7_i315_3_lut_rep_795 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n29468)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_7_i315_3_lut_rep_795.init = 16'h3838;
    LUT4 mux_196_Mux_8_i475_3_lut_4_lut (.A(n26996), .B(index_i[2]), .C(index_i[3]), 
         .D(n26875), .Z(n475_adj_2491)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_8_i475_3_lut_4_lut.init = 16'hf101;
    LUT4 mux_197_Mux_1_i700_3_lut_4_lut (.A(n26973), .B(index_q[3]), .C(index_q[4]), 
         .D(n684_adj_2318), .Z(n700_adj_2492)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_1_i700_3_lut_4_lut.init = 16'hefe0;
    LUT4 i19945_2_lut (.A(index_q[3]), .B(index_q[5]), .Z(n22401)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19945_2_lut.init = 16'h8888;
    LUT4 i20734_3_lut_4_lut (.A(n26836), .B(index_i[3]), .C(index_i[4]), 
         .D(n46), .Z(n23190)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20734_3_lut_4_lut.init = 16'h8f80;
    LUT4 index_q_1__bdd_4_lut_26349 (.A(index_q[1]), .B(index_q[3]), .C(index_q[0]), 
         .D(index_q[2]), .Z(n28805)) /* synthesis lut_function=(A (B (C+(D))+!B (C (D)))+!A !(B (C)+!B !(C+(D)))) */ ;
    defparam index_q_1__bdd_4_lut_26349.init = 16'hbd94;
    LUT4 n28805_bdd_3_lut (.A(n28805), .B(index_q[1]), .C(index_q[4]), 
         .Z(n28806)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n28805_bdd_3_lut.init = 16'hcaca;
    LUT4 n730_bdd_3_lut_23428 (.A(n27032), .B(n26991), .C(index_i[3]), 
         .Z(n24962)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n730_bdd_3_lut_23428.init = 16'hcaca;
    PFUMX mux_197_Mux_7_i190 (.BLUT(n22113), .ALUT(n173_adj_2493), .C0(index_q[5]), 
          .Z(n190)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 mux_197_Mux_5_i891_3_lut (.A(n875_adj_2494), .B(n890_adj_2376), 
         .C(index_q[4]), .Z(n891_adj_2495)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_5_i891_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_5_i860_3_lut (.A(n15_adj_2496), .B(n859_adj_2497), 
         .C(index_q[4]), .Z(n860_adj_2498)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_5_i860_3_lut.init = 16'hcaca;
    LUT4 i21646_3_lut (.A(n21397), .B(n21398), .C(index_q[4]), .Z(n21399)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21646_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_5_i636_4_lut (.A(n157_adj_2499), .B(n26892), .C(index_q[4]), 
         .D(index_q[3]), .Z(n636_adj_2500)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_5_i636_4_lut.init = 16'h3aca;
    LUT4 mux_196_Mux_3_i796_3_lut (.A(index_i[2]), .B(n731_adj_2501), .C(index_i[4]), 
         .Z(n796_adj_2502)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_3_i796_3_lut.init = 16'hacac;
    LUT4 mux_196_Mux_6_i731_3_lut (.A(n26928), .B(n29468), .C(index_i[3]), 
         .Z(n731_adj_2501)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_6_i731_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_0_i781_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n781)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A (B (C)+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i781_4_lut_4_lut_4_lut.init = 16'h0cb4;
    LUT4 n21595_bdd_4_lut_23769 (.A(n27035), .B(n763_adj_2414), .C(index_i[5]), 
         .D(index_i[4]), .Z(n24617)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam n21595_bdd_4_lut_23769.init = 16'hcfca;
    PFUMX i20281 (.BLUT(n669_adj_2503), .ALUT(n700_adj_2504), .C0(index_i[5]), 
          .Z(n22737));
    LUT4 i21649_3_lut (.A(n17786), .B(n17787), .C(index_q[4]), .Z(n17788)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21649_3_lut.init = 16'hcaca;
    PFUMX i19529 (.BLUT(n21964), .ALUT(n21965), .C0(index_i[4]), .Z(n21966));
    PFUMX i20282 (.BLUT(n22002), .ALUT(n763_adj_2356), .C0(index_i[5]), 
          .Z(n22738));
    PFUMX i20283 (.BLUT(n22005), .ALUT(n828_adj_2505), .C0(index_i[5]), 
          .Z(n22739));
    LUT4 mux_196_Mux_5_i124_3_lut (.A(n26900), .B(n27026), .C(index_i[3]), 
         .Z(n124_adj_2506)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_5_i124_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_5_i507_3_lut (.A(n491_adj_2507), .B(n506_adj_2445), 
         .C(index_q[4]), .Z(n507_adj_2508)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_5_i507_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_5_i476_3_lut (.A(n460_adj_2509), .B(n475), .C(index_q[4]), 
         .Z(n476_adj_2510)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_5_i476_3_lut.init = 16'hcaca;
    PFUMX i20284 (.BLUT(n860_adj_2511), .ALUT(n22008), .C0(index_i[5]), 
          .Z(n22740));
    LUT4 mux_197_Mux_5_i413_3_lut (.A(n397_adj_2512), .B(n251_adj_2371), 
         .C(index_q[4]), .Z(n413_adj_2513)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_5_i413_3_lut.init = 16'hcaca;
    PFUMX i19535 (.BLUT(n21970), .ALUT(n21971), .C0(index_i[4]), .Z(n21972));
    LUT4 n197_bdd_3_lut_23227 (.A(n26991), .B(index_i[3]), .C(n27023), 
         .Z(n24959)) /* synthesis lut_function=(A (B+(C))+!A !(B+!(C))) */ ;
    defparam n197_bdd_3_lut_23227.init = 16'hb8b8;
    LUT4 i15560_3_lut (.A(n17822), .B(n17823), .C(index_q[4]), .Z(n17824)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15560_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_5_i125_3_lut (.A(n109_adj_2514), .B(n124_adj_2515), 
         .C(index_q[4]), .Z(n125_adj_2516)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_5_i125_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_5_i797_3_lut_4_lut (.A(index_q[4]), .B(index_q[3]), 
         .C(n27131), .D(n27099), .Z(n797_adj_2517)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_5_i797_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_197_Mux_5_i94_3_lut (.A(n653_adj_2253), .B(n635_adj_2419), 
         .C(index_q[4]), .Z(n94_adj_2518)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_5_i94_3_lut.init = 16'hcaca;
    LUT4 n404_bdd_3_lut_23234 (.A(n404), .B(n26934), .C(index_i[3]), .Z(n24965)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n404_bdd_3_lut_23234.init = 16'hcaca;
    LUT4 n404_bdd_3_lut_23731 (.A(index_i[3]), .B(n27027), .C(n27028), 
         .Z(n24966)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam n404_bdd_3_lut_23731.init = 16'he4e4;
    LUT4 mux_197_Mux_5_i31_3_lut (.A(n15_adj_2496), .B(n30_adj_2519), .C(index_q[4]), 
         .Z(n31_adj_2520)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_5_i31_3_lut.init = 16'hcaca;
    LUT4 n470_bdd_3_lut (.A(n26989), .B(n29487), .C(index_i[3]), .Z(n24969)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n470_bdd_3_lut.init = 16'hacac;
    PFUMX i21011 (.BLUT(n557_adj_2521), .ALUT(n572_adj_2522), .C0(index_i[4]), 
          .Z(n23467));
    LUT4 i15570_4_lut (.A(index_q[0]), .B(index_q[4]), .C(index_q[1]), 
         .D(n26994), .Z(n286_adj_2523)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i15570_4_lut.init = 16'hccc8;
    LUT4 index_q_5__bdd_3_lut (.A(index_q[5]), .B(n29040), .C(index_q[3]), 
         .Z(n29041)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam index_q_5__bdd_3_lut.init = 16'hcaca;
    LUT4 index_q_6__bdd_4_lut_26157 (.A(index_q[6]), .B(index_q[5]), .C(index_q[1]), 
         .D(index_q[0]), .Z(n29039)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C))+!A (B (C)+!B !(C)))) */ ;
    defparam index_q_6__bdd_4_lut_26157.init = 16'h3cbc;
    LUT4 i20728_4_lut_4_lut (.A(n26767), .B(n26872), .C(index_q[5]), .D(index_q[4]), 
         .Z(n23184)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C+(D))+!B !(C (D)+!C !(D)))) */ ;
    defparam i20728_4_lut_4_lut.init = 16'hcf50;
    LUT4 index_q_6__bdd_1_lut (.A(index_q[5]), .Z(n29038)) /* synthesis lut_function=(!(A)) */ ;
    defparam index_q_6__bdd_1_lut.init = 16'h5555;
    LUT4 n27101_bdd_3_lut_26398 (.A(n26871), .B(index_q[6]), .C(index_q[5]), 
         .Z(n29042)) /* synthesis lut_function=(!(A (B)+!A (C))) */ ;
    defparam n27101_bdd_3_lut_26398.init = 16'h2727;
    PFUMX i21012 (.BLUT(n589_adj_2524), .ALUT(n604_adj_2317), .C0(index_i[4]), 
          .Z(n23468));
    LUT4 n27101_bdd_4_lut (.A(n27101), .B(index_q[6]), .C(index_q[2]), 
         .D(index_q[5]), .Z(n29043)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A !(B (C+(D))+!B (D)))) */ ;
    defparam n27101_bdd_4_lut.init = 16'h5fe0;
    LUT4 n29044_bdd_3_lut (.A(n29044), .B(n29041), .C(index_q[4]), .Z(n29045)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n29044_bdd_3_lut.init = 16'hcaca;
    PFUMX i20098 (.BLUT(n221), .ALUT(n252_adj_2307), .C0(index_q[5]), 
          .Z(n22554));
    PFUMX i20303 (.BLUT(n94_adj_2525), .ALUT(n125_adj_2526), .C0(index_i[5]), 
          .Z(n22759));
    CCU2D add_377_11 (.A0(quarter_wave_sample_register_q[10]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_q[11]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17575), .COUT(n17576), 
          .S0(o_val_pipeline_q_0__15__N_2189[10]), .S1(o_val_pipeline_q_0__15__N_2189[11]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(80[29:60])
    defparam add_377_11.INIT0 = 16'hf555;
    defparam add_377_11.INIT1 = 16'hf555;
    defparam add_377_11.INJECT1_0 = "NO";
    defparam add_377_11.INJECT1_1 = "NO";
    LUT4 mux_197_Mux_1_i924_3_lut (.A(n316_adj_2527), .B(n923_adj_2528), 
         .C(index_q[4]), .Z(n924_adj_2529)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_1_i924_3_lut.init = 16'hcaca;
    PFUMX i20304 (.BLUT(n158_adj_2530), .ALUT(n189_adj_2286), .C0(index_i[5]), 
          .Z(n22760));
    PFUMX i24769 (.BLUT(n27186), .ALUT(n27187), .C0(index_q[0]), .Z(n27188));
    LUT4 n24973_bdd_3_lut (.A(n24973), .B(n157_adj_2531), .C(index_i[4]), 
         .Z(n24974)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n24973_bdd_3_lut.init = 16'hcaca;
    LUT4 i21674_3_lut (.A(n21766), .B(n21767), .C(index_q[4]), .Z(n21768)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21674_3_lut.init = 16'hcaca;
    PFUMX i20305 (.BLUT(n221_adj_2489), .ALUT(n252_adj_2284), .C0(index_i[5]), 
          .Z(n22761));
    LUT4 mux_197_Mux_6_i285_3_lut_4_lut (.A(n27064), .B(index_q[2]), .C(index_q[3]), 
         .D(n27083), .Z(n285_adj_2422)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_6_i285_3_lut_4_lut.init = 16'hf606;
    LUT4 i18958_3_lut_4_lut (.A(n27064), .B(index_q[2]), .C(index_q[3]), 
         .D(n29474), .Z(n21395)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18958_3_lut_4_lut.init = 16'h6f60;
    LUT4 index_q_7__bdd_4_lut_24900 (.A(index_q[7]), .B(n125_adj_2532), 
         .C(n24748), .D(index_q[5]), .Z(n26706)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(B (C+(D))+!B !((D)+!C)))) */ ;
    defparam index_q_7__bdd_4_lut_24900.init = 16'h66f0;
    LUT4 index_i_7__bdd_4_lut_24924 (.A(index_i[7]), .B(n15124), .C(n24731), 
         .D(index_i[5]), .Z(n26707)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(B (C+(D))+!B !((D)+!C)))) */ ;
    defparam index_i_7__bdd_4_lut_24924.init = 16'h66f0;
    LUT4 index_i_6__bdd_4_lut_26215 (.A(index_i[6]), .B(index_i[5]), .C(index_i[1]), 
         .D(index_i[0]), .Z(n29159)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C))+!A (B (C)+!B !(C)))) */ ;
    defparam index_i_6__bdd_4_lut_26215.init = 16'h3cbc;
    LUT4 i19696_3_lut_4_lut (.A(n27064), .B(index_q[2]), .C(index_q[3]), 
         .D(n27098), .Z(n22133)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19696_3_lut_4_lut.init = 16'hf606;
    LUT4 index_i_6__bdd_1_lut (.A(index_i[5]), .Z(n29158)) /* synthesis lut_function=(!(A)) */ ;
    defparam index_i_6__bdd_1_lut.init = 16'h5555;
    LUT4 n187_bdd_4_lut_24157 (.A(n26836), .B(index_i[6]), .C(index_i[5]), 
         .D(n27003), .Z(n24994)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(D))+!A !(B (C+(D))+!B (D)))) */ ;
    defparam n187_bdd_4_lut_24157.init = 16'h7f40;
    LUT4 mux_197_Mux_3_i460_3_lut_4_lut (.A(n27064), .B(index_q[2]), .C(index_q[3]), 
         .D(n29493), .Z(n460_adj_2430)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_3_i460_3_lut_4_lut.init = 16'h6f60;
    LUT4 index_i_5__bdd_3_lut (.A(index_i[5]), .B(n29160), .C(index_i[3]), 
         .Z(n29161)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam index_i_5__bdd_3_lut.init = 16'hcaca;
    LUT4 n26927_bdd_3_lut (.A(n26876), .B(index_i[6]), .C(index_i[5]), 
         .Z(n29162)) /* synthesis lut_function=(!(A (B)+!A (C))) */ ;
    defparam n26927_bdd_3_lut.init = 16'h2727;
    LUT4 n26927_bdd_4_lut (.A(n26927), .B(index_i[6]), .C(index_i[2]), 
         .D(index_i[5]), .Z(n29163)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A !(B (C+(D))+!B (D)))) */ ;
    defparam n26927_bdd_4_lut.init = 16'h5fe0;
    LUT4 n29164_bdd_3_lut (.A(n29164), .B(n29161), .C(index_i[4]), .Z(n29165)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n29164_bdd_3_lut.init = 16'hcaca;
    PFUMX i20306 (.BLUT(n286_adj_2533), .ALUT(n22017), .C0(index_i[5]), 
          .Z(n22762));
    LUT4 n24997_bdd_3_lut (.A(n27211), .B(n24994), .C(index_i[4]), .Z(n24998)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n24997_bdd_3_lut.init = 16'hcaca;
    LUT4 i19666_3_lut_4_lut_4_lut (.A(n26927), .B(n26934), .C(index_i[3]), 
         .D(index_i[2]), .Z(n22103)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B+(C))) */ ;
    defparam i19666_3_lut_4_lut_4_lut.init = 16'hfc5c;
    LUT4 mux_197_Mux_1_i763_3_lut_4_lut (.A(index_q[4]), .B(index_q[3]), 
         .C(n27145), .D(n27099), .Z(n763_adj_2391)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_1_i763_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_197_Mux_1_i301_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n301)) /* synthesis lut_function=(A (B (C+(D))+!B !(D))+!A !(B (C+(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_1_i301_3_lut_4_lut_4_lut.init = 16'h99b6;
    LUT4 n25000_bdd_3_lut (.A(n25000), .B(n24998), .C(index_i[3]), .Z(n25001)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n25000_bdd_3_lut.init = 16'hcaca;
    PFUMX i20307 (.BLUT(n349_adj_2534), .ALUT(n22020), .C0(index_i[5]), 
          .Z(n22763));
    LUT4 i12055_2_lut_rep_590 (.A(index_q[2]), .B(index_q[0]), .Z(n26913)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12055_2_lut_rep_590.init = 16'h8888;
    PFUMX i21013 (.BLUT(n620_adj_2535), .ALUT(n635_adj_2536), .C0(index_i[4]), 
          .Z(n23469));
    LUT4 index_q_4__bdd_4_lut_25375 (.A(index_q[4]), .B(n26772), .C(n24488), 
         .D(index_q[5]), .Z(n26709)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (B (C (D))+!B (C+!(D)))) */ ;
    defparam index_q_4__bdd_4_lut_25375.init = 16'hf099;
    LUT4 mux_197_Mux_1_i349_3_lut (.A(n541), .B(n348), .C(index_q[4]), 
         .Z(n349_adj_2537)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_1_i349_3_lut.init = 16'hcaca;
    LUT4 i19603_3_lut_4_lut (.A(n26927), .B(index_i[2]), .C(index_i[3]), 
         .D(n308), .Z(n22040)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19603_3_lut_4_lut.init = 16'hf202;
    PFUMX i20308 (.BLUT(n413_adj_2538), .ALUT(n444_adj_2389), .C0(index_i[5]), 
          .Z(n22764));
    LUT4 mux_196_Mux_7_i506_3_lut_4_lut (.A(n26927), .B(index_i[2]), .C(index_i[3]), 
         .D(n29491), .Z(n506_adj_2359)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_7_i506_3_lut_4_lut.init = 16'h2f20;
    LUT4 i21692_3_lut (.A(n22147), .B(n22148), .C(index_q[4]), .Z(n22149)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21692_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_2_i189_3_lut_3_lut_4_lut (.A(index_i[1]), .B(n27035), 
         .C(n173), .D(index_i[4]), .Z(n189_adj_2539)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(C+(D)))) */ ;
    defparam mux_196_Mux_2_i189_3_lut_3_lut_4_lut.init = 16'h77f0;
    PFUMX i20309 (.BLUT(n476_adj_2540), .ALUT(n507_adj_2541), .C0(index_i[5]), 
          .Z(n22765));
    PFUMX i20310 (.BLUT(n22023), .ALUT(n573_adj_2393), .C0(index_i[5]), 
          .Z(n22766));
    LUT4 i11413_2_lut_3_lut_4_lut (.A(index_i[1]), .B(n27035), .C(index_i[5]), 
         .D(index_i[4]), .Z(n508_adj_2542)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;
    defparam i11413_2_lut_3_lut_4_lut.init = 16'hf080;
    PFUMX i19550 (.BLUT(n21985), .ALUT(n21986), .C0(index_q[4]), .Z(n21987));
    LUT4 i20875_3_lut_4_lut_4_lut (.A(n26821), .B(index_i[4]), .C(index_i[5]), 
         .D(n26842), .Z(n23331)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C)+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20875_3_lut_4_lut_4_lut.init = 16'h0434;
    PFUMX i20311 (.BLUT(n12091), .ALUT(n22026), .C0(index_i[5]), .Z(n22767));
    LUT4 mux_196_Mux_8_i892_3_lut_4_lut (.A(n26821), .B(index_i[4]), .C(index_i[5]), 
         .D(n860_adj_2278), .Z(n892_adj_2543)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_8_i892_3_lut_4_lut.init = 16'h4f40;
    PFUMX i20312 (.BLUT(n669_adj_2544), .ALUT(n700_adj_2545), .C0(index_i[5]), 
          .Z(n22768));
    L6MUX21 i20313 (.D0(n22029), .D1(n763), .SD(index_i[5]), .Z(n22769));
    PFUMX i20315 (.BLUT(n860_adj_2546), .ALUT(n891_adj_2547), .C0(index_i[5]), 
          .Z(n22771));
    LUT4 n269_bdd_3_lut_23599_4_lut (.A(n27068), .B(index_q[2]), .C(index_q[3]), 
         .D(n27066), .Z(n25209)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n269_bdd_3_lut_23599_4_lut.init = 16'hf606;
    PFUMX mux_197_Mux_1_i636 (.BLUT(n620_adj_2548), .ALUT(n635_adj_2549), 
          .C0(index_q[4]), .Z(n636_adj_2550)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 mux_197_Mux_3_i890_3_lut_4_lut (.A(n27068), .B(index_q[2]), .C(index_q[3]), 
         .D(n356), .Z(n890_adj_2425)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_3_i890_3_lut_4_lut.init = 16'h6f60;
    PFUMX i20316 (.BLUT(n924_adj_2551), .ALUT(n22032), .C0(index_i[5]), 
          .Z(n22772));
    LUT4 i19318_3_lut_4_lut (.A(n27068), .B(index_q[2]), .C(index_q[3]), 
         .D(n27083), .Z(n21755)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19318_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_197_Mux_1_i94_3_lut (.A(index_q[0]), .B(n93_adj_2552), .C(index_q[4]), 
         .Z(n94_adj_2553)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_1_i94_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_0_i348_3_lut_4_lut (.A(n27068), .B(index_q[2]), .C(index_q[3]), 
         .D(n29477), .Z(n348_adj_2554)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i348_3_lut_4_lut.init = 16'h6f60;
    LUT4 i9455_3_lut (.A(n12015), .B(n27082), .C(index_q[3]), .Z(n12016)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9455_3_lut.init = 16'hcaca;
    PFUMX i20317 (.BLUT(n22035), .ALUT(n1018), .C0(index_i[5]), .Z(n22773));
    PFUMX i21014 (.BLUT(n653_adj_2555), .ALUT(n668_adj_2556), .C0(index_i[4]), 
          .Z(n23470));
    PFUMX mux_197_Mux_8_i764 (.BLUT(n716_adj_2557), .ALUT(n732_adj_2558), 
          .C0(n22399), .Z(n764)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 mux_197_Mux_5_i124_3_lut (.A(n26887), .B(n27103), .C(index_q[3]), 
         .Z(n124_adj_2515)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_5_i124_3_lut.init = 16'hcaca;
    LUT4 i19480_3_lut_4_lut (.A(n27101), .B(index_q[2]), .C(index_q[3]), 
         .D(n27058), .Z(n21917)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19480_3_lut_4_lut.init = 16'h6f60;
    PFUMX i21015 (.BLUT(n684_adj_2338), .ALUT(n699_adj_2559), .C0(index_i[4]), 
          .Z(n23471));
    LUT4 i19300_3_lut_4_lut_4_lut_4_lut (.A(n27101), .B(index_q[2]), .C(index_q[3]), 
         .D(index_q[4]), .Z(n21737)) /* synthesis lut_function=(A (B)+!A (B (C (D))+!B !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19300_3_lut_4_lut_4_lut_4_lut.init = 16'hc999;
    LUT4 mux_197_Mux_2_i684_3_lut_4_lut (.A(n27101), .B(index_q[2]), .C(index_q[3]), 
         .D(n29477), .Z(n684_adj_2560)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_2_i684_3_lut_4_lut.init = 16'h6f60;
    LUT4 n254_bdd_4_lut (.A(index_q[5]), .B(index_q[3]), .C(index_q[6]), 
         .D(index_q[4]), .Z(n26215)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;
    defparam n254_bdd_4_lut.init = 16'hf8f0;
    LUT4 mux_196_Mux_8_i732_3_lut (.A(index_i[3]), .B(n15106), .C(index_i[5]), 
         .Z(n732_adj_2561)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_8_i732_3_lut.init = 16'h3a3a;
    LUT4 mux_197_Mux_0_i851_3_lut_3_lut_rep_802 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n29475)) /* synthesis lut_function=(A (B+(C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i851_3_lut_3_lut_rep_802.init = 16'hadad;
    LUT4 i20608_3_lut (.A(n27086), .B(n27105), .C(index_q[3]), .Z(n23064)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20608_3_lut.init = 16'hcaca;
    PFUMX i20335 (.BLUT(n158_adj_2562), .ALUT(n189_adj_2539), .C0(index_i[5]), 
          .Z(n22791));
    L6MUX21 i24611 (.D0(n26564), .D1(n26561), .SD(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_2141[4]));
    LUT4 i21723_3_lut (.A(n21922), .B(n21923), .C(index_i[4]), .Z(n21924)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i21723_3_lut.init = 16'hcaca;
    PFUMX i19553 (.BLUT(n21988), .ALUT(n21989), .C0(index_q[4]), .Z(n21990));
    LUT4 n26220_bdd_3_lut (.A(n27202), .B(n26216), .C(index_q[7]), .Z(n26221)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n26220_bdd_3_lut.init = 16'hcaca;
    PFUMX i20336 (.BLUT(n221_adj_2563), .ALUT(n22041), .C0(index_i[5]), 
          .Z(n22792));
    LUT4 mux_197_Mux_7_i475_3_lut_4_lut (.A(n27101), .B(index_q[2]), .C(index_q[3]), 
         .D(n27086), .Z(n475_adj_2564)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_7_i475_3_lut_4_lut.init = 16'h9f90;
    LUT4 n254_bdd_4_lut_adj_84 (.A(index_i[5]), .B(index_i[3]), .C(index_i[6]), 
         .D(index_i[4]), .Z(n26223)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;
    defparam n254_bdd_4_lut_adj_84.init = 16'hf8f0;
    PFUMX i20337 (.BLUT(n286_adj_2565), .ALUT(n317_adj_2566), .C0(index_i[5]), 
          .Z(n22793));
    PFUMX i21016 (.BLUT(n716_adj_2567), .ALUT(n731_adj_2348), .C0(index_i[4]), 
          .Z(n23472));
    LUT4 mux_197_Mux_6_i891_3_lut (.A(n78), .B(n890_adj_2311), .C(index_q[4]), 
         .Z(n891_adj_2568)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_6_i891_3_lut.init = 16'hcaca;
    PFUMX i24609 (.BLUT(n26563), .ALUT(n26562), .C0(index_q[8]), .Z(n26564));
    LUT4 mux_197_Mux_7_i653_3_lut_4_lut (.A(n27101), .B(index_q[2]), .C(index_q[3]), 
         .D(n27088), .Z(n653_adj_2569)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_7_i653_3_lut_4_lut.init = 16'hf606;
    PFUMX i20338 (.BLUT(n349_adj_2570), .ALUT(n22044), .C0(index_i[5]), 
          .Z(n22794));
    LUT4 i19302_4_lut_4_lut_4_lut (.A(n27101), .B(index_q[2]), .C(index_q[4]), 
         .D(index_q[3]), .Z(n21739)) /* synthesis lut_function=(A (B)+!A !(B (C+(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19302_4_lut_4_lut_4_lut.init = 16'h999c;
    LUT4 mux_197_Mux_0_i796_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n796)) /* synthesis lut_function=(A (B (C+(D))+!B (C (D)))+!A !(B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i796_3_lut_4_lut_4_lut.init = 16'hadc0;
    PFUMX i20339 (.BLUT(n413_adj_2571), .ALUT(n22047), .C0(index_i[5]), 
          .Z(n22795));
    LUT4 n26228_bdd_3_lut (.A(n27199), .B(n26224), .C(index_i[7]), .Z(n26229)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n26228_bdd_3_lut.init = 16'hcaca;
    PFUMX i20340 (.BLUT(n22050), .ALUT(n507_adj_2572), .C0(index_i[5]), 
          .Z(n22796));
    LUT4 mux_197_Mux_6_i828_4_lut (.A(n812), .B(n13909), .C(index_q[4]), 
         .D(index_q[2]), .Z(n828_adj_2573)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_6_i828_4_lut.init = 16'hfaca;
    LUT4 mux_197_Mux_6_i797_3_lut (.A(n653_adj_2464), .B(n26719), .C(index_q[4]), 
         .Z(n797_adj_2574)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_6_i797_3_lut.init = 16'hcaca;
    PFUMX i20341 (.BLUT(n22053), .ALUT(n573), .C0(index_i[5]), .Z(n22797));
    PFUMX i20342 (.BLUT(n605_adj_2575), .ALUT(n22056), .C0(index_i[5]), 
          .Z(n22798));
    PFUMX i20343 (.BLUT(n669_adj_2576), .ALUT(n700_adj_2470), .C0(index_i[5]), 
          .Z(n22799));
    LUT4 mux_197_Mux_6_i669_3_lut (.A(n653_adj_2253), .B(n668_adj_2254), 
         .C(index_q[4]), .Z(n669_adj_2577)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_6_i669_3_lut.init = 16'hcaca;
    PFUMX i20344 (.BLUT(n732_adj_2578), .ALUT(n763_adj_2579), .C0(index_i[5]), 
          .Z(n22800));
    L6MUX21 i22940 (.D0(n24624), .D1(n26700), .SD(index_i[6]), .Z(n24625));
    PFUMX i21017 (.BLUT(n747_adj_2580), .ALUT(n762_adj_2351), .C0(index_i[4]), 
          .Z(n23473));
    PFUMX i22938 (.BLUT(n24623), .ALUT(n24622), .C0(index_i[5]), .Z(n24624));
    L6MUX21 i20346 (.D0(n860_adj_2266), .D1(n891), .SD(index_i[5]), .Z(n22802));
    PFUMX i24606 (.BLUT(n26560), .ALUT(n22624), .C0(index_q[8]), .Z(n26561));
    PFUMX i19559 (.BLUT(n21994), .ALUT(n21995), .C0(index_i[4]), .Z(n476));
    CCU2D add_377_9 (.A0(quarter_wave_sample_register_q[8]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_q[9]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17574), .COUT(n17575), 
          .S0(o_val_pipeline_q_0__15__N_2189[8]), .S1(o_val_pipeline_q_0__15__N_2189[9]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(80[29:60])
    defparam add_377_9.INIT0 = 16'hf555;
    defparam add_377_9.INIT1 = 16'hf555;
    defparam add_377_9.INJECT1_0 = "NO";
    defparam add_377_9.INJECT1_1 = "NO";
    LUT4 mux_197_Mux_6_i542_3_lut (.A(n812_adj_2581), .B(n541_adj_2424), 
         .C(index_q[4]), .Z(n542_adj_2582)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_6_i542_3_lut.init = 16'hcaca;
    PFUMX mux_197_Mux_8_i574 (.BLUT(n542_adj_2344), .ALUT(n12119), .C0(index_q[5]), 
          .Z(n574)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 mux_197_Mux_6_i252_4_lut (.A(index_q[2]), .B(n251_adj_2371), .C(index_q[4]), 
         .D(n11119), .Z(n252_adj_2583)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_6_i252_4_lut.init = 16'hc5ca;
    LUT4 i20607_3_lut (.A(n1001), .B(n27061), .C(index_q[3]), .Z(n23063)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20607_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_2_i452_3_lut_3_lut_rep_763 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n27086)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_2_i452_3_lut_3_lut_rep_763.init = 16'hc7c7;
    LUT4 i22175_3_lut (.A(n25900), .B(n252_adj_2583), .C(index_q[5]), 
         .Z(n22471)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22175_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_4_lut (.A(n26737), .B(index_q[5]), .C(index_q[8]), .D(n19798), 
         .Z(n20197)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_3_lut_4_lut.init = 16'hfff8;
    PFUMX i20365 (.BLUT(n94_adj_2584), .ALUT(n22062), .C0(index_i[5]), 
          .Z(n22821));
    L6MUX21 i20366 (.D0(n22065), .D1(n22068), .SD(index_i[5]), .Z(n22822));
    PFUMX i20368 (.BLUT(n22071), .ALUT(n317_adj_2585), .C0(index_i[5]), 
          .Z(n22824));
    LUT4 i15573_4_lut (.A(index_i[0]), .B(index_i[4]), .C(index_i[1]), 
         .D(n26898), .Z(n286_adj_2586)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i15573_4_lut.init = 16'hccc8;
    LUT4 n21568_bdd_3_lut (.A(n26716), .B(n701), .C(index_i[6]), .Z(n26246)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n21568_bdd_3_lut.init = 16'hacac;
    PFUMX i20369 (.BLUT(n349_adj_2587), .ALUT(n22074), .C0(index_i[5]), 
          .Z(n22825));
    L6MUX21 i20370 (.D0(n22077), .D1(n22080), .SD(index_i[5]), .Z(n22826));
    L6MUX21 i20371 (.D0(n22083), .D1(n22086), .SD(index_i[5]), .Z(n22827));
    LUT4 n26249_bdd_3_lut (.A(n28559), .B(n23334), .C(index_i[8]), .Z(n26250)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n26249_bdd_3_lut.init = 16'hcaca;
    CCU2D add_377_7 (.A0(quarter_wave_sample_register_q[6]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_q[7]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17573), .COUT(n17574), 
          .S1(o_val_pipeline_q_0__15__N_2189[7]));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(80[29:60])
    defparam add_377_7.INIT0 = 16'hf555;
    defparam add_377_7.INIT1 = 16'hf555;
    defparam add_377_7.INJECT1_0 = "NO";
    defparam add_377_7.INJECT1_1 = "NO";
    L6MUX21 i20373 (.D0(n22092), .D1(n636), .SD(index_i[5]), .Z(n22829));
    LUT4 n21577_bdd_3_lut (.A(n26717), .B(n701_adj_2588), .C(index_q[6]), 
         .Z(n26261)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n21577_bdd_3_lut.init = 16'hacac;
    PFUMX i20374 (.BLUT(n22095), .ALUT(n700_adj_2345), .C0(index_i[5]), 
          .Z(n22830));
    LUT4 n26264_bdd_3_lut (.A(n28537), .B(n23181), .C(index_q[8]), .Z(n26265)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n26264_bdd_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_1_i620_3_lut_4_lut (.A(n27092), .B(index_q[1]), .C(index_q[3]), 
         .D(n27082), .Z(n620_adj_2548)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_1_i620_3_lut_4_lut.init = 16'hdfd0;
    L6MUX21 i20376 (.D0(n22098), .D1(n22101), .SD(index_i[5]), .Z(n22832));
    PFUMX i20378 (.BLUT(n924_adj_2589), .ALUT(n22107), .C0(index_i[5]), 
          .Z(n22834));
    LUT4 i19549_3_lut_4_lut (.A(n27092), .B(index_q[1]), .C(index_q[3]), 
         .D(n498), .Z(n21986)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19549_3_lut_4_lut.init = 16'hdfd0;
    LUT4 mux_197_Mux_7_i892_3_lut (.A(n62_adj_2590), .B(n891_adj_2277), 
         .C(index_q[5]), .Z(n892_adj_2312)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_7_i892_3_lut.init = 16'hcaca;
    LUT4 i19309_3_lut (.A(n747_adj_2591), .B(n908_adj_2592), .C(index_q[4]), 
         .Z(n21746)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19309_3_lut.init = 16'hcaca;
    LUT4 i19308_3_lut (.A(n716_adj_2416), .B(n14928), .C(index_q[4]), 
         .Z(n21745)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19308_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_0_i173_3_lut_4_lut (.A(n27092), .B(index_q[1]), .C(index_q[3]), 
         .D(n27080), .Z(n173_adj_2593)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i173_3_lut_4_lut.init = 16'hdfd0;
    LUT4 i20864_3_lut_4_lut (.A(n26766), .B(n26770), .C(index_i[5]), .D(index_i[6]), 
         .Z(n23320)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (B+((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20864_3_lut_4_lut.init = 16'hffc5;
    LUT4 i19306_3_lut (.A(n93_adj_2594), .B(n699_adj_2313), .C(index_q[4]), 
         .Z(n21743)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19306_3_lut.init = 16'hcaca;
    PFUMX i20379 (.BLUT(n987), .ALUT(n22110), .C0(index_i[5]), .Z(n22835));
    LUT4 i19305_3_lut (.A(n653_adj_2569), .B(n26747), .C(index_q[4]), 
         .Z(n21742)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19305_3_lut.init = 16'hcaca;
    LUT4 i19299_3_lut (.A(n526_adj_2595), .B(n15_adj_2413), .C(index_q[4]), 
         .Z(n21736)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19299_3_lut.init = 16'hcaca;
    PFUMX i19577 (.BLUT(n22012), .ALUT(n22013), .C0(index_i[4]), .Z(n22014));
    LUT4 i19296_3_lut (.A(n397_adj_2596), .B(n475_adj_2564), .C(index_q[4]), 
         .Z(n21733)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19296_3_lut.init = 16'hcaca;
    PFUMX i21018 (.BLUT(n781_adj_2597), .ALUT(n796_adj_2368), .C0(index_i[4]), 
          .Z(n23474));
    LUT4 i19294_3_lut (.A(n348_adj_2598), .B(n443_adj_2599), .C(index_q[4]), 
         .Z(n21731)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19294_3_lut.init = 16'hcaca;
    LUT4 i19293_3_lut (.A(n397_adj_2596), .B(n781_adj_2600), .C(index_q[4]), 
         .Z(n21730)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19293_3_lut.init = 16'hcaca;
    LUT4 n22745_bdd_3_lut_24404 (.A(n22745), .B(n24869), .C(index_i[7]), 
         .Z(n26296)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n22745_bdd_3_lut_24404.init = 16'hcaca;
    LUT4 i19291_3_lut (.A(n364_adj_2362), .B(n890_adj_2376), .C(index_q[4]), 
         .Z(n21728)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19291_3_lut.init = 16'hcaca;
    PFUMX i21019 (.BLUT(n812_adj_2360), .ALUT(n12109), .C0(index_i[4]), 
          .Z(n23475));
    LUT4 i19290_3_lut (.A(n333_adj_2601), .B(n348_adj_2598), .C(index_q[4]), 
         .Z(n21727)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19290_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_3_i251_3_lut_4_lut (.A(n27101), .B(index_q[2]), .C(index_q[3]), 
         .D(n26893), .Z(n14814)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_3_i251_3_lut_4_lut.init = 16'h8f80;
    LUT4 n22747_bdd_3_lut (.A(n22747), .B(n22748), .C(index_i[7]), .Z(n26294)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n22747_bdd_3_lut.init = 16'hcaca;
    PFUMX i20811 (.BLUT(n23251), .ALUT(n23252), .C0(index_q[5]), .Z(n23267));
    CCU2D add_377_5 (.A0(quarter_wave_sample_register_q[4]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_q[5]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17572), .COUT(n17573));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(80[29:60])
    defparam add_377_5.INIT0 = 16'hf555;
    defparam add_377_5.INIT1 = 16'hf555;
    defparam add_377_5.INJECT1_0 = "NO";
    defparam add_377_5.INJECT1_1 = "NO";
    LUT4 index_q_0__bdd_4_lut_24742 (.A(index_q[0]), .B(index_q[3]), .C(index_q[1]), 
         .D(index_q[2]), .Z(n27122)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C))+!A (B (C (D)+!C !(D))+!B !(C+!(D))))) */ ;
    defparam index_q_0__bdd_4_lut_24742.init = 16'h16d3;
    LUT4 index_q_1__bdd_4_lut_24774 (.A(index_q[1]), .B(index_q[0]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n27174)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A !(B ((D)+!C)+!B (D))) */ ;
    defparam index_q_1__bdd_4_lut_24774.init = 16'h8a51;
    LUT4 mux_197_Mux_6_i939_3_lut_rep_397_3_lut_4_lut (.A(n27101), .B(index_q[2]), 
         .C(index_q[3]), .D(n26871), .Z(n26720)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_6_i939_3_lut_rep_397_3_lut_4_lut.init = 16'h08f8;
    LUT4 n22745_bdd_3_lut (.A(n22744), .B(n22743), .C(index_i[7]), .Z(n26297)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n22745_bdd_3_lut.init = 16'hacac;
    PFUMX i24767 (.BLUT(n27182), .ALUT(n27183), .C0(index_q[1]), .Z(n27184));
    PFUMX i20812 (.BLUT(n23253), .ALUT(n23254), .C0(index_q[5]), .Z(n23268));
    LUT4 mux_196_Mux_0_i188_3_lut (.A(n27002), .B(n931_adj_2602), .C(index_i[3]), 
         .Z(n188_adj_2603)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_0_i188_3_lut.init = 16'hcaca;
    PFUMX i24562 (.BLUT(n26513), .ALUT(n26512), .C0(index_q[4]), .Z(n26514));
    LUT4 i21784_3_lut (.A(n716_adj_2411), .B(n731_adj_2604), .C(index_q[4]), 
         .Z(n732_adj_2605)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21784_3_lut.init = 16'hcaca;
    LUT4 i22707_2_lut_rep_410_3_lut_4_lut (.A(n27101), .B(index_q[2]), .C(index_q[5]), 
         .D(n26967), .Z(n26733)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i22707_2_lut_rep_410_3_lut_4_lut.init = 16'h0f7f;
    LUT4 i11251_3_lut (.A(index_q[3]), .B(index_q[1]), .C(index_q[0]), 
         .Z(n13925)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11251_3_lut.init = 16'hecec;
    LUT4 mux_197_Mux_8_i78_3_lut_4_lut (.A(n27101), .B(index_q[2]), .C(index_q[3]), 
         .D(n27088), .Z(n78)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_8_i78_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_197_Mux_2_i669_3_lut (.A(n653_adj_2606), .B(n475_adj_2377), 
         .C(index_q[4]), .Z(n669_adj_2607)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_2_i669_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_5_i939_3_lut_3_lut_4_lut (.A(n27101), .B(index_q[2]), 
         .C(n954_adj_2608), .D(index_q[4]), .Z(n939_adj_2296)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_5_i939_3_lut_3_lut_4_lut.init = 16'hf077;
    LUT4 mux_197_Mux_9_i364_3_lut_3_lut_4_lut (.A(n27101), .B(index_q[2]), 
         .C(n26893), .D(index_q[3]), .Z(n364)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_9_i364_3_lut_3_lut_4_lut.init = 16'h77f0;
    L6MUX21 i20813 (.D0(n23255), .D1(n23256), .SD(index_q[5]), .Z(n23269));
    LUT4 mux_197_Mux_2_i605_3_lut (.A(n142_adj_2436), .B(n604_adj_2609), 
         .C(index_q[4]), .Z(n605_adj_2610)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_2_i605_3_lut.init = 16'hcaca;
    LUT4 i21791_3_lut (.A(n27141), .B(n21479), .C(index_q[4]), .Z(n21480)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21791_3_lut.init = 16'hcaca;
    PFUMX i20814 (.BLUT(n23257), .ALUT(n23258), .C0(index_q[5]), .Z(n23270));
    LUT4 i21711_3_lut (.A(n27193), .B(n22133), .C(index_q[4]), .Z(n22134)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21711_3_lut.init = 16'hcaca;
    LUT4 i21795_3_lut (.A(n21475), .B(n21476), .C(index_q[4]), .Z(n21477)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21795_3_lut.init = 16'hcaca;
    PFUMX i19592 (.BLUT(n22027), .ALUT(n22028), .C0(index_i[4]), .Z(n22029));
    LUT4 mux_197_Mux_2_i413_3_lut (.A(n397_adj_2611), .B(n954_adj_2608), 
         .C(index_q[4]), .Z(n413_adj_2612)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_2_i413_3_lut.init = 16'hcaca;
    LUT4 i20258_3_lut (.A(n25736), .B(n23060), .C(index_q[6]), .Z(n22714)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20258_3_lut.init = 16'hcaca;
    L6MUX21 i20816 (.D0(n23261), .D1(n23262), .SD(index_q[5]), .Z(n23272));
    LUT4 i22045_3_lut (.A(n27192), .B(n124_adj_2613), .C(index_i[4]), 
         .Z(n23192)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22045_3_lut.init = 16'hcaca;
    LUT4 i22678_2_lut (.A(index_i[3]), .B(index_i[2]), .Z(n22374)) /* synthesis lut_function=(A+!(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i22678_2_lut.init = 16'hbbbb;
    LUT4 mux_197_Mux_2_i317_3_lut (.A(n668_adj_2428), .B(n316_adj_2614), 
         .C(index_q[4]), .Z(n317_adj_2615)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_2_i317_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_2_i286_3_lut (.A(n270_adj_2616), .B(n653_adj_2268), 
         .C(index_q[4]), .Z(n286_adj_2617)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_2_i286_3_lut.init = 16'hcaca;
    LUT4 i19329_3_lut_3_lut_4_lut (.A(n27101), .B(index_q[2]), .C(n1001), 
         .D(index_q[3]), .Z(n21766)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19329_3_lut_3_lut_4_lut.init = 16'hf077;
    L6MUX21 i20817 (.D0(n23263), .D1(n23264), .SD(index_q[5]), .Z(n23273));
    LUT4 n572_bdd_3_lut_24262_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n26011)) /* synthesis lut_function=(A (B (C+(D)))+!A (B ((D)+!C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n572_bdd_3_lut_24262_4_lut.init = 16'hcc94;
    LUT4 i21805_3_lut (.A(n142_adj_2412), .B(n13947), .C(index_q[4]), 
         .Z(n158_adj_2618)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21805_3_lut.init = 16'hcaca;
    LUT4 i11449_2_lut_rep_390_3_lut_4_lut (.A(n26767), .B(index_q[4]), .C(index_q[6]), 
         .D(index_q[5]), .Z(n26713)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11449_2_lut_rep_390_3_lut_4_lut.init = 16'hf080;
    L6MUX21 i20818 (.D0(n23265), .D1(n23266), .SD(index_q[5]), .Z(n23274));
    LUT4 i19562_then_4_lut (.A(index_i[2]), .B(index_i[1]), .C(index_i[4]), 
         .D(index_i[3]), .Z(n27176)) /* synthesis lut_function=(A (B (C+(D))+!B !(C))+!A !(B (C+(D))+!B !(C+!(D)))) */ ;
    defparam i19562_then_4_lut.init = 16'h9a97;
    LUT4 mux_197_Mux_1_i986_3_lut (.A(n27102), .B(n27081), .C(index_q[3]), 
         .Z(n986_adj_2619)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_1_i986_3_lut.init = 16'hcaca;
    L6MUX21 i20827 (.D0(n21933), .D1(n21936), .SD(index_i[5]), .Z(n23283));
    LUT4 mux_197_Mux_3_i700_3_lut_4_lut (.A(index_q[4]), .B(index_q[3]), 
         .C(n684_adj_2620), .D(n27094), .Z(n700_adj_2621)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_3_i700_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i20263_3_lut_4_lut (.A(n26768), .B(n26769), .C(index_q[5]), .D(index_q[6]), 
         .Z(n22719)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (B+((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20263_3_lut_4_lut.init = 16'hffc5;
    LUT4 i19678_3_lut (.A(n27102), .B(n851), .C(index_q[3]), .Z(n22115)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19678_3_lut.init = 16'hcaca;
    PFUMX mux_197_Mux_2_i891 (.BLUT(n875_adj_2622), .ALUT(n890_adj_2623), 
          .C0(index_q[4]), .Z(n891_adj_2624)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 i19677_3_lut (.A(n27078), .B(n27062), .C(index_q[3]), .Z(n22114)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19677_3_lut.init = 16'hcaca;
    LUT4 i12392_2_lut_3_lut_4_lut (.A(n26772), .B(index_q[4]), .C(index_q[6]), 
         .D(index_q[5]), .Z(n15088)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12392_2_lut_3_lut_4_lut.init = 16'hfef0;
    LUT4 i19675_3_lut (.A(n27102), .B(n26887), .C(index_q[3]), .Z(n22112)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19675_3_lut.init = 16'hcaca;
    LUT4 i19674_3_lut (.A(n27105), .B(n851), .C(index_q[3]), .Z(n22111)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19674_3_lut.init = 16'hcaca;
    PFUMX mux_197_Mux_2_i860 (.BLUT(n844_adj_2625), .ALUT(n859_adj_2626), 
          .C0(index_q[4]), .Z(n860_adj_2627)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 i19539_3_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[0]), 
         .D(index_i[3]), .Z(n21976)) /* synthesis lut_function=(A (B (C (D))+!B !(C (D)+!C !(D)))+!A (B (C)+!B !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19539_3_lut_4_lut_4_lut.init = 16'hc371;
    LUT4 i20758_3_lut (.A(n23207), .B(n28254), .C(index_i[6]), .Z(n23214)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20758_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_7_i173_3_lut (.A(n27078), .B(n26887), .C(index_q[3]), 
         .Z(n173_adj_2493)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_7_i173_3_lut.init = 16'hcaca;
    LUT4 i20759_3_lut (.A(n25495), .B(n23210), .C(index_i[6]), .Z(n23215)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20759_3_lut.init = 16'hcaca;
    LUT4 i19671_3_lut (.A(n26977), .B(n27029), .C(index_i[3]), .Z(n22108)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19671_3_lut.init = 16'hcaca;
    PFUMX i20409 (.BLUT(n956_adj_2628), .ALUT(n20333), .C0(index_q[6]), 
          .Z(n22865));
    LUT4 i21925_3_lut (.A(n22108), .B(n22109), .C(index_i[4]), .Z(n22110)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21925_3_lut.init = 16'hcaca;
    LUT4 i19282_3_lut (.A(n491_adj_2629), .B(n541), .C(index_q[4]), .Z(n21719)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19282_3_lut.init = 16'hcaca;
    PFUMX i19220 (.BLUT(n21655), .ALUT(n21656), .C0(index_i[5]), .Z(n21657));
    LUT4 i19281_3_lut (.A(n397), .B(n475_adj_2630), .C(index_q[4]), .Z(n21718)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19281_3_lut.init = 16'hcaca;
    LUT4 n25213_bdd_3_lut_24446 (.A(n22474), .B(n25238), .C(index_q[6]), 
         .Z(n26351)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n25213_bdd_3_lut_24446.init = 16'hcaca;
    LUT4 i19668_3_lut (.A(n38), .B(n773), .C(index_i[3]), .Z(n22105)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19668_3_lut.init = 16'hcaca;
    LUT4 i21928_3_lut (.A(n22105), .B(n22106), .C(index_i[4]), .Z(n22107)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21928_3_lut.init = 16'hcaca;
    L6MUX21 i20831 (.D0(n21942), .D1(n17813), .SD(index_i[5]), .Z(n23287));
    PFUMX i19223 (.BLUT(n21658), .ALUT(n21659), .C0(index_i[5]), .Z(n21660));
    LUT4 i19279_3_lut (.A(n251_adj_2314), .B(n443_adj_2309), .C(index_q[4]), 
         .Z(n21716)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19279_3_lut.init = 16'hcaca;
    LUT4 i19278_3_lut (.A(n397), .B(n14928), .C(index_q[4]), .Z(n21715)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;
    defparam i19278_3_lut.init = 16'h3a3a;
    L6MUX21 i20832 (.D0(n21945), .D1(n12055), .SD(index_i[5]), .Z(n23288));
    LUT4 i19660_3_lut (.A(n27025), .B(n26934), .C(index_i[3]), .Z(n22097)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19660_3_lut.init = 16'hcaca;
    PFUMX i20834 (.BLUT(n542_adj_2631), .ALUT(n573_adj_2632), .C0(index_i[5]), 
          .Z(n23290));
    LUT4 mux_197_Mux_3_i781_3_lut (.A(n27062), .B(n27058), .C(index_q[3]), 
         .Z(n781_adj_2600)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_3_i781_3_lut.init = 16'hcaca;
    PFUMX i20835 (.BLUT(n605), .ALUT(n636_adj_2633), .C0(index_i[5]), 
          .Z(n23291));
    LUT4 n25213_bdd_3_lut_25670 (.A(n25213), .B(n22473), .C(index_q[6]), 
         .Z(n26352)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n25213_bdd_3_lut_25670.init = 16'hcaca;
    PFUMX i20836 (.BLUT(n669_adj_2634), .ALUT(n700_adj_2635), .C0(index_i[5]), 
          .Z(n23292));
    LUT4 mux_197_Mux_10_i574_4_lut_4_lut (.A(n26772), .B(index_q[4]), .C(index_q[5]), 
         .D(n26753), .Z(n574_adj_2401)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_10_i574_4_lut_4_lut.init = 16'h1f1c;
    LUT4 i19512_3_lut_3_lut_4_lut (.A(index_i[2]), .B(n26996), .C(n26928), 
         .D(index_i[3]), .Z(n21949)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (B (C (D))+!B (C+!(D)))) */ ;
    defparam i19512_3_lut_3_lut_4_lut.init = 16'hf099;
    LUT4 i19645_3_lut (.A(n29470), .B(n27023), .C(index_i[3]), .Z(n22082)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19645_3_lut.init = 16'hcaca;
    LUT4 n476_bdd_3_lut_23143_4_lut (.A(index_i[2]), .B(n26996), .C(index_i[4]), 
         .D(n491_adj_2636), .Z(n24864)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+(D)))) */ ;
    defparam n476_bdd_3_lut_23143_4_lut.init = 16'h9f90;
    LUT4 i19587_3_lut_3_lut_4_lut (.A(index_i[2]), .B(n26996), .C(n26900), 
         .D(index_i[3]), .Z(n22024)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (B (C (D))+!B (C+!(D)))) */ ;
    defparam i19587_3_lut_3_lut_4_lut.init = 16'hf099;
    LUT4 i19638_3_lut (.A(n27025), .B(n29471), .C(index_i[3]), .Z(n22075)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19638_3_lut.init = 16'hcaca;
    PFUMX i20837 (.BLUT(n732_adj_2637), .ALUT(n21951), .C0(index_i[5]), 
          .Z(n23293));
    LUT4 n25449_bdd_3_lut (.A(n25449), .B(n22469), .C(index_q[6]), .Z(n26354)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n25449_bdd_3_lut.init = 16'hcaca;
    PFUMX i20838 (.BLUT(n797_adj_2638), .ALUT(n828_adj_2639), .C0(index_i[5]), 
          .Z(n23294));
    LUT4 i21938_3_lut (.A(n22072), .B(n22073), .C(index_i[4]), .Z(n22074)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21938_3_lut.init = 16'hcaca;
    PFUMX i20839 (.BLUT(n860), .ALUT(n891_adj_2640), .C0(index_i[5]), 
          .Z(n23295));
    LUT4 mux_197_Mux_5_i731_3_lut (.A(n29473), .B(n29474), .C(index_q[3]), 
         .Z(n731_adj_2641)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_5_i731_3_lut.init = 16'hcaca;
    LUT4 i22310_3_lut (.A(n27188), .B(n27191), .C(index_q[5]), .Z(n21711)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22310_3_lut.init = 16'hcaca;
    LUT4 n25096_bdd_3_lut (.A(n25096), .B(n476_adj_2423), .C(index_q[5]), 
         .Z(n25097)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n25096_bdd_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_6_i653_3_lut (.A(n26933), .B(n619), .C(index_i[3]), 
         .Z(n653_adj_2642)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_6_i653_3_lut.init = 16'hcaca;
    LUT4 i19269_3_lut (.A(n78), .B(n93_adj_2594), .C(index_q[4]), .Z(n21706)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19269_3_lut.init = 16'hcaca;
    LUT4 i12368_2_lut_3_lut_4_lut (.A(n26775), .B(index_i[4]), .C(index_i[6]), 
         .D(index_i[5]), .Z(n15064)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i12368_2_lut_3_lut_4_lut.init = 16'hfef0;
    LUT4 mux_196_Mux_5_i397_3_lut (.A(n26993), .B(n204), .C(index_i[3]), 
         .Z(n397_adj_2643)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_5_i397_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_10_i574_4_lut_4_lut (.A(n26775), .B(index_i[4]), .C(index_i[5]), 
         .D(n26759), .Z(n574_adj_2403)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_10_i574_4_lut_4_lut.init = 16'h1f1c;
    LUT4 mux_196_Mux_0_i986_3_lut (.A(n27027), .B(n985_adj_2644), .C(index_i[3]), 
         .Z(n986_adj_2645)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_0_i986_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_0_i971_3_lut (.A(n27028), .B(n27000), .C(index_i[3]), 
         .Z(n971_adj_2646)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_0_i971_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_3_i860_3_lut_4_lut (.A(index_i[2]), .B(n26996), .C(index_i[4]), 
         .D(n859_adj_2647), .Z(n860_adj_2546)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam mux_196_Mux_3_i860_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_197_Mux_0_i676_3_lut_4_lut_3_lut_rep_764 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n27087)) /* synthesis lut_function=(A (B)+!A !(B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i676_3_lut_4_lut_3_lut_rep_764.init = 16'h9898;
    LUT4 i19266_3_lut (.A(n15), .B(n526_adj_2417), .C(index_q[4]), .Z(n21703)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19266_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_1_i317_3_lut (.A(n301_adj_2648), .B(n908_adj_2358), 
         .C(index_i[4]), .Z(n317_adj_2585)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_1_i317_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_5_i506_3_lut (.A(n26977), .B(n29470), .C(index_i[3]), 
         .Z(n506_adj_2649)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_5_i506_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_0_i939_4_lut (.A(n773), .B(n26848), .C(index_i[3]), 
         .D(index_i[2]), .Z(n939_adj_2650)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_0_i939_4_lut.init = 16'hfaca;
    LUT4 mux_196_Mux_7_i892_3_lut (.A(n62), .B(n891_adj_2292), .C(index_i[5]), 
         .Z(n892)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_7_i892_3_lut.init = 16'hcaca;
    PFUMX i24503 (.BLUT(n26416), .ALUT(n29485), .C0(index_q[3]), .Z(n26417));
    LUT4 mux_196_Mux_0_i923_3_lut (.A(n26928), .B(n26999), .C(index_i[3]), 
         .Z(n923_adj_2651)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_0_i923_3_lut.init = 16'hcaca;
    LUT4 i19261_3_lut (.A(n747_adj_2297), .B(n762_adj_2298), .C(index_i[4]), 
         .Z(n21698)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19261_3_lut.init = 16'hcaca;
    LUT4 i19260_3_lut (.A(n716_adj_2267), .B(n14858), .C(index_i[4]), 
         .Z(n21697)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19260_3_lut.init = 16'hcaca;
    LUT4 i19258_3_lut (.A(n93_adj_2652), .B(n699_adj_2336), .C(index_i[4]), 
         .Z(n21695)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19258_3_lut.init = 16'hcaca;
    LUT4 i19257_3_lut (.A(n653_adj_2385), .B(n26748), .C(index_i[4]), 
         .Z(n21694)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19257_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_7_i443_3_lut_4_lut (.A(index_i[2]), .B(n26996), .C(index_i[3]), 
         .D(n26928), .Z(n443_adj_2653)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;
    defparam mux_196_Mux_7_i443_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_196_Mux_0_i30_3_lut (.A(n29492), .B(n27003), .C(index_i[3]), 
         .Z(n30_adj_2654)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_0_i30_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_4_i158_3_lut (.A(n142_adj_2655), .B(n157_adj_2499), 
         .C(index_q[4]), .Z(n158_adj_2656)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_4_i158_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_5_i15_3_lut (.A(n26932), .B(n29472), .C(index_i[3]), 
         .Z(n15_adj_2471)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_5_i15_3_lut.init = 16'hcaca;
    PFUMX i24765 (.BLUT(n27178), .ALUT(n27179), .C0(index_q[0]), .Z(n27180));
    LUT4 mux_196_Mux_5_i859_3_lut (.A(n308), .B(n26932), .C(index_i[3]), 
         .Z(n859_adj_2657)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_5_i859_3_lut.init = 16'hcaca;
    PFUMX i19232 (.BLUT(n21667), .ALUT(n21668), .C0(index_i[5]), .Z(n21669));
    CCU2D add_377_3 (.A0(quarter_wave_sample_register_q[2]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(quarter_wave_sample_register_q[3]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n17571), .COUT(n17572));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(80[29:60])
    defparam add_377_3.INIT0 = 16'hf555;
    defparam add_377_3.INIT1 = 16'hf555;
    defparam add_377_3.INJECT1_0 = "NO";
    defparam add_377_3.INJECT1_1 = "NO";
    LUT4 mux_196_Mux_5_i875_3_lut (.A(n26900), .B(n29491), .C(index_i[3]), 
         .Z(n875_adj_2658)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_5_i875_3_lut.init = 16'hcaca;
    PFUMX i19235 (.BLUT(n21670), .ALUT(n21671), .C0(index_i[5]), .Z(n21672));
    LUT4 i19626_3_lut (.A(n723), .B(n26934), .C(index_i[3]), .Z(n22063)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19626_3_lut.init = 16'hcaca;
    LUT4 i21945_3_lut (.A(n27185), .B(n22061), .C(index_i[4]), .Z(n22062)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21945_3_lut.init = 16'hcaca;
    LUT4 i19251_3_lut (.A(n526_adj_2659), .B(n541_adj_2660), .C(index_i[4]), 
         .Z(n21688)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19251_3_lut.init = 16'hcaca;
    LUT4 i19479_3_lut_3_lut_4_lut (.A(n27085), .B(index_q[2]), .C(n27062), 
         .D(index_q[3]), .Z(n21916)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (B (C (D))+!B (C+!(D)))) */ ;
    defparam i19479_3_lut_3_lut_4_lut.init = 16'hf099;
    LUT4 i19014_3_lut_3_lut_4_lut (.A(n27085), .B(index_q[2]), .C(n26887), 
         .D(index_q[3]), .Z(n21451)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (B (C (D))+!B (C+!(D)))) */ ;
    defparam i19014_3_lut_3_lut_4_lut.init = 16'hf099;
    LUT4 mux_197_Mux_2_i653_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n653_adj_2606)) /* synthesis lut_function=(A (B (C+!(D))+!B !(D))+!A !(B (C+!(D))+!B !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_2_i653_3_lut_4_lut.init = 16'h94aa;
    LUT4 i20722_3_lut_4_lut_4_lut (.A(n26817), .B(index_q[4]), .C(index_q[5]), 
         .D(n26796), .Z(n23178)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C)+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20722_3_lut_4_lut_4_lut.init = 16'h0434;
    LUT4 i19562_else_4_lut (.A(index_i[2]), .B(index_i[1]), .C(index_i[4]), 
         .D(index_i[3]), .Z(n27175)) /* synthesis lut_function=(!(A (B (C)+!B (C+(D)))+!A !(B (C (D)+!C !(D))+!B (C+!(D))))) */ ;
    defparam i19562_else_4_lut.init = 16'h581f;
    LUT4 i19248_3_lut (.A(n397_adj_2661), .B(n475_adj_2384), .C(index_i[4]), 
         .Z(n21685)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19248_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_8_i892_3_lut_4_lut (.A(n26817), .B(index_q[4]), .C(index_q[5]), 
         .D(n860_adj_2662), .Z(n892_adj_2663)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_8_i892_3_lut_4_lut.init = 16'h4f40;
    LUT4 n476_bdd_3_lut_23642_4_lut (.A(n27085), .B(index_q[2]), .C(index_q[4]), 
         .D(n491_adj_2664), .Z(n25408)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+(D)))) */ ;
    defparam n476_bdd_3_lut_23642_4_lut.init = 16'h9f90;
    LUT4 mux_197_Mux_3_i860_3_lut_4_lut (.A(n27085), .B(index_q[2]), .C(index_q[4]), 
         .D(n859_adj_2665), .Z(n860_adj_2666)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam mux_197_Mux_3_i860_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_197_Mux_6_i860_3_lut_3_lut (.A(n26747), .B(index_q[4]), .C(n844_adj_2667), 
         .Z(n860_adj_2668)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam mux_197_Mux_6_i860_3_lut_3_lut.init = 16'h7474;
    PFUMX i19238 (.BLUT(n21673), .ALUT(n21674), .C0(index_i[5]), .Z(n21675));
    LUT4 mux_197_Mux_7_i443_3_lut_4_lut (.A(n27085), .B(index_q[2]), .C(index_q[3]), 
         .D(n27062), .Z(n443_adj_2599)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;
    defparam mux_197_Mux_7_i443_3_lut_4_lut.init = 16'h6f60;
    LUT4 i19617_3_lut (.A(n404), .B(n26991), .C(index_i[3]), .Z(n22054)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19617_3_lut.init = 16'hcaca;
    LUT4 i19246_3_lut (.A(n348_adj_2669), .B(n443_adj_2653), .C(index_i[4]), 
         .Z(n21683)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19246_3_lut.init = 16'hcaca;
    LUT4 i21960_3_lut (.A(n22054), .B(n22055), .C(index_i[4]), .Z(n22056)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21960_3_lut.init = 16'hcaca;
    PFUMX i19241 (.BLUT(n21676), .ALUT(n21677), .C0(index_i[5]), .Z(n21678));
    LUT4 i19245_3_lut (.A(n397_adj_2661), .B(n731_adj_2501), .C(index_i[4]), 
         .Z(n21682)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19245_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_3_i1018_3_lut_4_lut (.A(index_q[1]), .B(n26994), .C(index_q[4]), 
         .D(n19855), .Z(n1018_adj_2670)) /* synthesis lut_function=(A (C+!(D))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_3_i1018_3_lut_4_lut.init = 16'he0ef;
    LUT4 i19243_3_lut (.A(n364_adj_2323), .B(n379_adj_2327), .C(index_i[4]), 
         .Z(n21680)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19243_3_lut.init = 16'hcaca;
    PFUMX i20442 (.BLUT(n22894), .ALUT(n22895), .C0(index_i[5]), .Z(n22898));
    LUT4 i19242_3_lut (.A(n333_adj_2671), .B(n348_adj_2669), .C(index_i[4]), 
         .Z(n21679)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19242_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_2_i700_3_lut_4_lut (.A(index_q[1]), .B(n26994), .C(index_q[4]), 
         .D(n684_adj_2560), .Z(n700_adj_2672)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_2_i700_3_lut_4_lut.init = 16'hefe0;
    LUT4 mux_197_Mux_3_i747_3_lut (.A(n27099), .B(n498), .C(index_q[3]), 
         .Z(n747_adj_2673)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_3_i747_3_lut.init = 16'hcaca;
    PFUMX i20443 (.BLUT(n22896), .ALUT(n22897), .C0(index_i[5]), .Z(n22899));
    PFUMX i24763 (.BLUT(n27175), .ALUT(n27176), .C0(index_i[0]), .Z(n27177));
    LUT4 mux_196_Mux_4_i61_3_lut (.A(n27025), .B(n26978), .C(index_i[3]), 
         .Z(n61_adj_2475)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_4_i61_3_lut.init = 16'hcaca;
    LUT4 n25100_bdd_3_lut_23416 (.A(n27184), .B(n25098), .C(index_q[5]), 
         .Z(n25101)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n25100_bdd_3_lut_23416.init = 16'hcaca;
    LUT4 i19267_3_lut_3_lut (.A(n26747), .B(index_q[4]), .C(n109_adj_2349), 
         .Z(n21704)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam i19267_3_lut_3_lut.init = 16'h7474;
    LUT4 mux_196_Mux_4_i270_3_lut (.A(n29488), .B(n26977), .C(index_i[3]), 
         .Z(n270_adj_2674)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_4_i270_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_4_i15_3_lut (.A(n29470), .B(n773), .C(index_i[3]), 
         .Z(n15_adj_2478)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_4_i15_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_4_i348_3_lut (.A(n26983), .B(n29489), .C(index_i[3]), 
         .Z(n348_adj_2675)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_4_i348_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_2_i955_then_4_lut (.A(index_q[4]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n27179)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B (C+!(D))+!B !(C (D)))) */ ;
    defparam mux_197_Mux_2_i955_then_4_lut.init = 16'he95d;
    LUT4 i19612_3_lut (.A(n404), .B(n26989), .C(index_i[3]), .Z(n22049)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19612_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_2_i955_else_4_lut (.A(index_q[4]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n27178)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+(D)))+!A !(B (C+!(D))+!B !(C+!(D))))) */ ;
    defparam mux_197_Mux_2_i955_else_4_lut.init = 16'h49c6;
    LUT4 i18993_3_lut (.A(n588), .B(n29493), .C(index_q[3]), .Z(n21430)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18993_3_lut.init = 16'hcaca;
    PFUMX i20449 (.BLUT(n22901), .ALUT(n22902), .C0(index_i[5]), .Z(n22905));
    LUT4 i11372_2_lut_rep_391_3_lut_4_lut (.A(n26781), .B(index_i[4]), .C(index_i[6]), 
         .D(index_i[5]), .Z(n26714)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11372_2_lut_rep_391_3_lut_4_lut.init = 16'hf080;
    LUT4 i20027_3_lut_4_lut_4_lut (.A(n26816), .B(index_q[5]), .C(index_q[4]), 
         .D(n26774), .Z(n22483)) /* synthesis lut_function=(A (B+(C (D)))+!A (B+((D)+!C))) */ ;
    defparam i20027_3_lut_4_lut_4_lut.init = 16'hfdcd;
    LUT4 i19234_3_lut (.A(n491_adj_2676), .B(n506), .C(index_i[4]), .Z(n21671)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19234_3_lut.init = 16'hcaca;
    LUT4 i19233_3_lut (.A(n397_adj_2392), .B(n475_adj_2491), .C(index_i[4]), 
         .Z(n21670)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19233_3_lut.init = 16'hcaca;
    LUT4 i19231_3_lut (.A(n251_adj_2306), .B(n443_adj_2308), .C(index_i[4]), 
         .Z(n21668)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19231_3_lut.init = 16'hcaca;
    LUT4 i19230_3_lut (.A(n397_adj_2392), .B(n14858), .C(index_i[4]), 
         .Z(n21667)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;
    defparam i19230_3_lut.init = 16'h3a3a;
    PFUMX i23366 (.BLUT(n25101), .ALUT(n25097), .C0(index_q[6]), .Z(n25102));
    PFUMX i21021 (.BLUT(n875_adj_2677), .ALUT(n890_adj_2337), .C0(index_i[4]), 
          .Z(n23477));
    LUT4 i21968_3_lut (.A(n22045), .B(n22046), .C(index_i[4]), .Z(n22047)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21968_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_4_i684_3_lut (.A(n619), .B(n108), .C(index_i[3]), 
         .Z(n684_adj_2678)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_4_i684_3_lut.init = 16'hcaca;
    LUT4 i19606_3_lut (.A(n26989), .B(n27026), .C(index_i[3]), .Z(n22043)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19606_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_3_i93_3_lut_4_lut (.A(n27085), .B(index_q[2]), .C(index_q[3]), 
         .D(n27088), .Z(n93_adj_2434)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_3_i93_3_lut_4_lut.init = 16'hefe0;
    LUT4 index_i_0__bdd_4_lut_24773 (.A(index_i[0]), .B(index_i[3]), .C(index_i[1]), 
         .D(index_i[2]), .Z(n27181)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C))+!A (B (C (D)+!C !(D))+!B !(C+!(D))))) */ ;
    defparam index_i_0__bdd_4_lut_24773.init = 16'h16d3;
    LUT4 mux_197_Mux_9_i124_3_lut_3_lut_4_lut (.A(n27085), .B(index_q[2]), 
         .C(n26893), .D(index_q[3]), .Z(n124_adj_2402)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_9_i124_3_lut_3_lut_4_lut.init = 16'h11f0;
    LUT4 i21970_3_lut (.A(n22042), .B(n22043), .C(index_i[4]), .Z(n22044)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21970_3_lut.init = 16'hcaca;
    PFUMX i20450 (.BLUT(n22903), .ALUT(n22904), .C0(index_i[5]), .Z(n22906));
    LUT4 mux_197_Mux_5_i15_3_lut (.A(n27078), .B(n29477), .C(index_q[3]), 
         .Z(n15_adj_2496)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_5_i15_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_8_i475_3_lut_3_lut_4_lut (.A(n27085), .B(index_q[2]), 
         .C(n26893), .D(index_q[3]), .Z(n475_adj_2630)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_8_i475_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 mux_197_Mux_0_i1002_3_lut_3_lut_4_lut (.A(n27085), .B(index_q[2]), 
         .C(n1001), .D(index_q[3]), .Z(n1002)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i1002_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 mux_197_Mux_7_i890_3_lut_3_lut_4_lut (.A(n27085), .B(index_q[2]), 
         .C(n26871), .D(index_q[3]), .Z(n890_adj_2276)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_7_i890_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 i21974_3_lut (.A(n22039), .B(n22040), .C(index_i[4]), .Z(n22041)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21974_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_6_i891_3_lut (.A(n301_adj_2679), .B(n890_adj_2490), 
         .C(index_i[4]), .Z(n891_adj_2640)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_6_i891_3_lut.init = 16'hcaca;
    PFUMX mux_197_Mux_3_i763 (.BLUT(n747_adj_2673), .ALUT(n762_adj_2305), 
          .C0(index_q[4]), .Z(n763_adj_2680)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 mux_196_Mux_6_i828_4_lut (.A(n812_adj_2681), .B(n14178), .C(index_i[4]), 
         .D(index_i[2]), .Z(n828_adj_2639)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_6_i828_4_lut.init = 16'hfaca;
    LUT4 mux_196_Mux_6_i797_3_lut (.A(n781_adj_2260), .B(n26809), .C(index_i[4]), 
         .Z(n797_adj_2638)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_6_i797_3_lut.init = 16'hcaca;
    LUT4 i23364_then_3_lut (.A(index_q[0]), .B(index_q[4]), .C(index_q[3]), 
         .Z(n27183)) /* synthesis lut_function=(A (B)+!A (B (C)+!B !(C))) */ ;
    defparam i23364_then_3_lut.init = 16'hc9c9;
    LUT4 i22487_3_lut_4_lut (.A(n26874), .B(n19801), .C(index_i[8]), .D(n766), 
         .Z(n21533)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i22487_3_lut_4_lut.init = 16'hefe0;
    LUT4 i22485_3_lut_4_lut (.A(n26870), .B(n19798), .C(index_q[8]), .D(n766_adj_2682), 
         .Z(n21539)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i22485_3_lut_4_lut.init = 16'hefe0;
    PFUMX i19244 (.BLUT(n21679), .ALUT(n21680), .C0(index_i[5]), .Z(n21681));
    LUT4 i23364_else_3_lut (.A(index_q[0]), .B(index_q[2]), .C(index_q[4]), 
         .D(index_q[3]), .Z(n27182)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C (D)+!C !(D))+!B !(C)))) */ ;
    defparam i23364_else_3_lut.init = 16'h1e58;
    PFUMX i19247 (.BLUT(n21682), .ALUT(n21683), .C0(index_i[5]), .Z(n21684));
    LUT4 mux_196_Mux_6_i669_3_lut (.A(n653_adj_2642), .B(n668_adj_2683), 
         .C(index_i[4]), .Z(n669_adj_2634)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_6_i669_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_6_i542_3_lut (.A(n526), .B(n541_adj_2684), .C(index_i[4]), 
         .Z(n542_adj_2631)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_6_i542_3_lut.init = 16'hcaca;
    LUT4 i19221_3_lut (.A(n301_adj_2679), .B(n93_adj_2652), .C(index_i[4]), 
         .Z(n21658)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19221_3_lut.init = 16'hcaca;
    LUT4 i19594_3_lut (.A(n396), .B(n26934), .C(index_i[3]), .Z(n22031)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19594_3_lut.init = 16'hcaca;
    LUT4 i12189_3_lut (.A(index_i[3]), .B(index_i[1]), .C(index_i[0]), 
         .Z(n14875)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i12189_3_lut.init = 16'hc8c8;
    LUT4 i21985_3_lut (.A(n22030), .B(n22031), .C(index_i[4]), .Z(n22032)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21985_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_3_i348_3_lut (.A(n29487), .B(n26934), .C(index_i[3]), 
         .Z(n348_adj_2685)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_3_i348_3_lut.init = 16'hcaca;
    LUT4 i19218_3_lut (.A(n15_adj_2686), .B(n30), .C(index_i[4]), .Z(n21655)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19218_3_lut.init = 16'hcaca;
    PFUMX i19250 (.BLUT(n21685), .ALUT(n21686), .C0(index_i[5]), .Z(n21687));
    LUT4 mux_196_Mux_6_i252_4_lut (.A(index_i[2]), .B(n251_adj_2687), .C(index_i[4]), 
         .D(n11274), .Z(n252_adj_2688)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_6_i252_4_lut.init = 16'hc5ca;
    LUT4 i22254_3_lut (.A(n25653), .B(n252_adj_2688), .C(index_i[5]), 
         .Z(n23285)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22254_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_3_i684_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[4]), .Z(n684_adj_2620)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A !(B ((D)+!C)+!B (C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_3_i684_3_lut_3_lut_4_lut.init = 16'h5594;
    LUT4 mux_197_Mux_0_i908_3_lut_4_lut (.A(index_q[0]), .B(n27090), .C(index_q[3]), 
         .D(n27087), .Z(n908)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (C+!(D)))) */ ;
    defparam mux_197_Mux_0_i908_3_lut_4_lut.init = 16'h2f20;
    LUT4 i19591_3_lut (.A(n26988), .B(n27032), .C(index_i[3]), .Z(n22028)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19591_3_lut.init = 16'hcaca;
    PFUMX i19253 (.BLUT(n21688), .ALUT(n21689), .C0(index_i[5]), .Z(n21690));
    LUT4 mux_196_Mux_3_i908_3_lut (.A(n27029), .B(n26978), .C(index_i[3]), 
         .Z(n908_adj_2689)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_3_i908_3_lut.init = 16'hcaca;
    LUT4 i20802_3_lut (.A(n236), .B(n251), .C(index_q[4]), .Z(n23258)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20802_3_lut.init = 16'hcaca;
    LUT4 i21990_3_lut (.A(n22024), .B(n22025), .C(index_i[4]), .Z(n22026)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21990_3_lut.init = 16'hcaca;
    LUT4 i22669_2_lut (.A(index_q[5]), .B(index_q[4]), .Z(n22399)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i22669_2_lut.init = 16'heeee;
    PFUMX i20463 (.BLUT(n22915), .ALUT(n22916), .C0(index_q[5]), .Z(n22919));
    LUT4 n986_bdd_4_lut_4_lut_4_lut (.A(index_q[0]), .B(n27090), .C(index_q[4]), 
         .D(index_q[3]), .Z(n24708)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (D))+!A (B (C (D)+!C !(D))+!B (D)))) */ ;
    defparam n986_bdd_4_lut_4_lut_4_lut.init = 16'h0c73;
    LUT4 i19582_3_lut (.A(n29471), .B(n26977), .C(index_i[3]), .Z(n22019)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19582_3_lut.init = 16'hcaca;
    PFUMX i19628 (.BLUT(n22063), .ALUT(n22064), .C0(index_i[4]), .Z(n22065));
    LUT4 i19581_3_lut (.A(n27028), .B(n26993), .C(index_i[3]), .Z(n22018)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19581_3_lut.init = 16'hcaca;
    LUT4 i21997_3_lut (.A(n22018), .B(n22019), .C(index_i[4]), .Z(n22020)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21997_3_lut.init = 16'hcaca;
    LUT4 i20795_3_lut (.A(n15_adj_2413), .B(n27174), .C(index_q[4]), .Z(n23251)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20795_3_lut.init = 16'hcaca;
    PFUMX i19631 (.BLUT(n22066), .ALUT(n22067), .C0(index_i[4]), .Z(n22068));
    LUT4 n715_bdd_3_lut (.A(n27087), .B(n652), .C(index_q[3]), .Z(n26513)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n715_bdd_3_lut.init = 16'hcaca;
    PFUMX i22933 (.BLUT(n21595), .ALUT(n24617), .C0(index_i[6]), .Z(n24618));
    CCU2D add_377_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(quarter_wave_sample_register_q[0]), .B1(quarter_wave_sample_register_q[1]), 
          .C1(GND_net), .D1(GND_net), .COUT(n17571));   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(80[29:60])
    defparam add_377_1.INIT0 = 16'hF000;
    defparam add_377_1.INIT1 = 16'ha666;
    defparam add_377_1.INJECT1_0 = "NO";
    defparam add_377_1.INJECT1_1 = "NO";
    LUT4 i19035_3_lut_3_lut_4_lut (.A(index_q[0]), .B(n27090), .C(n26893), 
         .D(index_q[3]), .Z(n21472)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(C+(D)))) */ ;
    defparam i19035_3_lut_3_lut_4_lut.init = 16'h77f0;
    PFUMX i20464 (.BLUT(n22917), .ALUT(n22918), .C0(index_q[5]), .Z(n22920));
    LUT4 i19579_3_lut (.A(n29497), .B(n26933), .C(index_i[3]), .Z(n22016)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19579_3_lut.init = 16'hcaca;
    LUT4 i19578_3_lut (.A(n27001), .B(n619), .C(index_i[3]), .Z(n22015)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19578_3_lut.init = 16'hcaca;
    LUT4 index_i_1__bdd_4_lut_25572 (.A(index_i[1]), .B(index_i[0]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n27185)) /* synthesis lut_function=(!(A (B (D)+!B (C+!(D)))+!A !(B (C (D)+!C !(D))+!B !((D)+!C)))) */ ;
    defparam index_i_1__bdd_4_lut_25572.init = 16'h429c;
    PFUMX i20470 (.BLUT(n22922), .ALUT(n22923), .C0(index_q[5]), .Z(n22926));
    LUT4 mux_196_Mux_2_i270_3_lut (.A(n26932), .B(n29490), .C(index_i[3]), 
         .Z(n270_adj_2690)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_2_i270_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_2_i316_3_lut (.A(n26988), .B(n27025), .C(index_i[3]), 
         .Z(n316_adj_2691)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_2_i316_3_lut.init = 16'hcaca;
    PFUMX i20143 (.BLUT(n158_adj_2656), .ALUT(n189_adj_2692), .C0(index_q[5]), 
          .Z(n22599));
    LUT4 i21999_3_lut (.A(n22015), .B(n22016), .C(index_i[4]), .Z(n22017)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21999_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_2_i397_3_lut (.A(n29497), .B(n26928), .C(index_i[3]), 
         .Z(n397_adj_2693)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_2_i397_3_lut.init = 16'hcaca;
    PFUMX i20471 (.BLUT(n22924), .ALUT(n22925), .C0(index_q[5]), .Z(n22927));
    PFUMX i21022 (.BLUT(n908_adj_2694), .ALUT(n923_adj_2651), .C0(index_i[4]), 
          .Z(n23478));
    PFUMX i19256 (.BLUT(n21691), .ALUT(n21692), .C0(index_i[5]), .Z(n21693));
    PFUMX i19259 (.BLUT(n21694), .ALUT(n21695), .C0(index_i[5]), .Z(n21696));
    LUT4 i11478_3_lut_4_lut (.A(index_q[0]), .B(n27090), .C(n26967), .D(index_q[5]), 
         .Z(n318)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (C (D))) */ ;
    defparam i11478_3_lut_4_lut.init = 16'hf800;
    LUT4 i19722_3_lut_3_lut_4_lut (.A(index_q[0]), .B(n27090), .C(index_q[3]), 
         .D(n26893), .Z(n22159)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A !(C+(D))) */ ;
    defparam i19722_3_lut_3_lut_4_lut.init = 16'h808f;
    PFUMX i19262 (.BLUT(n21697), .ALUT(n21698), .C0(index_i[5]), .Z(n21699));
    LUT4 i20298_3_lut (.A(n22749), .B(n22750), .C(index_i[7]), .Z(n22754)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20298_3_lut.init = 16'hcaca;
    PFUMX i21023 (.BLUT(n939_adj_2650), .ALUT(n954_adj_2695), .C0(index_i[4]), 
          .Z(n23479));
    LUT4 mux_196_Mux_1_i924_3_lut (.A(n908_adj_2282), .B(n412_adj_2320), 
         .C(index_i[4]), .Z(n924_adj_2589)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_1_i924_3_lut.init = 16'hcaca;
    LUT4 n62_bdd_3_lut_24483_4_lut (.A(n27063), .B(index_q[3]), .C(index_q[4]), 
         .D(n30_adj_2696), .Z(n24807)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n62_bdd_3_lut_24483_4_lut.init = 16'hf808;
    LUT4 i19570_3_lut (.A(n27032), .B(n396), .C(index_i[3]), .Z(n22007)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19570_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_adj_85 (.A(index_q[0]), .B(index_q[4]), .C(index_q[2]), 
         .Z(n20689)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_3_lut_adj_85.init = 16'hfefe;
    LUT4 i21931_3_lut (.A(n22093), .B(n22094), .C(index_i[4]), .Z(n22095)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21931_3_lut.init = 16'hcaca;
    LUT4 i19287_3_lut_4_lut_4_lut (.A(n26871), .B(index_q[4]), .C(index_q[3]), 
         .D(n26854), .Z(n21724)) /* synthesis lut_function=(A (B (C)+!B !(C+!(D)))+!A (B (C)+!B (C+(D)))) */ ;
    defparam i19287_3_lut_4_lut_4_lut.init = 16'hd3d0;
    LUT4 i22011_3_lut (.A(n22006), .B(n22007), .C(index_i[4]), .Z(n22008)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22011_3_lut.init = 16'hcaca;
    PFUMX i19268 (.BLUT(n21703), .ALUT(n21704), .C0(index_q[5]), .Z(n21705));
    PFUMX i21024 (.BLUT(n971_adj_2646), .ALUT(n986_adj_2645), .C0(index_i[4]), 
          .Z(n23480));
    L6MUX21 i24451 (.D0(n26355), .D1(n26353), .SD(index_q[8]), .Z(n26356));
    LUT4 i20461_3_lut_3_lut_4_lut_4_lut (.A(n27063), .B(index_q[3]), .C(index_q[4]), 
         .D(n26854), .Z(n22917)) /* synthesis lut_function=(!(A (B (C)+!B ((D)+!C))+!A (B+((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20461_3_lut_3_lut_4_lut_4_lut.init = 16'h0838;
    PFUMX i21025 (.BLUT(n1002_adj_2484), .ALUT(n1017_adj_2697), .C0(index_i[4]), 
          .Z(n23481));
    LUT4 i19566_3_lut (.A(n773), .B(n27025), .C(index_i[3]), .Z(n22003)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19566_3_lut.init = 16'hcaca;
    LUT4 i19564_3_lut (.A(n723), .B(n396), .C(index_i[3]), .Z(n22001)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19564_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_1_i349_3_lut (.A(n506), .B(n348_adj_2698), .C(index_i[4]), 
         .Z(n349_adj_2587)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_1_i349_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_1_i986_3_lut (.A(n29491), .B(n29487), .C(index_i[3]), 
         .Z(n986_adj_2699)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_1_i986_3_lut.init = 16'hcaca;
    LUT4 i21940_3_lut (.A(n22069), .B(n22070), .C(index_i[4]), .Z(n22071)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21940_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_2_i955_then_4_lut (.A(index_i[4]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n27124)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B (C+!(D))+!B !(C (D)))) */ ;
    defparam mux_196_Mux_2_i955_then_4_lut.init = 16'he95d;
    LUT4 i9558_3_lut_4_lut_4_lut (.A(n27063), .B(index_q[3]), .C(index_q[5]), 
         .D(n26871), .Z(n12120)) /* synthesis lut_function=(A (B+(C (D)))+!A (B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9558_3_lut_4_lut_4_lut.init = 16'hf8c8;
    LUT4 index_q_3__bdd_3_lut_24675_4_lut_4_lut (.A(n27063), .B(index_q[3]), 
         .C(index_q[4]), .D(n26861), .Z(n24492)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C))+!A !(B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam index_q_3__bdd_3_lut_24675_4_lut_4_lut.init = 16'h838f;
    LUT4 mux_196_Mux_1_i94_3_lut (.A(index_i[0]), .B(n93_adj_2397), .C(index_i[4]), 
         .Z(n94_adj_2584)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_1_i94_3_lut.init = 16'hcaca;
    PFUMX mux_197_Mux_5_i732 (.BLUT(n11958), .ALUT(n731_adj_2641), .C0(index_q[4]), 
          .Z(n732_adj_2700)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 n123_bdd_3_lut_23671_4_lut (.A(n27093), .B(index_q[2]), .C(n27065), 
         .D(index_q[3]), .Z(n25443)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (B (C+!(D))+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n123_bdd_3_lut_23671_4_lut.init = 16'hf066;
    PFUMX i19271 (.BLUT(n21706), .ALUT(n21707), .C0(index_q[5]), .Z(n21708));
    PFUMX i24449 (.BLUT(n26354), .ALUT(n22485), .C0(index_q[7]), .Z(n26355));
    LUT4 i19272_3_lut_then_4_lut (.A(index_q[4]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n27187)) /* synthesis lut_function=(A (B (C)+!B !(C (D)+!C !(D)))+!A !(B (C)+!B !(C (D)+!C !(D)))) */ ;
    defparam i19272_3_lut_then_4_lut.init = 16'h96a5;
    LUT4 i22475_3_lut (.A(n24626), .B(n22662), .C(index_i[8]), .Z(n22664)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22475_3_lut.init = 16'hcaca;
    LUT4 i19557_3_lut (.A(n29497), .B(n29472), .C(index_i[3]), .Z(n21994)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19557_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_3_i668_3_lut_4_lut (.A(n27093), .B(index_q[2]), .C(index_q[3]), 
         .D(n27080), .Z(n668_adj_2428)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_3_i668_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_197_Mux_4_i763_3_lut_4_lut (.A(n27093), .B(index_q[2]), .C(index_q[4]), 
         .D(n747_adj_2367), .Z(n763_adj_2701)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_4_i763_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_196_Mux_9_i364_3_lut_3_lut_4_lut (.A(n26937), .B(index_i[1]), 
         .C(index_i[3]), .D(n26882), .Z(n364_adj_2279)) /* synthesis lut_function=(!(A (C (D))+!A (B (C (D))+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_9_i364_3_lut_3_lut_4_lut.init = 16'h0efe;
    LUT4 n22624_bdd_3_lut (.A(n22617), .B(n22618), .C(index_q[7]), .Z(n26560)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n22624_bdd_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_0_i572_3_lut_4_lut (.A(n26937), .B(index_i[1]), .C(index_i[3]), 
         .D(n27028), .Z(n572_adj_2522)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_0_i572_3_lut_4_lut.init = 16'hefe0;
    PFUMX i19640 (.BLUT(n22075), .ALUT(n22076), .C0(index_i[4]), .Z(n22077));
    LUT4 i21956_3_lut (.A(n716_adj_2275), .B(n731_adj_2702), .C(index_i[4]), 
         .Z(n732_adj_2578)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21956_3_lut.init = 16'hcaca;
    PFUMX i19643 (.BLUT(n22078), .ALUT(n22079), .C0(index_i[4]), .Z(n22080));
    LUT4 i19641_3_lut_3_lut_4_lut (.A(n26937), .B(index_i[1]), .C(n26876), 
         .D(index_i[3]), .Z(n22078)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19641_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 i19608_3_lut_3_lut_4_lut (.A(n26937), .B(index_i[1]), .C(index_i[3]), 
         .D(n26876), .Z(n22045)) /* synthesis lut_function=(!(A (C (D))+!A (B (C (D))+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19608_3_lut_3_lut_4_lut.init = 16'h0efe;
    PFUMX i19646 (.BLUT(n22081), .ALUT(n22082), .C0(index_i[4]), .Z(n22083));
    LUT4 index_i_3__bdd_3_lut_22937_3_lut_4_lut (.A(n26937), .B(index_i[1]), 
         .C(index_i[4]), .D(index_i[3]), .Z(n24622)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam index_i_3__bdd_3_lut_22937_3_lut_4_lut.init = 16'hf10f;
    LUT4 n24625_bdd_3_lut_26342 (.A(n24625), .B(n24618), .C(index_i[7]), 
         .Z(n24626)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n24625_bdd_3_lut_26342.init = 16'hcaca;
    PFUMX i19649 (.BLUT(n22084), .ALUT(n22085), .C0(index_i[4]), .Z(n22086));
    LUT4 mux_196_Mux_2_i669_3_lut (.A(n653_adj_2703), .B(n475_adj_2704), 
         .C(index_i[4]), .Z(n669_adj_2576)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_2_i669_3_lut.init = 16'hcaca;
    LUT4 n25413_bdd_3_lut_24608 (.A(n25413), .B(n22615), .C(index_q[7]), 
         .Z(n26562)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n25413_bdd_3_lut_24608.init = 16'hacac;
    LUT4 mux_197_Mux_0_i220_3_lut (.A(n27058), .B(n27081), .C(index_q[3]), 
         .Z(n220)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i220_3_lut.init = 16'hcaca;
    LUT4 n25413_bdd_3_lut_25592 (.A(n22613), .B(n22614), .C(index_q[7]), 
         .Z(n26563)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n25413_bdd_3_lut_25592.init = 16'hcaca;
    LUT4 mux_196_Mux_2_i605_3_lut (.A(n142_adj_2705), .B(n604_adj_2361), 
         .C(index_i[4]), .Z(n605_adj_2575)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_2_i605_3_lut.init = 16'hcaca;
    LUT4 i21964_3_lut (.A(n29500), .B(n22052), .C(index_i[4]), .Z(n22053)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21964_3_lut.init = 16'hcaca;
    LUT4 i11613_3_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .Z(n11274)) /* synthesis lut_function=(!((B (C))+!A)) */ ;
    defparam i11613_3_lut.init = 16'h2a2a;
    LUT4 i21966_3_lut (.A(n22048), .B(n22049), .C(index_i[4]), .Z(n22050)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21966_3_lut.init = 16'hcaca;
    PFUMX i24447 (.BLUT(n26352), .ALUT(n26351), .C0(index_q[7]), .Z(n26353));
    LUT4 mux_196_Mux_2_i413_3_lut (.A(n397_adj_2693), .B(n954_adj_2706), 
         .C(index_i[4]), .Z(n413_adj_2571)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_2_i413_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_2_i317_3_lut (.A(n668_adj_2354), .B(n316_adj_2691), 
         .C(index_i[4]), .Z(n317_adj_2566)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_2_i317_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_3_i251_3_lut_4_lut (.A(n26937), .B(index_i[1]), .C(index_i[3]), 
         .D(n26882), .Z(n15108)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_3_i251_3_lut_4_lut.init = 16'hfe0e;
    LUT4 mux_196_Mux_2_i286_3_lut (.A(n270_adj_2690), .B(n653_adj_2707), 
         .C(index_i[4]), .Z(n286_adj_2565)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_2_i286_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_0_i716_3_lut (.A(n27033), .B(n26978), .C(index_i[3]), 
         .Z(n716_adj_2567)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_0_i716_3_lut.init = 16'hcaca;
    LUT4 i19552_3_lut (.A(n27100), .B(n29494), .C(index_q[3]), .Z(n21989)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19552_3_lut.init = 16'hcaca;
    LUT4 i21976_3_lut (.A(n142), .B(n14203), .C(index_i[4]), .Z(n158_adj_2562)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21976_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_6_i668_3_lut (.A(n108), .B(n27002), .C(index_i[3]), 
         .Z(n668_adj_2683)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_6_i668_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_6_i684_3_lut (.A(n26900), .B(n29497), .C(index_i[3]), 
         .Z(n684_adj_2708)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_6_i684_3_lut.init = 16'hcaca;
    LUT4 i9485_4_lut_4_lut (.A(n26937), .B(index_i[1]), .C(index_i[3]), 
         .D(n20693), .Z(n12046)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A (B (C)+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9485_4_lut_4_lut.init = 16'h0e3e;
    PFUMX i19655 (.BLUT(n22090), .ALUT(n22091), .C0(index_i[4]), .Z(n22092));
    LUT4 mux_196_Mux_0_i653_3_lut (.A(n26900), .B(n26977), .C(index_i[3]), 
         .Z(n653_adj_2555)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_0_i653_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_8_i732_3_lut (.A(index_q[3]), .B(n15132), .C(index_q[5]), 
         .Z(n732_adj_2558)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_8_i732_3_lut.init = 16'h3a3a;
    LUT4 i21983_3_lut (.A(n22033), .B(n27181), .C(index_i[4]), .Z(n22035)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21983_3_lut.init = 16'hcaca;
    LUT4 i11355_2_lut_rep_415_3_lut_4_lut (.A(n26937), .B(index_i[1]), .C(index_i[4]), 
         .D(index_i[3]), .Z(n26738)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11355_2_lut_rep_415_3_lut_4_lut.init = 16'hfef0;
    LUT4 i19236_4_lut_4_lut_3_lut_4_lut (.A(n26937), .B(index_i[1]), .C(index_i[4]), 
         .D(index_i[3]), .Z(n21673)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19236_4_lut_4_lut_3_lut_4_lut.init = 16'h11ef;
    LUT4 mux_196_Mux_3_i924_3_lut (.A(n908_adj_2689), .B(index_i[0]), .C(index_i[4]), 
         .Z(n924_adj_2551)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_3_i924_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_3_i891_3_lut (.A(n541_adj_2684), .B(n890_adj_2709), 
         .C(index_i[4]), .Z(n891_adj_2547)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_3_i891_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_3_i669_3_lut (.A(n653_adj_2707), .B(n668_adj_2354), 
         .C(index_i[4]), .Z(n669_adj_2544)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_3_i669_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_2_i955_else_4_lut (.A(index_i[4]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n27123)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C+(D)))+!A !(B (C+!(D))+!B !(C+!(D))))) */ ;
    defparam mux_196_Mux_2_i955_else_4_lut.init = 16'h49c6;
    LUT4 mux_196_Mux_7_i333_3_lut (.A(n27001), .B(n26900), .C(index_i[3]), 
         .Z(n333_adj_2671)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_7_i333_3_lut.init = 16'hcaca;
    PFUMX i19661 (.BLUT(n22096), .ALUT(n22097), .C0(index_i[4]), .Z(n22098));
    LUT4 i9530_4_lut (.A(n27046), .B(n26836), .C(index_i[3]), .D(index_i[4]), 
         .Z(n12091)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B ((D)+!C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9530_4_lut.init = 16'h3afa;
    LUT4 mux_196_Mux_7_i348_3_lut (.A(n29491), .B(n26999), .C(index_i[3]), 
         .Z(n348_adj_2669)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_7_i348_3_lut.init = 16'hcaca;
    LUT4 i19548_3_lut (.A(n27099), .B(n29494), .C(index_q[3]), .Z(n21985)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19548_3_lut.init = 16'hcaca;
    LUT4 i19272_3_lut_else_4_lut (.A(index_q[4]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n27186)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C+!(D)))+!A !(B ((D)+!C)+!B (C (D)+!C !(D))))) */ ;
    defparam i19272_3_lut_else_4_lut.init = 16'h5685;
    PFUMX i19664 (.BLUT(n22099), .ALUT(n22100), .C0(index_i[4]), .Z(n22101));
    LUT4 i21992_3_lut (.A(n22021), .B(n22022), .C(index_i[4]), .Z(n22023)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21992_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_7_i397_3_lut (.A(n29491), .B(n27001), .C(index_i[3]), 
         .Z(n397_adj_2661)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_7_i397_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_3_i476_3_lut (.A(n460_adj_2379), .B(n285_adj_2380), 
         .C(index_i[4]), .Z(n476_adj_2540)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_3_i476_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_8_i653_3_lut_rep_398_3_lut_4_lut (.A(index_i[0]), .B(n27046), 
         .C(n26882), .D(index_i[3]), .Z(n26721)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(C+(D)))) */ ;
    defparam mux_196_Mux_8_i653_3_lut_rep_398_3_lut_4_lut.init = 16'h77f0;
    PFUMX i19280 (.BLUT(n21715), .ALUT(n21716), .C0(index_q[5]), .Z(n21717));
    LUT4 mux_196_Mux_11_i638_4_lut_4_lut (.A(n26738), .B(index_i[5]), .C(index_i[6]), 
         .D(n26777), .Z(n638_adj_2710)) /* synthesis lut_function=(A (B (C (D))+!B !(C))+!A (B ((D)+!C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_11_i638_4_lut_4_lut.init = 16'hc707;
    PFUMX i19667 (.BLUT(n22102), .ALUT(n22103), .C0(index_i[4]), .Z(n22104));
    LUT4 mux_196_Mux_3_i413_3_lut (.A(n397_adj_2711), .B(n26976), .C(index_i[4]), 
         .Z(n413_adj_2538)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_3_i413_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_0_i620_3_lut (.A(n29491), .B(n29488), .C(index_i[3]), 
         .Z(n620_adj_2535)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_0_i620_3_lut.init = 16'hcaca;
    LUT4 i19546_3_lut (.A(n27103), .B(n29485), .C(index_q[3]), .Z(n21983)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19546_3_lut.init = 16'hcaca;
    LUT4 i11409_3_lut_4_lut (.A(index_i[0]), .B(n27046), .C(n26995), .D(index_i[5]), 
         .Z(n318_adj_2418)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (C (D))) */ ;
    defparam i11409_3_lut_4_lut.init = 16'hf800;
    PFUMX i19283 (.BLUT(n21718), .ALUT(n21719), .C0(index_q[5]), .Z(n21720));
    LUT4 mux_196_Mux_3_i286_4_lut (.A(n93_adj_2487), .B(index_i[2]), .C(index_i[4]), 
         .D(n14875), .Z(n286_adj_2533)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_3_i286_4_lut.init = 16'h3aca;
    PFUMX i19286 (.BLUT(n21721), .ALUT(n21722), .C0(index_q[5]), .Z(n21723));
    LUT4 i21658_3_lut (.A(n21982), .B(n21983), .C(index_q[4]), .Z(n21984)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21658_3_lut.init = 16'hcaca;
    LUT4 i19543_3_lut (.A(n29489), .B(n27024), .C(index_i[3]), .Z(n21980)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19543_3_lut.init = 16'hcaca;
    LUT4 i19542_3_lut (.A(n26991), .B(n396), .C(index_i[3]), .Z(n21979)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19542_3_lut.init = 16'hcaca;
    L6MUX21 i20514 (.D0(n22968), .D1(n22969), .SD(index_i[5]), .Z(n22970));
    LUT4 i22023_3_lut (.A(n21979), .B(n21980), .C(index_i[4]), .Z(n21981)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22023_3_lut.init = 16'hcaca;
    LUT4 i19540_3_lut (.A(n27031), .B(n26977), .C(index_i[3]), .Z(n21977)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19540_3_lut.init = 16'hcaca;
    LUT4 i22025_3_lut (.A(n21976), .B(n21977), .C(index_i[4]), .Z(n21978)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22025_3_lut.init = 16'hcaca;
    LUT4 n699_bdd_4_lut_4_lut_4_lut (.A(index_i[0]), .B(n27046), .C(index_i[4]), 
         .D(index_i[3]), .Z(n24639)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (D))+!A (B (C (D)+!C !(D))+!B (D)))) */ ;
    defparam n699_bdd_4_lut_4_lut_4_lut.init = 16'h0c73;
    PFUMX mux_196_Mux_1_i891 (.BLUT(n882), .ALUT(n890_adj_2712), .C0(n26925), 
          .Z(n891_adj_2301)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 n62_bdd_3_lut_4_lut (.A(n27048), .B(index_i[3]), .C(index_i[4]), 
         .D(n30_adj_2713), .Z(n24785)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n62_bdd_3_lut_4_lut.init = 16'hf808;
    LUT4 mux_196_Mux_3_i158_3_lut (.A(n142_adj_2705), .B(n157_adj_2319), 
         .C(index_i[4]), .Z(n158_adj_2530)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_3_i158_3_lut.init = 16'hcaca;
    PFUMX i19289 (.BLUT(n21724), .ALUT(n21725), .C0(index_q[5]), .Z(n21726));
    LUT4 mux_196_Mux_3_i125_3_lut (.A(n46_adj_2714), .B(n30), .C(index_i[4]), 
         .Z(n125_adj_2526)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_3_i125_3_lut.init = 16'hcaca;
    LUT4 i20440_3_lut_3_lut_4_lut_4_lut (.A(n27048), .B(index_i[3]), .C(index_i[4]), 
         .D(n26882), .Z(n22896)) /* synthesis lut_function=(!(A (B (C)+!B ((D)+!C))+!A (B+((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20440_3_lut_3_lut_4_lut_4_lut.init = 16'h0838;
    LUT4 i9486_3_lut_4_lut_4_lut (.A(n27048), .B(index_i[3]), .C(index_i[5]), 
         .D(n26876), .Z(n12047)) /* synthesis lut_function=(A (B+(C (D)))+!A (B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9486_3_lut_4_lut_4_lut.init = 16'hf8c8;
    LUT4 mux_196_Mux_0_i589_3_lut (.A(n26999), .B(n773), .C(index_i[3]), 
         .Z(n589_adj_2524)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_0_i589_3_lut.init = 16'hcaca;
    LUT4 index_i_3__bdd_3_lut_23776_4_lut_4_lut (.A(n27048), .B(index_i[3]), 
         .C(index_i[4]), .D(n26836), .Z(n24623)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C))+!A !(B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam index_i_3__bdd_3_lut_23776_4_lut_4_lut.init = 16'h838f;
    LUT4 i19273_3_lut_then_4_lut (.A(index_q[4]), .B(index_q[1]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n27190)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)+!C !(D)))+!A !(B (C+!(D))+!B (C (D)+!C !(D))))) */ ;
    defparam i19273_3_lut_then_4_lut.init = 16'h5a65;
    PFUMX i19679 (.BLUT(n22114), .ALUT(n22115), .C0(index_q[4]), .Z(n22116));
    LUT4 i22031_3_lut (.A(n21973), .B(n21974), .C(index_i[4]), .Z(n21975)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22031_3_lut.init = 16'hcaca;
    LUT4 i20286_4_lut (.A(n22014), .B(n1002_adj_2715), .C(index_i[5]), 
         .D(index_i[4]), .Z(n22742)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;
    defparam i20286_4_lut.init = 16'hfaca;
    LUT4 i19533_3_lut (.A(n27024), .B(n29471), .C(index_i[3]), .Z(n21970)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19533_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_4_i860_3_lut (.A(n506_adj_2649), .B(n25320), .C(index_i[4]), 
         .Z(n860_adj_2511)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_4_i860_3_lut.init = 16'hcaca;
    LUT4 i22013_3_lut (.A(n22003), .B(n22004), .C(index_i[4]), .Z(n22005)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22013_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_5_i700_3_lut (.A(n460_adj_2716), .B(n27022), .C(index_i[4]), 
         .Z(n700_adj_2454)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_5_i700_3_lut.init = 16'hcaca;
    LUT4 i11420_2_lut_3_lut_4_lut (.A(n26854), .B(n26967), .C(index_q[6]), 
         .D(index_q[5]), .Z(n254_adj_2717)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11420_2_lut_3_lut_4_lut.init = 16'hfef0;
    LUT4 i22015_3_lut (.A(n22000), .B(n22001), .C(index_i[4]), .Z(n22002)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22015_3_lut.init = 16'hcaca;
    LUT4 i19527_3_lut (.A(n396), .B(n29471), .C(index_i[3]), .Z(n21964)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19527_3_lut.init = 16'hcaca;
    LUT4 i19273_3_lut_else_4_lut (.A(index_q[4]), .B(index_q[1]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n27189)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A !(B (C+!(D))+!B ((D)+!C)))) */ ;
    defparam i19273_3_lut_else_4_lut.init = 16'h59e5;
    LUT4 mux_196_Mux_4_i700_3_lut (.A(n684_adj_2678), .B(index_i[1]), .C(index_i[4]), 
         .Z(n700_adj_2504)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_4_i700_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_4_i669_3_lut (.A(n781_adj_2260), .B(n668_adj_2326), 
         .C(index_i[4]), .Z(n669_adj_2503)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_4_i669_3_lut.init = 16'hcaca;
    PFUMX i20517 (.BLUT(n158_adj_2618), .ALUT(n189_adj_2353), .C0(index_q[5]), 
          .Z(n22973));
    LUT4 mux_196_Mux_4_i542_3_lut (.A(n30), .B(n506), .C(index_i[4]), 
         .Z(n542_adj_2718)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_4_i542_3_lut.init = 16'hcaca;
    LUT4 i20280_4_lut (.A(n26813), .B(n27177), .C(index_i[5]), .D(index_i[4]), 
         .Z(n22736)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam i20280_4_lut.init = 16'hc5ca;
    PFUMX i20518 (.BLUT(n221_adj_2719), .ALUT(n21468), .C0(index_q[5]), 
          .Z(n22974));
    LUT4 i22019_3_lut (.A(n22111), .B(n22112), .C(index_q[4]), .Z(n22113)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i22019_3_lut.init = 16'hcaca;
    PFUMX i20519 (.BLUT(n286_adj_2617), .ALUT(n317_adj_2615), .C0(index_q[5]), 
          .Z(n22975));
    PFUMX i20520 (.BLUT(n349_adj_2720), .ALUT(n21471), .C0(index_q[5]), 
          .Z(n22976));
    LUT4 i18991_3_lut (.A(n900), .B(n356), .C(index_q[3]), .Z(n21428)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18991_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_2_i270_3_lut (.A(n27078), .B(n27061), .C(index_q[3]), 
         .Z(n270_adj_2616)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_2_i270_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_2_i316_3_lut (.A(n27096), .B(n29493), .C(index_q[3]), 
         .Z(n316_adj_2614)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_2_i316_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_2_i397_3_lut (.A(n29485), .B(n27062), .C(index_q[3]), 
         .Z(n397_adj_2611)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_2_i397_3_lut.init = 16'hcaca;
    PFUMX i20521 (.BLUT(n413_adj_2612), .ALUT(n21474), .C0(index_q[5]), 
          .Z(n22977));
    LUT4 i19525_3_lut (.A(n26993), .B(n27032), .C(index_i[3]), .Z(n21962)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19525_3_lut.init = 16'hcaca;
    LUT4 i19524_3_lut (.A(n26934), .B(n27028), .C(index_i[3]), .Z(n21961)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19524_3_lut.init = 16'hcaca;
    LUT4 i19522_3_lut (.A(n26989), .B(n27028), .C(index_i[3]), .Z(n21959)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19522_3_lut.init = 16'hcaca;
    PFUMX i20737 (.BLUT(n142_adj_2721), .ALUT(n157_adj_2722), .C0(index_i[4]), 
          .Z(n23193));
    LUT4 mux_196_Mux_4_i286_3_lut (.A(n270_adj_2674), .B(n15_adj_2478), 
         .C(index_i[4]), .Z(n286_adj_2488)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_4_i286_3_lut.init = 16'hcaca;
    PFUMX i20522 (.BLUT(n21477), .ALUT(n507_adj_2723), .C0(index_q[5]), 
          .Z(n22978));
    LUT4 i19518_3_lut (.A(n27024), .B(n27028), .C(index_i[3]), .Z(n21955)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19518_3_lut.init = 16'hcaca;
    LUT4 i22425_3_lut_rep_393_4_lut (.A(n26860), .B(index_i[5]), .C(index_i[8]), 
         .D(n1021), .Z(n26716)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i22425_3_lut_rep_393_4_lut.init = 16'hf808;
    LUT4 mux_197_Mux_7_i333_3_lut (.A(n27104), .B(n26887), .C(index_q[3]), 
         .Z(n333_adj_2601)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_7_i333_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_7_i348_3_lut (.A(n27102), .B(n27086), .C(index_q[3]), 
         .Z(n348_adj_2598)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_7_i348_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_4_i94_3_lut (.A(n61_adj_2475), .B(n26979), .C(index_i[4]), 
         .Z(n94_adj_2483)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_4_i94_3_lut.init = 16'hcaca;
    PFUMX i20523 (.BLUT(n21480), .ALUT(n573_adj_2405), .C0(index_q[5]), 
          .Z(n22979));
    LUT4 i11344_2_lut_3_lut_4_lut (.A(n26882), .B(n26995), .C(index_i[6]), 
         .D(index_i[5]), .Z(n254_adj_2350)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i11344_2_lut_3_lut_4_lut.init = 16'hfef0;
    PFUMX i20524 (.BLUT(n605_adj_2610), .ALUT(n21483), .C0(index_q[5]), 
          .Z(n22980));
    LUT4 mux_197_Mux_3_i262_rep_765 (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .Z(n27088)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_3_i262_rep_765.init = 16'h7c7c;
    LUT4 mux_196_Mux_7_i123_3_lut_3_lut_rep_676 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26999)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_7_i123_3_lut_3_lut_rep_676.init = 16'hc7c7;
    LUT4 mux_197_Mux_7_i397_3_lut (.A(n27102), .B(n27104), .C(index_q[3]), 
         .Z(n397_adj_2596)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_7_i397_3_lut.init = 16'hcaca;
    PFUMX i20525 (.BLUT(n669_adj_2607), .ALUT(n700_adj_2672), .C0(index_q[5]), 
          .Z(n22981));
    PFUMX i20738 (.BLUT(n173_adj_2407), .ALUT(n188_adj_2603), .C0(index_i[4]), 
          .Z(n23194));
    L6MUX21 i24407 (.D0(n26298), .D1(n26295), .SD(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2126[4]));
    LUT4 i19516_3_lut (.A(n27026), .B(n29497), .C(index_i[3]), .Z(n21953)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19516_3_lut.init = 16'hcaca;
    PFUMX i20526 (.BLUT(n732_adj_2605), .ALUT(n763_adj_2724), .C0(index_q[5]), 
          .Z(n22982));
    LUT4 i21610_3_lut (.A(n21952), .B(n21953), .C(index_i[4]), .Z(n21954)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21610_3_lut.init = 16'hcaca;
    LUT4 i22423_3_lut_rep_394_4_lut (.A(n26840), .B(index_q[5]), .C(index_q[8]), 
         .D(n1021_adj_2725), .Z(n26717)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i22423_3_lut_rep_394_4_lut.init = 16'hf808;
    LUT4 i21890_3_lut (.A(n21949), .B(n21950), .C(index_i[4]), .Z(n21951)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21890_3_lut.init = 16'hcaca;
    PFUMX i24405 (.BLUT(n26297), .ALUT(n26296), .C0(index_i[8]), .Z(n26298));
    LUT4 n21321_bdd_3_lut_23674 (.A(n27094), .B(n27083), .C(index_q[3]), 
         .Z(n25446)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n21321_bdd_3_lut_23674.init = 16'hcaca;
    LUT4 mux_197_Mux_6_i732_3_lut_4_lut (.A(n27104), .B(index_q[3]), .C(index_q[4]), 
         .D(n781_adj_2600), .Z(n732_adj_2726)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_6_i732_3_lut_4_lut.init = 16'hf909;
    LUT4 i19507_3_lut (.A(n404), .B(n26990), .C(index_i[3]), .Z(n21944)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19507_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_5_i891_3_lut (.A(n875_adj_2658), .B(n379_adj_2327), 
         .C(index_i[4]), .Z(n891_adj_2461)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_5_i891_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_5_i860_3_lut (.A(n15_adj_2471), .B(n859_adj_2657), 
         .C(index_i[4]), .Z(n860_adj_2460)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_5_i860_3_lut.init = 16'hcaca;
    LUT4 i20733_3_lut (.A(n541_adj_2660), .B(n30_adj_2654), .C(index_i[4]), 
         .Z(n23189)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20733_3_lut.init = 16'hcaca;
    LUT4 i19506_3_lut (.A(n29489), .B(n396), .C(index_i[3]), .Z(n21943)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19506_3_lut.init = 16'hcaca;
    L6MUX21 i20528 (.D0(n860_adj_2627), .D1(n891_adj_2624), .SD(index_q[5]), 
            .Z(n22984));
    LUT4 mux_196_Mux_6_i844_3_lut_4_lut (.A(n26927), .B(index_i[2]), .C(index_i[3]), 
         .D(n29492), .Z(n844_adj_2259)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_6_i844_3_lut_4_lut.init = 16'hf808;
    LUT4 i22051_3_lut (.A(n21967), .B(n21968), .C(index_i[4]), .Z(n21969)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22051_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_8_i301_3_lut_4_lut (.A(n26927), .B(index_i[2]), .C(index_i[3]), 
         .D(n70), .Z(n301_adj_2679)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_8_i301_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_196_Mux_5_i636_4_lut (.A(n157_adj_2396), .B(n26794), .C(index_i[4]), 
         .D(index_i[3]), .Z(n636_adj_2453)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A (B ((D)+!C)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_5_i636_4_lut.init = 16'h3aca;
    LUT4 i15548_3_lut (.A(n26990), .B(n26993), .C(index_i[3]), .Z(n17812)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15548_3_lut.init = 16'hcaca;
    PFUMX i19292 (.BLUT(n21727), .ALUT(n21728), .C0(index_q[5]), .Z(n21729));
    LUT4 i15547_3_lut (.A(n26993), .B(n29489), .C(index_i[3]), .Z(n17811)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15547_3_lut.init = 16'hcaca;
    LUT4 i22054_3_lut (.A(n17814), .B(n17815), .C(index_i[4]), .Z(n17816)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22054_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_5_i507_3_lut (.A(n491_adj_2727), .B(n506_adj_2649), 
         .C(index_i[4]), .Z(n507)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_5_i507_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_5_i476_3_lut (.A(n460_adj_2716), .B(n475_adj_2728), 
         .C(index_i[4]), .Z(n476_adj_2449)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_5_i476_3_lut.init = 16'hcaca;
    PFUMX i24402 (.BLUT(n26294), .ALUT(n22754), .C0(index_i[8]), .Z(n26295));
    LUT4 mux_196_Mux_5_i413_3_lut (.A(n397_adj_2643), .B(n251_adj_2687), 
         .C(index_i[4]), .Z(n413_adj_2447)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_5_i413_3_lut.init = 16'hcaca;
    PFUMX i24728 (.BLUT(n27119), .ALUT(n27120), .C0(index_q[3]), .Z(n62_adj_2590));
    LUT4 i15566_3_lut (.A(n17828), .B(n17829), .C(index_i[4]), .Z(n17830)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15566_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_5_i125_3_lut (.A(n109_adj_2729), .B(n124_adj_2506), 
         .C(index_i[4]), .Z(n125_adj_2444)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_5_i125_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_5_i94_3_lut (.A(n653_adj_2642), .B(n635_adj_2730), 
         .C(index_i[4]), .Z(n94)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_5_i94_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_6_i700_3_lut_4_lut (.A(n27104), .B(index_q[3]), .C(index_q[4]), 
         .D(n684_adj_2256), .Z(n700_adj_2731)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_6_i700_3_lut_4_lut.init = 16'h9f90;
    L6MUX21 i20552 (.D0(n23006), .D1(n23007), .SD(index_i[5]), .Z(n23008));
    LUT4 mux_197_Mux_5_i397_3_lut (.A(n27098), .B(n204_adj_2732), .C(index_q[3]), 
         .Z(n397_adj_2512)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_5_i397_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut (.A(index_i[6]), .B(n26849), .C(index_i[5]), .D(index_i[4]), 
         .Z(n20362)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i1_4_lut.init = 16'hfffe;
    LUT4 i17578_4_lut (.A(n27045), .B(n892_adj_2451), .C(index_i[6]), 
         .D(index_i[5]), .Z(n19870)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D))))) */ ;
    defparam i17578_4_lut.init = 16'h3a35;
    PFUMX i19295 (.BLUT(n21730), .ALUT(n21731), .C0(index_q[5]), .Z(n21732));
    LUT4 i22420_3_lut (.A(n19870), .B(n20362), .C(index_i[7]), .Z(n22662)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22420_3_lut.init = 16'hcaca;
    L6MUX21 i20964 (.D0(n23404), .D1(n23405), .SD(index_q[5]), .Z(n23420));
    L6MUX21 i20965 (.D0(n23406), .D1(n23407), .SD(index_q[5]), .Z(n23421));
    L6MUX21 i20966 (.D0(n23408), .D1(n23409), .SD(index_q[5]), .Z(n23422));
    L6MUX21 i20967 (.D0(n23410), .D1(n23411), .SD(index_q[5]), .Z(n23423));
    LUT4 i1_3_lut_4_lut_adj_86 (.A(n26738), .B(index_i[5]), .C(index_i[8]), 
         .D(n19801), .Z(n20198)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i1_3_lut_4_lut_adj_86.init = 16'hfff8;
    PFUMX i19298 (.BLUT(n21733), .ALUT(n21734), .C0(index_q[5]), .Z(n21735));
    PFUMX i19301 (.BLUT(n21736), .ALUT(n21737), .C0(index_q[5]), .Z(n21738));
    LUT4 i19504_3_lut (.A(n29489), .B(n26990), .C(index_i[3]), .Z(n21941)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19504_3_lut.init = 16'hcaca;
    LUT4 i19503_3_lut (.A(n396), .B(n204), .C(index_i[3]), .Z(n21940)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19503_3_lut.init = 16'hcaca;
    L6MUX21 i20559 (.D0(n23013), .D1(n23014), .SD(index_i[5]), .Z(n23015));
    L6MUX21 i20968 (.D0(n23412), .D1(n23413), .SD(index_q[5]), .Z(n23424));
    PFUMX i19304 (.BLUT(n21739), .ALUT(n21740), .C0(index_q[5]), .Z(n21741));
    LUT4 index_i_0__bdd_4_lut_25303 (.A(index_i[0]), .B(index_i[3]), .C(index_i[1]), 
         .D(index_i[2]), .Z(n27192)) /* synthesis lut_function=(A (B (C)+!B !(C+!(D)))+!A !(B ((D)+!C)+!B !(C (D)+!C !(D)))) */ ;
    defparam index_i_0__bdd_4_lut_25303.init = 16'h92c1;
    PFUMX i19307 (.BLUT(n21742), .ALUT(n21743), .C0(index_q[5]), .Z(n21744));
    LUT4 index_i_4__bdd_2_lut_3_lut_4_lut (.A(n26927), .B(index_i[2]), .C(index_i[5]), 
         .D(n26995), .Z(n24733)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam index_i_4__bdd_2_lut_3_lut_4_lut.init = 16'h0f7f;
    LUT4 mux_196_Mux_8_i15_3_lut_4_lut (.A(n26927), .B(index_i[2]), .C(index_i[3]), 
         .D(n27003), .Z(n15_adj_2686)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_8_i15_3_lut_4_lut.init = 16'hf808;
    L6MUX21 i20969 (.D0(n23414), .D1(n23415), .SD(index_q[5]), .Z(n23425));
    PFUMX i19310 (.BLUT(n21745), .ALUT(n21746), .C0(index_q[5]), .Z(n21747));
    LUT4 mux_197_Mux_14_i511_4_lut_4_lut (.A(n26713), .B(index_q[7]), .C(index_q[8]), 
         .D(n254_adj_2717), .Z(n511_adj_2733)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (B (C+!(D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_14_i511_4_lut_4_lut.init = 16'h1c10;
    LUT4 index_q_1__bdd_4_lut_25966 (.A(index_q[1]), .B(index_q[0]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n27193)) /* synthesis lut_function=(!(A (B (D)+!B (C+!(D)))+!A !(B (C (D)+!C !(D))+!B !((D)+!C)))) */ ;
    defparam index_q_1__bdd_4_lut_25966.init = 16'h429c;
    LUT4 mux_197_Mux_5_i30_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n30_adj_2519)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A (B+!(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_5_i30_3_lut_4_lut.init = 16'hcc67;
    LUT4 mux_197_Mux_5_i506_3_lut (.A(n27072), .B(n29475), .C(index_q[3]), 
         .Z(n506_adj_2445)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_5_i506_3_lut.init = 16'hcaca;
    L6MUX21 i20970 (.D0(n23416), .D1(n23417), .SD(index_q[5]), .Z(n23426));
    LUT4 i22082_3_lut (.A(n286_adj_2523), .B(n317), .C(index_q[5]), .Z(n23175)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22082_3_lut.init = 16'hcaca;
    L6MUX21 i20566 (.D0(n23020), .D1(n23021), .SD(index_i[5]), .Z(n23022));
    LUT4 i19656_3_lut_3_lut_4_lut (.A(n26927), .B(index_i[2]), .C(n38), 
         .D(index_i[3]), .Z(n22093)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19656_3_lut_3_lut_4_lut.init = 16'hf077;
    LUT4 mux_196_Mux_8_i173_3_lut_3_lut_4_lut (.A(n26927), .B(index_i[2]), 
         .C(n954_adj_2706), .D(index_i[4]), .Z(n173_adj_2734)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C+!(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_8_i173_3_lut_3_lut_4_lut.init = 16'hf077;
    L6MUX21 i20971 (.D0(n23418), .D1(n23419), .SD(index_q[5]), .Z(n23427));
    PFUMX i24382 (.BLUT(n26265), .ALUT(n26263), .C0(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_2141[10]));
    LUT4 mux_197_Mux_5_i859_3_lut (.A(n851), .B(n27078), .C(index_q[3]), 
         .Z(n859_adj_2497)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_5_i859_3_lut.init = 16'hcaca;
    LUT4 i19489_3_lut (.A(n29491), .B(n308), .C(index_i[3]), .Z(n21926)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19489_3_lut.init = 16'hcaca;
    LUT4 i19488_3_lut (.A(n26932), .B(n26928), .C(index_i[3]), .Z(n21925)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19488_3_lut.init = 16'hcaca;
    LUT4 i11249_3_lut_3_lut_3_lut_rep_804 (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[0]), .Z(n29477)) /* synthesis lut_function=(!(A+!(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11249_3_lut_3_lut_3_lut_rep_804.init = 16'h4545;
    LUT4 i19740_3_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[2]), .C(index_q[0]), 
         .D(index_q[3]), .Z(n22177)) /* synthesis lut_function=(!(A ((D)+!B)+!A !(B (D)+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19740_3_lut_4_lut_4_lut.init = 16'h4588;
    LUT4 i9419_3_lut_4_lut_4_lut (.A(index_q[3]), .B(index_q[2]), .C(index_q[0]), 
         .D(index_q[1]), .Z(n844_adj_2625)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9419_3_lut_4_lut_4_lut.init = 16'hf00e;
    LUT4 i19486_3_lut (.A(n29491), .B(n26900), .C(index_i[3]), .Z(n21923)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19486_3_lut.init = 16'hcaca;
    LUT4 i19485_3_lut (.A(n27002), .B(n308), .C(index_i[3]), .Z(n21922)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19485_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_7_i173_3_lut (.A(n26932), .B(n26900), .C(index_i[3]), 
         .Z(n173_adj_2735)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_7_i173_3_lut.init = 16'hcaca;
    LUT4 i11625_3_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[3]), 
         .Z(n11119)) /* synthesis lut_function=(!((B (C))+!A)) */ ;
    defparam i11625_3_lut.init = 16'h2a2a;
    LUT4 i22097_3_lut (.A(n28806), .B(n26514), .C(index_q[5]), .Z(n22611)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22097_3_lut.init = 16'hcaca;
    PFUMX i24380 (.BLUT(n21577), .ALUT(n26261), .C0(index_q[7]), .Z(n26262));
    LUT4 i22101_3_lut (.A(n542_adj_2466), .B(n573_adj_2406), .C(index_q[5]), 
         .Z(n22605)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22101_3_lut.init = 16'hcaca;
    PFUMX i24371 (.BLUT(n26250), .ALUT(n26248), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2126[10]));
    LUT4 i21731_3_lut (.A(n21916), .B(n21917), .C(index_q[4]), .Z(n21918)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21731_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_5_i875_3_lut (.A(n26887), .B(n27102), .C(index_q[3]), 
         .Z(n875_adj_2494)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_5_i875_3_lut.init = 16'hcaca;
    LUT4 i15545_3_lut (.A(n27097), .B(n27098), .C(index_q[3]), .Z(n17809)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15545_3_lut.init = 16'hcaca;
    LUT4 i15544_3_lut (.A(n27098), .B(n27080), .C(index_q[3]), .Z(n17808)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i15544_3_lut.init = 16'hcaca;
    LUT4 i19477_3_lut (.A(n498), .B(n27077), .C(index_q[3]), .Z(n21914)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19477_3_lut.init = 16'hcaca;
    LUT4 i18984_3_lut (.A(n29485), .B(n29477), .C(index_q[3]), .Z(n21421)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18984_3_lut.init = 16'hcaca;
    LUT4 i19474_3_lut (.A(n498), .B(n27097), .C(index_q[3]), .Z(n21911)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19474_3_lut.init = 16'hcaca;
    LUT4 n269_bdd_3_lut_23453 (.A(n27095), .B(index_q[3]), .C(n27079), 
         .Z(n25208)) /* synthesis lut_function=(A (B+(C))+!A !(B+!(C))) */ ;
    defparam n269_bdd_3_lut_23453.init = 16'hb8b8;
    LUT4 i19473_3_lut (.A(n27080), .B(n356), .C(index_q[3]), .Z(n21910)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19473_3_lut.init = 16'hcaca;
    L6MUX21 i20013 (.D0(n21756), .D1(n21759), .SD(index_q[5]), .Z(n22469));
    LUT4 n285_bdd_3_lut (.A(n27095), .B(n29474), .C(index_q[3]), .Z(n25211)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n285_bdd_3_lut.init = 16'hacac;
    PFUMX i24369 (.BLUT(n21568), .ALUT(n26246), .C0(index_i[7]), .Z(n26247));
    LUT4 i20605_3_lut (.A(n27105), .B(n26887), .C(index_q[3]), .Z(n23061)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20605_3_lut.init = 16'hcaca;
    LUT4 i19494_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[2]), .C(index_i[1]), 
         .D(index_i[3]), .Z(n21931)) /* synthesis lut_function=(!(A (B+!((D)+!C))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19494_3_lut_4_lut_4_lut.init = 16'h6646;
    LUT4 mux_196_Mux_6_i636_4_lut_4_lut (.A(index_i[1]), .B(index_i[4]), 
         .C(n635_adj_2730), .D(n14441), .Z(n636_adj_2633)) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_6_i636_4_lut_4_lut.init = 16'hf3d1;
    L6MUX21 i20017 (.D0(n21765), .D1(n17810), .SD(index_q[5]), .Z(n22473));
    L6MUX21 i20018 (.D0(n21912), .D1(n11929), .SD(index_q[5]), .Z(n22474));
    PFUMX i20020 (.BLUT(n542_adj_2582), .ALUT(n573_adj_2736), .C0(index_q[5]), 
          .Z(n22476));
    PFUMX i20021 (.BLUT(n605_adj_2737), .ALUT(n636_adj_2738), .C0(index_q[5]), 
          .Z(n22477));
    LUT4 mux_197_Mux_0_i762_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n762)) /* synthesis lut_function=(A (B+!((D)+!C))+!A !(B (D)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i762_3_lut_4_lut_4_lut.init = 16'h98fc;
    LUT4 mux_197_Mux_2_i859_3_lut_4_lut (.A(index_q[0]), .B(n27063), .C(index_q[3]), 
         .D(n27095), .Z(n859_adj_2626)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_2_i859_3_lut_4_lut.init = 16'h4f40;
    LUT4 n21914_bdd_3_lut_23535 (.A(n29495), .B(n29494), .C(index_q[3]), 
         .Z(n25233)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n21914_bdd_3_lut_23535.init = 16'hcaca;
    LUT4 i19219_3_lut_3_lut (.A(n26748), .B(index_i[4]), .C(n46_adj_2714), 
         .Z(n21656)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;
    defparam i19219_3_lut_3_lut.init = 16'h7474;
    LUT4 n459_bdd_3_lut_23538 (.A(n27100), .B(n27081), .C(index_q[3]), 
         .Z(n25236)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n459_bdd_3_lut_23538.init = 16'hacac;
    LUT4 mux_197_Mux_0_i684_3_lut_4_lut (.A(index_q[0]), .B(n27063), .C(index_q[3]), 
         .D(n27087), .Z(n684)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i684_3_lut_4_lut.init = 16'h4f40;
    PFUMX i20022 (.BLUT(n669_adj_2577), .ALUT(n700_adj_2731), .C0(index_q[5]), 
          .Z(n22478));
    LUT4 mux_197_Mux_4_i61_3_lut (.A(n29493), .B(n27076), .C(index_q[3]), 
         .Z(n61)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_4_i61_3_lut.init = 16'hcaca;
    LUT4 i19020_3_lut_4_lut (.A(index_q[0]), .B(n27063), .C(index_q[3]), 
         .D(n27070), .Z(n21457)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19020_3_lut_4_lut.init = 16'hf404;
    PFUMX i20023 (.BLUT(n732_adj_2726), .ALUT(n21918), .C0(index_q[5]), 
          .Z(n22479));
    LUT4 mux_197_Mux_3_i62_3_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[4]), .D(n812), .Z(n62_adj_2739)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_3_i62_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_197_Mux_3_i94_3_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[4]), .D(n93_adj_2434), .Z(n94_adj_2740)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_3_i94_3_lut_4_lut.init = 16'hf606;
    PFUMX i24356 (.BLUT(n26229), .ALUT(n1022_adj_2357), .C0(index_i[9]), 
          .Z(quarter_wave_sample_register_i_15__N_2126[12]));
    PFUMX i20024 (.BLUT(n797_adj_2574), .ALUT(n828_adj_2573), .C0(index_q[5]), 
          .Z(n22480));
    LUT4 mux_197_Mux_4_i270_3_lut (.A(n27082), .B(n27072), .C(index_q[3]), 
         .Z(n270)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_4_i270_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_4_i15_3_lut (.A(n29475), .B(n588), .C(index_q[3]), 
         .Z(n15_adj_2456)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_4_i15_3_lut.init = 16'hcaca;
    PFUMX i20025 (.BLUT(n860_adj_2668), .ALUT(n891_adj_2568), .C0(index_q[5]), 
          .Z(n22481));
    LUT4 mux_197_Mux_4_i348_3_lut (.A(n27066), .B(n27080), .C(index_q[3]), 
         .Z(n348_adj_2741)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_4_i348_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_4_i684_3_lut (.A(n652), .B(n660), .C(index_q[3]), 
         .Z(n684_adj_2462)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_4_i684_3_lut.init = 16'hcaca;
    LUT4 i3507_2_lut_rep_595 (.A(index_q[0]), .B(index_q[1]), .Z(n26918)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i3507_2_lut_rep_595.init = 16'h6666;
    PFUMX i24352 (.BLUT(n254), .ALUT(n26223), .C0(index_i[8]), .Z(n26224));
    LUT4 mux_197_Mux_1_i732_3_lut (.A(n716_adj_2332), .B(n491_adj_2507), 
         .C(index_q[4]), .Z(n732_adj_2390)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_1_i732_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_3_i619_3_lut_rep_564_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n26887)) /* synthesis lut_function=(!(A (B)+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_3_i619_3_lut_rep_564_3_lut.init = 16'h6363;
    PFUMX i24350 (.BLUT(n26221), .ALUT(n1022), .C0(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_2141[12]));
    LUT4 mux_196_Mux_4_i205_3_lut_4_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[1]), .D(index_i[3]), .Z(n205)) /* synthesis lut_function=(!(A (B (D)+!B (C (D)))+!A !(B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_4_i205_3_lut_4_lut.init = 16'h46aa;
    LUT4 mux_197_Mux_1_i882_3_lut_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n882_adj_2742)) /* synthesis lut_function=(A ((C)+!B)+!A !((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_1_i882_3_lut_3_lut.init = 16'ha6a6;
    L6MUX21 i20604 (.D0(n23058), .D1(n23059), .SD(index_q[5]), .Z(n23060));
    L6MUX21 mux_196_Mux_7_i253 (.D0(n12050), .D1(n21927), .SD(index_i[5]), 
            .Z(n253_adj_2743)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    L6MUX21 i20611 (.D0(n23065), .D1(n23066), .SD(index_q[5]), .Z(n23067));
    PFUMX mux_196_Mux_7_i190 (.BLUT(n21924), .ALUT(n173_adj_2735), .C0(index_i[5]), 
          .Z(n190_adj_2744)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 mux_197_Mux_8_i124_3_lut_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n124)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C+!(D)))+!A (B (C (D)+!C !(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_8_i124_3_lut_3_lut_4_lut_4_lut.init = 16'h07c1;
    PFUMX mux_196_Mux_8_i764 (.BLUT(n716_adj_2280), .ALUT(n732_adj_2561), 
          .C0(n22372), .Z(n764_adj_2333)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 mux_197_Mux_0_i939_4_lut (.A(n588), .B(n27071), .C(index_q[3]), 
         .D(index_q[2]), .Z(n939)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i939_4_lut.init = 16'hfaca;
    LUT4 mux_197_Mux_0_i739_3_lut_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n588)) /* synthesis lut_function=(!(A (B+(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i739_3_lut_3_lut.init = 16'h5656;
    PFUMX mux_196_Mux_8_i574 (.BLUT(n542), .ALUT(n12046), .C0(index_i[5]), 
          .Z(n574_adj_2328)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 i21614_3_lut (.A(n21409), .B(n21410), .C(index_q[4]), .Z(n21411)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21614_3_lut.init = 16'hcaca;
    LUT4 i11267_3_lut (.A(index_q[3]), .B(index_q[1]), .C(index_q[0]), 
         .Z(n13941)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11267_3_lut.init = 16'hc8c8;
    LUT4 mux_197_Mux_3_i348_3_lut (.A(n27081), .B(n27077), .C(index_q[3]), 
         .Z(n348_adj_2745)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_3_i348_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_5_i828_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[4]), .D(n26994), .Z(n828_adj_2746)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_5_i828_4_lut_4_lut.init = 16'hc66c;
    LUT4 i22170_3_lut (.A(n924_adj_2747), .B(n955_adj_2339), .C(index_q[5]), 
         .Z(n22482)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22170_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_6_i844_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n844_adj_2667)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (B (C)+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_6_i844_3_lut_4_lut_4_lut.init = 16'hc1e0;
    L6MUX21 i20618 (.D0(n23072), .D1(n23073), .SD(index_q[5]), .Z(n23074));
    LUT4 i9600_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n12165)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B ((D)+!C)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9600_3_lut_4_lut_4_lut.init = 16'h6c3c;
    LUT4 mux_197_Mux_3_i908_3_lut (.A(n27070), .B(n27076), .C(index_q[3]), 
         .Z(n908_adj_2420)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_3_i908_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_6_i660_3_lut_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n660)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_6_i660_3_lut_3_lut.init = 16'hc6c6;
    LUT4 mux_197_Mux_3_i507_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[4]), .D(n491_adj_2365), .Z(n507_adj_2748)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_3_i507_3_lut_4_lut.init = 16'h6f60;
    L6MUX21 i20625 (.D0(n23079), .D1(n23080), .SD(index_q[5]), .Z(n23081));
    LUT4 i22446_3_lut (.A(n25271), .B(n22471), .C(index_q[6]), .Z(n22485)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22446_3_lut.init = 16'hcaca;
    LUT4 i20328_3_lut (.A(n22778), .B(n22779), .C(index_i[7]), .Z(n22784)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20328_3_lut.init = 16'hcaca;
    LUT4 i20323_3_lut (.A(n22768), .B(n22769), .C(index_i[6]), .Z(n22779)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20323_3_lut.init = 16'hcaca;
    PFUMX i20626 (.BLUT(n12016), .ALUT(n62_adj_2749), .C0(index_q[5]), 
          .Z(n23082));
    LUT4 i20388_3_lut (.A(n22836), .B(n22837), .C(index_i[7]), .Z(n22844)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20388_3_lut.init = 16'hcaca;
    LUT4 i20381_3_lut (.A(n22822), .B(n25607), .C(index_i[6]), .Z(n22837)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20381_3_lut.init = 16'hcaca;
    LUT4 i20390_3_lut (.A(n22840), .B(n22841), .C(index_i[7]), .Z(n22846)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20390_3_lut.init = 16'hcaca;
    LUT4 i20384_3_lut (.A(n25613), .B(n22829), .C(index_i[6]), .Z(n22840)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20384_3_lut.init = 16'hcaca;
    PFUMX i20627 (.BLUT(n94_adj_2553), .ALUT(n22134), .C0(index_q[5]), 
          .Z(n23083));
    LUT4 i20650_3_lut (.A(n23098), .B(n23099), .C(index_q[7]), .Z(n23106)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20650_3_lut.init = 16'hcaca;
    LUT4 i20643_3_lut (.A(n23084), .B(n25970), .C(index_q[6]), .Z(n23099)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20643_3_lut.init = 16'hcaca;
    LUT4 i20652_3_lut (.A(n23102), .B(n23103), .C(index_q[7]), .Z(n23108)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20652_3_lut.init = 16'hcaca;
    LUT4 i20646_3_lut (.A(n26016), .B(n23091), .C(index_q[6]), .Z(n23102)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20646_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_6_i732_3_lut_4_lut (.A(n27001), .B(index_i[3]), .C(index_i[4]), 
         .D(n731_adj_2501), .Z(n732_adj_2637)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_6_i732_3_lut_4_lut.init = 16'hf909;
    LUT4 i20198_3_lut (.A(n22648), .B(n22649), .C(index_q[7]), .Z(n22654)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20198_3_lut.init = 16'hcaca;
    LUT4 i20193_3_lut (.A(n22638), .B(n22639), .C(index_q[6]), .Z(n22649)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20193_3_lut.init = 16'hcaca;
    LUT4 i20246_3_lut (.A(n22691), .B(n22692), .C(index_i[6]), .Z(n22702)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20246_3_lut.init = 16'hcaca;
    LUT4 i20357_3_lut (.A(n24908), .B(n22806), .C(index_i[7]), .Z(n22813)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20357_3_lut.init = 16'hcaca;
    LUT4 i8814_4_lut_4_lut (.A(index_i[3]), .B(index_i[0]), .C(index_i[1]), 
         .D(index_i[2]), .Z(n11334)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (D)+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i8814_4_lut_4_lut.init = 16'h0bf4;
    LUT4 i20395_3_lut (.A(n24809), .B(n29045), .C(index_q[7]), .Z(n22851)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20395_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_6_i700_3_lut_4_lut (.A(n27001), .B(index_i[3]), .C(index_i[4]), 
         .D(n684_adj_2708), .Z(n700_adj_2635)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(B (C+!(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_6_i700_3_lut_4_lut.init = 16'h9f90;
    LUT4 i11585_4_lut_4_lut (.A(index_i[3]), .B(index_i[2]), .C(index_i[0]), 
         .D(index_i[1]), .Z(n875_adj_2677)) /* synthesis lut_function=((B (C)+!B (D))+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11585_4_lut_4_lut.init = 16'hf7d5;
    L6MUX21 i20628 (.D0(n22140), .D1(n22143), .SD(index_q[5]), .Z(n23084));
    LUT4 i22667_2_lut (.A(index_q[3]), .B(index_q[2]), .Z(n22413)) /* synthesis lut_function=(A+!(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i22667_2_lut.init = 16'hbbbb;
    LUT4 i20539_3_lut (.A(n25102), .B(n22988), .C(index_q[7]), .Z(n22995)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20539_3_lut.init = 16'hcaca;
    LUT4 i21039_3_lut (.A(n23492), .B(n23493), .C(index_i[7]), .Z(n23495)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21039_3_lut.init = 16'hcaca;
    LUT4 i20446_3_lut_4_lut_3_lut (.A(index_i[3]), .B(index_i[4]), .C(n26836), 
         .Z(n22902)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20446_3_lut_4_lut_3_lut.init = 16'h6464;
    LUT4 mux_196_Mux_1_i987_3_lut_4_lut_4_lut (.A(index_i[3]), .B(n986_adj_2699), 
         .C(index_i[4]), .D(n29468), .Z(n987)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_1_i987_3_lut_4_lut_4_lut.init = 16'hc5c0;
    LUT4 mux_197_Mux_0_i923_3_lut (.A(n27062), .B(n27086), .C(index_q[3]), 
         .Z(n923)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i923_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_6_i251_3_lut_4_lut (.A(n26848), .B(index_i[2]), .C(index_i[3]), 
         .D(n27023), .Z(n251_adj_2687)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_6_i251_3_lut_4_lut.init = 16'hf606;
    PFUMX i24345 (.BLUT(n254_adj_2255), .ALUT(n26215), .C0(index_q[8]), 
          .Z(n26216));
    LUT4 i19264_4_lut_3_lut (.A(index_i[3]), .B(index_i[4]), .C(n26876), 
         .Z(n21701)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19264_4_lut_3_lut.init = 16'h6565;
    LUT4 i19644_3_lut_4_lut (.A(index_i[0]), .B(index_i[2]), .C(index_i[1]), 
         .D(index_i[3]), .Z(n22081)) /* synthesis lut_function=(A (B (D)+!B (C+(D)))+!A !(B (D)+!B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19644_3_lut_4_lut.init = 16'haa65;
    PFUMX i20630 (.BLUT(n22149), .ALUT(n317_adj_2409), .C0(index_q[5]), 
          .Z(n23086));
    LUT4 i19330_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21767)) /* synthesis lut_function=(!(A ((D)+!C)+!A !(B ((D)+!C)+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19330_3_lut_3_lut_4_lut.init = 16'h55a4;
    PFUMX i20631 (.BLUT(n349_adj_2537), .ALUT(n22152), .C0(index_q[5]), 
          .Z(n23087));
    LUT4 mux_196_Mux_2_i221_4_lut_4_lut (.A(index_i[3]), .B(index_i[4]), 
         .C(n26876), .D(n26759), .Z(n221_adj_2563)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (B+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_2_i221_4_lut_4_lut.init = 16'hf7c4;
    LUT4 i9487_3_lut_3_lut (.A(index_i[3]), .B(index_i[4]), .C(n12047), 
         .Z(n12048)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9487_3_lut_3_lut.init = 16'h7474;
    LUT4 i5940_2_lut_rep_599 (.A(index_i[0]), .B(index_i[2]), .Z(n26922)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i5940_2_lut_rep_599.init = 16'h6666;
    LUT4 i22379_3_lut (.A(n22985), .B(n25817), .C(index_q[6]), .Z(n22994)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22379_3_lut.init = 16'hcaca;
    LUT4 i20116_3_lut (.A(n22561), .B(n22562), .C(index_q[6]), .Z(n22572)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20116_3_lut.init = 16'hcaca;
    LUT4 i9512_3_lut_4_lut (.A(n26848), .B(index_i[2]), .C(n27045), .D(n27023), 
         .Z(n444_adj_2448)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9512_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_196_Mux_6_i157_3_lut_4_lut (.A(n26848), .B(index_i[2]), .C(index_i[3]), 
         .D(n26977), .Z(n157_adj_2531)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_6_i157_3_lut_4_lut.init = 16'hf606;
    LUT4 i19030_3_lut_4_lut (.A(n27101), .B(index_q[2]), .C(index_q[3]), 
         .D(n851), .Z(n21467)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19030_3_lut_4_lut.init = 16'hf202;
    LUT4 i19038_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21475)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+(D)))+!A !(B (D)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19038_3_lut_4_lut_4_lut.init = 16'h99c7;
    LUT4 i15551_3_lut_3_lut (.A(index_i[0]), .B(index_i[2]), .C(index_i[3]), 
         .Z(n17815)) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i15551_3_lut_3_lut.init = 16'h6a6a;
    LUT4 mux_196_Mux_4_i349_3_lut_4_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[4]), .D(n348_adj_2675), .Z(n349)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_4_i349_3_lut_4_lut.init = 16'hf606;
    PFUMX i23263 (.BLUT(n24999), .ALUT(n26882), .C0(index_i[4]), .Z(n25000));
    LUT4 mux_196_Mux_4_i828_3_lut_4_lut (.A(index_i[4]), .B(index_i[3]), 
         .C(n812_adj_2273), .D(n26992), .Z(n828_adj_2505)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_4_i828_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_197_Mux_7_i506_3_lut_4_lut (.A(n27101), .B(index_q[2]), .C(index_q[3]), 
         .D(n27102), .Z(n506_adj_2750)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_7_i506_3_lut_4_lut.init = 16'h2f20;
    PFUMX i26204 (.BLUT(n29163), .ALUT(n29162), .C0(index_i[3]), .Z(n29164));
    LUT4 mux_196_Mux_5_i797_3_lut_4_lut (.A(index_i[4]), .B(index_i[3]), 
         .C(n27137), .D(n27024), .Z(n797_adj_2458)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_5_i797_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n389_bdd_3_lut_24616_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n25635)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C))+!A (B (C (D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n389_bdd_3_lut_24616_3_lut_4_lut.init = 16'h0fc7;
    LUT4 mux_197_Mux_0_i653_3_lut (.A(n26887), .B(n27072), .C(index_q[3]), 
         .Z(n653)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i653_3_lut.init = 16'hcaca;
    PFUMX i26201 (.BLUT(n29159), .ALUT(n29158), .C0(index_i[2]), .Z(n29160));
    LUT4 mux_196_Mux_1_i763_3_lut_4_lut (.A(index_i[4]), .B(index_i[3]), 
         .C(n27208), .D(n27024), .Z(n763_adj_2300)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_1_i763_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i12190_2_lut_rep_600 (.A(index_i[2]), .B(index_i[0]), .Z(n26923)) /* synthesis lut_function=(A (B)) */ ;
    defparam i12190_2_lut_rep_600.init = 16'h8888;
    LUT4 index_i_8__bdd_3_lut_24659_then_4_lut (.A(index_i[4]), .B(index_i[6]), 
         .C(index_i[5]), .D(n26781), .Z(n27198)) /* synthesis lut_function=(!(A (B (C+(D)))+!A (B (C)))) */ ;
    defparam index_i_8__bdd_3_lut_24659_then_4_lut.init = 16'h373f;
    LUT4 mux_196_Mux_4_i747_3_lut_4_lut (.A(n26848), .B(index_i[2]), .C(index_i[3]), 
         .D(n27032), .Z(n747_adj_2355)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_4_i747_3_lut_4_lut.init = 16'hf606;
    LUT4 i20203_3_lut (.A(n24787), .B(n29165), .C(index_i[7]), .Z(n22659)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20203_3_lut.init = 16'hcaca;
    LUT4 i20211_3_lut (.A(n190_adj_2744), .B(n253_adj_2743), .C(index_i[6]), 
         .Z(n22667)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20211_3_lut.init = 16'hcaca;
    LUT4 i20212_3_lut (.A(n23022), .B(n21681), .C(index_i[6]), .Z(n22668)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20212_3_lut.init = 16'hcaca;
    L6MUX21 i20632 (.D0(n22158), .D1(n22161), .SD(index_q[5]), .Z(n23088));
    L6MUX21 i20633 (.D0(n22167), .D1(n22170), .SD(index_q[5]), .Z(n23089));
    LUT4 i18960_3_lut_4_lut (.A(index_q[0]), .B(n27090), .C(index_q[3]), 
         .D(n29493), .Z(n21397)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A ((D)+!C)) */ ;
    defparam i18960_3_lut_4_lut.init = 16'hfd0d;
    L6MUX21 i20635 (.D0(n22179), .D1(n636_adj_2550), .SD(index_q[5]), 
            .Z(n23091));
    PFUMX i20636 (.BLUT(n21768), .ALUT(n700_adj_2492), .C0(index_q[5]), 
          .Z(n23092));
    LUT4 i20347_4_lut_4_lut (.A(index_i[4]), .B(index_i[5]), .C(n27125), 
         .D(n908_adj_2358), .Z(n22803)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam i20347_4_lut_4_lut.init = 16'hd1c0;
    PFUMX i23244 (.BLUT(n24974), .ALUT(n26922), .C0(index_i[5]), .Z(n24975));
    PFUMX i23242 (.BLUT(n27021), .ALUT(n24972), .C0(index_i[2]), .Z(n24973));
    L6MUX21 i23240 (.D0(n24970), .D1(n24967), .SD(index_i[5]), .Z(n24971));
    LUT4 index_i_8__bdd_3_lut_24659_else_4_lut (.A(n26835), .B(index_i[4]), 
         .C(index_i[6]), .D(index_i[5]), .Z(n27197)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;
    defparam index_i_8__bdd_3_lut_24659_else_4_lut.init = 16'hf080;
    L6MUX21 i20638 (.D0(n21771), .D1(n21774), .SD(index_q[5]), .Z(n23094));
    PFUMX i23238 (.BLUT(n24969), .ALUT(n475_adj_2704), .C0(index_i[4]), 
          .Z(n24970));
    PFUMX i20640 (.BLUT(n924_adj_2529), .ALUT(n21780), .C0(index_q[5]), 
          .Z(n23096));
    PFUMX i20641 (.BLUT(n987_adj_2751), .ALUT(n21783), .C0(index_q[5]), 
          .Z(n23097));
    PFUMX i26117 (.BLUT(n29043), .ALUT(n29042), .C0(index_q[3]), .Z(n29044));
    LUT4 i22672_2_lut_rep_602 (.A(index_i[4]), .B(index_i[3]), .Z(n26925)) /* synthesis lut_function=((B)+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i22672_2_lut_rep_602.init = 16'hdddd;
    PFUMX i26115 (.BLUT(n29039), .ALUT(n29038), .C0(index_q[2]), .Z(n29040));
    LUT4 mux_196_Mux_3_i797_3_lut_4_lut (.A(index_i[4]), .B(index_i[3]), 
         .C(n796_adj_2502), .D(n70), .Z(n797)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_3_i797_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i20873_3_lut_4_lut_4_lut (.A(n26849), .B(index_i[4]), .C(index_i[5]), 
         .D(n26781), .Z(n23329)) /* synthesis lut_function=(A ((C+!(D))+!B)+!A (B (C+!(D))+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20873_3_lut_4_lut_4_lut.init = 16'he3ef;
    LUT4 i11263_2_lut_rep_767 (.A(index_q[1]), .B(index_q[2]), .Z(n27090)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11263_2_lut_rep_767.init = 16'h8888;
    LUT4 i21038_3_lut (.A(n23490), .B(n23491), .C(index_i[7]), .Z(n23494)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21038_3_lut.init = 16'hcaca;
    PFUMX i20095 (.BLUT(n31_adj_2520), .ALUT(n21984), .C0(index_q[5]), 
          .Z(n22551));
    LUT4 i9557_4_lut_4_lut (.A(n27092), .B(index_q[1]), .C(index_q[3]), 
         .D(n20689), .Z(n12119)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A (B (C)+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9557_4_lut_4_lut.init = 16'h0e3e;
    PFUMX i23235 (.BLUT(n24966), .ALUT(n24965), .C0(index_i[4]), .Z(n24967));
    LUT4 mux_197_Mux_5_i491_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n491_adj_2507)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A !(B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_5_i491_3_lut_4_lut_4_lut.init = 16'ha54a;
    PFUMX i20096 (.BLUT(n94_adj_2518), .ALUT(n125_adj_2516), .C0(index_q[5]), 
          .Z(n22552));
    LUT4 n25269_bdd_3_lut (.A(n25269), .B(n157_adj_2752), .C(index_q[4]), 
         .Z(n25270)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n25269_bdd_3_lut.init = 16'hcaca;
    L6MUX21 i23232 (.D0(n24963), .D1(n24961), .SD(index_i[5]), .Z(n24964));
    PFUMX i20097 (.BLUT(n17824), .ALUT(n14460), .C0(index_q[5]), .Z(n22553));
    PFUMX i23230 (.BLUT(n24962), .ALUT(n285_adj_2380), .C0(index_i[4]), 
          .Z(n24963));
    LUT4 index_q_8__bdd_3_lut_then_4_lut (.A(index_q[4]), .B(index_q[6]), 
         .C(index_q[5]), .D(n26767), .Z(n27201)) /* synthesis lut_function=(!(A (B (C+(D)))+!A (B (C)))) */ ;
    defparam index_q_8__bdd_3_lut_then_4_lut.init = 16'h373f;
    LUT4 mux_196_Mux_1_i62_3_lut_4_lut (.A(index_i[0]), .B(index_i[3]), 
         .C(index_i[2]), .D(index_i[4]), .Z(n62_adj_2753)) /* synthesis lut_function=(A (B (D)+!B ((D)+!C))+!A !(B (D)+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_1_i62_3_lut_4_lut.init = 16'haa56;
    L6MUX21 i20099 (.D0(n21987), .D1(n21990), .SD(index_q[5]), .Z(n22555));
    LUT4 mux_197_Mux_0_i572_3_lut_4_lut (.A(n27092), .B(index_q[1]), .C(index_q[3]), 
         .D(n29494), .Z(n572)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i572_3_lut_4_lut.init = 16'hefe0;
    L6MUX21 i20100 (.D0(n21393), .D1(n21396), .SD(index_q[5]), .Z(n22556));
    PFUMX i20101 (.BLUT(n413_adj_2513), .ALUT(n444_adj_2369), .C0(index_q[5]), 
          .Z(n22557));
    PFUMX i20102 (.BLUT(n476_adj_2510), .ALUT(n507_adj_2508), .C0(index_q[5]), 
          .Z(n22558));
    LUT4 mux_196_Mux_4_i252_4_lut_4_lut (.A(index_i[0]), .B(index_i[3]), 
         .C(n27048), .D(index_i[4]), .Z(n252_adj_2486)) /* synthesis lut_function=(!(A (B (D)+!B !(D))+!A !(B ((D)+!C)+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_4_i252_4_lut_4_lut.init = 16'h669d;
    PFUMX mux_197_Mux_1_i891 (.BLUT(n882_adj_2742), .ALUT(n890_adj_2754), 
          .C0(n26911), .Z(n891_adj_2394)) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 index_q_3__bdd_3_lut_22851_3_lut_4_lut (.A(n27092), .B(index_q[1]), 
         .C(index_q[4]), .D(index_q[3]), .Z(n24491)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam index_q_3__bdd_3_lut_22851_3_lut_4_lut.init = 16'hf10f;
    LUT4 i20168_3_lut (.A(n22619), .B(n22620), .C(index_q[7]), .Z(n22624)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20168_3_lut.init = 16'hcaca;
    PFUMX i20103 (.BLUT(n17788), .ALUT(n573_adj_2755), .C0(index_q[5]), 
          .Z(n22559));
    LUT4 i11475_2_lut_rep_414_3_lut_4_lut (.A(n27092), .B(index_q[1]), .C(index_q[4]), 
         .D(index_q[3]), .Z(n26737)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11475_2_lut_rep_414_3_lut_4_lut.init = 16'hfef0;
    LUT4 i19284_4_lut_4_lut_3_lut_4_lut (.A(n27092), .B(index_q[1]), .C(index_q[4]), 
         .D(index_q[3]), .Z(n21721)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19284_4_lut_4_lut_3_lut_4_lut.init = 16'h11ef;
    LUT4 i11498_2_lut_rep_659 (.A(index_i[0]), .B(index_i[1]), .Z(n26982)) /* synthesis lut_function=((B)+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11498_2_lut_rep_659.init = 16'hdddd;
    PFUMX i23228 (.BLUT(n24960), .ALUT(n24959), .C0(index_i[4]), .Z(n24961));
    LUT4 n400_bdd_3_lut_24707_4_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .Z(n25491)) /* synthesis lut_function=(!(A (B)+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n400_bdd_3_lut_24707_4_lut_3_lut.init = 16'h6262;
    LUT4 mux_196_Mux_0_i908_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n908_adj_2694)) /* synthesis lut_function=(!(A (B (C (D))+!B !(D))+!A (B+((D)+!C)))) */ ;
    defparam mux_196_Mux_0_i908_3_lut_4_lut_4_lut.init = 16'h2a98;
    PFUMX i20104 (.BLUT(n605_adj_2756), .ALUT(n636_adj_2500), .C0(index_q[5]), 
          .Z(n22560));
    LUT4 i11629_2_lut_rep_548_3_lut (.A(index_q[1]), .B(index_q[2]), .C(index_q[0]), 
         .Z(n26871)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11629_2_lut_rep_548_3_lut.init = 16'h8080;
    PFUMX i20105 (.BLUT(n21399), .ALUT(n700_adj_2757), .C0(index_q[5]), 
          .Z(n22561));
    LUT4 mux_197_Mux_3_i796_3_lut_3_lut (.A(index_q[4]), .B(n781_adj_2600), 
         .C(index_q[2]), .Z(n796_adj_2372)) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam mux_197_Mux_3_i796_3_lut_3_lut.init = 16'he4e4;
    LUT4 i9554_4_lut_4_lut (.A(index_q[4]), .B(n22401), .C(n27214), .D(n27088), 
         .Z(n12116)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam i9554_4_lut_4_lut.init = 16'hf4b0;
    LUT4 i20468_3_lut_4_lut (.A(n26854), .B(index_q[3]), .C(index_q[4]), 
         .D(n26817), .Z(n22924)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20468_3_lut_4_lut.init = 16'hfe0e;
    LUT4 i20529_4_lut_4_lut (.A(index_q[4]), .B(index_q[5]), .C(n27180), 
         .D(n908_adj_2408), .Z(n22985)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(49[8] 89[6])
    defparam i20529_4_lut_4_lut.init = 16'hd1c0;
    LUT4 i12208_2_lut_rep_604 (.A(index_i[0]), .B(index_i[1]), .Z(n26927)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i12208_2_lut_rep_604.init = 16'heeee;
    L6MUX21 i20106 (.D0(n732_adj_2700), .D1(n21402), .SD(index_q[5]), 
            .Z(n22562));
    PFUMX i20107 (.BLUT(n797_adj_2517), .ALUT(n828_adj_2746), .C0(index_q[5]), 
          .Z(n22563));
    LUT4 index_q_8__bdd_3_lut_else_4_lut (.A(n26859), .B(index_q[4]), .C(index_q[6]), 
         .D(index_q[5]), .Z(n27200)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;
    defparam index_q_8__bdd_3_lut_else_4_lut.init = 16'hf080;
    PFUMX i20108 (.BLUT(n860_adj_2498), .ALUT(n891_adj_2495), .C0(index_q[5]), 
          .Z(n22564));
    LUT4 n173_bdd_4_lut (.A(n173_adj_2734), .B(n70), .C(index_i[4]), .D(index_i[3]), 
         .Z(n24641)) /* synthesis lut_function=(A (B+(C+!(D)))+!A !((C+!(D))+!B)) */ ;
    defparam n173_bdd_4_lut.init = 16'hacaa;
    LUT4 i20549_3_lut (.A(n26999), .B(n27002), .C(index_i[3]), .Z(n23005)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20549_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_7_i691_3_lut_rep_677 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27000)) /* synthesis lut_function=(!(A (B (C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_7_i691_3_lut_rep_677.init = 16'h7e7e;
    LUT4 i11245_2_lut_rep_778 (.A(index_q[0]), .B(index_q[1]), .Z(n27101)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11245_2_lut_rep_778.init = 16'heeee;
    LUT4 mux_196_Mux_7_i572_3_lut_3_lut_rep_486_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n26809)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)+!C !(D)))) */ ;
    defparam mux_196_Mux_7_i572_3_lut_3_lut_rep_486_4_lut.init = 16'hfe01;
    LUT4 i11369_2_lut_rep_458_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n26781)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i11369_2_lut_rep_458_3_lut_4_lut.init = 16'hfef0;
    LUT4 n26247_bdd_3_lut_3_lut (.A(n1021), .B(index_i[8]), .C(n26247), 
         .Z(n26248)) /* synthesis lut_function=(A (B+(C))+!A !(B+!(C))) */ ;
    defparam n26247_bdd_3_lut_3_lut.init = 16'hb8b8;
    LUT4 mux_197_Mux_3_i828_3_lut_3_lut_4_lut (.A(n26854), .B(index_q[3]), 
         .C(n157_adj_2437), .D(index_q[4]), .Z(n828_adj_2429)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_3_i828_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 mux_196_Mux_7_i924_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[4]), .D(n27035), .Z(n924_adj_2758)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B ((D)+!C))) */ ;
    defparam mux_196_Mux_7_i924_3_lut_3_lut_4_lut.init = 16'hf10f;
    LUT4 mux_196_Mux_2_i931_3_lut_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n931_adj_2602)) /* synthesis lut_function=(!(A (B (C))+!A (B (C)+!B !(C)))) */ ;
    defparam mux_196_Mux_2_i931_3_lut_3_lut_3_lut.init = 16'h3e3e;
    LUT4 index_i_5__bdd_3_lut_23860_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n25577)) /* synthesis lut_function=(A (B (C)+!B (C+(D)))+!A (B (C)+!B !(C (D)+!C !(D)))) */ ;
    defparam index_i_5__bdd_3_lut_23860_4_lut_4_lut_4_lut.init = 16'he3f0;
    LUT4 i11470_2_lut_rep_559_3_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .Z(n26882)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i11470_2_lut_rep_559_3_lut.init = 16'he0e0;
    LUT4 i20548_3_lut (.A(n38), .B(n29490), .C(index_i[3]), .Z(n23004)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20548_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_8_i397_3_lut_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n397_adj_2392)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B ((D)+!C))) */ ;
    defparam mux_196_Mux_8_i397_3_lut_3_lut_3_lut_4_lut.init = 16'hf10f;
    LUT4 i5810_2_lut_rep_698 (.A(index_i[0]), .B(index_i[1]), .Z(n27021)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i5810_2_lut_rep_698.init = 16'h6666;
    LUT4 i11435_2_lut_rep_443_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[4]), .D(n27035), .Z(n26766)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i11435_2_lut_rep_443_3_lut_4_lut.init = 16'hfef0;
    LUT4 n526_bdd_3_lut_24373_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n25605)) /* synthesis lut_function=(!(A (B)+!A !(B (C+(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n526_bdd_3_lut_24373_4_lut_4_lut_4_lut.init = 16'h6663;
    LUT4 mux_196_Mux_3_i30_3_lut_3_lut_4_lut_4_lut_3_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[2]), .D(index_i[3]), .Z(n30_adj_2481)) /* synthesis lut_function=(A (C)+!A (B (C)+!B ((D)+!C))) */ ;
    defparam mux_196_Mux_3_i30_3_lut_3_lut_4_lut_4_lut_3_lut_4_lut.init = 16'hf1e1;
    LUT4 i12375_1_lut_rep_408_2_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n26731)) /* synthesis lut_function=(!(A (C+(D))+!A (B (C+(D))+!B (C)))) */ ;
    defparam i12375_1_lut_rep_408_2_lut_3_lut_4_lut.init = 16'h010f;
    LUT4 mux_196_Mux_1_i882_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n882)) /* synthesis lut_function=(A ((C)+!B)+!A !((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_1_i882_3_lut_3_lut.init = 16'ha6a6;
    LUT4 mux_196_Mux_8_i46_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n46_adj_2714)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (B (C)+!B !(C (D)+!C !(D)))) */ ;
    defparam mux_196_Mux_8_i46_3_lut_4_lut_4_lut_4_lut.init = 16'hc1f0;
    LUT4 mux_197_Mux_0_i14_3_lut_rep_739_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n27062)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i14_3_lut_rep_739_3_lut.init = 16'he3e3;
    LUT4 mux_196_Mux_0_i333_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n333_adj_2759)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B (D))) */ ;
    defparam mux_196_Mux_0_i333_3_lut_3_lut_4_lut.init = 16'hf10e;
    LUT4 i19602_3_lut_3_lut_4_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n22039)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B !((D)+!C)))) */ ;
    defparam i19602_3_lut_3_lut_4_lut_3_lut_4_lut.init = 16'h11ef;
    LUT4 i9510_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(n27035), .D(index_i[4]), .Z(n221_adj_2760)) /* synthesis lut_function=(!(A (B)+!A (B (C+(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9510_3_lut_4_lut_4_lut_4_lut.init = 16'h3336;
    LUT4 mux_197_Mux_9_i30_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[0]), .D(index_q[3]), .Z(n30_adj_2696)) /* synthesis lut_function=(A (B (C (D))+!B !(D))+!A !(B+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_9_i30_3_lut_4_lut_4_lut_4_lut.init = 16'h8033;
    LUT4 i9593_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n12158)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B ((D)+!C)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9593_3_lut_4_lut_4_lut.init = 16'h6c3c;
    LUT4 mux_196_Mux_2_i731_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n731_adj_2702)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_2_i731_3_lut_4_lut_4_lut.init = 16'h6cc6;
    LUT4 mux_196_Mux_3_i157_3_lut_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n157_adj_2319)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B !(C+(D))))) */ ;
    defparam mux_196_Mux_3_i157_3_lut_3_lut_3_lut_4_lut.init = 16'h1ff0;
    LUT4 mux_196_Mux_5_i356_3_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n396)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_5_i356_3_lut_4_lut_3_lut.init = 16'h6d6d;
    LUT4 i19639_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n22076)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (B (C+!(D))+!B (D))) */ ;
    defparam i19639_3_lut_4_lut_4_lut_4_lut.init = 16'hf1cc;
    LUT4 i11556_2_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n635)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A (B (C+!(D))+!B (C+(D)))) */ ;
    defparam i11556_2_lut_4_lut_4_lut.init = 16'hf1fc;
    LUT4 i9496_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n526)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+(D)))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9496_3_lut_4_lut_4_lut.init = 16'h666c;
    LUT4 i19629_3_lut_4_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n22066)) /* synthesis lut_function=(A (B (D)+!B ((D)+!C))+!A (B (D)+!B (C+!(D)))) */ ;
    defparam i19629_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'hfe13;
    LUT4 mux_196_Mux_7_i29_3_lut_rep_678 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27001)) /* synthesis lut_function=(A (B+!(C))+!A !((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_7_i29_3_lut_rep_678.init = 16'h8e8e;
    LUT4 i11427_2_lut_rep_575 (.A(index_i[2]), .B(index_i[3]), .Z(n26898)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11427_2_lut_rep_575.init = 16'heeee;
    LUT4 n21326_bdd_3_lut_23555 (.A(n26992), .B(n27022), .C(index_i[3]), 
         .Z(n25319)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n21326_bdd_3_lut_23555.init = 16'hcaca;
    LUT4 i18973_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .D(index_q[0]), .Z(n21410)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C (D)+!C !(D)))+!A !(B (D)+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18973_3_lut_4_lut_4_lut_4_lut.init = 16'h7c03;
    LUT4 mux_196_Mux_7_i235_3_lut_rep_605 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26928)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C)+!B !(C))) */ ;
    defparam mux_196_Mux_7_i235_3_lut_rep_605.init = 16'he3e3;
    LUT4 i19662_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n22099)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C (D)))+!A (B (C+(D))+!B !(C)))) */ ;
    defparam i19662_4_lut_4_lut_4_lut.init = 16'h301c;
    LUT4 mux_196_Mux_0_i699_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n699_adj_2559)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (D))+!A (B (C+!(D))+!B !(C+!(D))))) */ ;
    defparam mux_196_Mux_0_i699_3_lut_3_lut_4_lut.init = 16'h1c33;
    LUT4 mux_196_Mux_7_i541_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n541_adj_2660)) /* synthesis lut_function=(A (B (C)+!B ((D)+!C))+!A (B (C)+!B !(C))) */ ;
    defparam mux_196_Mux_7_i541_3_lut_4_lut_4_lut.init = 16'he3c3;
    LUT4 mux_196_Mux_7_i60_3_lut_4_lut_3_lut_rep_679 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27002)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_7_i60_3_lut_4_lut_3_lut_rep_679.init = 16'h1818;
    LUT4 i22235_3_lut (.A(n286_adj_2586), .B(n317_adj_2288), .C(index_i[5]), 
         .Z(n23328)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22235_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_0_i747_3_lut_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n747_adj_2580)) /* synthesis lut_function=(!(A (B+!(C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_0_i747_3_lut_3_lut_4_lut_4_lut.init = 16'h6556;
    LUT4 mux_196_Mux_7_i156_3_lut_3_lut_rep_577_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26900)) /* synthesis lut_function=(!(A (B)+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_7_i156_3_lut_3_lut_rep_577_3_lut.init = 16'h6363;
    LUT4 mux_196_Mux_3_i507_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[4]), .D(n491_adj_2382), .Z(n507_adj_2541)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_3_i507_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_196_Mux_6_i573_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[4]), .D(n572_adj_2761), .Z(n573_adj_2632)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_6_i573_3_lut_4_lut.init = 16'hf909;
    LUT4 mux_196_Mux_6_i660_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n108)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_6_i660_3_lut_3_lut.init = 16'hc6c6;
    LUT4 n521_bdd_3_lut_24221_4_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .Z(n24972)) /* synthesis lut_function=(A (B)+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n521_bdd_3_lut_24221_4_lut_3_lut.init = 16'hd9d9;
    LUT4 mux_196_Mux_4_i773_3_lut_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n773)) /* synthesis lut_function=(!(A (B+(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_4_i773_3_lut_3_lut_3_lut.init = 16'h5656;
    LUT4 mux_196_Mux_5_i828_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[4]), .D(n26898), .Z(n828_adj_2459)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D)))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_5_i828_4_lut_4_lut.init = 16'hc66c;
    LUT4 i20269_3_lut (.A(n22722), .B(n22723), .C(index_q[8]), .Z(n22725)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20269_3_lut.init = 16'hcaca;
    LUT4 i9595_3_lut_4_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[4]), .Z(n12160)) /* synthesis lut_function=(!(A (B)+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9595_3_lut_4_lut_4_lut_3_lut.init = 16'h6262;
    PFUMX i20364 (.BLUT(n12104), .ALUT(n62_adj_2753), .C0(index_i[5]), 
          .Z(n22820));
    LUT4 mux_196_Mux_6_i92_3_lut_4_lut_3_lut_rep_699 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27022)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_6_i92_3_lut_4_lut_3_lut_rep_699.init = 16'h6969;
    LUT4 mux_196_Mux_6_i250_3_lut_4_lut_3_lut_rep_700 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27023)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_6_i250_3_lut_4_lut_3_lut_rep_700.init = 16'h9696;
    LUT4 mux_196_Mux_5_i739_rep_701 (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .Z(n27024)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_5_i739_rep_701.init = 16'h6464;
    LUT4 mux_196_Mux_4_i70_3_lut_3_lut_rep_702 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27025)) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_4_i70_3_lut_3_lut_rep_702.init = 16'h6a6a;
    LUT4 mux_196_Mux_6_i627_3_lut_4_lut_3_lut_rep_703 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27026)) /* synthesis lut_function=(A ((C)+!B)+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_6_i627_3_lut_4_lut_3_lut_rep_703.init = 16'he6e6;
    LUT4 mux_196_Mux_6_i518_3_lut_3_lut_rep_704 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27027)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_6_i518_3_lut_3_lut_rep_704.init = 16'h6c6c;
    LUT4 mux_196_Mux_6_i467_3_lut_3_lut_3_lut_rep_705 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27028)) /* synthesis lut_function=(!(A (B)+!A (B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_6_i467_3_lut_3_lut_3_lut_rep_705.init = 16'h3636;
    LUT4 mux_196_Mux_5_i683_3_lut_4_lut_4_lut_3_lut_rep_706 (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[2]), .Z(n27029)) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_5_i683_3_lut_4_lut_4_lut_3_lut_rep_706.init = 16'h6b6b;
    PFUMX i20302 (.BLUT(n31_adj_2482), .ALUT(n62_adj_2762), .C0(index_i[5]), 
          .Z(n22758));
    LUT4 mux_197_Mux_10_i413_3_lut_3_lut_4_lut (.A(n26854), .B(index_q[3]), 
         .C(n26796), .D(index_q[4]), .Z(n413_adj_2763)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_10_i413_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 mux_196_Mux_5_i109_3_lut_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .Z(n109_adj_2729)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_5_i109_3_lut_3_lut_3_lut.init = 16'h3939;
    PFUMX i20142 (.BLUT(n94_adj_2480), .ALUT(n21411), .C0(index_q[5]), 
          .Z(n22598));
    LUT4 mux_196_Mux_6_i60_3_lut_4_lut_3_lut_rep_708 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27031)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_6_i60_3_lut_4_lut_3_lut_rep_708.init = 16'hd6d6;
    LUT4 mux_196_Mux_5_i371_3_lut_4_lut_4_lut_3_lut_rep_709 (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[2]), .Z(n27032)) /* synthesis lut_function=(A ((C)+!B)+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_5_i371_3_lut_4_lut_4_lut_3_lut_rep_709.init = 16'hb6b6;
    LUT4 mux_196_Mux_5_i754_3_lut_4_lut_4_lut_3_lut_rep_710 (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[2]), .Z(n27033)) /* synthesis lut_function=(!(A (B)+!A ((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_5_i754_3_lut_4_lut_4_lut_3_lut_rep_710.init = 16'h2626;
    LUT4 i19596_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n22033)) /* synthesis lut_function=(!(A (B)+!A (B (C+(D))+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19596_3_lut_3_lut_4_lut.init = 16'h3326;
    LUT4 mux_196_Mux_1_i301_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n301_adj_2648)) /* synthesis lut_function=(A (B (C+(D))+!B !(D))+!A !(B (C+(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_1_i301_3_lut_4_lut_4_lut.init = 16'h99b6;
    LUT4 n21326_bdd_3_lut_23728_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n25320)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C))+!A !(B (C+!(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n21326_bdd_3_lut_23728_4_lut_4_lut.init = 16'h5ad6;
    LUT4 i19531_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21968)) /* synthesis lut_function=(A (B (C)+!B !(C (D)+!C !(D)))+!A (B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19531_3_lut_4_lut_4_lut.init = 16'hd6a5;
    LUT4 mux_196_Mux_5_i30_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n30_adj_2472)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A (B+!(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_5_i30_3_lut_4_lut.init = 16'hcc67;
    LUT4 mux_196_Mux_5_i460_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n460_adj_2716)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A !(B (C)+!B !(C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_5_i460_3_lut_4_lut_4_lut.init = 16'h6b5a;
    PFUMX i20271 (.BLUT(n31_adj_2479), .ALUT(n62_adj_2476), .C0(index_i[5]), 
          .Z(n22727));
    LUT4 mux_196_Mux_6_i475_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n475_adj_2704)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A !(B (C+(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_6_i475_3_lut_4_lut_4_lut.init = 16'h9936;
    LUT4 mux_196_Mux_0_i124_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n124_adj_2613)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A !(B (D)+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_0_i124_3_lut_4_lut_4_lut.init = 16'h6c99;
    LUT4 mux_196_Mux_6_i635_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n635_adj_2730)) /* synthesis lut_function=(A (B (C+(D))+!B !(D))+!A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_6_i635_3_lut_4_lut.init = 16'hcce6;
    LUT4 mux_196_Mux_2_i491_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n491_adj_2764)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A !(B (C)+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_2_i491_3_lut_4_lut_4_lut.init = 16'h6a5a;
    PFUMX i23177 (.BLUT(n24907), .ALUT(n24903), .C0(index_i[6]), .Z(n24908));
    LUT4 i19563_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n22000)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19563_3_lut_4_lut.init = 16'h64cc;
    LUT4 i9518_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n12079)) /* synthesis lut_function=(!(A (B (D)+!B (C+!(D)))+!A !(B (D)+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9518_3_lut_4_lut_4_lut.init = 16'h4699;
    PFUMX i20144 (.BLUT(n221_adj_2765), .ALUT(n252_adj_2766), .C0(index_q[5]), 
          .Z(n22600));
    LUT4 n92_bdd_3_lut_23826_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n25610)) /* synthesis lut_function=(A (B (C+(D))+!B ((D)+!C))+!A !(B (C+(D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n92_bdd_3_lut_23826_4_lut.init = 16'haa96;
    LUT4 mux_196_Mux_0_i142_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n142_adj_2721)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C))+!A !(B (C (D)+!C !(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_0_i142_3_lut_4_lut_4_lut.init = 16'ha569;
    PFUMX i20225 (.BLUT(n31_adj_2473), .ALUT(n21954), .C0(index_i[5]), 
          .Z(n22681));
    LUT4 i9369_2_lut_rep_711 (.A(index_q[2]), .B(index_q[3]), .Z(n27034)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9369_2_lut_rep_711.init = 16'h8888;
    PFUMX i20145 (.BLUT(n286_adj_2469), .ALUT(n21414), .C0(index_q[5]), 
          .Z(n22601));
    LUT4 i11652_2_lut_rep_473_3_lut (.A(index_q[2]), .B(index_q[3]), .C(index_q[1]), 
         .Z(n26796)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11652_2_lut_rep_473_3_lut.init = 16'h8080;
    LUT4 i20469_3_lut_3_lut_3_lut_4_lut (.A(index_q[2]), .B(index_q[3]), 
         .C(index_q[4]), .D(index_q[1]), .Z(n22925)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20469_3_lut_3_lut_3_lut_4_lut.init = 16'h878f;
    LUT4 i11567_2_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n668_adj_2556)) /* synthesis lut_function=(!(A ((D)+!B)+!A (B ((D)+!C)+!B (C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11567_2_lut_4_lut_4_lut_4_lut.init = 16'h00c9;
    LUT4 i20466_3_lut_3_lut_4_lut (.A(n26854), .B(index_q[3]), .C(n923_adj_2528), 
         .D(index_q[4]), .Z(n22922)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20466_3_lut_3_lut_4_lut.init = 16'hf011;
    PFUMX i20172 (.BLUT(n31_adj_2468), .ALUT(n62_adj_2739), .C0(index_q[5]), 
          .Z(n22628));
    LUT4 i18963_3_lut (.A(n27099), .B(n29473), .C(index_q[3]), .Z(n21400)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18963_3_lut.init = 16'hcaca;
    LUT4 i19964_1_lut_2_lut (.A(index_q[2]), .B(index_q[3]), .Z(n22420)) /* synthesis lut_function=(!(A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19964_1_lut_2_lut.init = 16'h7777;
    PFUMX i20146 (.BLUT(n349_adj_2767), .ALUT(n21417), .C0(index_q[5]), 
          .Z(n22602));
    LUT4 i11597_2_lut_rep_445_3_lut_4_lut (.A(index_q[2]), .B(index_q[3]), 
         .C(index_q[4]), .D(n27101), .Z(n26768)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11597_2_lut_rep_445_3_lut_4_lut.init = 16'hf8f0;
    LUT4 mux_196_Mux_6_i498_3_lut_4_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n404)) /* synthesis lut_function=(A (B+!(C))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_6_i498_3_lut_4_lut_4_lut_3_lut.init = 16'h9b9b;
    LUT4 mux_197_Mux_7_i924_3_lut_3_lut_4_lut (.A(index_q[2]), .B(index_q[3]), 
         .C(index_q[4]), .D(n27101), .Z(n924_adj_2768)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_7_i924_3_lut_3_lut_4_lut.init = 16'h878f;
    LUT4 i11477_2_lut_rep_446_3_lut_4_lut (.A(index_q[2]), .B(index_q[3]), 
         .C(index_q[4]), .D(n27085), .Z(n26769)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11477_2_lut_rep_446_3_lut_4_lut.init = 16'hf8f0;
    LUT4 i11497_2_lut_rep_712 (.A(index_i[2]), .B(index_i[3]), .Z(n27035)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11497_2_lut_rep_712.init = 16'h8888;
    LUT4 i11766_2_lut_2_lut_3_lut (.A(index_i[2]), .B(index_i[3]), .C(index_i[0]), 
         .Z(n14441)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11766_2_lut_2_lut_3_lut.init = 16'h0808;
    LUT4 i15565_3_lut_3_lut_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n17829)) /* synthesis lut_function=(!(A (B (C)+!B !(C (D)+!C !(D)))+!A !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i15565_3_lut_3_lut_3_lut_4_lut.init = 16'h780f;
    LUT4 i11735_2_lut_rep_519_3_lut (.A(index_i[2]), .B(index_i[3]), .C(index_i[1]), 
         .Z(n26842)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11735_2_lut_rep_519_3_lut.init = 16'h8080;
    LUT4 i20448_3_lut_3_lut_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[4]), .D(index_i[1]), .Z(n22904)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20448_3_lut_3_lut_3_lut_4_lut.init = 16'h878f;
    LUT4 i8005_3_lut_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), .C(index_i[1]), 
         .D(index_i[0]), .Z(n157_adj_2396)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(D))+!A !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i8005_3_lut_3_lut_4_lut.init = 16'h7780;
    PFUMX i20151 (.BLUT(n669_adj_2465), .ALUT(n700_adj_2463), .C0(index_q[5]), 
          .Z(n22607));
    LUT4 i20546_3_lut (.A(n27002), .B(n26900), .C(index_i[3]), .Z(n23002)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20546_3_lut.init = 16'hcaca;
    PFUMX i20152 (.BLUT(n21429), .ALUT(n763_adj_2701), .C0(index_q[5]), 
          .Z(n22608));
    LUT4 i15564_3_lut_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), .C(index_i[1]), 
         .D(index_i[0]), .Z(n17828)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i15564_3_lut_3_lut_4_lut.init = 16'hf078;
    LUT4 i11693_2_lut_rep_526_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n26849)) /* synthesis lut_function=(A (B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11693_2_lut_rep_526_3_lut_4_lut.init = 16'h8880;
    LUT4 i9539_3_lut_4_lut_4_lut_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n875_adj_2263)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(D))+!A !(D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9539_3_lut_4_lut_4_lut_3_lut_4_lut.init = 16'h887f;
    LUT4 i9498_3_lut_3_lut_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n541_adj_2684)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9498_3_lut_3_lut_3_lut_4_lut.init = 16'h870f;
    LUT4 mux_197_Mux_5_i700_3_lut (.A(n460_adj_2509), .B(n27083), .C(index_q[4]), 
         .Z(n700_adj_2757)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_5_i700_3_lut.init = 16'hcaca;
    LUT4 i22248_3_lut (.A(n924_adj_2769), .B(n955), .C(index_i[5]), .Z(n23296)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22248_3_lut.init = 16'hcaca;
    LUT4 i11667_2_lut_rep_512_3_lut (.A(index_i[2]), .B(index_i[3]), .C(index_i[1]), 
         .Z(n26835)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11667_2_lut_rep_512_3_lut.init = 16'hfefe;
    L6MUX21 i21026 (.D0(n23466), .D1(n23467), .SD(index_i[5]), .Z(n23482));
    L6MUX21 i21027 (.D0(n23468), .D1(n23469), .SD(index_i[5]), .Z(n23483));
    LUT4 i9532_3_lut_3_lut_4_lut_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n762_adj_2270)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C (D)+!C !(D)))+!A !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9532_3_lut_3_lut_4_lut_3_lut_4_lut.init = 16'h700f;
    LUT4 mux_196_Mux_8_i14_3_lut_rep_680 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n27003)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_8_i14_3_lut_rep_680.init = 16'h8383;
    LUT4 i19950_1_lut_2_lut (.A(index_i[2]), .B(index_i[3]), .Z(n22406)) /* synthesis lut_function=(!(A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19950_1_lut_2_lut.init = 16'h7777;
    LUT4 i1_2_lut_rep_541_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), .C(index_i[1]), 
         .D(index_i[0]), .Z(n26864)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i1_2_lut_rep_541_3_lut_4_lut.init = 16'h8000;
    LUT4 mux_196_Mux_7_i77_3_lut_3_lut_rep_609 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26932)) /* synthesis lut_function=(A (B)+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_7_i77_3_lut_3_lut_rep_609.init = 16'h9c9c;
    LUT4 mux_196_Mux_5_i38_3_lut_3_lut_4_lut_3_lut_rep_610 (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[2]), .Z(n26933)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_5_i38_3_lut_3_lut_4_lut_3_lut_rep_610.init = 16'h1919;
    LUT4 mux_196_Mux_6_i505_3_lut_rep_611 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26934)) /* synthesis lut_function=(A (B)+!A (B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_6_i505_3_lut_rep_611.init = 16'hc9c9;
    LUT4 i11260_2_lut_rep_493_3_lut (.A(index_q[1]), .B(index_q[2]), .C(index_q[3]), 
         .Z(n26816)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11260_2_lut_rep_493_3_lut.init = 16'hf8f8;
    LUT4 i19659_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n22096)) /* synthesis lut_function=(A (B (C)+!B (C (D)+!C !(D)))+!A !(B (C+!(D))+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19659_3_lut_4_lut_4_lut.init = 16'ha593;
    L6MUX21 i24182 (.D0(n26015), .D1(n26012), .SD(index_q[5]), .Z(n26016));
    LUT4 mux_196_Mux_3_i397_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n397_adj_2711)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !(B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_3_i397_3_lut_4_lut_4_lut.init = 16'ha95a;
    PFUMX i20141 (.BLUT(n31), .ALUT(n62_adj_2455), .C0(index_q[5]), .Z(n22597));
    L6MUX21 i25790 (.D0(n28558), .D1(n28555), .SD(index_i[7]), .Z(n28559));
    PFUMX i25788 (.BLUT(n28557), .ALUT(n28556), .C0(index_i[5]), .Z(n28558));
    LUT4 i19669_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n22106)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C+(D)))+!A (B (C)+!B !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19669_3_lut_4_lut_4_lut.init = 16'hc95a;
    PFUMX i24180 (.BLUT(n26014), .ALUT(n26013), .C0(index_q[4]), .Z(n26015));
    LUT4 i19515_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n21952)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(D))+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19515_3_lut_3_lut_4_lut.init = 16'h3319;
    LUT4 mux_196_Mux_3_i859_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n859_adj_2647)) /* synthesis lut_function=(!(A (B (D)+!B !(D))+!A (B (C+(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_3_i859_3_lut_3_lut_4_lut.init = 16'h339c;
    L6MUX21 i21028 (.D0(n23470), .D1(n23471), .SD(index_i[5]), .Z(n23484));
    PFUMX i20153 (.BLUT(n21432), .ALUT(n828_adj_2457), .C0(index_q[5]), 
          .Z(n22609));
    LUT4 i19605_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n22042)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C))+!A !(B ((D)+!C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19605_3_lut_4_lut_4_lut.init = 16'h925a;
    PFUMX i25786 (.BLUT(n23337), .ALUT(n28554), .C0(index_i[6]), .Z(n28555));
    LUT4 i12180_2_lut_rep_614 (.A(index_i[2]), .B(index_i[0]), .Z(n26937)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i12180_2_lut_rep_614.init = 16'heeee;
    LUT4 n45_bdd_2_lut_3_lut_3_lut_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[1]), .D(index_i[3]), .Z(n25706)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B ((D)+!C)))) */ ;
    defparam n45_bdd_2_lut_3_lut_3_lut_4_lut.init = 16'h00fe;
    LUT4 mux_197_Mux_5_i781_3_lut_4_lut_4_lut_then_4_lut (.A(index_q[3]), 
         .B(index_q[0]), .C(index_q[4]), .D(index_q[2]), .Z(n27130)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_5_i781_3_lut_4_lut_4_lut_then_4_lut.init = 16'hece0;
    LUT4 i1_2_lut_rep_552_3_lut (.A(index_i[2]), .B(index_i[0]), .C(index_i[1]), 
         .Z(n26875)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_552_3_lut.init = 16'hfefe;
    LUT4 mux_196_Mux_5_i954_3_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[1]), .Z(n954_adj_2706)) /* synthesis lut_function=(!(A (C)+!A (B+((D)+!C)))) */ ;
    defparam mux_196_Mux_5_i954_3_lut_4_lut_4_lut.init = 16'h0a1a;
    PFUMX i24177 (.BLUT(n26011), .ALUT(n26746), .C0(index_q[4]), .Z(n26012));
    L6MUX21 i25770 (.D0(n28536), .D1(n28533), .SD(index_q[7]), .Z(n28537));
    PFUMX i20154 (.BLUT(n860_adj_2446), .ALUT(n21435), .C0(index_q[5]), 
          .Z(n22610));
    PFUMX i25768 (.BLUT(n28535), .ALUT(n28534), .C0(index_q[5]), .Z(n28536));
    LUT4 mux_196_Mux_9_i285_3_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[1]), .Z(n285_adj_2386)) /* synthesis lut_function=(A (C)+!A !(B+(C+(D)))) */ ;
    defparam mux_196_Mux_9_i285_3_lut_4_lut_4_lut.init = 16'ha0a1;
    LUT4 i11354_2_lut_rep_452_3_lut_4_lut (.A(index_i[2]), .B(index_i[0]), 
         .C(index_i[3]), .D(index_i[1]), .Z(n26775)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;
    defparam i11354_2_lut_rep_452_3_lut_4_lut.init = 16'hf0e0;
    LUT4 mux_196_Mux_3_i700_3_lut_4_lut (.A(index_i[4]), .B(index_i[3]), 
         .C(n684_adj_2770), .D(n26992), .Z(n700_adj_2545)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_3_i700_3_lut_4_lut.init = 16'hf4b0;
    LUT4 mux_197_Mux_5_i781_3_lut_4_lut_4_lut_else_4_lut (.A(index_q[3]), 
         .B(index_q[0]), .C(index_q[4]), .Z(n27129)) /* synthesis lut_function=(!(A (C)+!A (B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_5_i781_3_lut_4_lut_4_lut_else_4_lut.init = 16'h1f1f;
    LUT4 i22456_3_lut (.A(n24975), .B(n23285), .C(index_i[6]), .Z(n23299)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22456_3_lut.init = 16'hcaca;
    PFUMX i25766 (.BLUT(n23184), .ALUT(n28532), .C0(index_q[6]), .Z(n28533));
    LUT4 mux_196_Mux_0_i635_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n635_adj_2536)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_0_i635_3_lut_4_lut_4_lut.init = 16'hfd0a;
    LUT4 mux_197_Mux_8_i860_3_lut_4_lut (.A(n26893), .B(index_q[3]), .C(index_q[4]), 
         .D(n26856), .Z(n860_adj_2662)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_8_i860_3_lut_4_lut.init = 16'h08f8;
    PFUMX i24753 (.BLUT(n27159), .ALUT(n27160), .C0(index_q[1]), .Z(n27161));
    LUT4 i19497_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n21934)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (D))+!A !(D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19497_3_lut_4_lut_4_lut_4_lut.init = 16'ha25d;
    L6MUX21 i21029 (.D0(n23472), .D1(n23473), .SD(index_i[5]), .Z(n23485));
    LUT4 mux_197_Mux_3_i157_3_lut_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n157_adj_2437)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_3_i157_3_lut_3_lut_3_lut_4_lut.init = 16'h1ff0;
    LUT4 index_q_5__bdd_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n25801)) /* synthesis lut_function=(A (B (C)+!B (C+(D)))+!A (B (C)+!B !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam index_q_5__bdd_3_lut_4_lut_4_lut_4_lut.init = 16'he3f0;
    LUT4 i12163_1_lut_2_lut_3_lut_4_lut (.A(n26854), .B(index_q[3]), .C(index_q[5]), 
         .D(index_q[4]), .Z(n381_adj_2415)) /* synthesis lut_function=(!(A (C+(D))+!A (B (C+(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12163_1_lut_2_lut_3_lut_4_lut.init = 16'h010f;
    L6MUX21 i21030 (.D0(n23474), .D1(n23475), .SD(index_i[5]), .Z(n23486));
    LUT4 i15522_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .D(index_q[0]), .Z(n17786)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C (D)+!C !(D)))+!A !(B (D)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i15522_3_lut_4_lut_4_lut_4_lut.init = 16'h83fc;
    LUT4 i22258_3_lut (.A(n25830), .B(n21749), .C(index_q[5]), .Z(n21750)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22258_3_lut.init = 16'hcaca;
    L6MUX21 i21031 (.D0(n23476), .D1(n23477), .SD(index_i[5]), .Z(n23487));
    L6MUX21 i21032 (.D0(n23478), .D1(n23479), .SD(index_i[5]), .Z(n23488));
    PFUMX i20173 (.BLUT(n94_adj_2740), .ALUT(n125_adj_2440), .C0(index_q[5]), 
          .Z(n22629));
    PFUMX i20174 (.BLUT(n158_adj_2438), .ALUT(n189), .C0(index_q[5]), 
          .Z(n22630));
    LUT4 mux_196_Mux_1_i908_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n908_adj_2282)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+(D)))+!A (B (C+(D))+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_1_i908_3_lut_4_lut_4_lut_4_lut.init = 16'h332d;
    L6MUX21 i21033 (.D0(n23480), .D1(n23481), .SD(index_i[5]), .Z(n23489));
    PFUMX i20175 (.BLUT(n221_adj_2295), .ALUT(n252), .C0(index_q[5]), 
          .Z(n22631));
    LUT4 mux_197_Mux_4_i93_3_lut_4_lut_3_lut_rep_734_4_lut (.A(index_q[1]), 
         .B(index_q[2]), .C(index_q[3]), .D(index_q[0]), .Z(n27057)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_4_i93_3_lut_4_lut_3_lut_rep_734_4_lut.init = 16'h07f0;
    L6MUX21 i24152 (.D0(n25969), .D1(n25967), .SD(index_q[4]), .Z(n25970));
    LUT4 mux_197_Mux_10_i252_3_lut_4_lut_4_lut (.A(n26854), .B(index_q[3]), 
         .C(index_q[4]), .D(n26861), .Z(n252_adj_2442)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B (C (D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_10_i252_3_lut_4_lut_4_lut.init = 16'h3efe;
    LUT4 i11546_2_lut_rep_528_2_lut (.A(index_i[1]), .B(index_i[0]), .Z(n26851)) /* synthesis lut_function=((B)+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11546_2_lut_rep_528_2_lut.init = 16'hdddd;
    PFUMX i24150 (.BLUT(n26753), .ALUT(n25968), .C0(index_q[5]), .Z(n25969));
    LUT4 mux_196_Mux_4_i340_3_lut_rep_660 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26983)) /* synthesis lut_function=(A (B+!(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_4_i340_3_lut_rep_660.init = 16'hdada;
    LUT4 i9416_2_lut_3_lut (.A(index_q[1]), .B(index_q[2]), .C(index_q[3]), 
         .Z(n11977)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9416_2_lut_3_lut.init = 16'h8080;
    PFUMX i20176 (.BLUT(n286), .ALUT(n21444), .C0(index_q[5]), .Z(n22632));
    PFUMX i24148 (.BLUT(n25966), .ALUT(n25965), .C0(index_q[5]), .Z(n25967));
    LUT4 i18957_3_lut (.A(n356), .B(n29473), .C(index_q[3]), .Z(n21394)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18957_3_lut.init = 16'hcaca;
    LUT4 i18955_3_lut (.A(n27098), .B(n29474), .C(index_q[3]), .Z(n21392)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18955_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_87 (.A(index_q[6]), .B(n26856), .C(index_q[5]), 
         .D(index_q[4]), .Z(n20366)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_4_lut_adj_87.init = 16'hfffe;
    LUT4 i18954_3_lut (.A(n27077), .B(n29494), .C(index_q[3]), .Z(n21391)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i18954_3_lut.init = 16'hcaca;
    LUT4 i17611_4_lut (.A(n27044), .B(n892_adj_2441), .C(index_q[6]), 
         .D(index_q[5]), .Z(n19907)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D))))) */ ;
    defparam i17611_4_lut.init = 16'h3a35;
    LUT4 i22461_3_lut (.A(n19907), .B(n20366), .C(index_q[7]), .Z(n22854)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22461_3_lut.init = 16'hcaca;
    PFUMX i19129 (.BLUT(n445), .ALUT(n508_adj_2542), .C0(index_i[6]), 
          .Z(n21566));
    LUT4 mux_196_Mux_5_i761_3_lut_4_lut_3_lut_rep_663 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26986)) /* synthesis lut_function=(A (B)+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_5_i761_3_lut_4_lut_3_lut_rep_663.init = 16'hd9d9;
    PFUMX i20177 (.BLUT(n349_adj_2771), .ALUT(n21447), .C0(index_q[5]), 
          .Z(n22633));
    PFUMX i20178 (.BLUT(n413_adj_2433), .ALUT(n444_adj_2772), .C0(index_q[5]), 
          .Z(n22634));
    PFUMX i20179 (.BLUT(n476_adj_2431), .ALUT(n507_adj_2748), .C0(index_q[5]), 
          .Z(n22635));
    PFUMX i20180 (.BLUT(n21450), .ALUT(n573_adj_2398), .C0(index_q[5]), 
          .Z(n22636));
    LUT4 mux_196_Mux_6_i572_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n572_adj_2761)) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_6_i572_3_lut_4_lut.init = 16'hccd9;
    LUT4 n53_bdd_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n25317)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n53_bdd_3_lut_4_lut_4_lut.init = 16'ha5ad;
    LUT4 i19632_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n22069)) /* synthesis lut_function=(!(A (B (C (D))+!B (C (D)+!C !(D)))+!A !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19632_3_lut_4_lut_4_lut.init = 16'h5aad;
    PFUMX i20181 (.BLUT(n11973), .ALUT(n21453), .C0(index_q[5]), .Z(n22637));
    LUT4 mux_196_Mux_4_i723_3_lut_4_lut_3_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .Z(n723)) /* synthesis lut_function=(A (B (C))+!A (B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_4_i723_3_lut_4_lut_3_lut_3_lut.init = 16'hd4d4;
    LUT4 i19615_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n22052)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D))+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19615_3_lut_4_lut.init = 16'hccdb;
    LUT4 mux_197_Mux_3_i30_3_lut_3_lut_4_lut_3_lut_4_lut (.A(index_q[0]), 
         .B(index_q[1]), .C(index_q[3]), .D(index_q[2]), .Z(n30_adj_2467)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_3_i30_3_lut_3_lut_4_lut_3_lut_4_lut.init = 16'hfe11;
    PFUMX i20182 (.BLUT(n669), .ALUT(n700_adj_2621), .C0(index_q[5]), 
          .Z(n22638));
    LUT4 mux_196_Mux_1_i732_3_lut (.A(n716_adj_2330), .B(n491_adj_2727), 
         .C(index_i[4]), .Z(n732_adj_2299)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_1_i732_3_lut.init = 16'hcaca;
    L6MUX21 i20183 (.D0(n21456), .D1(n763_adj_2680), .SD(index_q[5]), 
            .Z(n22639));
    PFUMX i23146 (.BLUT(n24868), .ALUT(n24865), .C0(index_i[6]), .Z(n24869));
    PFUMX i20185 (.BLUT(n860_adj_2666), .ALUT(n891_adj_2426), .C0(index_q[5]), 
          .Z(n22641));
    LUT4 i7650_2_lut_rep_721 (.A(index_q[3]), .B(index_q[4]), .Z(n27044)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i7650_2_lut_rep_721.init = 16'h8888;
    LUT4 i1_2_lut_rep_547_3_lut (.A(index_q[3]), .B(index_q[4]), .C(index_q[5]), 
         .Z(n26870)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_2_lut_rep_547_3_lut.init = 16'hf8f8;
    LUT4 i1_2_lut_3_lut (.A(index_q[3]), .B(index_q[4]), .C(index_q[5]), 
         .Z(n20559)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_2_lut_3_lut.init = 16'h8080;
    LUT4 i22399_3_lut (.A(n22803), .B(n25588), .C(index_i[6]), .Z(n22812)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22399_3_lut.init = 16'hcaca;
    LUT4 i20721_3_lut_3_lut_4_lut (.A(index_q[3]), .B(index_q[4]), .C(n413_adj_2763), 
         .D(index_q[5]), .Z(n23177)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20721_3_lut_3_lut_4_lut.init = 16'h77f0;
    LUT4 i11689_2_lut_3_lut_4_lut (.A(index_q[3]), .B(index_q[4]), .C(index_q[2]), 
         .D(n27085), .Z(n125_adj_2532)) /* synthesis lut_function=(A (B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11689_2_lut_3_lut_4_lut.init = 16'h8880;
    PFUMX i20186 (.BLUT(n924_adj_2421), .ALUT(n21459), .C0(index_q[5]), 
          .Z(n22642));
    LUT4 mux_197_Mux_4_i491_3_lut_4_lut_4_lut (.A(index_q[2]), .B(n27102), 
         .C(index_q[3]), .D(n27085), .Z(n491_adj_2664)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_4_i491_3_lut_4_lut_4_lut.init = 16'hfc5c;
    LUT4 i12072_3_lut_3_lut (.A(index_q[2]), .B(index_q[0]), .C(index_q[1]), 
         .Z(n1001)) /* synthesis lut_function=(A (C)+!A (B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12072_3_lut_3_lut.init = 16'hf4f4;
    LUT4 mux_196_Mux_5_i731_3_lut (.A(n29471), .B(n27032), .C(index_i[3]), 
         .Z(n731_adj_2283)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_5_i731_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_0_i364_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n364_adj_2773)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A ((C+!(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_0_i364_3_lut_3_lut_4_lut.init = 16'hdb55;
    LUT4 n26262_bdd_3_lut_3_lut (.A(n1021_adj_2725), .B(index_q[8]), .C(n26262), 
         .Z(n26263)) /* synthesis lut_function=(A (B+(C))+!A !(B+!(C))) */ ;
    defparam n26262_bdd_3_lut_3_lut.init = 16'hb8b8;
    LUT4 mux_197_Mux_5_i924_4_lut_3_lut (.A(index_q[2]), .B(n13925), .C(index_q[4]), 
         .Z(n924_adj_2774)) /* synthesis lut_function=(!(A (B+(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_5_i924_4_lut_3_lut.init = 16'h5656;
    LUT4 mux_197_Mux_0_i620_3_lut (.A(n27102), .B(n27082), .C(index_q[3]), 
         .Z(n620_adj_2251)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i620_3_lut.init = 16'hcaca;
    LUT4 i11418_2_lut_rep_722 (.A(index_i[3]), .B(index_i[4]), .Z(n27045)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11418_2_lut_rep_722.init = 16'h8888;
    PFUMX i20187 (.BLUT(n21462), .ALUT(n1018_adj_2670), .C0(index_q[5]), 
          .Z(n22643));
    LUT4 mux_197_Mux_8_i412_3_lut_4_lut_3_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .Z(n14928)) /* synthesis lut_function=(A (B+!(C))+!A !((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_8_i412_3_lut_4_lut_3_lut.init = 16'h8e8e;
    LUT4 n18009_bdd_4_lut_then_4_lut (.A(index_i[3]), .B(index_i[4]), .C(index_i[1]), 
         .D(index_i[2]), .Z(n27207)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B+(C (D)+!C !(D)))) */ ;
    defparam n18009_bdd_4_lut_then_4_lut.init = 16'hf44f;
    LUT4 i9528_3_lut_3_lut_3_lut_4_lut (.A(index_i[3]), .B(index_i[4]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n444_adj_2427)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C))+!A (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9528_3_lut_3_lut_3_lut_4_lut.init = 16'h0f87;
    LUT4 i1_2_lut_rep_551_3_lut (.A(index_i[3]), .B(index_i[4]), .C(index_i[5]), 
         .Z(n26874)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i1_2_lut_rep_551_3_lut.init = 16'hf8f8;
    LUT4 i20720_3_lut_4_lut_4_lut (.A(n26856), .B(index_q[4]), .C(index_q[5]), 
         .D(n26767), .Z(n23176)) /* synthesis lut_function=(A ((C+!(D))+!B)+!A (B (C+!(D))+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20720_3_lut_4_lut_4_lut.init = 16'he3ef;
    LUT4 i19569_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n22006)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19569_3_lut_4_lut_4_lut.init = 16'hda5a;
    LUT4 i11782_2_lut_rep_569_3_lut (.A(index_q[1]), .B(index_q[2]), .C(index_q[0]), 
         .Z(n26892)) /* synthesis lut_function=(A (B+!(C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11782_2_lut_rep_569_3_lut.init = 16'h8f8f;
    LUT4 i19654_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n22091)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C))+!A !(B (C)+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19654_3_lut_4_lut_4_lut.init = 16'h5ad3;
    LUT4 i20874_3_lut_3_lut_4_lut (.A(index_i[3]), .B(index_i[4]), .C(n413), 
         .D(index_i[5]), .Z(n23330)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20874_3_lut_3_lut_4_lut.init = 16'h77f0;
    LUT4 i1_2_lut_3_lut_adj_88 (.A(index_i[3]), .B(index_i[4]), .C(index_i[5]), 
         .Z(n20555)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i1_2_lut_3_lut_adj_88.init = 16'h8080;
    LUT4 i22293_3_lut (.A(n28270), .B(n27232), .C(index_i[5]), .Z(n22741)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22293_3_lut.init = 16'hcaca;
    LUT4 i8234_2_lut_rep_723 (.A(index_i[1]), .B(index_i[2]), .Z(n27046)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i8234_2_lut_rep_723.init = 16'h8888;
    LUT4 mux_196_Mux_9_i30_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .D(index_i[3]), .Z(n30_adj_2713)) /* synthesis lut_function=(A (B (C (D))+!B !(D))+!A !(B+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_9_i30_3_lut_4_lut_4_lut_4_lut.init = 16'h8033;
    LUT4 i20797_3_lut_3_lut_4_lut (.A(n26861), .B(index_q[3]), .C(n93_adj_2775), 
         .D(index_q[4]), .Z(n23253)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C+!(D))) */ ;
    defparam i20797_3_lut_3_lut_4_lut.init = 16'hf077;
    LUT4 n18009_bdd_4_lut_else_4_lut (.A(index_i[3]), .B(index_i[4]), .C(index_i[1]), 
         .D(index_i[2]), .Z(n27206)) /* synthesis lut_function=(!(A (B (D)+!B ((D)+!C))+!A !(B+!((D)+!C)))) */ ;
    defparam n18009_bdd_4_lut_else_4_lut.init = 16'h44fc;
    LUT4 mux_196_Mux_3_i349_3_lut_3_lut (.A(index_i[1]), .B(index_i[4]), 
         .C(n348_adj_2685), .Z(n349_adj_2534)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_3_i349_3_lut_3_lut.init = 16'hd1d1;
    LUT4 mux_196_Mux_4_i93_3_lut_4_lut_3_lut_rep_656_4_lut (.A(index_i[1]), 
         .B(index_i[2]), .C(index_i[3]), .D(index_i[0]), .Z(n26979)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_4_i93_3_lut_4_lut_3_lut_rep_656_4_lut.init = 16'h07f0;
    LUT4 i9534_2_lut_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[3]), 
         .Z(n12095)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9534_2_lut_3_lut.init = 16'h8080;
    LUT4 i11659_2_lut_rep_553_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[0]), 
         .Z(n26876)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11659_2_lut_rep_553_3_lut.init = 16'h8080;
    LUT4 i23261_then_4_lut (.A(index_i[6]), .B(index_i[2]), .C(index_i[5]), 
         .D(index_i[0]), .Z(n27210)) /* synthesis lut_function=(A ((C+!(D))+!B)+!A !(B (C (D))+!B !(C+(D)))) */ ;
    defparam i23261_then_4_lut.init = 16'hb7fe;
    LUT4 i22297_3_lut (.A(n542_adj_2718), .B(n573_adj_2387), .C(index_i[5]), 
         .Z(n22735)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22297_3_lut.init = 16'hcaca;
    LUT4 i19609_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .D(index_i[3]), .Z(n22046)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(D))+!A (B+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19609_3_lut_4_lut_4_lut_4_lut.init = 16'h3380;
    PFUMX i19138 (.BLUT(n445_adj_2334), .ALUT(n508), .C0(index_q[6]), 
          .Z(n21575));
    L6MUX21 i25559 (.D0(n28253), .D1(n28250), .SD(index_i[5]), .Z(n28254));
    LUT4 i19537_3_lut_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n21974)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C (D)+!C !(D)))+!A !(B (D)+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19537_3_lut_4_lut_4_lut_4_lut.init = 16'h7c03;
    PFUMX i25557 (.BLUT(n28252), .ALUT(n28251), .C0(index_i[3]), .Z(n28253));
    PFUMX i25555 (.BLUT(n28249), .ALUT(n28248), .C0(index_i[3]), .Z(n28250));
    LUT4 i11763_2_lut_rep_471_2_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .Z(n26794)) /* synthesis lut_function=(A (B+!(C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11763_2_lut_rep_471_2_lut_3_lut.init = 16'h8f8f;
    LUT4 i19567_3_lut_4_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n22004)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19567_3_lut_4_lut_3_lut_4_lut.init = 16'hf80f;
    LUT4 i11429_2_lut_rep_490_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[3]), 
         .Z(n26813)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11429_2_lut_rep_490_3_lut.init = 16'hf8f8;
    PFUMX i20255 (.BLUT(n22709), .ALUT(n22710), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2126[5]));
    PFUMX i20743 (.BLUT(n333_adj_2759), .ALUT(n348_adj_2776), .C0(index_i[4]), 
          .Z(n23199));
    LUT4 i23261_else_4_lut (.A(index_i[2]), .Z(n27209)) /* synthesis lut_function=(A) */ ;
    defparam i23261_else_4_lut.init = 16'haaaa;
    PFUMX i20744 (.BLUT(n364_adj_2773), .ALUT(n379), .C0(index_i[4]), 
          .Z(n23200));
    LUT4 i11584_2_lut_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), .C(index_i[1]), 
         .D(index_i[0]), .Z(n844_adj_2262)) /* synthesis lut_function=(A ((C (D)+!C !(D))+!B)+!A (B+(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11584_2_lut_3_lut_4_lut.init = 16'hf66f;
    LUT4 i19044_3_lut (.A(n498), .B(n27095), .C(index_q[3]), .Z(n21481)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19044_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_3_i142_3_lut_3_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .Z(n142_adj_2705)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_3_i142_3_lut_3_lut_3_lut.init = 16'h3838;
    LUT4 i21789_3_lut (.A(n21481), .B(n21482), .C(index_q[4]), .Z(n21483)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21789_3_lut.init = 16'hcaca;
    PFUMX i20745 (.BLUT(n397_adj_2410), .ALUT(n412_adj_2335), .C0(index_i[4]), 
          .Z(n23201));
    PFUMX i20332 (.BLUT(n22786), .ALUT(n22787), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2126[3]));
    PFUMX i19706 (.BLUT(n22141), .ALUT(n22142), .C0(index_q[4]), .Z(n22143));
    LUT4 mux_196_Mux_6_i924_3_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[4]), .D(n762_adj_2298), .Z(n924_adj_2769)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_6_i924_3_lut_4_lut.init = 16'h6f60;
    LUT4 i11391_2_lut_rep_453_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n26776)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11391_2_lut_rep_453_3_lut_4_lut.init = 16'hf8f0;
    LUT4 mux_196_Mux_8_i491_3_lut_3_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n491_adj_2676)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_8_i491_3_lut_3_lut_3_lut_4_lut.init = 16'h7870;
    LUT4 i11658_2_lut_rep_724 (.A(index_i[1]), .B(index_i[2]), .C(index_i[0]), 
         .Z(n27047)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11658_2_lut_rep_724.init = 16'h7070;
    LUT4 mux_196_Mux_0_i1017_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[0]), .D(index_i[3]), .Z(n1017_adj_2697)) /* synthesis lut_function=(A (B (D)+!B !((D)+!C))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_0_i1017_4_lut_4_lut_4_lut.init = 16'hdd70;
    LUT4 i11560_2_lut_rep_725 (.A(index_i[1]), .B(index_i[2]), .Z(n27048)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11560_2_lut_rep_725.init = 16'heeee;
    LUT4 i19536_3_lut_4_lut_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .D(index_i[0]), .Z(n21973)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19536_3_lut_4_lut_3_lut_4_lut.init = 16'h0fe0;
    LUT4 i11287_2_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n635_adj_2549)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A (B (C+!(D))+!B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11287_2_lut_4_lut_4_lut.init = 16'hf1fc;
    LUT4 mux_196_Mux_9_i93_3_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .Z(n93_adj_2290)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_9_i93_3_lut_3_lut.init = 16'hc1c1;
    LUT4 i11661_2_lut_rep_469_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[0]), 
         .Z(n26792)) /* synthesis lut_function=(A (C)+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11661_2_lut_rep_469_3_lut.init = 16'hf1f1;
    LUT4 i9561_3_lut_then_4_lut (.A(index_q[4]), .B(index_q[0]), .C(index_q[1]), 
         .D(index_q[2]), .Z(n27213)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C+(D)))+!A (B (C+(D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9561_3_lut_then_4_lut.init = 16'hd54a;
    LUT4 mux_196_Mux_8_i412_3_lut_4_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .Z(n14858)) /* synthesis lut_function=(A (B+!(C))+!A !((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_8_i412_3_lut_4_lut_3_lut.init = 16'h8e8e;
    PFUMX i20394 (.BLUT(n22848), .ALUT(n22849), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2126[1]));
    LUT4 i11499_2_lut_rep_664 (.A(index_i[0]), .B(index_i[1]), .Z(n26987)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11499_2_lut_rep_664.init = 16'h4444;
    LUT4 i11240_2_lut_rep_451_3_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .D(index_q[0]), .Z(n26774)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11240_2_lut_rep_451_3_lut_4_lut.init = 16'hf8f0;
    PFUMX i20228 (.BLUT(n221_adj_2760), .ALUT(n252_adj_2329), .C0(index_i[5]), 
          .Z(n22684));
    LUT4 i19672_3_lut_3_lut_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[3]), 
         .Z(n22109)) /* synthesis lut_function=(A (C)+!A (B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19672_3_lut_3_lut_3_lut.init = 16'he5e5;
    LUT4 i11259_2_lut_rep_444_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n26767)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11259_2_lut_rep_444_3_lut_4_lut.init = 16'hfef0;
    LUT4 i11414_2_lut_rep_554_3_lut (.A(index_i[1]), .B(index_i[2]), .C(index_i[3]), 
         .Z(n26877)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11414_2_lut_rep_554_3_lut.init = 16'he0e0;
    LUT4 mux_196_Mux_4_i236_3_lut_4_lut_3_lut_rep_653_4_lut (.A(index_i[1]), 
         .B(index_i[2]), .C(index_i[3]), .D(index_i[0]), .Z(n26976)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_4_i236_3_lut_4_lut_3_lut_rep_653_4_lut.init = 16'hf01f;
    LUT4 i9561_3_lut_else_4_lut (.A(index_q[4]), .B(index_q[0]), .C(index_q[1]), 
         .D(index_q[2]), .Z(n27212)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A !(B (D)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9561_3_lut_else_4_lut.init = 16'ha955;
    LUT4 i20762_3_lut (.A(n23215), .B(n23216), .C(index_i[7]), .Z(n23218)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20762_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_0_i954_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n954_adj_2695)) /* synthesis lut_function=(A (D)+!A !(B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_0_i954_3_lut_4_lut_4_lut.init = 16'haf40;
    LUT4 n197_bdd_3_lut_23707_4_lut (.A(n26851), .B(index_i[2]), .C(index_i[3]), 
         .D(n26983), .Z(n24960)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n197_bdd_3_lut_23707_4_lut.init = 16'hf606;
    PFUMX i20746 (.BLUT(n428), .ALUT(n443_adj_2302), .C0(index_i[4]), 
          .Z(n23202));
    LUT4 mux_196_Mux_9_i412_3_lut_3_lut_4_lut_3_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[3]), .Z(n412_adj_2320)) /* synthesis lut_function=(!(A (B (C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_9_i412_3_lut_3_lut_4_lut_3_lut.init = 16'h7e7e;
    LUT4 mux_197_Mux_3_i142_3_lut_3_lut_3_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .Z(n142_adj_2436)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_3_i142_3_lut_3_lut_3_lut.init = 16'h3838;
    LUT4 i11415_2_lut_rep_454_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[4]), .D(index_i[3]), .Z(n26777)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11415_2_lut_rep_454_3_lut_4_lut.init = 16'hfef0;
    LUT4 n10476_bdd_3_lut_23772_4_lut_4_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[4]), .D(index_i[3]), .Z(n24619)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C+(D)))+!A (B (C (D)+!C !(D))+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n10476_bdd_3_lut_23772_4_lut_4_lut_4_lut.init = 16'hc10f;
    LUT4 mux_196_Mux_8_i93_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n93_adj_2652)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C))+!A (B (C+!(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_8_i93_3_lut_3_lut_4_lut.init = 16'h0f83;
    PFUMX i20747 (.BLUT(n460_adj_2321), .ALUT(n475_adj_2381), .C0(index_i[4]), 
          .Z(n23203));
    PFUMX i20656 (.BLUT(n23110), .ALUT(n23111), .C0(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_2141[1]));
    LUT4 i23175_then_3_lut (.A(index_i[0]), .B(index_i[4]), .C(index_i[3]), 
         .Z(n27216)) /* synthesis lut_function=(A (B)+!A (B (C)+!B !(C))) */ ;
    defparam i23175_then_3_lut.init = 16'hc9c9;
    LUT4 i23175_else_3_lut (.A(index_i[0]), .B(index_i[2]), .C(index_i[4]), 
         .D(index_i[3]), .Z(n27215)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C (D)+!C !(D))+!B !(C)))) */ ;
    defparam i23175_else_3_lut.init = 16'h1e58;
    PFUMX i20748 (.BLUT(n491_adj_2777), .ALUT(n11334), .C0(index_i[4]), 
          .Z(n23204));
    LUT4 mux_196_Mux_3_i676_3_lut_4_lut_3_lut_rep_665 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26988)) /* synthesis lut_function=(A (B (C))+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_3_i676_3_lut_4_lut_3_lut_rep_665.init = 16'h9494;
    LUT4 i23144_then_4_lut (.A(index_i[0]), .B(index_i[4]), .C(index_i[1]), 
         .D(index_i[3]), .Z(n27219)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B (C (D)+!C !(D))+!B !(C (D)+!C !(D))))) */ ;
    defparam i23144_then_4_lut.init = 16'h3c69;
    LUT4 i19039_3_lut (.A(n498), .B(n27100), .C(index_q[3]), .Z(n21476)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19039_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_6_i459_rep_666 (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .Z(n26989)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_6_i459_rep_666.init = 16'h4d4d;
    LUT4 i19239_3_lut_4_lut_4_lut (.A(n26876), .B(index_i[4]), .C(index_i[3]), 
         .D(n26882), .Z(n21676)) /* synthesis lut_function=(A (B (C)+!B !(C+!(D)))+!A (B (C)+!B (C+(D)))) */ ;
    defparam i19239_3_lut_4_lut_4_lut.init = 16'hd3d0;
    PFUMX i20125 (.BLUT(n22579), .ALUT(n22580), .C0(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_2141[5]));
    LUT4 mux_196_Mux_6_i371_3_lut_4_lut_4_lut_3_lut_rep_667 (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[2]), .Z(n26990)) /* synthesis lut_function=(!(A (B+!(C))+!A ((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_6_i371_3_lut_4_lut_4_lut_3_lut_rep_667.init = 16'h2424;
    LUT4 mux_197_Mux_5_i851_3_lut_4_lut_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n851)) /* synthesis lut_function=(A ((C)+!B)+!A (B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_5_i851_3_lut_4_lut_3_lut.init = 16'he7e7;
    LUT4 mux_197_Mux_6_i796_3_lut_rep_396_3_lut_3_lut_4_lut (.A(index_q[0]), 
         .B(index_q[1]), .C(index_q[3]), .D(index_q[2]), .Z(n26719)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_6_i796_3_lut_rep_396_3_lut_3_lut_4_lut.init = 16'hfe01;
    PFUMX i19721 (.BLUT(n22156), .ALUT(n22157), .C0(index_q[4]), .Z(n22158));
    LUT4 mux_197_Mux_8_i491_3_lut_3_lut_3_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .D(index_q[0]), .Z(n491_adj_2629)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_8_i491_3_lut_3_lut_3_lut_4_lut.init = 16'h7870;
    PFUMX i19724 (.BLUT(n22159), .ALUT(n22160), .C0(index_q[4]), .Z(n22161));
    LUT4 i19720_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n22157)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B ((D)+!C)+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19720_3_lut_4_lut_4_lut.init = 16'hfc1c;
    PFUMX i19730 (.BLUT(n22165), .ALUT(n22166), .C0(index_q[4]), .Z(n22167));
    PFUMX i20202 (.BLUT(n22656), .ALUT(n22657), .C0(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_2141[3]));
    LUT4 mux_196_Mux_6_i269_rep_668 (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .Z(n26991)) /* synthesis lut_function=(A (C)+!A !((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_6_i269_rep_668.init = 16'ha4a4;
    PFUMX i19733 (.BLUT(n22168), .ALUT(n22169), .C0(index_q[4]), .Z(n22170));
    LUT4 mux_196_Mux_6_i22_rep_669 (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .Z(n26992)) /* synthesis lut_function=(!(A (C)+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_6_i22_rep_669.init = 16'h4a4a;
    LUT4 i23144_else_4_lut (.A(index_i[0]), .B(index_i[4]), .C(index_i[1]), 
         .D(index_i[3]), .Z(n27218)) /* synthesis lut_function=(!(A (B (C)+!B !(C (D)+!C !(D)))+!A (B ((D)+!C)+!B !((D)+!C)))) */ ;
    defparam i23144_else_4_lut.init = 16'h394b;
    LUT4 i18994_3_lut_3_lut_4_lut (.A(index_q[1]), .B(index_q[2]), .C(index_q[3]), 
         .D(index_q[0]), .Z(n21431)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18994_3_lut_3_lut_4_lut.init = 16'hf80f;
    PFUMX i24086 (.BLUT(n25899), .ALUT(n26974), .C0(index_q[4]), .Z(n25900));
    LUT4 mux_196_Mux_6_i378_3_lut_4_lut_3_lut_rep_670 (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n26993)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_6_i378_3_lut_4_lut_3_lut_rep_670.init = 16'h4949;
    LUT4 i19036_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[0]), .D(index_q[3]), .Z(n21473)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(D))+!A (B+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19036_3_lut_4_lut_4_lut_4_lut.init = 16'h3380;
    PFUMX i20270 (.BLUT(n22724), .ALUT(n22725), .C0(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_2141[8]));
    PFUMX i19742 (.BLUT(n22177), .ALUT(n22178), .C0(index_q[4]), .Z(n22179));
    LUT4 mux_197_Mux_1_i923_3_lut_3_lut_4_lut_3_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .Z(n923_adj_2528)) /* synthesis lut_function=(!(A (B (C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_1_i923_3_lut_3_lut_4_lut_3_lut.init = 16'h7e7e;
    LUT4 i11728_2_lut_rep_768 (.A(index_q[1]), .B(index_q[2]), .C(index_q[0]), 
         .Z(n27091)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11728_2_lut_rep_768.init = 16'h7070;
    PFUMX i20363 (.BLUT(n22817), .ALUT(n22818), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2126[2]));
    LUT4 i21797_3_lut (.A(n21472), .B(n21473), .C(index_q[4]), .Z(n21474)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21797_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_0_i1017_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[0]), .D(index_q[3]), .Z(n1017)) /* synthesis lut_function=(A (B (D)+!B !((D)+!C))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i1017_4_lut_4_lut_4_lut.init = 16'hdd70;
    LUT4 i12067_2_lut_rep_769 (.A(index_q[2]), .B(index_q[0]), .Z(n27092)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12067_2_lut_rep_769.init = 16'heeee;
    PFUMX i20273 (.BLUT(n158), .ALUT(n189_adj_2366), .C0(index_i[5]), 
          .Z(n22729));
    LUT4 mux_197_Mux_2_i173_3_lut_4_lut_4_lut_4_lut (.A(index_q[2]), .B(index_q[0]), 
         .C(index_q[3]), .D(index_q[1]), .Z(n173_adj_2352)) /* synthesis lut_function=(!(A (C)+!A (B (C+!(D))+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_2_i173_3_lut_4_lut_4_lut_4_lut.init = 16'h0f1a;
    LUT4 mux_196_Mux_2_i890_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n890_adj_2264)) /* synthesis lut_function=(A (B (D)+!B !((D)+!C))+!A !(B (C+(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_2_i890_3_lut_4_lut_4_lut.init = 16'h9934;
    LUT4 i19635_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n22072)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (D))+!A !(B (C (D))+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19635_3_lut_3_lut_4_lut.init = 16'h4933;
    LUT4 i19704_3_lut_4_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n22141)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))+!A (B (C)+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19704_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'hf1e3;
    PFUMX i9368 (.BLUT(n12148), .ALUT(n12149), .C0(n22420), .Z(n11929));
    LUT4 i19701_3_lut (.A(n900), .B(n27077), .C(index_q[3]), .Z(n22138)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19701_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_5_i491_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n491_adj_2727)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A !(B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_5_i491_3_lut_4_lut_4_lut.init = 16'ha54a;
    LUT4 mux_197_Mux_2_i931_3_lut_3_lut_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n931)) /* synthesis lut_function=(!(A (B (C))+!A (B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_2_i931_3_lut_3_lut_3_lut.init = 16'h3e3e;
    LUT4 i22328_3_lut (.A(n25708), .B(n21701), .C(index_i[5]), .Z(n21702)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22328_3_lut.init = 16'hcaca;
    PFUMX i20401 (.BLUT(n22855), .ALUT(n22856), .C0(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_2141[9]));
    LUT4 i19657_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n22094)) /* synthesis lut_function=(!(A ((D)+!C)+!A !(B ((D)+!C)+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19657_3_lut_3_lut_4_lut.init = 16'h55a4;
    L6MUX21 i20854 (.D0(n23306), .D1(n23307), .SD(index_i[8]), .Z(n23310));
    PFUMX i20871 (.BLUT(n23325), .ALUT(n23326), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2126[8]));
    LUT4 mux_197_Mux_0_i589_3_lut (.A(n27086), .B(n588), .C(index_q[3]), 
         .Z(n589)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i589_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_0_i781_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n781_adj_2597)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A (B (C)+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_0_i781_4_lut_4_lut_4_lut.init = 16'h0cb4;
    PFUMX i9571 (.BLUT(n12164), .ALUT(n12165), .C0(n22413), .Z(n12134));
    PFUMX i20545 (.BLUT(n22999), .ALUT(n23000), .C0(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_2141[2]));
    PFUMX i9494 (.BLUT(n12160), .ALUT(n12161), .C0(n22406), .Z(n12055));
    LUT4 mux_196_Mux_0_i491_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n491_adj_2777)) /* synthesis lut_function=(!(A (B (D)+!B !(C+!(D)))+!A ((C+!(D))+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_0_i491_3_lut_4_lut.init = 16'h24aa;
    LUT4 i1_2_lut_rep_570_3_lut (.A(index_q[2]), .B(index_q[0]), .C(index_q[1]), 
         .Z(n26893)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_2_lut_rep_570_3_lut.init = 16'hfefe;
    LUT4 mux_197_Mux_5_i954_3_lut_4_lut_4_lut (.A(index_q[2]), .B(index_q[0]), 
         .C(index_q[3]), .D(index_q[1]), .Z(n954_adj_2608)) /* synthesis lut_function=(!(A (C)+!A (B+((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_5_i954_3_lut_4_lut_4_lut.init = 16'h0a1a;
    LUT4 mux_196_Mux_5_i781_3_lut_4_lut_4_lut_then_4_lut (.A(index_i[3]), 
         .B(index_i[0]), .C(index_i[4]), .D(index_i[2]), .Z(n27136)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_5_i781_3_lut_4_lut_4_lut_then_4_lut.init = 16'hece0;
    LUT4 n476_bdd_3_lut_23421_3_lut (.A(index_i[1]), .B(index_i[4]), .C(n124_adj_2506), 
         .Z(n24902)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n476_bdd_3_lut_23421_3_lut.init = 16'hd1d1;
    LUT4 mux_197_Mux_2_i731_3_lut_3_lut_4_lut (.A(index_q[2]), .B(index_q[3]), 
         .C(index_q[1]), .D(index_q[0]), .Z(n731_adj_2604)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(B (C)+!B !(C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_2_i731_3_lut_3_lut_4_lut.init = 16'h69f0;
    LUT4 n172_bdd_2_lut_3_lut_3_lut_4_lut (.A(index_q[2]), .B(index_q[0]), 
         .C(index_q[1]), .D(index_q[3]), .Z(n25828)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B ((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n172_bdd_2_lut_3_lut_3_lut_4_lut.init = 16'h00fe;
    LUT4 mux_196_Mux_5_i781_3_lut_4_lut_4_lut_else_4_lut (.A(index_i[3]), 
         .B(index_i[0]), .C(index_i[4]), .Z(n27135)) /* synthesis lut_function=(!(A (C)+!A (B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_5_i781_3_lut_4_lut_4_lut_else_4_lut.init = 16'h1f1f;
    LUT4 mux_197_Mux_6_i924_3_lut_4_lut (.A(index_q[2]), .B(index_q[3]), 
         .C(index_q[4]), .D(n908_adj_2592), .Z(n924_adj_2747)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_6_i924_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_197_Mux_2_i763_4_lut_4_lut (.A(index_q[0]), .B(n11977), .C(index_q[4]), 
         .D(n157_adj_2752), .Z(n763_adj_2724)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_2_i763_4_lut_4_lut.init = 16'hdfd0;
    LUT4 mux_196_Mux_3_i653_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n653_adj_2707)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A !(B (D)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_3_i653_3_lut_4_lut_4_lut.init = 16'h4d99;
    LUT4 mux_197_Mux_2_i349_3_lut_3_lut (.A(index_q[0]), .B(index_q[4]), 
         .C(n348_adj_2778), .Z(n349_adj_2720)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_2_i349_3_lut_3_lut.init = 16'hd1d1;
    LUT4 mux_197_Mux_2_i507_3_lut_3_lut (.A(index_q[0]), .B(index_q[4]), 
         .C(n491_adj_2374), .Z(n507_adj_2723)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_2_i507_3_lut_3_lut.init = 16'h7474;
    LUT4 i9393_3_lut_4_lut_4_lut (.A(index_q[0]), .B(n29493), .C(index_q[4]), 
         .D(index_q[3]), .Z(n605_adj_2756)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A !(B+(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9393_3_lut_4_lut_4_lut.init = 16'h555c;
    LUT4 mux_197_Mux_5_i573_3_lut_3_lut (.A(index_q[0]), .B(index_q[4]), 
         .C(n572_adj_2779), .Z(n573_adj_2755)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_5_i573_3_lut_3_lut.init = 16'hd1d1;
    LUT4 i11789_2_lut_3_lut_3_lut (.A(index_q[0]), .B(index_q[3]), .C(index_q[2]), 
         .Z(n14464)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11789_2_lut_3_lut_3_lut.init = 16'h4040;
    LUT4 mux_196_Mux_5_i475_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n475_adj_2728)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_5_i475_3_lut_4_lut_4_lut.init = 16'hd4a5;
    PFUMX mux_197_Mux_14_i1023 (.BLUT(n511_adj_2733), .ALUT(n20197), .C0(index_q[9]), 
          .Z(quarter_wave_sample_register_q_15__N_2141[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 i11633_4_lut (.A(n26870), .B(index_q[7]), .C(n892_adj_2441), 
         .D(index_q[6]), .Z(n1021_adj_2725)) /* synthesis lut_function=(A (B+(C (D)))+!A (B+(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11633_4_lut.init = 16'hfcdd;
    LUT4 mux_197_Mux_4_i142_3_lut_4_lut_3_lut (.A(index_q[0]), .B(index_q[3]), 
         .C(index_q[2]), .Z(n142_adj_2655)) /* synthesis lut_function=(A (B (C))+!A !(B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_4_i142_3_lut_4_lut_3_lut.init = 16'h9595;
    LUT4 mux_196_Mux_0_i157_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n157_adj_2722)) /* synthesis lut_function=(A (B (C+!(D))+!B !(D))+!A (B (D)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_0_i157_3_lut_4_lut.init = 16'hd4aa;
    LUT4 mux_197_Mux_6_i908_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), 
         .B(index_q[1]), .C(index_q[3]), .D(index_q[2]), .Z(n908_adj_2592)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A (B (C (D)+!C !(D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_6_i908_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h1cf0;
    LUT4 mux_197_Mux_4_i221_3_lut_3_lut (.A(index_q[0]), .B(index_q[4]), 
         .C(n205_adj_2780), .Z(n221_adj_2765)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_4_i221_3_lut_3_lut.init = 16'h7474;
    LUT4 i19167_3_lut_3_lut_4_lut (.A(n26863), .B(index_q[4]), .C(n700), 
         .D(index_q[5]), .Z(n21604)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19167_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 mux_196_Mux_0_i557_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n557_adj_2521)) /* synthesis lut_function=(A ((D)+!C)+!A !((D)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_0_i557_3_lut_4_lut.init = 16'haa4e;
    LUT4 i19344_3_lut (.A(n27072), .B(n27070), .C(index_q[3]), .Z(n21781)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19344_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_3_i444_3_lut_4_lut (.A(index_q[0]), .B(index_q[3]), 
         .C(n27090), .D(index_q[4]), .Z(n444_adj_2772)) /* synthesis lut_function=(!(A (B (D)+!B (C (D)))+!A !(B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_3_i444_3_lut_4_lut.init = 16'h46aa;
    LUT4 n572_bdd_3_lut_24632_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .D(index_i[3]), .Z(n25608)) /* synthesis lut_function=(A (B (C+(D)))+!A (B ((D)+!C)+!B !((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n572_bdd_3_lut_24632_4_lut.init = 16'hcc94;
    LUT4 i21663_3_lut (.A(n21781), .B(n21782), .C(index_q[4]), .Z(n21783)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21663_3_lut.init = 16'hcaca;
    LUT4 n476_bdd_3_lut_23890 (.A(n476_adj_2423), .B(n25408), .C(index_q[5]), 
         .Z(n25409)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n476_bdd_3_lut_23890.init = 16'hcaca;
    LUT4 mux_197_Mux_4_i252_4_lut_4_lut (.A(index_q[0]), .B(index_q[3]), 
         .C(n27063), .D(index_q[4]), .Z(n252_adj_2766)) /* synthesis lut_function=(!(A (B (D)+!B !(D))+!A !(B ((D)+!C)+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_4_i252_4_lut_4_lut.init = 16'h669d;
    LUT4 mux_197_Mux_1_i62_3_lut_4_lut (.A(index_q[0]), .B(index_q[3]), 
         .C(index_q[2]), .D(index_q[4]), .Z(n62_adj_2749)) /* synthesis lut_function=(A (B (D)+!B ((D)+!C))+!A !(B (D)+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_1_i62_3_lut_4_lut.init = 16'haa56;
    LUT4 mux_197_Mux_10_i701_4_lut_4_lut (.A(n26863), .B(index_q[4]), .C(index_q[5]), 
         .D(n26774), .Z(n701_adj_2588)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B (C (D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_10_i701_4_lut_4_lut.init = 16'h3efe;
    L6MUX21 i12912362_i1 (.D0(n23281), .D1(n23434), .SD(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_2141[0]));
    LUT4 i19341_3_lut (.A(n1001), .B(n588), .C(index_q[3]), .Z(n21778)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19341_3_lut.init = 16'hcaca;
    L6MUX21 i12900356_i1 (.D0(n23219), .D1(n23496), .SD(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2126[0]));
    PFUMX i24027 (.BLUT(n25829), .ALUT(n25828), .C0(index_q[4]), .Z(n25830));
    PFUMX mux_196_Mux_14_i1023 (.BLUT(n511), .ALUT(n20198), .C0(index_i[9]), 
          .Z(quarter_wave_sample_register_i_15__N_2126[13])) /* synthesis LSE_LINE_FILE_ID=3, LSE_LCOL=70, LSE_RCOL=134, LSE_LLINE=21, LSE_RLINE=21 */ ;
    LUT4 i21665_3_lut (.A(n21778), .B(n21779), .C(index_q[4]), .Z(n21780)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21665_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_2_i653_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n653_adj_2703)) /* synthesis lut_function=(A (B (C+!(D))+!B !(D))+!A !(B (C+!(D))+!B !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_2_i653_3_lut_4_lut.init = 16'h94aa;
    LUT4 mux_196_Mux_3_i684_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[4]), .Z(n684_adj_2770)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A !(B ((D)+!C)+!B (C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_3_i684_3_lut_3_lut_4_lut.init = 16'h5594;
    LUT4 i11446_4_lut (.A(n26874), .B(index_i[7]), .C(n892_adj_2451), 
         .D(index_i[6]), .Z(n1021)) /* synthesis lut_function=(A (B+(C (D)))+!A (B+(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11446_4_lut.init = 16'hfcdd;
    L6MUX21 i23092 (.D0(n24808), .D1(n24806), .SD(index_q[6]), .Z(n24809));
    L6MUX21 i24014 (.D0(n25816), .D1(n25814), .SD(index_q[5]), .Z(n25817));
    LUT4 mux_196_Mux_3_i747_3_lut (.A(n27024), .B(n404), .C(index_i[3]), 
         .Z(n747_adj_2269)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_3_i747_3_lut.init = 16'hcaca;
    PFUMX i24012 (.BLUT(n572_adj_2779), .ALUT(n25815), .C0(index_q[4]), 
          .Z(n25816));
    PFUMX i24010 (.BLUT(n25813), .ALUT(n25812), .C0(index_q[4]), .Z(n25814));
    PFUMX i23090 (.BLUT(n24807), .ALUT(n62_adj_2590), .C0(index_q[5]), 
          .Z(n24808));
    LUT4 n476_bdd_3_lut_23415_3_lut (.A(index_q[1]), .B(index_q[4]), .C(n124_adj_2515), 
         .Z(n25096)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n476_bdd_3_lut_23415_3_lut.init = 16'hd1d1;
    LUT4 mux_197_Mux_7_i956_3_lut_3_lut_4_lut (.A(n26863), .B(index_q[4]), 
         .C(n924_adj_2768), .D(index_q[5]), .Z(n956_adj_2628)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_7_i956_3_lut_3_lut_4_lut.init = 16'h11f0;
    LUT4 mux_197_Mux_6_i636_4_lut_4_lut (.A(index_q[1]), .B(index_q[4]), 
         .C(n635_adj_2419), .D(n14464), .Z(n636_adj_2738)) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_6_i636_4_lut_4_lut.init = 16'hf3d1;
    L6MUX21 i24003 (.D0(n25805), .D1(n25803), .SD(index_q[4]), .Z(n25806));
    PFUMX i24001 (.BLUT(n25804), .ALUT(n26732), .C0(index_q[5]), .Z(n25805));
    LUT4 i1_2_lut_rep_671 (.A(index_q[3]), .B(index_q[2]), .Z(n26994)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_2_lut_rep_671.init = 16'heeee;
    PFUMX i23088 (.BLUT(n24805), .ALUT(n24804), .C0(index_q[5]), .Z(n24806));
    LUT4 i19333_3_lut (.A(n29493), .B(n27077), .C(index_q[3]), .Z(n21770)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19333_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_11_i766_3_lut (.A(n638), .B(n765), .C(index_q[7]), 
         .Z(n766_adj_2682)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_11_i766_3_lut.init = 16'h3a3a;
    LUT4 mux_197_Mux_0_i46_3_lut_4_lut_4_lut_4_lut (.A(index_q[2]), .B(index_q[0]), 
         .C(index_q[1]), .D(index_q[3]), .Z(n46_adj_2304)) /* synthesis lut_function=(A (D)+!A (B+(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i46_3_lut_4_lut_4_lut_4_lut.init = 16'hfe55;
    LUT4 i11247_3_lut_3_lut_3_lut (.A(index_q[1]), .B(index_q[2]), .C(index_q[0]), 
         .Z(n652)) /* synthesis lut_function=(!(A ((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11247_3_lut_3_lut_3_lut.init = 16'h5d5d;
    LUT4 mux_197_Mux_9_i285_3_lut_4_lut_4_lut (.A(index_q[2]), .B(index_q[0]), 
         .C(index_q[3]), .D(index_q[1]), .Z(n285_adj_2399)) /* synthesis lut_function=(A (C)+!A !(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_9_i285_3_lut_4_lut_4_lut.init = 16'ha0a1;
    LUT4 i11697_2_lut_rep_536_3_lut (.A(index_q[3]), .B(index_q[2]), .C(index_q[1]), 
         .Z(n26859)) /* synthesis lut_function=(A+(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11697_2_lut_rep_536_3_lut.init = 16'hfefe;
    LUT4 i7656_2_lut_rep_644 (.A(index_q[3]), .B(index_q[4]), .Z(n26967)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i7656_2_lut_rep_644.init = 16'heeee;
    LUT4 i9372_3_lut_4_lut (.A(index_q[3]), .B(index_q[4]), .C(n27075), 
         .D(n29485), .Z(n605_adj_2737)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9372_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i9399_3_lut_3_lut_4_lut (.A(index_q[3]), .B(index_q[2]), .C(index_q[1]), 
         .D(index_q[0]), .Z(n812_adj_2581)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9399_3_lut_3_lut_4_lut.init = 16'h1ef0;
    LUT4 i1_3_lut_rep_517_4_lut (.A(index_q[3]), .B(index_q[4]), .C(index_q[2]), 
         .D(n27085), .Z(n26840)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_3_lut_rep_517_4_lut.init = 16'hfffe;
    LUT4 i1_3_lut_4_lut_adj_89 (.A(index_q[3]), .B(index_q[4]), .C(index_q[5]), 
         .D(n27090), .Z(n20333)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i1_3_lut_4_lut_adj_89.init = 16'hfffe;
    LUT4 n21464_bdd_3_lut_3_lut (.A(index_q[1]), .B(n812_adj_2581), .C(index_q[4]), 
         .Z(n25098)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n21464_bdd_3_lut_3_lut.init = 16'h5c5c;
    LUT4 mux_196_Mux_4_i491_3_lut_4_lut_4_lut (.A(index_i[2]), .B(n29491), 
         .C(index_i[3]), .D(n26996), .Z(n491_adj_2636)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_4_i491_3_lut_4_lut_4_lut.init = 16'hfc5c;
    PFUMX i20799 (.BLUT(n142_adj_2781), .ALUT(n157), .C0(index_q[4]), 
          .Z(n23255));
    LUT4 i19327_3_lut (.A(n27080), .B(n27097), .C(index_q[3]), .Z(n21764)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19327_3_lut.init = 16'hcaca;
    PFUMX i23999 (.BLUT(n25802), .ALUT(n25801), .C0(index_q[5]), .Z(n25803));
    LUT4 i19326_3_lut (.A(n356), .B(n204_adj_2732), .C(index_q[3]), .Z(n21763)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19326_3_lut.init = 16'hcaca;
    LUT4 index_i_6__bdd_4_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[6]), 
         .C(index_i[5]), .D(n26882), .Z(n24999)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (D))+!A (B (C (D))+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam index_i_6__bdd_4_lut_4_lut_4_lut.init = 16'h04f7;
    LUT4 mux_197_Mux_3_i349_3_lut_3_lut (.A(index_q[1]), .B(index_q[4]), 
         .C(n348_adj_2745), .Z(n349_adj_2771)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_3_i349_3_lut_3_lut.init = 16'hd1d1;
    LUT4 i11264_2_lut_rep_449_3_lut_4_lut (.A(index_q[2]), .B(index_q[0]), 
         .C(index_q[3]), .D(index_q[1]), .Z(n26772)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11264_2_lut_rep_449_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i11528_3_lut_3_lut_4_lut_4_lut (.A(index_i[2]), .B(index_i[3]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n14203)) /* synthesis lut_function=(!(A ((C+(D))+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11528_3_lut_3_lut_4_lut_4_lut.init = 16'h555d;
    LUT4 i23837_then_4_lut (.A(index_i[0]), .B(index_i[4]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n27231)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)+!C !(D))+!B (C (D)))) */ ;
    defparam i23837_then_4_lut.init = 16'hda0e;
    LUT4 i11785_3_lut_4_lut_4_lut_4_lut (.A(index_q[1]), .B(n27034), .C(index_q[4]), 
         .D(index_q[0]), .Z(n14460)) /* synthesis lut_function=(!(A (((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11785_3_lut_4_lut_4_lut_4_lut.init = 16'h55d5;
    LUT4 i23837_else_4_lut (.A(index_i[0]), .B(index_i[4]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n27230)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C))+!A (B (C)+!B (C+(D)))) */ ;
    defparam i23837_else_4_lut.init = 16'hf178;
    LUT4 mux_196_Mux_11_i766_3_lut (.A(n638_adj_2710), .B(n765_adj_2289), 
         .C(index_i[7]), .Z(n766)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_11_i766_3_lut.init = 16'h3a3a;
    LUT4 mux_197_Mux_8_i716_3_lut_4_lut_4_lut_4_lut (.A(index_q[2]), .B(index_q[0]), 
         .C(index_q[1]), .D(index_q[3]), .Z(n716_adj_2557)) /* synthesis lut_function=(!(A (D)+!A !(B+(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_8_i716_3_lut_4_lut_4_lut_4_lut.init = 16'h55fe;
    LUT4 i11036_2_lut_rep_770 (.A(index_q[0]), .B(index_q[1]), .Z(n27093)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11036_2_lut_rep_770.init = 16'h4444;
    PFUMX i20800 (.BLUT(n173_adj_2593), .ALUT(n188), .C0(index_q[4]), 
          .Z(n23256));
    LUT4 i19158_3_lut_3_lut_4_lut (.A(n26864), .B(index_i[4]), .C(n700_adj_2293), 
         .D(index_i[5]), .Z(n21595)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19158_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 mux_196_Mux_5_i924_4_lut_3_lut (.A(index_i[2]), .B(n14871), .C(index_i[4]), 
         .Z(n924)) /* synthesis lut_function=(!(A (B+(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_5_i924_4_lut_3_lut.init = 16'h5656;
    LUT4 i20563_3_lut (.A(n308), .B(n29468), .C(index_i[3]), .Z(n23019)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20563_3_lut.init = 16'hcaca;
    LUT4 i7503_2_lut_rep_672 (.A(index_i[3]), .B(index_i[4]), .Z(n26995)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i7503_2_lut_rep_672.init = 16'heeee;
    LUT4 mux_197_Mux_2_i908_3_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[0]), .D(index_q[3]), .Z(n908_adj_2408)) /* synthesis lut_function=(!(A (B+!(D))+!A !(B+!(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_2_i908_3_lut_4_lut_4_lut.init = 16'h6645;
    LUT4 i20562_3_lut (.A(n619), .B(n29491), .C(index_i[3]), .Z(n23018)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20562_3_lut.init = 16'hcaca;
    LUT4 i6529_2_lut_rep_740 (.A(index_q[1]), .B(index_q[2]), .Z(n27063)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i6529_2_lut_rep_740.init = 16'heeee;
    LUT4 mux_196_Mux_10_i701_4_lut_4_lut (.A(n26864), .B(index_i[4]), .C(index_i[5]), 
         .D(n26776), .Z(n701)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B (C (D))+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_10_i701_4_lut_4_lut.init = 16'h3efe;
    LUT4 i11729_2_lut_rep_511_3_lut (.A(index_q[1]), .B(index_q[2]), .C(index_q[0]), 
         .Z(n26834)) /* synthesis lut_function=(A (C)+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11729_2_lut_rep_511_3_lut.init = 16'hf1f1;
    LUT4 i11530_2_lut_rep_525_2_lut (.A(index_i[1]), .B(index_i[0]), .Z(n26848)) /* synthesis lut_function=(!(A+!(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11530_2_lut_rep_525_2_lut.init = 16'h4444;
    LUT4 i20561_3_lut (.A(n29472), .B(n27001), .C(index_i[3]), .Z(n23017)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20561_3_lut.init = 16'hcaca;
    LUT4 i20560_3_lut (.A(n29468), .B(n26999), .C(index_i[3]), .Z(n23016)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20560_3_lut.init = 16'hcaca;
    PFUMX i24726 (.BLUT(n27116), .ALUT(n27117), .C0(index_q[2]), .Z(n27118));
    LUT4 i1_3_lut_rep_537_4_lut (.A(index_i[3]), .B(index_i[4]), .C(index_i[2]), 
         .D(n26996), .Z(n26860)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i1_3_lut_rep_537_4_lut.init = 16'hfffe;
    L6MUX21 i23076 (.D0(n24786), .D1(n24784), .SD(index_i[6]), .Z(n24787));
    LUT4 mux_197_Mux_4_i236_3_lut_4_lut_3_lut_rep_733_4_lut (.A(index_q[1]), 
         .B(index_q[2]), .C(index_q[3]), .D(index_q[0]), .Z(n27056)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_4_i236_3_lut_4_lut_3_lut_rep_733_4_lut.init = 16'hf01f;
    LUT4 mux_196_Mux_7_i956_3_lut_3_lut_4_lut (.A(n26864), .B(index_i[4]), 
         .C(n924_adj_2758), .D(index_i[5]), .Z(n956)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_7_i956_3_lut_3_lut_4_lut.init = 16'h11f0;
    LUT4 i9514_3_lut_3_lut_4_lut (.A(index_i[3]), .B(index_i[4]), .C(n27025), 
         .D(index_i[0]), .Z(n605_adj_2452)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9514_3_lut_3_lut_4_lut.init = 16'h10fe;
    LUT4 mux_197_Mux_9_i93_3_lut_3_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .Z(n93_adj_2274)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_9_i93_3_lut_3_lut.init = 16'hc1c1;
    LUT4 n10942_bdd_3_lut_24671_4_lut_4_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[4]), .D(index_q[3]), .Z(n24488)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C+(D)))+!A (B (C (D)+!C !(D))+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n10942_bdd_3_lut_24671_4_lut_4_lut_4_lut.init = 16'hc10f;
    PFUMX i23074 (.BLUT(n24785), .ALUT(n62), .C0(index_i[5]), .Z(n24786));
    LUT4 i11482_2_lut_rep_549_3_lut (.A(index_q[1]), .B(index_q[2]), .C(index_q[3]), 
         .Z(n26872)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11482_2_lut_rep_549_3_lut.init = 16'he0e0;
    PFUMX i19097 (.BLUT(n21532), .ALUT(n21533), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2126[11]));
    LUT4 i1_3_lut_4_lut_adj_90 (.A(index_i[3]), .B(index_i[4]), .C(index_i[5]), 
         .D(n27046), .Z(n20334)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i1_3_lut_4_lut_adj_90.init = 16'hfffe;
    PFUMX i23072 (.BLUT(n24783), .ALUT(n24782), .C0(index_i[5]), .Z(n24784));
    PFUMX i20805 (.BLUT(n333), .ALUT(n348_adj_2554), .C0(index_q[4]), 
          .Z(n23261));
    LUT4 i11550_2_lut_rep_673 (.A(index_i[0]), .B(index_i[1]), .Z(n26996)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11550_2_lut_rep_673.init = 16'h8888;
    LUT4 i11483_2_lut_rep_450_3_lut_4_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[4]), .D(index_q[3]), .Z(n26773)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11483_2_lut_rep_450_3_lut_4_lut.init = 16'hfef0;
    LUT4 i9592_3_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[4]), 
         .Z(n12157)) /* synthesis lut_function=(A (B)+!A !(B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9592_3_lut_4_lut_3_lut.init = 16'h9898;
    LUT4 i18972_3_lut_3_lut_4_lut (.A(index_q[1]), .B(index_q[2]), .C(index_q[3]), 
         .D(index_q[0]), .Z(n21409)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18972_3_lut_3_lut_4_lut.init = 16'h0fe0;
    PFUMX i20806 (.BLUT(n364_adj_2782), .ALUT(n379_adj_2310), .C0(index_q[4]), 
          .Z(n23262));
    LUT4 i19345_3_lut_3_lut_3_lut (.A(index_q[1]), .B(index_q[2]), .C(index_q[3]), 
         .Z(n21782)) /* synthesis lut_function=(A (C)+!A (B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19345_3_lut_3_lut_3_lut.init = 16'he5e5;
    LUT4 mux_197_Mux_1_i890_4_lut_4_lut_4_lut_4_lut (.A(index_q[3]), .B(index_q[4]), 
         .C(n26887), .D(index_q[0]), .Z(n890_adj_2754)) /* synthesis lut_function=(!(A (B (D)+!B !(C))+!A (B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_1_i890_4_lut_4_lut_4_lut_4_lut.init = 16'h31fd;
    LUT4 i20537_3_lut (.A(n25806), .B(n22984), .C(index_q[6]), .Z(n22993)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20537_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_0_i954_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n954)) /* synthesis lut_function=(A (D)+!A !(B (C (D)+!C !(D))+!B (C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i954_3_lut_4_lut_4_lut.init = 16'haf40;
    LUT4 i20467_3_lut_4_lut_3_lut (.A(index_q[3]), .B(index_q[4]), .C(n26861), 
         .Z(n22923)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20467_3_lut_4_lut_3_lut.init = 16'h6464;
    PFUMX i20807 (.BLUT(n397_adj_2370), .ALUT(n412), .C0(index_q[4]), 
          .Z(n23263));
    LUT4 i21765_3_lut (.A(n620_adj_2783), .B(n14525), .C(index_q[4]), 
         .Z(n21740)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21765_3_lut.init = 16'hcaca;
    LUT4 i19033_3_lut (.A(n27100), .B(n27103), .C(index_q[3]), .Z(n21470)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i19033_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_1_i987_3_lut_4_lut_4_lut (.A(index_q[3]), .B(n986_adj_2619), 
         .C(index_q[4]), .D(n27058), .Z(n987_adj_2751)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_1_i987_3_lut_4_lut_4_lut.init = 16'hc5c0;
    PFUMX i19103 (.BLUT(n21538), .ALUT(n21539), .C0(index_q[9]), .Z(quarter_wave_sample_register_q_15__N_2141[11]));
    LUT4 i8831_4_lut_4_lut (.A(index_q[3]), .B(index_q[0]), .C(index_q[1]), 
         .D(index_q[2]), .Z(n11354)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (D)+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i8831_4_lut_4_lut.init = 16'h0bf4;
    L6MUX21 i23937 (.D0(n25735), .D1(n25732), .SD(index_q[5]), .Z(n25736));
    LUT4 i11079_4_lut_4_lut (.A(index_q[3]), .B(index_q[2]), .C(index_q[0]), 
         .D(index_q[1]), .Z(n875)) /* synthesis lut_function=((B (C)+!B (D))+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11079_4_lut_4_lut.init = 16'hf7d5;
    LUT4 i21800_3_lut (.A(n21469), .B(n21470), .C(index_q[4]), .Z(n21471)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21800_3_lut.init = 16'hcaca;
    PFUMX i23935 (.BLUT(n25734), .ALUT(n25733), .C0(index_q[4]), .Z(n25735));
    LUT4 i19312_4_lut_3_lut (.A(index_q[3]), .B(index_q[4]), .C(n26871), 
         .Z(n21749)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19312_4_lut_3_lut.init = 16'h6565;
    LUT4 mux_197_Mux_2_i221_4_lut_4_lut (.A(index_q[3]), .B(index_q[4]), 
         .C(n26871), .D(n26753), .Z(n221_adj_2719)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (B+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_2_i221_4_lut_4_lut.init = 16'hf7c4;
    LUT4 mux_196_Mux_3_i1002_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n19881)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (D))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_3_i1002_3_lut_3_lut_4_lut.init = 16'hf708;
    LUT4 i9559_3_lut_3_lut (.A(index_q[3]), .B(index_q[4]), .C(n12120), 
         .Z(n12121)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9559_3_lut_3_lut.init = 16'h7474;
    PFUMX i20808 (.BLUT(n428_adj_2303), .ALUT(n443), .C0(index_q[4]), 
          .Z(n23264));
    LUT4 i11048_2_lut_rep_741 (.A(index_q[0]), .B(index_q[1]), .Z(n27064)) /* synthesis lut_function=((B)+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11048_2_lut_rep_741.init = 16'hdddd;
    LUT4 i11496_3_lut_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n14171)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (D))+!A (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11496_3_lut_3_lut_3_lut_4_lut.init = 16'h00f7;
    LUT4 i11503_2_lut_2_lut_3_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .Z(n14178)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11503_2_lut_2_lut_3_lut.init = 16'h0808;
    PFUMX i20809 (.BLUT(n460), .ALUT(n475_adj_2364), .C0(index_q[4]), 
          .Z(n23265));
    LUT4 i7137_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n157_adj_2499)) /* synthesis lut_function=(!(A (C (D))+!A !(B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i7137_3_lut_4_lut_4_lut.init = 16'h4aaa;
    PFUMX i20810 (.BLUT(n491_adj_2477), .ALUT(n11354), .C0(index_q[4]), 
          .Z(n23266));
    LUT4 mux_196_Mux_8_i635_3_lut_4_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n635_adj_2341)) /* synthesis lut_function=(!(A (B (C (D))+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_8_i635_3_lut_4_lut_3_lut_4_lut.init = 16'h0ff8;
    LUT4 i22732_2_lut_rep_498_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n26821)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i22732_2_lut_rep_498_3_lut_4_lut.init = 16'h0007;
    LUT4 i19320_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n21757)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (D))+!A !(D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19320_3_lut_4_lut_4_lut_4_lut.init = 16'ha25d;
    LUT4 mux_197_Mux_0_i635_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n635_adj_2252)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i635_3_lut_4_lut_4_lut.init = 16'hfd0a;
    LUT4 mux_196_Mux_4_i1002_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n1002_adj_2715)) /* synthesis lut_function=(A (B (C (D))+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_4_i1002_3_lut_3_lut_4_lut.init = 16'hf007;
    LUT4 mux_197_Mux_6_i396_3_lut_4_lut_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n356)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_6_i396_3_lut_4_lut_3_lut.init = 16'h6d6d;
    LUT4 i12422_2_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(n27045), 
         .D(index_i[2]), .Z(n15124)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i12422_2_lut_3_lut_4_lut.init = 16'hf080;
    LUT4 mux_197_Mux_0_i316_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n316_adj_2527)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+(D)))+!A (B (C+(D))+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i316_3_lut_4_lut_4_lut_4_lut.init = 16'h332d;
    PFUMX i23932 (.BLUT(n78), .ALUT(n25731), .C0(index_q[4]), .Z(n25732));
    LUT4 i19647_3_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[3]), 
         .D(index_i[2]), .Z(n22084)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A (B (C)+!B !(C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19647_3_lut_4_lut_4_lut.init = 16'h3c8c;
    LUT4 mux_197_Mux_6_i60_3_lut_4_lut_3_lut_rep_742 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n27065)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_6_i60_3_lut_4_lut_3_lut_rep_742.init = 16'hd6d6;
    LUT4 mux_197_Mux_2_i773_3_lut_rep_743 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n27066)) /* synthesis lut_function=(A (B+!(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_2_i773_3_lut_rep_743.init = 16'hdada;
    LUT4 n123_bdd_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n25444)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !(C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n123_bdd_3_lut_4_lut_4_lut.init = 16'ha5ad;
    LUT4 i19710_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n22147)) /* synthesis lut_function=(!(A (B (C (D))+!B (C (D)+!C !(D)))+!A !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19710_3_lut_4_lut_4_lut.init = 16'h5aad;
    LUT4 i18996_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21433)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18996_3_lut_4_lut_4_lut.init = 16'hda5a;
    LUT4 i19741_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n22178)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C))+!A !(B (C)+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19741_3_lut_4_lut_4_lut.init = 16'h5ad3;
    LUT4 i18961_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21398)) /* synthesis lut_function=(A (B (C)+!B !(C (D)+!C !(D)))+!A (B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18961_3_lut_4_lut_4_lut.init = 16'hd6a5;
    LUT4 n21321_bdd_3_lut_23996_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n25447)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C))+!A !(B (C+!(D))+!B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n21321_bdd_3_lut_23996_4_lut_4_lut.init = 16'h5ad6;
    LUT4 i11316_2_lut_rep_745 (.A(index_q[0]), .B(index_q[1]), .Z(n27068)) /* synthesis lut_function=(A+!(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11316_2_lut_rep_745.init = 16'hbbbb;
    LUT4 i19045_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n21482)) /* synthesis lut_function=(A (C+(D))+!A !(B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19045_3_lut_4_lut_4_lut.init = 16'haba5;
    LUT4 index_q_0__bdd_4_lut_25125 (.A(index_q[0]), .B(index_q[3]), .C(index_q[1]), 
         .D(index_q[2]), .Z(n27141)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (C (D)))+!A !(B (C+!(D))+!B !(C+(D))))) */ ;
    defparam index_q_0__bdd_4_lut_25125.init = 16'h4ae7;
    LUT4 n642_bdd_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n25899)) /* synthesis lut_function=(!(A (D)+!A !(B (D)+!B (C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n642_bdd_4_lut_4_lut_4_lut.init = 16'h54bb;
    LUT4 i21803_3_lut (.A(n21466), .B(n21467), .C(index_q[4]), .Z(n21468)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21803_3_lut.init = 16'hcaca;
    LUT4 i22389_3_lut (.A(n12048), .B(n892_adj_2543), .C(index_i[6]), 
         .Z(n23319)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22389_3_lut.init = 16'hcaca;
    LUT4 i9421_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n875_adj_2622)) /* synthesis lut_function=(A (C (D))+!A !(B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9421_3_lut_4_lut_4_lut_4_lut.init = 16'hb555;
    LUT4 mux_197_Mux_6_i204_3_lut_3_lut_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n204_adj_2732)) /* synthesis lut_function=(!(A (C)+!A !((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_6_i204_3_lut_3_lut_3_lut.init = 16'h5b5b;
    LUT4 i20556_3_lut (.A(n29490), .B(n26999), .C(index_i[3]), .Z(n23012)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20556_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_1_i348_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n348_adj_2698)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A (B ((D)+!C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_1_i348_3_lut_4_lut_4_lut_4_lut.init = 16'h38f0;
    LUT4 i20555_3_lut (.A(n29472), .B(n108), .C(index_i[3]), .Z(n23011)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20555_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_0_i236_3_lut_3_lut (.A(index_q[0]), .B(index_q[2]), 
         .C(index_q[3]), .Z(n236)) /* synthesis lut_function=(A (B+(C))+!A !(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i236_3_lut_3_lut.init = 16'ha9a9;
    LUT4 mux_197_Mux_5_i459_3_lut_4_lut_3_lut_rep_747 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n27070)) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_5_i459_3_lut_4_lut_3_lut_rep_747.init = 16'h6b6b;
    LUT4 mux_197_Mux_5_i460_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n460_adj_2509)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A !(B (C)+!B !(C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_5_i460_3_lut_4_lut_4_lut.init = 16'h6b5a;
    LUT4 i20554_3_lut (.A(n619), .B(n27001), .C(index_i[3]), .Z(n23010)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20554_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_0_i364_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n364_adj_2782)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A ((C+!(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i364_3_lut_3_lut_4_lut.init = 16'hdb55;
    LUT4 i20553_3_lut (.A(n26900), .B(n26932), .C(index_i[3]), .Z(n23009)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20553_3_lut.init = 16'hcaca;
    LUT4 i19042_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21479)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D))+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19042_3_lut_4_lut.init = 16'hccdb;
    LUT4 i11314_2_lut_rep_748 (.A(index_q[0]), .B(index_q[1]), .Z(n27071)) /* synthesis lut_function=(!((B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11314_2_lut_rep_748.init = 16'h2222;
    LUT4 mux_197_Mux_4_i900_3_lut_4_lut_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n900)) /* synthesis lut_function=(A ((C)+!B)+!A !(B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_4_i900_3_lut_4_lut_3_lut.init = 16'hb2b2;
    PFUMX i19004 (.BLUT(n21439), .ALUT(n21440), .C0(index_q[4]), .Z(n21441));
    LUT4 mux_197_Mux_6_i157_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n157_adj_2752)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (D))+!A !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_6_i157_3_lut_4_lut_4_lut_4_lut.init = 16'h5d22;
    LUT4 mux_197_Mux_4_i205_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n205_adj_2780)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_4_i205_3_lut_4_lut_4_lut.init = 16'h5a2a;
    LUT4 index_q_4__bdd_3_lut_23048_4_lut (.A(n26893), .B(index_q[3]), .C(index_q[5]), 
         .D(index_q[4]), .Z(n24751)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam index_q_4__bdd_3_lut_23048_4_lut.init = 16'hf080;
    LUT4 mux_197_Mux_0_i985_3_lut_3_lut_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n985)) /* synthesis lut_function=(!(A (B+!(C))+!A (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i985_3_lut_3_lut_3_lut.init = 16'h2525;
    PFUMX i23908 (.BLUT(n25707), .ALUT(n25706), .C0(index_i[4]), .Z(n25708));
    LUT4 i9583_3_lut_4_lut_3_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[4]), 
         .Z(n12148)) /* synthesis lut_function=(!(A (B)+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9583_3_lut_4_lut_3_lut.init = 16'h6262;
    LUT4 mux_196_Mux_6_i812_3_lut_4_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n812_adj_2681)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(D))+!A !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_6_i812_3_lut_4_lut_3_lut_4_lut.init = 16'h7780;
    LUT4 mux_197_Mux_0_i652_3_lut_rep_749 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n27072)) /* synthesis lut_function=(!(A (B+(C))+!A !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i652_3_lut_rep_749.init = 16'h5252;
    LUT4 mux_197_Mux_0_i708_3_lut_4_lut_3_lut_rep_750 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n27073)) /* synthesis lut_function=(!(A (B)+!A ((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i708_3_lut_4_lut_3_lut_rep_750.init = 16'h2626;
    LUT4 mux_196_Mux_7_i526_3_lut_3_lut_4_lut_4_lut_3_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[3]), .D(index_i[2]), .Z(n526_adj_2659)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(D))+!A !(D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_7_i526_3_lut_3_lut_4_lut_4_lut_3_lut_4_lut.init = 16'h887f;
    LUT4 mux_196_Mux_8_i526_3_lut_3_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n526_adj_2340)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_8_i526_3_lut_3_lut_3_lut_4_lut.init = 16'h0f70;
    LUT4 i20355_3_lut (.A(n25582), .B(n22802), .C(index_i[6]), .Z(n22811)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20355_3_lut.init = 16'hcaca;
    LUT4 i18975_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21412)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C+!(D)))+!A !(B (C+!(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i18975_3_lut_4_lut_4_lut.init = 16'ha52b;
    LUT4 i20761_3_lut (.A(n23213), .B(n23214), .C(index_i[7]), .Z(n23217)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20761_3_lut.init = 16'hcaca;
    LUT4 i19023_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21460)) /* synthesis lut_function=(!(A (B)+!A (B (C+(D))+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19023_3_lut_3_lut_4_lut.init = 16'h3326;
    LUT4 n316_bdd_3_lut_24613_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n25632)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A !(B ((D)+!C)+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n316_bdd_3_lut_24613_3_lut_4_lut.init = 16'h552c;
    LUT4 i19317_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21754)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C))+!A !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19317_3_lut_4_lut_4_lut.init = 16'h5a52;
    LUT4 mux_197_Mux_2_i348_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n348_adj_2778)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_2_i348_3_lut_4_lut_4_lut.init = 16'h52a5;
    LUT4 i11407_2_lut_rep_513_3_lut (.A(index_i[0]), .B(index_i[1]), .C(index_i[2]), 
         .Z(n26836)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11407_2_lut_rep_513_3_lut.init = 16'hf8f8;
    LUT4 i22560_2_lut_rep_752 (.A(index_q[0]), .B(index_q[1]), .Z(n27075)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i22560_2_lut_rep_752.init = 16'h9999;
    LUT4 mux_196_Mux_8_i172_rep_34_3_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n70)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_8_i172_rep_34_3_lut_3_lut.init = 16'h7c7c;
    LUT4 mux_196_Mux_7_i491_3_lut_4_lut_4_lut_4_lut_4_lut (.A(index_i[0]), 
         .B(index_i[1]), .C(index_i[2]), .D(index_i[3]), .Z(n491)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A (B ((D)+!C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_7_i491_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'h3870;
    LUT4 i22558_2_lut_rep_650 (.A(index_q[1]), .B(index_q[2]), .Z(n26973)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i22558_2_lut_rep_650.init = 16'h9999;
    LUT4 i9370_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n541_adj_2424)) /* synthesis lut_function=(A (B (C (D))+!B !(C (D)))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9370_3_lut_4_lut_4_lut_4_lut.init = 16'h9333;
    LUT4 n442_bdd_2_lut_24016_3_lut (.A(index_q[1]), .B(index_q[2]), .C(index_q[3]), 
         .Z(n25812)) /* synthesis lut_function=(A (B+(C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n442_bdd_2_lut_24016_3_lut.init = 16'hf9f9;
    LUT4 i11073_2_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n668)) /* synthesis lut_function=(!(A ((D)+!B)+!A (B ((D)+!C)+!B (C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11073_2_lut_4_lut_4_lut_4_lut.init = 16'h00c9;
    LUT4 i15559_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n17823)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)))+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i15559_3_lut_4_lut_4_lut_4_lut.init = 16'h3999;
    LUT4 mux_197_Mux_0_i93_3_lut_3_lut (.A(index_q[1]), .B(index_q[2]), 
         .C(index_q[3]), .Z(n93_adj_2775)) /* synthesis lut_function=(A (B)+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i93_3_lut_3_lut.init = 16'h9c9c;
    LUT4 i3596_2_lut_rep_651 (.A(index_q[0]), .B(index_q[2]), .Z(n26974)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i3596_2_lut_rep_651.init = 16'h6666;
    LUT4 mux_196_Mux_7_i308_3_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .Z(n308)) /* synthesis lut_function=(A ((C)+!B)+!A (B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_7_i308_3_lut_4_lut_3_lut.init = 16'he7e7;
    LUT4 mux_197_Mux_5_i483_rep_771 (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .Z(n27094)) /* synthesis lut_function=(!(A (C)+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_5_i483_rep_771.init = 16'h4a4a;
    LUT4 i15558_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n17822)) /* synthesis lut_function=(A (B)+!A !(B (C (D))+!B !(C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i15558_3_lut_4_lut_4_lut.init = 16'h9ccc;
    LUT4 mux_197_Mux_2_i269_3_lut_3_lut_rep_738_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n27061)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_2_i269_3_lut_3_lut_rep_738_3_lut.init = 16'h3939;
    L6MUX21 i23046 (.D0(n24752), .D1(n26706), .SD(index_q[6]), .Z(n24753));
    LUT4 mux_197_Mux_6_i315_rep_772 (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .Z(n27095)) /* synthesis lut_function=(A (C)+!A !((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_6_i315_rep_772.init = 16'ha4a4;
    LUT4 i19728_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n22165)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !(B (C+!(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19728_3_lut_4_lut_4_lut.init = 16'ha5a9;
    LUT4 i9408_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(n27034), .D(index_q[4]), .Z(n189_adj_2692)) /* synthesis lut_function=(A (B (C (D)))+!A !(B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i9408_3_lut_4_lut_4_lut_4_lut.init = 16'h9555;
    PFUMX i23044 (.BLUT(n24751), .ALUT(n26733), .C0(index_q[7]), .Z(n24752));
    LUT4 mux_197_Mux_5_i572_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n572_adj_2779)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A !(B (C+(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_5_i572_3_lut_4_lut_4_lut.init = 16'ha9a5;
    L6MUX21 i23888 (.D0(n25671), .D1(n25668), .SD(index_i[5]), .Z(n25672));
    LUT4 i20039_3_lut (.A(n22490), .B(n22491), .C(index_q[7]), .Z(n22495)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20039_3_lut.init = 16'hcaca;
    PFUMX i23886 (.BLUT(n25670), .ALUT(n25669), .C0(index_i[4]), .Z(n25671));
    LUT4 i15523_3_lut_3_lut (.A(index_q[0]), .B(index_q[2]), .C(index_q[3]), 
         .Z(n17787)) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i15523_3_lut_3_lut.init = 16'h6a6a;
    LUT4 mux_196_Mux_3_i890_3_lut_4_lut (.A(n26851), .B(index_i[2]), .C(index_i[3]), 
         .D(n396), .Z(n890_adj_2709)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_3_i890_3_lut_4_lut.init = 16'h6f60;
    LUT4 n28_bdd_3_lut_24024_4_lut_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .Z(n25268)) /* synthesis lut_function=(A (B)+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n28_bdd_3_lut_24024_4_lut_3_lut.init = 16'hd9d9;
    LUT4 mux_197_Mux_5_i109_3_lut_3_lut_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .Z(n109_adj_2514)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_5_i109_3_lut_3_lut_3_lut.init = 16'h3939;
    LUT4 mux_197_Mux_2_i604_3_lut_4_lut_4_lut_4_lut_4_lut (.A(index_q[0]), 
         .B(index_q[1]), .C(index_q[3]), .D(index_q[2]), .Z(n604_adj_2609)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C (D)+!C !(D)))+!A (B (C)+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_2_i604_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'h3c9f;
    LUT4 i19495_3_lut_4_lut (.A(n26851), .B(index_i[2]), .C(index_i[3]), 
         .D(n27022), .Z(n21932)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19495_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_197_Mux_4_i349_3_lut_4_lut (.A(index_q[0]), .B(index_q[2]), 
         .C(index_q[4]), .D(n348_adj_2741), .Z(n349_adj_2767)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_4_i349_3_lut_4_lut.init = 16'hf606;
    LUT4 i19642_3_lut_4_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n22079)) /* synthesis lut_function=(!(A (B (C)+!B !(C+!(D)))+!A (B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19642_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'h383f;
    PFUMX i23883 (.BLUT(n301_adj_2679), .ALUT(n25667), .C0(index_i[4]), 
          .Z(n25668));
    LUT4 i11077_2_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[3]), 
         .D(index_q[2]), .Z(n844)) /* synthesis lut_function=(A (B+!(C (D)+!C !(D)))+!A !(B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11077_2_lut_3_lut_4_lut.init = 16'h9ff9;
    LUT4 mux_197_Mux_6_i573_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[4]), .D(n572_adj_2784), .Z(n573_adj_2736)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (B (C (D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_6_i573_3_lut_4_lut.init = 16'hf909;
    LUT4 mux_197_Mux_6_i498_3_lut_4_lut_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n498)) /* synthesis lut_function=(A (B+!(C))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_6_i498_3_lut_4_lut_3_lut.init = 16'h9b9b;
    LUT4 mux_197_Mux_4_i77_3_lut_rep_753 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n27076)) /* synthesis lut_function=(A (B (C))+!A !(B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_4_i77_3_lut_rep_753.init = 16'h9595;
    LUT4 i11472_2_lut_rep_436_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n26759)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11472_2_lut_rep_436_3_lut_4_lut.init = 16'hf080;
    LUT4 mux_196_Mux_3_i94_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[4]), .D(n93_adj_2487), .Z(n94_adj_2525)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_3_i94_3_lut_4_lut.init = 16'hf606;
    LUT4 mux_197_Mux_0_i660_3_lut_rep_754 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n27077)) /* synthesis lut_function=(A (B)+!A (B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i660_3_lut_rep_754.init = 16'hc9c9;
    LUT4 mux_197_Mux_2_i262_3_lut_3_lut_rep_755 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n27078)) /* synthesis lut_function=(A (B)+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_2_i262_3_lut_3_lut_rep_755.init = 16'h9c9c;
    LUT4 mux_197_Mux_6_i308_3_lut_4_lut_3_lut_rep_756 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n27079)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_6_i308_3_lut_4_lut_3_lut_rep_756.init = 16'h9696;
    LUT4 mux_196_Mux_3_i62_3_lut_4_lut (.A(index_i[1]), .B(index_i[2]), 
         .C(index_i[4]), .D(n812_adj_2681), .Z(n62_adj_2762)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_3_i62_3_lut_4_lut.init = 16'h6f60;
    LUT4 n518_bdd_3_lut_4_lut_4_lut_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[3]), .D(index_i[2]), .Z(n25603)) /* synthesis lut_function=(A (B (C)+!B !(D))+!A !(D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam n518_bdd_3_lut_4_lut_4_lut_3_lut_4_lut.init = 16'h80f7;
    LUT4 mux_197_Mux_6_i340_3_lut_4_lut_3_lut_rep_757 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n27080)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_6_i340_3_lut_4_lut_3_lut_rep_757.init = 16'h9292;
    LUT4 i5753_1_lut_rep_652 (.A(index_i[0]), .Z(n26975)) /* synthesis lut_function=(!(A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i5753_1_lut_rep_652.init = 16'h5555;
    LUT4 mux_197_Mux_2_i308_3_lut_4_lut_3_lut_rep_773 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n27096)) /* synthesis lut_function=(A (B (C))+!A !(B (C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_2_i308_3_lut_4_lut_3_lut_rep_773.init = 16'h9494;
    LUT4 mux_196_Mux_4_i221_3_lut_3_lut (.A(index_i[0]), .B(index_i[4]), 
         .C(n205), .Z(n221_adj_2485)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_4_i221_3_lut_3_lut.init = 16'h7474;
    LUT4 mux_197_Mux_6_i540_3_lut_3_lut_3_lut_rep_758 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n27081)) /* synthesis lut_function=(A (B (C)+!B !(C))+!A !(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_6_i540_3_lut_3_lut_3_lut_rep_758.init = 16'h9393;
    LUT4 mux_197_Mux_4_i262_3_lut_3_lut_rep_759 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n27082)) /* synthesis lut_function=(A (B+(C))+!A !(B+(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_4_i262_3_lut_3_lut_rep_759.init = 16'ha9a9;
    LUT4 mux_197_Mux_0_i134_3_lut_4_lut_3_lut_rep_760 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n27083)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i134_3_lut_4_lut_3_lut_rep_760.init = 16'h6969;
    LUT4 i9542_3_lut_4_lut_4_lut (.A(index_i[0]), .B(n773), .C(index_i[4]), 
         .D(n27048), .Z(n12103)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B ((D)+!C)+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i9542_3_lut_4_lut_4_lut.init = 16'h5c0c;
    LUT4 mux_197_Mux_5_i761_3_lut_4_lut_3_lut_rep_761 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n27084)) /* synthesis lut_function=(A (B)+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_5_i761_3_lut_4_lut_3_lut_rep_761.init = 16'hd9d9;
    LUT4 mux_197_Mux_6_i572_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n572_adj_2784)) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_6_i572_3_lut_4_lut.init = 16'hccd9;
    PFUMX i23869 (.BLUT(n25652), .ALUT(n26922), .C0(index_i[4]), .Z(n25653));
    LUT4 mux_197_Mux_0_i142_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n142_adj_2781)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C))+!A !(B (C (D)+!C !(D))+!B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i142_3_lut_4_lut_4_lut.init = 16'ha569;
    LUT4 mux_196_Mux_0_i985_3_lut_4_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[1]), .Z(n985_adj_2644)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_0_i985_3_lut_4_lut_4_lut_3_lut.init = 16'h1919;
    LUT4 mux_197_Mux_3_i397_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n397_adj_2432)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)+!C !(D)))+!A !(B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_3_i397_3_lut_4_lut_4_lut.init = 16'ha95a;
    LUT4 i19017_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21454)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A !(B (D)+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19017_3_lut_3_lut_4_lut.init = 16'ha955;
    LUT4 i19551_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21988)) /* synthesis lut_function=(A (B (C (D))+!B !(C (D)))+!A !(B (D)+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19551_3_lut_4_lut_4_lut.init = 16'h9366;
    LUT4 mux_197_Mux_6_i347_3_lut_4_lut_3_lut_rep_774 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n27097)) /* synthesis lut_function=(!(A (B+!(C))+!A ((C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_6_i347_3_lut_4_lut_3_lut_rep_774.init = 16'h2424;
    L6MUX21 i23853 (.D0(n25636), .D1(n25633), .SD(index_q[5]), .Z(n25637));
    LUT4 i19332_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21769)) /* synthesis lut_function=(A (B (C)+!B (C (D)+!C !(D)))+!A !(B (C+!(D))+!B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19332_3_lut_4_lut_4_lut.init = 16'ha593;
    LUT4 mux_196_Mux_6_i204_3_lut_4_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[2]), 
         .C(index_i[1]), .Z(n204)) /* synthesis lut_function=(!(A (B)+!A !(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_6_i204_3_lut_4_lut_4_lut_3_lut.init = 16'h6767;
    LUT4 mux_196_Mux_9_i62_3_lut_4_lut_then_4_lut (.A(index_i[4]), .B(index_i[2]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n27237)) /* synthesis lut_function=(!(A (B (C+(D)))+!A (B+(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_9_i62_3_lut_4_lut_then_4_lut.init = 16'h222b;
    L6MUX21 i23031 (.D0(n24735), .D1(n26707), .SD(index_i[6]), .Z(n24736));
    LUT4 i19032_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21469)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C))+!A !(B ((D)+!C)+!B !(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19032_3_lut_4_lut_4_lut.init = 16'h925a;
    PFUMX i23851 (.BLUT(n25635), .ALUT(n25634), .C0(index_q[4]), .Z(n25636));
    LUT4 mux_197_Mux_0_i812_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n812_adj_2257)) /* synthesis lut_function=(A (B (C+(D))+!B !(C))+!A (B (D)+!B !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i812_3_lut_4_lut_4_lut_4_lut.init = 16'hcf92;
    LUT4 n715_bdd_3_lut_24179_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n26013)) /* synthesis lut_function=(A (B (C+(D))+!B ((D)+!C))+!A !(B (C+(D))+!B ((D)+!C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n715_bdd_3_lut_24179_4_lut.init = 16'haa96;
    LUT4 mux_197_Mux_6_i378_3_lut_4_lut_3_lut_rep_775 (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n27098)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)+!B !(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_6_i378_3_lut_4_lut_3_lut_rep_775.init = 16'h4949;
    LUT4 mux_196_Mux_9_i62_3_lut_4_lut_else_4_lut (.A(index_i[4]), .B(index_i[2]), 
         .C(index_i[1]), .D(index_i[0]), .Z(n27236)) /* synthesis lut_function=((B+(C (D)))+!A) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_9_i62_3_lut_4_lut_else_4_lut.init = 16'hfddd;
    LUT4 mux_197_Mux_3_i859_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n859_adj_2665)) /* synthesis lut_function=(!(A (B (D)+!B !(D))+!A (B (C+(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_3_i859_3_lut_3_lut_4_lut.init = 16'h339c;
    LUT4 i22408_3_lut (.A(n12121), .B(n892_adj_2663), .C(index_q[6]), 
         .Z(n22718)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i22408_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_5_i739_rep_776 (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .Z(n27099)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_5_i739_rep_776.init = 16'h6464;
    PFUMX i23029 (.BLUT(n24734), .ALUT(n24733), .C0(index_i[7]), .Z(n24735));
    LUT4 i21770_3_lut (.A(n491_adj_2439), .B(n506_adj_2750), .C(index_q[4]), 
         .Z(n21734)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i21770_3_lut.init = 16'hcaca;
    LUT4 i19342_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .D(index_q[3]), .Z(n21779)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C+(D)))+!A (B (C)+!B !(C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19342_3_lut_4_lut_4_lut.init = 16'hc95a;
    PFUMX i21010 (.BLUT(n526_adj_2347), .ALUT(n541_adj_2346), .C0(index_i[4]), 
          .Z(n23466));
    LUT4 mux_197_Mux_1_i93_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n93_adj_2552)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B !(C+(D)))+!A !(B (C (D)+!C !(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_1_i93_3_lut_4_lut_4_lut.init = 16'h955a;
    LUT4 mux_196_Mux_0_i348_3_lut_4_lut (.A(n26851), .B(index_i[2]), .C(index_i[3]), 
         .D(n29472), .Z(n348_adj_2776)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_0_i348_3_lut_4_lut.init = 16'h6f60;
    LUT4 mux_197_Mux_6_i459_rep_777 (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .Z(n27100)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_6_i459_rep_777.init = 16'h4d4d;
    LUT4 mux_196_Mux_4_i142_3_lut_4_lut_3_lut (.A(index_i[0]), .B(index_i[3]), 
         .C(index_i[2]), .Z(n142_adj_2395)) /* synthesis lut_function=(A (B (C))+!A !(B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_4_i142_3_lut_4_lut_3_lut.init = 16'h9595;
    LUT4 i11408_2_lut_rep_447_3_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[4]), .D(n27035), .Z(n26770)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11408_2_lut_rep_447_3_lut_4_lut.init = 16'hf8f0;
    PFUMX i23848 (.BLUT(n25632), .ALUT(n316_adj_2527), .C0(index_q[4]), 
          .Z(n25633));
    LUT4 i11233_2_lut_rep_762 (.A(index_q[0]), .B(index_q[1]), .Z(n27085)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11233_2_lut_rep_762.init = 16'h8888;
    LUT4 i11235_2_lut_2_lut_3_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[3]), 
         .Z(n13909)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11235_2_lut_2_lut_3_lut.init = 16'h0808;
    LUT4 i12330_2_lut_rep_430_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n26753)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i12330_2_lut_rep_430_3_lut_4_lut.init = 16'hf080;
    LUT4 i11037_2_lut_rep_538_3_lut (.A(index_q[0]), .B(index_q[1]), .C(index_q[2]), 
         .Z(n26861)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11037_2_lut_rep_538_3_lut.init = 16'hf8f8;
    LUT4 i20820_3_lut (.A(n23269), .B(n23270), .C(index_q[6]), .Z(n23276)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20820_3_lut.init = 16'hcaca;
    LUT4 i22743_2_lut_rep_494_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n26817)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A (C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i22743_2_lut_rep_494_3_lut_4_lut.init = 16'h0007;
    LUT4 mux_196_Mux_2_i349_3_lut_3_lut (.A(index_i[0]), .B(index_i[4]), 
         .C(n348_adj_2474), .Z(n349_adj_2570)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_2_i349_3_lut_3_lut.init = 16'hd1d1;
    LUT4 i20821_3_lut (.A(n25637), .B(n23272), .C(index_q[6]), .Z(n23277)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20821_3_lut.init = 16'hcaca;
    LUT4 i20508_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n22964)) /* synthesis lut_function=(A (B (C)+!B !(C (D)+!C !(D)))+!A !(B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i20508_3_lut_4_lut_4_lut_4_lut.init = 16'h83f0;
    LUT4 mux_197_Mux_7_i526_3_lut_3_lut_4_lut_4_lut_3_lut_4_lut (.A(index_q[0]), 
         .B(index_q[1]), .C(index_q[3]), .D(index_q[2]), .Z(n526_adj_2595)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(D))+!A !(D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_7_i526_3_lut_3_lut_4_lut_4_lut_3_lut_4_lut.init = 16'h887f;
    LUT4 i19530_3_lut_4_lut_4_lut (.A(index_i[0]), .B(n27025), .C(index_i[3]), 
         .D(n27046), .Z(n21967)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19530_3_lut_4_lut_4_lut.init = 16'hcfc5;
    LUT4 n172_bdd_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n25829)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)+!C !(D)))+!A (B (C+!(D))+!B (C (D)+!C !(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n172_bdd_3_lut_4_lut_4_lut_4_lut.init = 16'h0f38;
    LUT4 i20977_3_lut (.A(n23430), .B(n23431), .C(index_q[7]), .Z(n23433)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20977_3_lut.init = 16'hcaca;
    LUT4 mux_196_Mux_1_i890_4_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[3]), 
         .C(n26900), .D(index_i[4]), .Z(n890_adj_2712)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (D))+!A !((C+(D))+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_1_i890_4_lut_4_lut_4_lut_4_lut.init = 16'h55f3;
    LUT4 mux_197_Mux_8_i635_3_lut_4_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n635_adj_2342)) /* synthesis lut_function=(!(A (B (C (D))+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_8_i635_3_lut_4_lut_3_lut_4_lut.init = 16'h0ff8;
    LUT4 i20976_3_lut (.A(n23428), .B(n23429), .C(index_q[7]), .Z(n23432)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i20976_3_lut.init = 16'hcaca;
    LUT4 mux_197_Mux_7_i747_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), 
         .B(index_q[1]), .C(index_q[3]), .D(index_q[2]), .Z(n747_adj_2591)) /* synthesis lut_function=(A (B (C)+!B (C (D)+!C !(D)))+!A (B (C+!(D))+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_7_i747_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hf0c7;
    LUT4 mux_197_Mux_7_i620_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n620_adj_2783)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A !(B (C+!(D))+!B (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_7_i620_3_lut_4_lut_4_lut_4_lut.init = 16'h8c33;
    L6MUX21 i23829 (.D0(n25612), .D1(n25609), .SD(index_i[5]), .Z(n25613));
    LUT4 mux_196_Mux_2_i507_3_lut_3_lut (.A(index_i[0]), .B(index_i[4]), 
         .C(n491_adj_2764), .Z(n507_adj_2572)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B+(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_2_i507_3_lut_3_lut.init = 16'h7474;
    PFUMX i23827 (.BLUT(n25611), .ALUT(n25610), .C0(index_i[4]), .Z(n25612));
    PFUMX i20209 (.BLUT(n22663), .ALUT(n22664), .C0(index_i[9]), .Z(quarter_wave_sample_register_i_15__N_2126[9]));
    LUT4 mux_196_Mux_5_i573_3_lut_3_lut (.A(index_i[0]), .B(index_i[4]), 
         .C(n572_adj_2435), .Z(n573_adj_2450)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_5_i573_3_lut_3_lut.init = 16'hd1d1;
    LUT4 i11554_2_lut_rep_426_4_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[1]), 
         .C(index_i[2]), .D(index_i[3]), .Z(n26749)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A (B+((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11554_2_lut_rep_426_4_lut_4_lut_4_lut_4_lut.init = 16'h0038;
    LUT4 mux_197_Mux_6_i730_3_lut_rep_735_3_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .Z(n27058)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_6_i730_3_lut_rep_735_3_lut.init = 16'h3838;
    PFUMX i23824 (.BLUT(n25608), .ALUT(n26749), .C0(index_i[4]), .Z(n25609));
    LUT4 n77_bdd_3_lut_24283_3_lut_4_lut_4_lut_3_lut_4_lut (.A(index_q[0]), 
         .B(index_q[1]), .C(index_q[3]), .D(index_q[2]), .Z(n25966)) /* synthesis lut_function=(A (B (C)+!B !(D))+!A !(D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam n77_bdd_3_lut_24283_3_lut_4_lut_4_lut_3_lut_4_lut.init = 16'h80f7;
    LUT4 mux_197_Mux_8_i93_3_lut_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n93_adj_2594)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B (D))+!A (B ((D)+!C)+!B (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_8_i93_3_lut_3_lut_4_lut_4_lut.init = 16'h08f3;
    LUT4 i19723_3_lut_4_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n22160)) /* synthesis lut_function=(!(A (B (D)+!B !((D)+!C))+!A (B (C+(D))+!B !((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i19723_3_lut_4_lut_4_lut_4_lut_4_lut.init = 16'h338f;
    LUT4 i11501_3_lut_3_lut_3_lut (.A(index_i[0]), .B(index_i[2]), .C(index_i[1]), 
         .Z(n619)) /* synthesis lut_function=(!(A (C)+!A !(B+!(C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11501_3_lut_3_lut_3_lut.init = 16'h4f4f;
    L6MUX21 i23822 (.D0(n25606), .D1(n25604), .SD(index_i[4]), .Z(n25607));
    PFUMX i23820 (.BLUT(n26759), .ALUT(n25605), .C0(index_i[5]), .Z(n25606));
    LUT4 mux_197_Mux_4_i653_3_lut_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), 
         .B(index_q[1]), .C(index_q[3]), .D(index_q[2]), .Z(n653_adj_2464)) /* synthesis lut_function=(A (B (D)+!B !(D))+!A (B (C (D)+!C !(D))+!B !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_4_i653_3_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hc837;
    LUT4 i20598_3_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n23054)) /* synthesis lut_function=(A (B (C)+!B !(C (D)+!C !(D)))+!A !(B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i20598_3_lut_4_lut_4_lut_4_lut.init = 16'h83f0;
    PFUMX i23818 (.BLUT(n25603), .ALUT(n25602), .C0(index_i[5]), .Z(n25604));
    LUT4 mux_197_Mux_4_i1002_3_lut_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n1002_adj_2443)) /* synthesis lut_function=(A (B (C (D))+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_4_i1002_3_lut_3_lut_3_lut_4_lut.init = 16'hf007;
    LUT4 mux_196_Mux_2_i763_4_lut_4_lut (.A(index_i[0]), .B(n12095), .C(index_i[4]), 
         .D(n157_adj_2531), .Z(n763_adj_2579)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C+(D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_2_i763_4_lut_4_lut.init = 16'hdfd0;
    LUT4 n25411_bdd_3_lut (.A(n27118), .B(n444), .C(index_q[5]), .Z(n25412)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n25411_bdd_3_lut.init = 16'hcaca;
    LUT4 n17993_bdd_4_lut_then_4_lut (.A(index_q[3]), .B(index_q[4]), .C(index_q[1]), 
         .D(index_q[2]), .Z(n27144)) /* synthesis lut_function=(A (C (D)+!C !(D))+!A (B+(C (D)+!C !(D)))) */ ;
    defparam n17993_bdd_4_lut_then_4_lut.init = 16'hf44f;
    LUT4 i11765_3_lut_4_lut_4_lut_4_lut (.A(index_i[0]), .B(index_i[4]), 
         .C(n27035), .D(index_i[1]), .Z(n14440)) /* synthesis lut_function=(!(A (D)+!A !(B (C+!(D))+!B !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i11765_3_lut_4_lut_4_lut_4_lut.init = 16'h40ff;
    LUT4 mux_197_Mux_8_i526_3_lut_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n526_adj_2343)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)+!C !(D)))+!A (C (D)+!C !(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_8_i526_3_lut_3_lut_3_lut_4_lut.init = 16'h0f70;
    L6MUX21 i23801 (.D0(n25587), .D1(n25585), .SD(index_i[5]), .Z(n25588));
    PFUMX i23799 (.BLUT(n572_adj_2435), .ALUT(n25586), .C0(index_i[4]), 
          .Z(n25587));
    PFUMX i23797 (.BLUT(n25584), .ALUT(n25583), .C0(index_i[4]), .Z(n25585));
    L6MUX21 i23795 (.D0(n25581), .D1(n25579), .SD(index_i[4]), .Z(n25582));
    PFUMX i23793 (.BLUT(n25580), .ALUT(n26731), .C0(index_i[5]), .Z(n25581));
    PFUMX i20222 (.BLUT(n22674), .ALUT(n22675), .C0(index_i[8]), .Z(n22678));
    PFUMX i23791 (.BLUT(n25578), .ALUT(n25577), .C0(index_i[5]), .Z(n25579));
    PFUMX i20948 (.BLUT(n526_adj_2325), .ALUT(n541_adj_2324), .C0(index_q[4]), 
          .Z(n23404));
    LUT4 mux_197_Mux_2_i890_3_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n890_adj_2623)) /* synthesis lut_function=(A (B (D)+!B !((D)+!C))+!A !(B (C+(D))+!B !(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_2_i890_3_lut_4_lut_4_lut.init = 16'h9934;
    L6MUX21 i22854 (.D0(n24493), .D1(n26709), .SD(index_q[6]), .Z(n24494));
    PFUMX i22852 (.BLUT(n24492), .ALUT(n24491), .C0(index_q[5]), .Z(n24493));
    PFUMX i22847 (.BLUT(n21604), .ALUT(n24486), .C0(index_q[6]), .Z(n24487));
    L6MUX21 i23010 (.D0(n24711), .D1(n24709), .SD(index_q[6]), .Z(n24712));
    LUT4 i19593_3_lut_4_lut_4_lut (.A(index_i[0]), .B(n27029), .C(index_i[3]), 
         .D(n27048), .Z(n22030)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam i19593_3_lut_4_lut_4_lut.init = 16'hc5c0;
    PFUMX i23008 (.BLUT(n924_adj_2774), .ALUT(n24710), .C0(index_q[5]), 
          .Z(n24711));
    L6MUX21 i20223 (.D0(n22676), .D1(n22677), .SD(index_i[8]), .Z(n22679));
    LUT4 mux_196_Mux_2_i859_3_lut_4_lut_4_lut (.A(index_i[0]), .B(n26991), 
         .C(index_i[3]), .D(n27048), .Z(n859)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B ((D)+!C)+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(67[46:73])
    defparam mux_196_Mux_2_i859_3_lut_4_lut_4_lut.init = 16'h5c0c;
    LUT4 i11286_2_lut_rep_423_4_lut_4_lut_4_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[2]), .D(index_q[3]), .Z(n26746)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A (B+((D)+!C)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11286_2_lut_rep_423_4_lut_4_lut_4_lut_4_lut.init = 16'h0038;
    LUT4 i11850_3_lut_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n14525)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (D))+!A (D))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam i11850_3_lut_3_lut_3_lut_4_lut.init = 16'h00f7;
    PFUMX i19019 (.BLUT(n21454), .ALUT(n21455), .C0(index_q[4]), .Z(n21456));
    PFUMX i23703 (.BLUT(n25494), .ALUT(n25490), .C0(index_i[4]), .Z(n25495));
    PFUMX i23006 (.BLUT(n24708), .ALUT(n26840), .C0(index_q[5]), .Z(n24709));
    PFUMX i20512 (.BLUT(n22964), .ALUT(n22965), .C0(index_i[4]), .Z(n22968));
    PFUMX i23701 (.BLUT(n25491), .ALUT(n26975), .C0(index_i[3]), .Z(n25492));
    LUT4 mux_197_Mux_3_i1002_3_lut_3_lut_4_lut (.A(index_q[0]), .B(index_q[1]), 
         .C(index_q[3]), .D(index_q[2]), .Z(n19855)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (D))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_3_i1002_3_lut_3_lut_4_lut.init = 16'hf708;
    LUT4 mux_197_Mux_0_i716_3_lut (.A(n27073), .B(n27076), .C(index_q[3]), 
         .Z(n716)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/quarter_wave_sine_lookup.v(68[46:73])
    defparam mux_197_Mux_0_i716_3_lut.init = 16'hcaca;
    L6MUX21 i23677 (.D0(n25448), .D1(n25445), .SD(index_q[5]), .Z(n25449));
    PFUMX i20513 (.BLUT(n22966), .ALUT(n22967), .C0(index_i[4]), .Z(n22969));
    PFUMX i23675 (.BLUT(n25447), .ALUT(n25446), .C0(index_q[4]), .Z(n25448));
    
endmodule
//
// Verilog Description of module \nco(OW=12)_U1 
//

module \nco(OW=12)_U1  (increment, o_phase, GND_net, dac_clk_p_c, i_resetb_N_301) /* synthesis syn_module_defined=1 */ ;
    input [30:0]increment;
    output [11:0]o_phase;
    input GND_net;
    input dac_clk_p_c;
    input i_resetb_N_301;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(28[49:58])
    
    wire n17726;
    wire [31:0]n133;
    
    wire n17725, n17724, n17723, n17722, n17721, n17720;
    wire [31:0]n233;
    
    wire n17719, n17718, n17717, n17716, n17715, n17714, n17713, 
        n17712;
    
    CCU2D phase_register_547_add_4_32 (.A0(increment[30]), .B0(o_phase[10]), 
          .C0(GND_net), .D0(GND_net), .A1(o_phase[11]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n17726), .S0(n133[30]), .S1(n133[31]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547_add_4_32.INIT0 = 16'h5666;
    defparam phase_register_547_add_4_32.INIT1 = 16'hfaaa;
    defparam phase_register_547_add_4_32.INJECT1_0 = "NO";
    defparam phase_register_547_add_4_32.INJECT1_1 = "NO";
    CCU2D phase_register_547_add_4_30 (.A0(increment[28]), .B0(o_phase[8]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[29]), .B1(o_phase[9]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17725), .COUT(n17726), .S0(n133[28]), 
          .S1(n133[29]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547_add_4_30.INIT0 = 16'h5666;
    defparam phase_register_547_add_4_30.INIT1 = 16'h5666;
    defparam phase_register_547_add_4_30.INJECT1_0 = "NO";
    defparam phase_register_547_add_4_30.INJECT1_1 = "NO";
    CCU2D phase_register_547_add_4_28 (.A0(increment[26]), .B0(o_phase[6]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[27]), .B1(o_phase[7]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17724), .COUT(n17725), .S0(n133[26]), 
          .S1(n133[27]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547_add_4_28.INIT0 = 16'h5666;
    defparam phase_register_547_add_4_28.INIT1 = 16'h5666;
    defparam phase_register_547_add_4_28.INJECT1_0 = "NO";
    defparam phase_register_547_add_4_28.INJECT1_1 = "NO";
    CCU2D phase_register_547_add_4_26 (.A0(increment[24]), .B0(o_phase[4]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[25]), .B1(o_phase[5]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17723), .COUT(n17724), .S0(n133[24]), 
          .S1(n133[25]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547_add_4_26.INIT0 = 16'h5666;
    defparam phase_register_547_add_4_26.INIT1 = 16'h5666;
    defparam phase_register_547_add_4_26.INJECT1_0 = "NO";
    defparam phase_register_547_add_4_26.INJECT1_1 = "NO";
    CCU2D phase_register_547_add_4_24 (.A0(increment[22]), .B0(o_phase[2]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[23]), .B1(o_phase[3]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17722), .COUT(n17723), .S0(n133[22]), 
          .S1(n133[23]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547_add_4_24.INIT0 = 16'h5666;
    defparam phase_register_547_add_4_24.INIT1 = 16'h5666;
    defparam phase_register_547_add_4_24.INJECT1_0 = "NO";
    defparam phase_register_547_add_4_24.INJECT1_1 = "NO";
    CCU2D phase_register_547_add_4_22 (.A0(increment[20]), .B0(o_phase[0]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[21]), .B1(o_phase[1]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17721), .COUT(n17722), .S0(n133[20]), 
          .S1(n133[21]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547_add_4_22.INIT0 = 16'h5666;
    defparam phase_register_547_add_4_22.INIT1 = 16'h5666;
    defparam phase_register_547_add_4_22.INJECT1_0 = "NO";
    defparam phase_register_547_add_4_22.INJECT1_1 = "NO";
    CCU2D phase_register_547_add_4_20 (.A0(increment[18]), .B0(n233[18]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[19]), .B1(n233[19]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17720), .COUT(n17721), .S0(n133[18]), 
          .S1(n133[19]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547_add_4_20.INIT0 = 16'h5666;
    defparam phase_register_547_add_4_20.INIT1 = 16'h5666;
    defparam phase_register_547_add_4_20.INJECT1_0 = "NO";
    defparam phase_register_547_add_4_20.INJECT1_1 = "NO";
    CCU2D phase_register_547_add_4_18 (.A0(increment[16]), .B0(n233[16]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[17]), .B1(n233[17]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17719), .COUT(n17720), .S0(n133[16]), 
          .S1(n133[17]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547_add_4_18.INIT0 = 16'h5666;
    defparam phase_register_547_add_4_18.INIT1 = 16'h5666;
    defparam phase_register_547_add_4_18.INJECT1_0 = "NO";
    defparam phase_register_547_add_4_18.INJECT1_1 = "NO";
    CCU2D phase_register_547_add_4_16 (.A0(increment[14]), .B0(n233[14]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[15]), .B1(n233[15]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17718), .COUT(n17719), .S0(n133[14]), 
          .S1(n133[15]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547_add_4_16.INIT0 = 16'h5666;
    defparam phase_register_547_add_4_16.INIT1 = 16'h5666;
    defparam phase_register_547_add_4_16.INJECT1_0 = "NO";
    defparam phase_register_547_add_4_16.INJECT1_1 = "NO";
    CCU2D phase_register_547_add_4_14 (.A0(increment[12]), .B0(n233[12]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[13]), .B1(n233[13]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17717), .COUT(n17718), .S0(n133[12]), 
          .S1(n133[13]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547_add_4_14.INIT0 = 16'h5666;
    defparam phase_register_547_add_4_14.INIT1 = 16'h5666;
    defparam phase_register_547_add_4_14.INJECT1_0 = "NO";
    defparam phase_register_547_add_4_14.INJECT1_1 = "NO";
    CCU2D phase_register_547_add_4_12 (.A0(increment[10]), .B0(n233[10]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[11]), .B1(n233[11]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17716), .COUT(n17717), .S0(n133[10]), 
          .S1(n133[11]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547_add_4_12.INIT0 = 16'h5666;
    defparam phase_register_547_add_4_12.INIT1 = 16'h5666;
    defparam phase_register_547_add_4_12.INJECT1_0 = "NO";
    defparam phase_register_547_add_4_12.INJECT1_1 = "NO";
    CCU2D phase_register_547_add_4_10 (.A0(increment[8]), .B0(n233[8]), 
          .C0(GND_net), .D0(GND_net), .A1(increment[9]), .B1(n233[9]), 
          .C1(GND_net), .D1(GND_net), .CIN(n17715), .COUT(n17716), .S0(n133[8]), 
          .S1(n133[9]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547_add_4_10.INIT0 = 16'h5666;
    defparam phase_register_547_add_4_10.INIT1 = 16'h5666;
    defparam phase_register_547_add_4_10.INJECT1_0 = "NO";
    defparam phase_register_547_add_4_10.INJECT1_1 = "NO";
    CCU2D phase_register_547_add_4_8 (.A0(increment[6]), .B0(n233[6]), .C0(GND_net), 
          .D0(GND_net), .A1(increment[7]), .B1(n233[7]), .C1(GND_net), 
          .D1(GND_net), .CIN(n17714), .COUT(n17715), .S0(n133[6]), .S1(n133[7]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547_add_4_8.INIT0 = 16'h5666;
    defparam phase_register_547_add_4_8.INIT1 = 16'h5666;
    defparam phase_register_547_add_4_8.INJECT1_0 = "NO";
    defparam phase_register_547_add_4_8.INJECT1_1 = "NO";
    CCU2D phase_register_547_add_4_6 (.A0(increment[4]), .B0(n233[4]), .C0(GND_net), 
          .D0(GND_net), .A1(increment[5]), .B1(n233[5]), .C1(GND_net), 
          .D1(GND_net), .CIN(n17713), .COUT(n17714), .S0(n133[4]), .S1(n133[5]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547_add_4_6.INIT0 = 16'h5666;
    defparam phase_register_547_add_4_6.INIT1 = 16'h5666;
    defparam phase_register_547_add_4_6.INJECT1_0 = "NO";
    defparam phase_register_547_add_4_6.INJECT1_1 = "NO";
    CCU2D phase_register_547_add_4_4 (.A0(increment[2]), .B0(n233[2]), .C0(GND_net), 
          .D0(GND_net), .A1(increment[3]), .B1(n233[3]), .C1(GND_net), 
          .D1(GND_net), .CIN(n17712), .COUT(n17713), .S0(n133[2]), .S1(n133[3]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547_add_4_4.INIT0 = 16'h5666;
    defparam phase_register_547_add_4_4.INIT1 = 16'h5666;
    defparam phase_register_547_add_4_4.INJECT1_0 = "NO";
    defparam phase_register_547_add_4_4.INJECT1_1 = "NO";
    CCU2D phase_register_547_add_4_2 (.A0(increment[0]), .B0(n233[0]), .C0(GND_net), 
          .D0(GND_net), .A1(increment[1]), .B1(n233[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n17712), .S1(n133[1]));   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547_add_4_2.INIT0 = 16'h7000;
    defparam phase_register_547_add_4_2.INIT1 = 16'h5666;
    defparam phase_register_547_add_4_2.INJECT1_0 = "NO";
    defparam phase_register_547_add_4_2.INJECT1_1 = "NO";
    LUT4 i15482_2_lut (.A(increment[0]), .B(n233[0]), .Z(n133[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i15482_2_lut.init = 16'h6666;
    FD1S3DX phase_register_547__i31 (.D(n133[31]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(o_phase[11])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i31.GSR = "DISABLED";
    FD1S3DX phase_register_547__i30 (.D(n133[30]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(o_phase[10])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i30.GSR = "DISABLED";
    FD1S3DX phase_register_547__i29 (.D(n133[29]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(o_phase[9])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i29.GSR = "DISABLED";
    FD1S3DX phase_register_547__i28 (.D(n133[28]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(o_phase[8])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i28.GSR = "DISABLED";
    FD1S3DX phase_register_547__i27 (.D(n133[27]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(o_phase[7])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i27.GSR = "DISABLED";
    FD1S3DX phase_register_547__i26 (.D(n133[26]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(o_phase[6])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i26.GSR = "DISABLED";
    FD1S3DX phase_register_547__i25 (.D(n133[25]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(o_phase[5])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i25.GSR = "DISABLED";
    FD1S3DX phase_register_547__i24 (.D(n133[24]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(o_phase[4])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i24.GSR = "DISABLED";
    FD1S3DX phase_register_547__i23 (.D(n133[23]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(o_phase[3])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i23.GSR = "DISABLED";
    FD1S3DX phase_register_547__i22 (.D(n133[22]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(o_phase[2])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i22.GSR = "DISABLED";
    FD1S3DX phase_register_547__i21 (.D(n133[21]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(o_phase[1])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i21.GSR = "DISABLED";
    FD1S3DX phase_register_547__i20 (.D(n133[20]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(o_phase[0])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i20.GSR = "DISABLED";
    FD1S3DX phase_register_547__i19 (.D(n133[19]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(n233[19])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i19.GSR = "DISABLED";
    FD1S3DX phase_register_547__i18 (.D(n133[18]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(n233[18])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i18.GSR = "DISABLED";
    FD1S3DX phase_register_547__i17 (.D(n133[17]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(n233[17])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i17.GSR = "DISABLED";
    FD1S3DX phase_register_547__i16 (.D(n133[16]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(n233[16])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i16.GSR = "DISABLED";
    FD1S3DX phase_register_547__i15 (.D(n133[15]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(n233[15])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i15.GSR = "DISABLED";
    FD1S3DX phase_register_547__i14 (.D(n133[14]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(n233[14])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i14.GSR = "DISABLED";
    FD1S3DX phase_register_547__i13 (.D(n133[13]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(n233[13])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i13.GSR = "DISABLED";
    FD1S3DX phase_register_547__i12 (.D(n133[12]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(n233[12])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i12.GSR = "DISABLED";
    FD1S3DX phase_register_547__i11 (.D(n133[11]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(n233[11])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i11.GSR = "DISABLED";
    FD1S3DX phase_register_547__i10 (.D(n133[10]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(n233[10])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i10.GSR = "DISABLED";
    FD1S3DX phase_register_547__i9 (.D(n133[9]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(n233[9])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i9.GSR = "DISABLED";
    FD1S3DX phase_register_547__i8 (.D(n133[8]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(n233[8])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i8.GSR = "DISABLED";
    FD1S3DX phase_register_547__i7 (.D(n133[7]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(n233[7])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i7.GSR = "DISABLED";
    FD1S3DX phase_register_547__i6 (.D(n133[6]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(n233[6])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i6.GSR = "DISABLED";
    FD1S3DX phase_register_547__i5 (.D(n133[5]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(n233[5])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i5.GSR = "DISABLED";
    FD1S3DX phase_register_547__i4 (.D(n133[4]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(n233[4])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i4.GSR = "DISABLED";
    FD1S3DX phase_register_547__i3 (.D(n133[3]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(n233[3])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i3.GSR = "DISABLED";
    FD1S3DX phase_register_547__i2 (.D(n133[2]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(n233[2])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i2.GSR = "DISABLED";
    FD1S3DX phase_register_547__i1 (.D(n133[1]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(n233[1])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i1.GSR = "DISABLED";
    FD1S3DX phase_register_547__i0 (.D(n133[0]), .CK(dac_clk_p_c), .CD(i_resetb_N_301), 
            .Q(n233[0])) /* synthesis syn_use_carry_chain=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/nco.v(25[22:50])
    defparam phase_register_547__i0.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module TSALL
// module not written out since it is a black-box. 
//

//
// Verilog Description of module efb_inst
//

module efb_inst (dac_clk_p_c, i_resetb_N_301, wb_cyc, wb_lo_data_7__N_96, 
            wb_we, \wb_addr[7] , \wb_addr[6] , \wb_addr[5] , \wb_addr[4] , 
            \wb_addr[3] , \wb_addr[2] , \wb_addr[1] , \wb_addr[0] , 
            \wb_odata[7] , \wb_odata[6] , \wb_odata[5] , \wb_odata[4] , 
            \wb_odata[3] , \wb_odata[2] , \wb_odata[1] , \wb_odata[0] , 
            pll_data_o, pll_ack, wb_lo_data, wb_lo_ack, pll_clk, pll_rst, 
            pll_stb, pll_we, pll_addr, pll_data_i, GND_net, VCC_net) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;
    input dac_clk_p_c;
    input i_resetb_N_301;
    input wb_cyc;
    input wb_lo_data_7__N_96;
    input wb_we;
    input \wb_addr[7] ;
    input \wb_addr[6] ;
    input \wb_addr[5] ;
    input \wb_addr[4] ;
    input \wb_addr[3] ;
    input \wb_addr[2] ;
    input \wb_addr[1] ;
    input \wb_addr[0] ;
    input \wb_odata[7] ;
    input \wb_odata[6] ;
    input \wb_odata[5] ;
    input \wb_odata[4] ;
    input \wb_odata[3] ;
    input \wb_odata[2] ;
    input \wb_odata[1] ;
    input \wb_odata[0] ;
    input [7:0]pll_data_o;
    input pll_ack;
    output [7:0]wb_lo_data;
    output wb_lo_ack;
    output pll_clk;
    output pll_rst;
    output pll_stb;
    output pll_we;
    output [4:0]pll_addr;
    output [7:0]pll_data_i;
    input GND_net;
    input VCC_net;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(28[49:58])
    
    EFB EFBInst_0 (.WBCLKI(dac_clk_p_c), .WBRSTI(i_resetb_N_301), .WBCYCI(wb_cyc), 
        .WBSTBI(wb_lo_data_7__N_96), .WBWEI(wb_we), .WBADRI0(\wb_addr[0] ), 
        .WBADRI1(\wb_addr[1] ), .WBADRI2(\wb_addr[2] ), .WBADRI3(\wb_addr[3] ), 
        .WBADRI4(\wb_addr[4] ), .WBADRI5(\wb_addr[5] ), .WBADRI6(\wb_addr[6] ), 
        .WBADRI7(\wb_addr[7] ), .WBDATI0(\wb_odata[0] ), .WBDATI1(\wb_odata[1] ), 
        .WBDATI2(\wb_odata[2] ), .WBDATI3(\wb_odata[3] ), .WBDATI4(\wb_odata[4] ), 
        .WBDATI5(\wb_odata[5] ), .WBDATI6(\wb_odata[6] ), .WBDATI7(\wb_odata[7] ), 
        .I2C1SCLI(GND_net), .I2C1SDAI(GND_net), .I2C2SCLI(GND_net), .I2C2SDAI(GND_net), 
        .SPISCKI(GND_net), .SPIMISOI(GND_net), .SPIMOSII(GND_net), .SPISCSN(GND_net), 
        .TCCLKI(GND_net), .TCRSTN(GND_net), .TCIC(GND_net), .UFMSN(VCC_net), 
        .PLL0DATI0(pll_data_o[0]), .PLL0DATI1(pll_data_o[1]), .PLL0DATI2(pll_data_o[2]), 
        .PLL0DATI3(pll_data_o[3]), .PLL0DATI4(pll_data_o[4]), .PLL0DATI5(pll_data_o[5]), 
        .PLL0DATI6(pll_data_o[6]), .PLL0DATI7(pll_data_o[7]), .PLL0ACKI(pll_ack), 
        .PLL1DATI0(GND_net), .PLL1DATI1(GND_net), .PLL1DATI2(GND_net), 
        .PLL1DATI3(GND_net), .PLL1DATI4(GND_net), .PLL1DATI5(GND_net), 
        .PLL1DATI6(GND_net), .PLL1DATI7(GND_net), .PLL1ACKI(GND_net), 
        .WBDATO0(wb_lo_data[0]), .WBDATO1(wb_lo_data[1]), .WBDATO2(wb_lo_data[2]), 
        .WBDATO3(wb_lo_data[3]), .WBDATO4(wb_lo_data[4]), .WBDATO5(wb_lo_data[5]), 
        .WBDATO6(wb_lo_data[6]), .WBDATO7(wb_lo_data[7]), .WBACKO(wb_lo_ack), 
        .PLLCLKO(pll_clk), .PLLRSTO(pll_rst), .PLL0STBO(pll_stb), .PLLWEO(pll_we), 
        .PLLADRO0(pll_addr[0]), .PLLADRO1(pll_addr[1]), .PLLADRO2(pll_addr[2]), 
        .PLLADRO3(pll_addr[3]), .PLLADRO4(pll_addr[4]), .PLLDATO0(pll_data_i[0]), 
        .PLLDATO1(pll_data_i[1]), .PLLDATO2(pll_data_i[2]), .PLLDATO3(pll_data_i[3]), 
        .PLLDATO4(pll_data_i[4]), .PLLDATO5(pll_data_i[5]), .PLLDATO6(pll_data_i[6]), 
        .PLLDATO7(pll_data_i[7])) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=8, LSE_LCOL=10, LSE_RCOL=3, LSE_LLINE=180, LSE_RLINE=192 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(180[10] 192[3])
    defparam EFBInst_0.EFB_I2C1 = "DISABLED";
    defparam EFBInst_0.EFB_I2C2 = "DISABLED";
    defparam EFBInst_0.EFB_SPI = "DISABLED";
    defparam EFBInst_0.EFB_TC = "DISABLED";
    defparam EFBInst_0.EFB_TC_PORTMODE = "WB";
    defparam EFBInst_0.EFB_UFM = "DISABLED";
    defparam EFBInst_0.EFB_WB_CLK_FREQ = "50.0";
    defparam EFBInst_0.DEV_DENSITY = "6900L";
    defparam EFBInst_0.UFM_INIT_PAGES = 0;
    defparam EFBInst_0.UFM_INIT_START_PAGE = 0;
    defparam EFBInst_0.UFM_INIT_ALL_ZEROS = "ENABLED";
    defparam EFBInst_0.UFM_INIT_FILE_NAME = "NONE";
    defparam EFBInst_0.UFM_INIT_FILE_FORMAT = "HEX";
    defparam EFBInst_0.I2C1_ADDRESSING = "7BIT";
    defparam EFBInst_0.I2C2_ADDRESSING = "7BIT";
    defparam EFBInst_0.I2C1_SLAVE_ADDR = "0b1000001";
    defparam EFBInst_0.I2C2_SLAVE_ADDR = "0b1000010";
    defparam EFBInst_0.I2C1_BUS_PERF = "100kHz";
    defparam EFBInst_0.I2C2_BUS_PERF = "100kHz";
    defparam EFBInst_0.I2C1_CLK_DIVIDER = 1;
    defparam EFBInst_0.I2C2_CLK_DIVIDER = 1;
    defparam EFBInst_0.I2C1_GEN_CALL = "DISABLED";
    defparam EFBInst_0.I2C2_GEN_CALL = "DISABLED";
    defparam EFBInst_0.I2C1_WAKEUP = "DISABLED";
    defparam EFBInst_0.I2C2_WAKEUP = "DISABLED";
    defparam EFBInst_0.SPI_MODE = "MASTER";
    defparam EFBInst_0.SPI_CLK_DIVIDER = 1;
    defparam EFBInst_0.SPI_LSB_FIRST = "DISABLED";
    defparam EFBInst_0.SPI_CLK_INV = "DISABLED";
    defparam EFBInst_0.SPI_PHASE_ADJ = "DISABLED";
    defparam EFBInst_0.SPI_SLAVE_HANDSHAKE = "DISABLED";
    defparam EFBInst_0.SPI_INTR_TXRDY = "DISABLED";
    defparam EFBInst_0.SPI_INTR_RXRDY = "DISABLED";
    defparam EFBInst_0.SPI_INTR_TXOVR = "DISABLED";
    defparam EFBInst_0.SPI_INTR_RXOVR = "DISABLED";
    defparam EFBInst_0.SPI_WAKEUP = "DISABLED";
    defparam EFBInst_0.TC_MODE = "CTCM";
    defparam EFBInst_0.TC_SCLK_SEL = "PCLOCK";
    defparam EFBInst_0.TC_CCLK_SEL = 1;
    defparam EFBInst_0.GSR = "ENABLED";
    defparam EFBInst_0.TC_TOP_SET = 65535;
    defparam EFBInst_0.TC_OCR_SET = 32767;
    defparam EFBInst_0.TC_OC_MODE = "TOGGLE";
    defparam EFBInst_0.TC_RESETN = "ENABLED";
    defparam EFBInst_0.TC_TOP_SEL = "OFF";
    defparam EFBInst_0.TC_OV_INT = "OFF";
    defparam EFBInst_0.TC_OCR_INT = "OFF";
    defparam EFBInst_0.TC_ICR_INT = "OFF";
    defparam EFBInst_0.TC_OVERFLOW = "DISABLED";
    defparam EFBInst_0.TC_ICAPTURE = "DISABLED";
    
endmodule
//
// Verilog Description of module clock_phase_shifter
//

module clock_phase_shifter (q_clk_p_c, i_clk_2f_N_2249, q_clk_n_c, i_clk_p_c, 
            lo_pll_out, i_clk_n_c) /* synthesis syn_module_defined=1 */ ;
    output q_clk_p_c;
    input i_clk_2f_N_2249;
    input q_clk_n_c;
    output i_clk_p_c;
    input lo_pll_out;
    input i_clk_n_c;
    
    wire i_clk_2f_N_2249 /* synthesis is_inv_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/clock_phase_shifter.v(11[21:28])
    wire lo_pll_out /* synthesis is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(160[6:16])
    
    FD1S3AX o_clk_q_10 (.D(q_clk_n_c), .CK(i_clk_2f_N_2249), .Q(q_clk_p_c)) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=21, LSE_RCOL=2, LSE_LLINE=161, LSE_RLINE=165 */ ;   // d:/documents/git_local/fm_modulator/rtl/clock_phase_shifter.v(17[8] 19[4])
    defparam o_clk_q_10.GSR = "DISABLED";
    FD1S3AX o_clk_i_9 (.D(i_clk_n_c), .CK(lo_pll_out), .Q(i_clk_p_c)) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=21, LSE_RCOL=2, LSE_LLINE=161, LSE_RLINE=165 */ ;   // d:/documents/git_local/fm_modulator/rtl/clock_phase_shifter.v(13[8] 15[4])
    defparam o_clk_i_9.GSR = "DISABLED";
    
endmodule
//
// Verilog Description of module sys_clk
//

module sys_clk (i_ref_clk_c, dac_clk_p_c, GND_net) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;
    input i_ref_clk_c;
    output dac_clk_p_c;
    input GND_net;
    
    wire i_ref_clk_c /* synthesis is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(22[12:21])
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(28[49:58])
    
    wire CLKFB_t;
    
    EHXPLLJ PLLInst_0 (.CLKI(i_ref_clk_c), .CLKFB(CLKFB_t), .PHASESEL0(GND_net), 
            .PHASESEL1(GND_net), .PHASEDIR(GND_net), .PHASESTEP(GND_net), 
            .LOADREG(GND_net), .STDBY(GND_net), .PLLWAKESYNC(GND_net), 
            .RST(GND_net), .RESETC(GND_net), .RESETD(GND_net), .RESETM(GND_net), 
            .ENCLKOP(GND_net), .ENCLKOS(GND_net), .ENCLKOS2(GND_net), 
            .ENCLKOS3(GND_net), .PLLCLK(GND_net), .PLLRST(GND_net), .PLLSTB(GND_net), 
            .PLLWE(GND_net), .PLLDATI0(GND_net), .PLLDATI1(GND_net), .PLLDATI2(GND_net), 
            .PLLDATI3(GND_net), .PLLDATI4(GND_net), .PLLDATI5(GND_net), 
            .PLLDATI6(GND_net), .PLLDATI7(GND_net), .PLLADDR0(GND_net), 
            .PLLADDR1(GND_net), .PLLADDR2(GND_net), .PLLADDR3(GND_net), 
            .PLLADDR4(GND_net), .CLKOP(dac_clk_p_c), .CLKINTFB(CLKFB_t)) /* synthesis FREQUENCY_PIN_CLKOP="96.000000", FREQUENCY_PIN_CLKI="12.000000", ICP_CURRENT="7", LPF_RESISTOR="8", syn_instantiated=1, LSE_LINE_FILE_ID=8, LSE_LCOL=10, LSE_RCOL=54, LSE_LLINE=37, LSE_RLINE=37 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(37[10:54])
    defparam PLLInst_0.CLKI_DIV = 1;
    defparam PLLInst_0.CLKFB_DIV = 8;
    defparam PLLInst_0.CLKOP_DIV = 5;
    defparam PLLInst_0.CLKOS_DIV = 1;
    defparam PLLInst_0.CLKOS2_DIV = 1;
    defparam PLLInst_0.CLKOS3_DIV = 1;
    defparam PLLInst_0.CLKOP_ENABLE = "ENABLED";
    defparam PLLInst_0.CLKOS_ENABLE = "DISABLED";
    defparam PLLInst_0.CLKOS2_ENABLE = "DISABLED";
    defparam PLLInst_0.CLKOS3_ENABLE = "DISABLED";
    defparam PLLInst_0.VCO_BYPASS_A0 = "DISABLED";
    defparam PLLInst_0.VCO_BYPASS_B0 = "DISABLED";
    defparam PLLInst_0.VCO_BYPASS_C0 = "DISABLED";
    defparam PLLInst_0.VCO_BYPASS_D0 = "DISABLED";
    defparam PLLInst_0.CLKOP_CPHASE = 4;
    defparam PLLInst_0.CLKOS_CPHASE = 0;
    defparam PLLInst_0.CLKOS2_CPHASE = 0;
    defparam PLLInst_0.CLKOS3_CPHASE = 0;
    defparam PLLInst_0.CLKOP_FPHASE = 0;
    defparam PLLInst_0.CLKOS_FPHASE = 0;
    defparam PLLInst_0.CLKOS2_FPHASE = 0;
    defparam PLLInst_0.CLKOS3_FPHASE = 0;
    defparam PLLInst_0.FEEDBK_PATH = "INT_DIVA";
    defparam PLLInst_0.FRACN_ENABLE = "DISABLED";
    defparam PLLInst_0.FRACN_DIV = 0;
    defparam PLLInst_0.CLKOP_TRIM_POL = "RISING";
    defparam PLLInst_0.CLKOP_TRIM_DELAY = 0;
    defparam PLLInst_0.CLKOS_TRIM_POL = "FALLING";
    defparam PLLInst_0.CLKOS_TRIM_DELAY = 0;
    defparam PLLInst_0.PLL_USE_WB = "DISABLED";
    defparam PLLInst_0.PREDIVIDER_MUXA1 = 0;
    defparam PLLInst_0.PREDIVIDER_MUXB1 = 0;
    defparam PLLInst_0.PREDIVIDER_MUXC1 = 0;
    defparam PLLInst_0.PREDIVIDER_MUXD1 = 0;
    defparam PLLInst_0.OUTDIVIDER_MUXA2 = "DIVA";
    defparam PLLInst_0.OUTDIVIDER_MUXB2 = "DIVB";
    defparam PLLInst_0.OUTDIVIDER_MUXC2 = "DIVC";
    defparam PLLInst_0.OUTDIVIDER_MUXD2 = "DIVD";
    defparam PLLInst_0.PLL_LOCK_MODE = 0;
    defparam PLLInst_0.STDBY_ENABLE = "DISABLED";
    defparam PLLInst_0.DPHASE_SOURCE = "DISABLED";
    defparam PLLInst_0.PLLRST_ENA = "DISABLED";
    defparam PLLInst_0.MRST_ENA = "DISABLED";
    defparam PLLInst_0.DCRST_ENA = "DISABLED";
    defparam PLLInst_0.DDRST_ENA = "DISABLED";
    defparam PLLInst_0.INTFB_WAKE = "DISABLED";
    
endmodule
//
// Verilog Description of module dynamic_pll
//

module dynamic_pll (i_clk_2f_N_2249, lo_pll_out, i_ref_clk_c, pll_clk, 
            pll_rst, pll_stb, pll_we, pll_data_i, pll_addr, pll_data_o, 
            pll_ack, GND_net) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;
    output i_clk_2f_N_2249;
    output lo_pll_out;
    input i_ref_clk_c;
    input pll_clk;
    input pll_rst;
    input pll_stb;
    input pll_we;
    input [7:0]pll_data_i;
    input [4:0]pll_addr;
    output [7:0]pll_data_o;
    output pll_ack;
    input GND_net;
    
    wire i_clk_2f_N_2249 /* synthesis is_inv_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/clock_phase_shifter.v(11[21:28])
    wire lo_pll_out /* synthesis is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(160[6:16])
    wire i_ref_clk_c /* synthesis is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(22[12:21])
    
    INV i26492 (.A(lo_pll_out), .Z(i_clk_2f_N_2249));
    EHXPLLJ PLLInst_0 (.CLKI(i_ref_clk_c), .CLKFB(lo_pll_out), .PHASESEL0(GND_net), 
            .PHASESEL1(GND_net), .PHASEDIR(GND_net), .PHASESTEP(GND_net), 
            .LOADREG(GND_net), .STDBY(GND_net), .PLLWAKESYNC(GND_net), 
            .RST(GND_net), .RESETC(GND_net), .RESETD(GND_net), .RESETM(GND_net), 
            .ENCLKOP(GND_net), .ENCLKOS(GND_net), .ENCLKOS2(GND_net), 
            .ENCLKOS3(GND_net), .PLLCLK(pll_clk), .PLLRST(pll_rst), .PLLSTB(pll_stb), 
            .PLLWE(pll_we), .PLLDATI0(pll_data_i[0]), .PLLDATI1(pll_data_i[1]), 
            .PLLDATI2(pll_data_i[2]), .PLLDATI3(pll_data_i[3]), .PLLDATI4(pll_data_i[4]), 
            .PLLDATI5(pll_data_i[5]), .PLLDATI6(pll_data_i[6]), .PLLDATI7(pll_data_i[7]), 
            .PLLADDR0(pll_addr[0]), .PLLADDR1(pll_addr[1]), .PLLADDR2(pll_addr[2]), 
            .PLLADDR3(pll_addr[3]), .PLLADDR4(pll_addr[4]), .CLKOP(lo_pll_out), 
            .PLLDATO0(pll_data_o[0]), .PLLDATO1(pll_data_o[1]), .PLLDATO2(pll_data_o[2]), 
            .PLLDATO3(pll_data_o[3]), .PLLDATO4(pll_data_o[4]), .PLLDATO5(pll_data_o[5]), 
            .PLLDATO6(pll_data_o[6]), .PLLDATO7(pll_data_o[7]), .PLLACK(pll_ack)) /* synthesis FREQUENCY_PIN_CLKOP="420.000000", FREQUENCY_PIN_CLKI="12.000000", ICP_CURRENT="6", LPF_RESISTOR="8", syn_instantiated=1, LSE_LINE_FILE_ID=8, LSE_LCOL=13, LSE_RCOL=5, LSE_LLINE=167, LSE_RLINE=178 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(167[13] 178[5])
    defparam PLLInst_0.CLKI_DIV = 1;
    defparam PLLInst_0.CLKFB_DIV = 35;
    defparam PLLInst_0.CLKOP_DIV = 1;
    defparam PLLInst_0.CLKOS_DIV = 1;
    defparam PLLInst_0.CLKOS2_DIV = 1;
    defparam PLLInst_0.CLKOS3_DIV = 1;
    defparam PLLInst_0.CLKOP_ENABLE = "ENABLED";
    defparam PLLInst_0.CLKOS_ENABLE = "DISABLED";
    defparam PLLInst_0.CLKOS2_ENABLE = "DISABLED";
    defparam PLLInst_0.CLKOS3_ENABLE = "DISABLED";
    defparam PLLInst_0.VCO_BYPASS_A0 = "DISABLED";
    defparam PLLInst_0.VCO_BYPASS_B0 = "DISABLED";
    defparam PLLInst_0.VCO_BYPASS_C0 = "DISABLED";
    defparam PLLInst_0.VCO_BYPASS_D0 = "DISABLED";
    defparam PLLInst_0.CLKOP_CPHASE = 0;
    defparam PLLInst_0.CLKOS_CPHASE = 0;
    defparam PLLInst_0.CLKOS2_CPHASE = 0;
    defparam PLLInst_0.CLKOS3_CPHASE = 0;
    defparam PLLInst_0.CLKOP_FPHASE = 0;
    defparam PLLInst_0.CLKOS_FPHASE = 0;
    defparam PLLInst_0.CLKOS2_FPHASE = 0;
    defparam PLLInst_0.CLKOS3_FPHASE = 0;
    defparam PLLInst_0.FEEDBK_PATH = "CLKOP";
    defparam PLLInst_0.FRACN_ENABLE = "ENABLED";
    defparam PLLInst_0.FRACN_DIV = 2731;
    defparam PLLInst_0.CLKOP_TRIM_POL = "RISING";
    defparam PLLInst_0.CLKOP_TRIM_DELAY = 0;
    defparam PLLInst_0.CLKOS_TRIM_POL = "FALLING";
    defparam PLLInst_0.CLKOS_TRIM_DELAY = 0;
    defparam PLLInst_0.PLL_USE_WB = "ENABLED";
    defparam PLLInst_0.PREDIVIDER_MUXA1 = 0;
    defparam PLLInst_0.PREDIVIDER_MUXB1 = 0;
    defparam PLLInst_0.PREDIVIDER_MUXC1 = 0;
    defparam PLLInst_0.PREDIVIDER_MUXD1 = 0;
    defparam PLLInst_0.OUTDIVIDER_MUXA2 = "DIVA";
    defparam PLLInst_0.OUTDIVIDER_MUXB2 = "DIVB";
    defparam PLLInst_0.OUTDIVIDER_MUXC2 = "DIVC";
    defparam PLLInst_0.OUTDIVIDER_MUXD2 = "DIVD";
    defparam PLLInst_0.PLL_LOCK_MODE = 0;
    defparam PLLInst_0.STDBY_ENABLE = "DISABLED";
    defparam PLLInst_0.DPHASE_SOURCE = "DISABLED";
    defparam PLLInst_0.PLLRST_ENA = "DISABLED";
    defparam PLLInst_0.MRST_ENA = "DISABLED";
    defparam PLLInst_0.DCRST_ENA = "DISABLED";
    defparam PLLInst_0.DDRST_ENA = "DISABLED";
    defparam PLLInst_0.INTFB_WAKE = "DISABLED";
    
endmodule
//
// Verilog Description of module \txuartlite(TIMING_BITS=24,CLOCKS_PER_BAUD=10000) 
//

module \txuartlite(TIMING_BITS=24,CLOCKS_PER_BAUD=10000)  (dac_clk_p_c, dac_clk_p_c_enable_322, 
            \lcl_data_7__N_511[0] , zero_baud_counter, o_wbu_uart_tx_c, 
            n26910, GND_net, \state[0] , \lcl_data[7] , n29502, \lcl_data[6] , 
            \lcl_data_7__N_511[6] , \lcl_data[5] , \lcl_data_7__N_511[5] , 
            \lcl_data[4] , \lcl_data_7__N_511[4] , \lcl_data[3] , \lcl_data_7__N_511[3] , 
            \lcl_data[2] , \lcl_data_7__N_511[2] , \lcl_data[1] , \lcl_data_7__N_511[1] , 
            o_busy_N_536, tx_busy, n17844) /* synthesis syn_module_defined=1 */ ;
    input dac_clk_p_c;
    input dac_clk_p_c_enable_322;
    input \lcl_data_7__N_511[0] ;
    output zero_baud_counter;
    output o_wbu_uart_tx_c;
    input n26910;
    input GND_net;
    output \state[0] ;
    output \lcl_data[7] ;
    input n29502;
    output \lcl_data[6] ;
    input \lcl_data_7__N_511[6] ;
    output \lcl_data[5] ;
    input \lcl_data_7__N_511[5] ;
    output \lcl_data[4] ;
    input \lcl_data_7__N_511[4] ;
    output \lcl_data[3] ;
    input \lcl_data_7__N_511[3] ;
    output \lcl_data[2] ;
    input \lcl_data_7__N_511[2] ;
    output \lcl_data[1] ;
    input \lcl_data_7__N_511[1] ;
    output o_busy_N_536;
    output tx_busy;
    input n17844;
    
    wire dac_clk_p_c /* synthesis SET_AS_NETWORK=dac_clk_p_c, is_clock=1 */ ;   // d:/documents/git_local/fm_modulator/rtl/top.v(28[49:58])
    wire [7:0]lcl_data;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(84[12:20])
    
    wire zero_baud_counter_N_525;
    wire [23:0]baud_counter;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(82[17:29])
    wire [23:0]baud_counter_23__N_483;
    
    wire n17655;
    wire [23:0]n108;
    
    wire n17654, n17653, n17652, n17651, n17650, n17649, n17648, 
        n17647, n17646, n17645, n17644;
    wire [3:0]state;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(83[12:17])
    
    wire n26907, n11532, n27154, n27153, n27157, n27156, n20311, 
        n26789, zero_baud_counter_N_528, n20839, n20847, n20845, n20837;
    wire [23:0]n133;
    
    wire n20823, n20833, n20835, n20825, n8997;
    wire [3:0]n27;
    
    wire n27158, n27155;
    
    FD1P3AY lcl_data_i0 (.D(\lcl_data_7__N_511[0] ), .SP(dac_clk_p_c_enable_322), 
            .CK(dac_clk_p_c), .Q(lcl_data[0])) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=62, LSE_RLINE=62 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(139[9] 143[40])
    defparam lcl_data_i0.GSR = "DISABLED";
    FD1S3AY zero_baud_counter_49 (.D(zero_baud_counter_N_525), .CK(dac_clk_p_c), 
            .Q(zero_baud_counter)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=62, LSE_RLINE=62 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam zero_baud_counter_49.GSR = "DISABLED";
    FD1S3AX baud_counter_i0 (.D(baud_counter_23__N_483[0]), .CK(dac_clk_p_c), 
            .Q(baud_counter[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=62, LSE_RLINE=62 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i0.GSR = "DISABLED";
    FD1P3IX o_uart_tx_48 (.D(lcl_data[0]), .SP(dac_clk_p_c_enable_322), 
            .CD(n26910), .CK(dac_clk_p_c), .Q(o_wbu_uart_tx_c)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=62, LSE_RLINE=62 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(154[9] 158[29])
    defparam o_uart_tx_48.GSR = "DISABLED";
    CCU2D sub_36_add_2_25 (.A0(baud_counter[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n17655), .S0(n108[23]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_25.INIT0 = 16'h5555;
    defparam sub_36_add_2_25.INIT1 = 16'h0000;
    defparam sub_36_add_2_25.INJECT1_0 = "NO";
    defparam sub_36_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_36_add_2_23 (.A0(baud_counter[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17654), .COUT(n17655), .S0(n108[21]), 
          .S1(n108[22]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_23.INIT0 = 16'h5555;
    defparam sub_36_add_2_23.INIT1 = 16'h5555;
    defparam sub_36_add_2_23.INJECT1_0 = "NO";
    defparam sub_36_add_2_23.INJECT1_1 = "NO";
    CCU2D sub_36_add_2_21 (.A0(baud_counter[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17653), .COUT(n17654), .S0(n108[19]), 
          .S1(n108[20]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_21.INIT0 = 16'h5555;
    defparam sub_36_add_2_21.INIT1 = 16'h5555;
    defparam sub_36_add_2_21.INJECT1_0 = "NO";
    defparam sub_36_add_2_21.INJECT1_1 = "NO";
    CCU2D sub_36_add_2_19 (.A0(baud_counter[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17652), .COUT(n17653), .S0(n108[17]), 
          .S1(n108[18]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_19.INIT0 = 16'h5555;
    defparam sub_36_add_2_19.INIT1 = 16'h5555;
    defparam sub_36_add_2_19.INJECT1_0 = "NO";
    defparam sub_36_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_36_add_2_17 (.A0(baud_counter[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17651), .COUT(n17652), .S0(n108[15]), 
          .S1(n108[16]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_17.INIT0 = 16'h5555;
    defparam sub_36_add_2_17.INIT1 = 16'h5555;
    defparam sub_36_add_2_17.INJECT1_0 = "NO";
    defparam sub_36_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_36_add_2_15 (.A0(baud_counter[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17650), .COUT(n17651), .S0(n108[13]), 
          .S1(n108[14]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_15.INIT0 = 16'h5555;
    defparam sub_36_add_2_15.INIT1 = 16'h5555;
    defparam sub_36_add_2_15.INJECT1_0 = "NO";
    defparam sub_36_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_36_add_2_13 (.A0(baud_counter[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17649), .COUT(n17650), .S0(n108[11]), 
          .S1(n108[12]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_13.INIT0 = 16'h5555;
    defparam sub_36_add_2_13.INIT1 = 16'h5555;
    defparam sub_36_add_2_13.INJECT1_0 = "NO";
    defparam sub_36_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_36_add_2_11 (.A0(baud_counter[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17648), .COUT(n17649), .S0(n108[9]), .S1(n108[10]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_11.INIT0 = 16'h5555;
    defparam sub_36_add_2_11.INIT1 = 16'h5555;
    defparam sub_36_add_2_11.INJECT1_0 = "NO";
    defparam sub_36_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_36_add_2_9 (.A0(baud_counter[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17647), .COUT(n17648), .S0(n108[7]), .S1(n108[8]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_9.INIT0 = 16'h5555;
    defparam sub_36_add_2_9.INIT1 = 16'h5555;
    defparam sub_36_add_2_9.INJECT1_0 = "NO";
    defparam sub_36_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_36_add_2_7 (.A0(baud_counter[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17646), .COUT(n17647), .S0(n108[5]), .S1(n108[6]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_7.INIT0 = 16'h5555;
    defparam sub_36_add_2_7.INIT1 = 16'h5555;
    defparam sub_36_add_2_7.INJECT1_0 = "NO";
    defparam sub_36_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_36_add_2_5 (.A0(baud_counter[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17645), .COUT(n17646), .S0(n108[3]), .S1(n108[4]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_5.INIT0 = 16'h5555;
    defparam sub_36_add_2_5.INIT1 = 16'h5555;
    defparam sub_36_add_2_5.INJECT1_0 = "NO";
    defparam sub_36_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_36_add_2_3 (.A0(baud_counter[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(baud_counter[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n17644), .COUT(n17645), .S0(n108[1]), .S1(n108[2]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_3.INIT0 = 16'h5555;
    defparam sub_36_add_2_3.INIT1 = 16'h5555;
    defparam sub_36_add_2_3.INJECT1_0 = "NO";
    defparam sub_36_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_36_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(baud_counter[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n17644), .S1(n108[0]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(222[20:39])
    defparam sub_36_add_2_1.INIT0 = 16'hF000;
    defparam sub_36_add_2_1.INIT1 = 16'h5555;
    defparam sub_36_add_2_1.INJECT1_0 = "NO";
    defparam sub_36_add_2_1.INJECT1_1 = "NO";
    LUT4 i1_2_lut_4_lut (.A(state[2]), .B(n26907), .C(state[1]), .D(zero_baud_counter), 
         .Z(n11532)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(110[14:26])
    defparam i1_2_lut_4_lut.init = 16'hff80;
    LUT4 state_546_mux_6_i3_4_lut_then_4_lut (.A(n26910), .B(\state[0] ), 
         .C(state[1]), .D(state[3]), .Z(n27154)) /* synthesis lut_function=(!(A (B (C+(D))+!B (D))+!A !(((D)+!C)+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(110[14:26])
    defparam state_546_mux_6_i3_4_lut_then_4_lut.init = 16'h553f;
    LUT4 state_546_mux_6_i3_4_lut_else_4_lut (.A(n26910), .B(\state[0] ), 
         .C(state[1]), .D(state[3]), .Z(n27153)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A !(B (C+(D))+!B (C (D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(110[14:26])
    defparam state_546_mux_6_i3_4_lut_else_4_lut.init = 16'h54c0;
    LUT4 state_546_mux_6_i4_4_lut_then_4_lut (.A(n26910), .B(state[2]), 
         .C(\state[0] ), .D(state[1]), .Z(n27157)) /* synthesis lut_function=(!(A (B+(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(110[14:26])
    defparam state_546_mux_6_i4_4_lut_then_4_lut.init = 16'h5557;
    LUT4 state_546_mux_6_i4_4_lut_else_4_lut (.A(state[2]), .B(\state[0] ), 
         .C(state[1]), .Z(n27156)) /* synthesis lut_function=(A (B (C))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(110[14:26])
    defparam state_546_mux_6_i4_4_lut_else_4_lut.init = 16'h8080;
    FD1S3IX baud_counter_i23 (.D(n108[23]), .CK(dac_clk_p_c), .CD(n11532), 
            .Q(baud_counter[23])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=62, LSE_RLINE=62 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i23.GSR = "DISABLED";
    FD1S3IX baud_counter_i22 (.D(n108[22]), .CK(dac_clk_p_c), .CD(n11532), 
            .Q(baud_counter[22])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=62, LSE_RLINE=62 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i22.GSR = "DISABLED";
    FD1S3IX baud_counter_i21 (.D(n108[21]), .CK(dac_clk_p_c), .CD(n11532), 
            .Q(baud_counter[21])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=62, LSE_RLINE=62 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i21.GSR = "DISABLED";
    FD1S3IX baud_counter_i20 (.D(n108[20]), .CK(dac_clk_p_c), .CD(n11532), 
            .Q(baud_counter[20])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=62, LSE_RLINE=62 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i20.GSR = "DISABLED";
    FD1S3IX baud_counter_i19 (.D(n108[19]), .CK(dac_clk_p_c), .CD(n11532), 
            .Q(baud_counter[19])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=62, LSE_RLINE=62 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i19.GSR = "DISABLED";
    FD1S3IX baud_counter_i18 (.D(n108[18]), .CK(dac_clk_p_c), .CD(n11532), 
            .Q(baud_counter[18])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=62, LSE_RLINE=62 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i18.GSR = "DISABLED";
    FD1S3IX baud_counter_i17 (.D(n108[17]), .CK(dac_clk_p_c), .CD(n11532), 
            .Q(baud_counter[17])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=62, LSE_RLINE=62 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i17.GSR = "DISABLED";
    FD1S3IX baud_counter_i16 (.D(n108[16]), .CK(dac_clk_p_c), .CD(n11532), 
            .Q(baud_counter[16])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=62, LSE_RLINE=62 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i16.GSR = "DISABLED";
    FD1S3IX baud_counter_i15 (.D(n108[15]), .CK(dac_clk_p_c), .CD(n11532), 
            .Q(baud_counter[15])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=62, LSE_RLINE=62 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i15.GSR = "DISABLED";
    FD1S3IX baud_counter_i14 (.D(n108[14]), .CK(dac_clk_p_c), .CD(n11532), 
            .Q(baud_counter[14])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=62, LSE_RLINE=62 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i14.GSR = "DISABLED";
    FD1S3AX baud_counter_i13 (.D(baud_counter_23__N_483[13]), .CK(dac_clk_p_c), 
            .Q(baud_counter[13])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=62, LSE_RLINE=62 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i13.GSR = "DISABLED";
    FD1S3IX baud_counter_i12 (.D(n108[12]), .CK(dac_clk_p_c), .CD(n11532), 
            .Q(baud_counter[12])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=62, LSE_RLINE=62 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i12.GSR = "DISABLED";
    FD1S3IX baud_counter_i11 (.D(n108[11]), .CK(dac_clk_p_c), .CD(n11532), 
            .Q(baud_counter[11])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=62, LSE_RLINE=62 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i11.GSR = "DISABLED";
    FD1S3AX baud_counter_i10 (.D(baud_counter_23__N_483[10]), .CK(dac_clk_p_c), 
            .Q(baud_counter[10])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=62, LSE_RLINE=62 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i10.GSR = "DISABLED";
    FD1S3AX baud_counter_i9 (.D(baud_counter_23__N_483[9]), .CK(dac_clk_p_c), 
            .Q(baud_counter[9])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=62, LSE_RLINE=62 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i9.GSR = "DISABLED";
    FD1S3AX baud_counter_i8 (.D(baud_counter_23__N_483[8]), .CK(dac_clk_p_c), 
            .Q(baud_counter[8])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=62, LSE_RLINE=62 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i8.GSR = "DISABLED";
    FD1S3IX baud_counter_i7 (.D(n108[7]), .CK(dac_clk_p_c), .CD(n11532), 
            .Q(baud_counter[7])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=62, LSE_RLINE=62 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i7.GSR = "DISABLED";
    FD1S3IX baud_counter_i6 (.D(n108[6]), .CK(dac_clk_p_c), .CD(n11532), 
            .Q(baud_counter[6])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=62, LSE_RLINE=62 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i6.GSR = "DISABLED";
    FD1S3IX baud_counter_i5 (.D(n108[5]), .CK(dac_clk_p_c), .CD(n11532), 
            .Q(baud_counter[5])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=62, LSE_RLINE=62 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i5.GSR = "DISABLED";
    FD1S3IX baud_counter_i4 (.D(n108[4]), .CK(dac_clk_p_c), .CD(n11532), 
            .Q(baud_counter[4])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=62, LSE_RLINE=62 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i4.GSR = "DISABLED";
    FD1S3AX baud_counter_i3 (.D(baud_counter_23__N_483[3]), .CK(dac_clk_p_c), 
            .Q(baud_counter[3])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=62, LSE_RLINE=62 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i3.GSR = "DISABLED";
    FD1S3AX baud_counter_i2 (.D(baud_counter_23__N_483[2]), .CK(dac_clk_p_c), 
            .Q(baud_counter[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=62, LSE_RLINE=62 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i2.GSR = "DISABLED";
    FD1S3AX baud_counter_i1 (.D(baud_counter_23__N_483[1]), .CK(dac_clk_p_c), 
            .Q(baud_counter[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=62, LSE_RLINE=62 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(205[9] 225[5])
    defparam baud_counter_i1.GSR = "DISABLED";
    FD1P3IX lcl_data_i7 (.D(n29502), .SP(zero_baud_counter), .CD(n26910), 
            .CK(dac_clk_p_c), .Q(\lcl_data[7] )) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=62, LSE_RLINE=62 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(139[9] 143[40])
    defparam lcl_data_i7.GSR = "DISABLED";
    LUT4 zero_baud_counter_I_0_51_4_lut (.A(n26910), .B(n20311), .C(n26789), 
         .D(zero_baud_counter_N_528), .Z(zero_baud_counter_N_525)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C))+!A !((C+(D))+!B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(217[12] 224[43])
    defparam zero_baud_counter_I_0_51_4_lut.init = 16'h5f53;
    LUT4 i1_4_lut (.A(n20839), .B(n20847), .C(n20845), .D(n20837), .Z(n20311)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(207[24:43])
    defparam i1_4_lut.init = 16'hfffe;
    FD1P3AY lcl_data_i6 (.D(\lcl_data_7__N_511[6] ), .SP(dac_clk_p_c_enable_322), 
            .CK(dac_clk_p_c), .Q(\lcl_data[6] )) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=62, LSE_RLINE=62 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(139[9] 143[40])
    defparam lcl_data_i6.GSR = "DISABLED";
    FD1P3AY lcl_data_i5 (.D(\lcl_data_7__N_511[5] ), .SP(dac_clk_p_c_enable_322), 
            .CK(dac_clk_p_c), .Q(\lcl_data[5] )) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=62, LSE_RLINE=62 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(139[9] 143[40])
    defparam lcl_data_i5.GSR = "DISABLED";
    FD1P3AY lcl_data_i4 (.D(\lcl_data_7__N_511[4] ), .SP(dac_clk_p_c_enable_322), 
            .CK(dac_clk_p_c), .Q(\lcl_data[4] )) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=62, LSE_RLINE=62 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(139[9] 143[40])
    defparam lcl_data_i4.GSR = "DISABLED";
    FD1P3AY lcl_data_i3 (.D(\lcl_data_7__N_511[3] ), .SP(dac_clk_p_c_enable_322), 
            .CK(dac_clk_p_c), .Q(\lcl_data[3] )) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=62, LSE_RLINE=62 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(139[9] 143[40])
    defparam lcl_data_i3.GSR = "DISABLED";
    FD1P3AY lcl_data_i2 (.D(\lcl_data_7__N_511[2] ), .SP(dac_clk_p_c_enable_322), 
            .CK(dac_clk_p_c), .Q(\lcl_data[2] )) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=62, LSE_RLINE=62 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(139[9] 143[40])
    defparam lcl_data_i2.GSR = "DISABLED";
    FD1P3AY lcl_data_i1 (.D(\lcl_data_7__N_511[1] ), .SP(dac_clk_p_c_enable_322), 
            .CK(dac_clk_p_c), .Q(\lcl_data[1] )) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=62, LSE_RLINE=62 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(139[9] 143[40])
    defparam lcl_data_i1.GSR = "DISABLED";
    LUT4 baud_counter_23__I_10_i14_4_lut (.A(n26910), .B(n133[13]), .C(n26789), 
         .D(zero_baud_counter_N_528), .Z(baud_counter_23__N_483[13])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((C+(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(217[12] 224[43])
    defparam baud_counter_23__I_10_i14_4_lut.init = 16'ha0ac;
    LUT4 i11518_2_lut (.A(n108[13]), .B(zero_baud_counter), .Z(n133[13])) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(224[4:43])
    defparam i11518_2_lut.init = 16'heeee;
    LUT4 baud_counter_23__I_10_i11_4_lut (.A(n26910), .B(n133[10]), .C(n26789), 
         .D(zero_baud_counter_N_528), .Z(baud_counter_23__N_483[10])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((C+(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(217[12] 224[43])
    defparam baud_counter_23__I_10_i11_4_lut.init = 16'ha0ac;
    LUT4 i11519_2_lut (.A(n108[10]), .B(zero_baud_counter), .Z(n133[10])) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(224[4:43])
    defparam i11519_2_lut.init = 16'heeee;
    LUT4 baud_counter_23__I_10_i10_4_lut (.A(n26910), .B(n133[9]), .C(n26789), 
         .D(zero_baud_counter_N_528), .Z(baud_counter_23__N_483[9])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((C+(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(217[12] 224[43])
    defparam baud_counter_23__I_10_i10_4_lut.init = 16'ha0ac;
    LUT4 i11520_2_lut (.A(n108[9]), .B(zero_baud_counter), .Z(n133[9])) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(224[4:43])
    defparam i11520_2_lut.init = 16'heeee;
    LUT4 baud_counter_23__I_10_i9_4_lut (.A(n26910), .B(n133[8]), .C(n26789), 
         .D(zero_baud_counter_N_528), .Z(baud_counter_23__N_483[8])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((C+(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(217[12] 224[43])
    defparam baud_counter_23__I_10_i9_4_lut.init = 16'ha0ac;
    LUT4 i11521_2_lut (.A(n108[8]), .B(zero_baud_counter), .Z(n133[8])) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(224[4:43])
    defparam i11521_2_lut.init = 16'heeee;
    LUT4 baud_counter_23__I_10_i4_4_lut (.A(n26910), .B(n133[3]), .C(n26789), 
         .D(zero_baud_counter_N_528), .Z(baud_counter_23__N_483[3])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((C+(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(217[12] 224[43])
    defparam baud_counter_23__I_10_i4_4_lut.init = 16'ha0ac;
    LUT4 i11522_2_lut (.A(n108[3]), .B(zero_baud_counter), .Z(n133[3])) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(224[4:43])
    defparam i11522_2_lut.init = 16'heeee;
    LUT4 baud_counter_23__I_10_i3_4_lut (.A(n26910), .B(n133[2]), .C(n26789), 
         .D(zero_baud_counter_N_528), .Z(baud_counter_23__N_483[2])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((C+(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(217[12] 224[43])
    defparam baud_counter_23__I_10_i3_4_lut.init = 16'ha0ac;
    LUT4 i11523_2_lut (.A(n108[2]), .B(zero_baud_counter), .Z(n133[2])) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(224[4:43])
    defparam i11523_2_lut.init = 16'heeee;
    LUT4 baud_counter_23__I_10_i2_4_lut (.A(n26910), .B(n133[1]), .C(n26789), 
         .D(zero_baud_counter_N_528), .Z(baud_counter_23__N_483[1])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((C+(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(217[12] 224[43])
    defparam baud_counter_23__I_10_i2_4_lut.init = 16'ha0ac;
    LUT4 i11524_2_lut (.A(n108[1]), .B(zero_baud_counter), .Z(n133[1])) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(224[4:43])
    defparam i11524_2_lut.init = 16'heeee;
    LUT4 i1_4_lut_adj_74 (.A(baud_counter[1]), .B(baud_counter[4]), .C(baud_counter[17]), 
         .D(baud_counter[5]), .Z(n20839)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(207[24:43])
    defparam i1_4_lut_adj_74.init = 16'hfffe;
    LUT4 i1_4_lut_adj_75 (.A(n20823), .B(baud_counter[0]), .C(n20833), 
         .D(baud_counter[19]), .Z(n20847)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(207[24:43])
    defparam i1_4_lut_adj_75.init = 16'hfffb;
    LUT4 i1_4_lut_adj_76 (.A(baud_counter[22]), .B(n20835), .C(n20825), 
         .D(baud_counter[12]), .Z(n20845)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(207[24:43])
    defparam i1_4_lut_adj_76.init = 16'hfffe;
    LUT4 i1_2_lut_rep_584 (.A(\state[0] ), .B(state[3]), .Z(n26907)) /* synthesis lut_function=(A (B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(110[14:26])
    defparam i1_2_lut_rep_584.init = 16'h8888;
    LUT4 i1_3_lut_rep_466_4_lut (.A(\state[0] ), .B(state[3]), .C(state[1]), 
         .D(state[2]), .Z(n26789)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(110[14:26])
    defparam i1_3_lut_rep_466_4_lut.init = 16'h8000;
    LUT4 i1_4_lut_adj_77 (.A(baud_counter[18]), .B(baud_counter[11]), .C(baud_counter[9]), 
         .D(baud_counter[20]), .Z(n20837)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(207[24:43])
    defparam i1_4_lut_adj_77.init = 16'hfffe;
    LUT4 i1_2_lut (.A(baud_counter[8]), .B(baud_counter[6]), .Z(n20823)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(207[24:43])
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i1_4_lut_adj_78 (.A(baud_counter[13]), .B(baud_counter[23]), .C(baud_counter[3]), 
         .D(baud_counter[16]), .Z(n20833)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(207[24:43])
    defparam i1_4_lut_adj_78.init = 16'hfffe;
    LUT4 i1_4_lut_adj_79 (.A(baud_counter[7]), .B(baud_counter[2]), .C(baud_counter[15]), 
         .D(baud_counter[14]), .Z(n20835)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(207[24:43])
    defparam i1_4_lut_adj_79.init = 16'hfffe;
    LUT4 i1_2_lut_adj_80 (.A(baud_counter[21]), .B(baud_counter[10]), .Z(n20825)) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(207[24:43])
    defparam i1_2_lut_adj_80.init = 16'heeee;
    LUT4 i1_4_lut_adj_81 (.A(state[1]), .B(n26907), .C(state[2]), .D(zero_baud_counter), 
         .Z(zero_baud_counter_N_528)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_adj_81.init = 16'h0400;
    LUT4 i22622_2_lut (.A(o_busy_N_536), .B(zero_baud_counter), .Z(n8997)) /* synthesis lut_function=(!(A (B))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(97[8] 113[6])
    defparam i22622_2_lut.init = 16'h7777;
    LUT4 i732_4_lut (.A(state[2]), .B(state[3]), .C(state[1]), .D(\state[0] ), 
         .Z(o_busy_N_536)) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;
    defparam i732_4_lut.init = 16'hccc8;
    LUT4 state_546_mux_6_i2_4_lut (.A(state[1]), .B(n26910), .C(o_busy_N_536), 
         .D(\state[0] ), .Z(n27[1])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(110[14:26])
    defparam state_546_mux_6_i2_4_lut.init = 16'h353a;
    LUT4 baud_counter_23__I_10_i1_4_lut (.A(n26910), .B(n133[0]), .C(n26789), 
         .D(zero_baud_counter_N_528), .Z(baud_counter_23__N_483[0])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((C+(D))+!B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(217[12] 224[43])
    defparam baud_counter_23__I_10_i1_4_lut.init = 16'ha0ac;
    LUT4 i11002_2_lut (.A(n108[0]), .B(zero_baud_counter), .Z(n133[0])) /* synthesis lut_function=(A+(B)) */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(224[4:43])
    defparam i11002_2_lut.init = 16'heeee;
    PFUMX i24751 (.BLUT(n27156), .ALUT(n27157), .C0(state[3]), .Z(n27158));
    PFUMX i24749 (.BLUT(n27153), .ALUT(n27154), .C0(state[2]), .Z(n27155));
    FD1S3JX r_busy_45 (.D(n8997), .CK(dac_clk_p_c), .PD(n26910), .Q(tx_busy)) /* synthesis lse_init_val=1, LSE_LINE_FILE_ID=8, LSE_LCOL=58, LSE_RCOL=115, LSE_LLINE=62, LSE_RLINE=62 */ ;   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(92[9] 114[5])
    defparam r_busy_45.GSR = "DISABLED";
    FD1P3AX state_546__i3 (.D(n27158), .SP(zero_baud_counter), .CK(dac_clk_p_c), 
            .Q(state[3]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(110[14:26])
    defparam state_546__i3.GSR = "DISABLED";
    FD1P3AX state_546__i2 (.D(n27155), .SP(zero_baud_counter), .CK(dac_clk_p_c), 
            .Q(state[2]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(110[14:26])
    defparam state_546__i2.GSR = "DISABLED";
    FD1P3AX state_546__i1 (.D(n27[1]), .SP(zero_baud_counter), .CK(dac_clk_p_c), 
            .Q(state[1]));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(110[14:26])
    defparam state_546__i1.GSR = "DISABLED";
    FD1P3AX state_546__i0 (.D(n17844), .SP(zero_baud_counter), .CK(dac_clk_p_c), 
            .Q(\state[0] ));   // d:/documents/git_local/fm_modulator/rtl/debug_bus/txuartlite.v(110[14:26])
    defparam state_546__i0.GSR = "DISABLED";
    
endmodule
